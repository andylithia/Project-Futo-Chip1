* NGSPICE file created from caparray_s1.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

.subckt caparray_s1 cap_series_gygyn cap_series_gygyp cap_series_gyn cap_series_gyp
+ cap_shunt_gyn cap_shunt_gyp cap_shunt_n cap_shunt_p tune_series_gy[0] tune_series_gy[1]
+ tune_series_gy[2] tune_series_gy[3] tune_series_gy[4] tune_series_gy[5] tune_series_gygy[0]
+ tune_series_gygy[1] tune_series_gygy[2] tune_series_gygy[3] tune_series_gygy[4]
+ tune_series_gygy[5] tune_shunt[0] tune_shunt[1] tune_shunt[2] tune_shunt[3] tune_shunt[4]
+ tune_shunt[5] tune_shunt[6] tune_shunt[7] tune_shunt_gy[0] tune_shunt_gy[1] tune_shunt_gy[2]
+ tune_shunt_gy[3] tune_shunt_gy[4] tune_shunt_gy[5] tune_shunt_gy[6] vdd vss
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g1\[12\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[12\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[72\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[72\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[117\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[117\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[7\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[7\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[61\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[61\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g8\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[0] gen_shunt_g8\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gy_g1\[3\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[3\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g11\[11\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[11\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g2\[3\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[3\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[88\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[88\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[114\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[114\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[37\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[37\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g1\[20\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[20\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[71\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[71\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[116\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[116\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[39\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[39\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[60\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[60\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[87\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[87\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[113\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[113\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[3\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[3\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[36\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[36\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[70\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[70\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[5\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[5\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[89\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[89\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[115\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[115\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[38\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[38\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[86\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[86\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[112\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[112\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[35\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[35\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[3\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[3\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[88\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[88\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g4\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[114\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[114\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[37\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[37\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[85\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[85\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[111\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[111\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[18\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[18\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[34\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[34\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[87\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[87\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[113\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[113\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[36\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[36\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[5\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[5\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g2\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[84\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[84\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g3\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[26\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[26\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[110\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[110\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[33\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[33\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[86\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[86\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[112\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[112\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[35\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[35\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[83\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[83\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[32\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[32\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[13\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[13\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g3\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[3]
+ gen_shunt_gygy_g3\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[85\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[85\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[18\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[18\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[111\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[111\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[34\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[34\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g11\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[12\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[12\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[82\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[82\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g3\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[127\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[127\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[21\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[21\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[84\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[84\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g3\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[26\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[26\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[110\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[110\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[39\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[39\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[33\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[33\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[81\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[81\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[126\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[126\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[49\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[49\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[83\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[83\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[32\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[32\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[38\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[38\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[6\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[6\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_series_gy_g1\[13\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[13\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g3\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[3]
+ gen_shunt_gygy_g3\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g3\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[80\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[80\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[99\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[99\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g7\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[1] gen_shunt_g7\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[125\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[125\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[48\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[48\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[12\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[12\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[82\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[82\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g3\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[37\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[37\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[127\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[127\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[21\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[21\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[6\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[6\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[98\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[98\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g3\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[39\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[39\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g7\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[1] gen_shunt_g7\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[124\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[124\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[47\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[47\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gygy_g2\[2\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[2\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[81\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[81\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[36\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[36\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[126\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[126\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[49\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[49\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[97\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[97\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[38\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[38\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[123\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[123\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[6\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[6\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[46\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[46\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[80\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[80\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[99\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[99\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[2\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[2\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g7\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[1] gen_shunt_g7\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[35\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[35\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[125\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[125\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[48\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[48\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[96\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[96\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[37\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[37\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[122\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[122\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[45\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[45\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[6\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[6\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g4\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[98\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[98\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g7\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[1] gen_shunt_g7\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[19\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[19\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[34\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[34\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[124\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[124\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[2\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[2\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[47\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[47\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gygy_g2\[2\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[2\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g3\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[2] gen_shunt_gy_g3\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[2]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[95\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[95\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[36\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[36\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[121\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[121\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[44\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[44\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g4\[0\].u_shunt_n cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[0] gen_shunt_gy_g4\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g3\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[97\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[97\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[27\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[27\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[33\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[33\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[123\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[123\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[46\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[46\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g4\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[2\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[2\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gy_g3\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[1] gen_shunt_gy_g3\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[94\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[94\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[35\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[35\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp2 cap_series_gygyp cap_series_gygyp tune_series_gygy[1]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[120\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[120\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[4\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[4\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[43\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[43\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g3\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g4\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[96\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[96\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[32\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[32\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[122\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[122\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[45\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[45\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[14\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[14\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[93\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[93\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[19\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[19\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[34\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[34\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g1\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[2\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[2\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[42\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[42\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g3\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[2] gen_shunt_gy_g3\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp3 cap_series_gygyp cap_series_gygyp tune_series_gygy[0]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp3/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[2]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[13\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[13\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[95\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[95\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g3\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g2\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[121\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[121\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[44\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[44\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[22\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[22\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g4\[0\].u_shunt_p cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[0] gen_shunt_gy_g4\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[92\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[92\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[27\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[27\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[33\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[33\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[41\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[41\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gy_g3\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[1] gen_shunt_gy_g3\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[94\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[94\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn2 cap_series_gygyn cap_series_gygyn tune_series_gygy[1]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[120\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[120\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[4\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[4\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[3\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[3\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[43\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[43\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[49\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[49\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[30\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[30\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[91\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[91\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[32\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[32\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[14\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[14\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[40\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[40\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[59\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[59\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[93\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[93\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g1\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[42\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[42\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[48\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[48\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g11\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn3 cap_series_gygyn cap_series_gygyn tune_series_gygy[0]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn3/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[13\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[13\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[3\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[3\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g4\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[90\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[90\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[22\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[22\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[58\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[58\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[92\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[92\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[41\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[41\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[47\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[47\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g6\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[3\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[3\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g2\[49\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[49\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[30\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[30\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[57\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[57\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g2\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[91\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[91\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g5\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[0]
+ gen_series_gy_g5\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[40\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[40\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[46\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[46\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[59\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[59\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g6\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[48\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[48\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[56\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[56\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g2\[3\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[3\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[90\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[90\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g1\[5\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[5\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[45\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[45\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[58\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[58\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g6\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[47\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[47\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[55\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[55\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g6\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[8\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[8\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[44\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[44\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[57\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[57\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g1\[5\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[5\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g6\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g5\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[0]
+ gen_series_gy_g5\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[28\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[28\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g2\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[46\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[46\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[54\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[54\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g6\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[43\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[43\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[56\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[56\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[5\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[5\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[45\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[45\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[15\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[15\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[7\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[7\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[53\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[53\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[8\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[8\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[42\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[42\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[55\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[55\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[14\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[14\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[8\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[8\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[44\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[44\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[23\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[23\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[5\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[5\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[52\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[52\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gy_g1\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[28\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[28\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g3\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[2] gen_shunt_gy_g3\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g2\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[41\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[41\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[54\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[54\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g3\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[43\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[43\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[31\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[31\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[51\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[51\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[10\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[10\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[40\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[40\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[15\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[15\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[7\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[7\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[53\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[53\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[59\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[59\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g3\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[1] gen_shunt_gy_g3\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g4\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[1]
+ gen_series_gy_g4\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[3\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[3\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g1\[8\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[8\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[42\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[42\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[50\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[50\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[69\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[69\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[14\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[14\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[23\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[23\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[52\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[52\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[58\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[58\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gy_g3\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[2] gen_shunt_gy_g3\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[41\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[41\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[68\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[68\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[31\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[31\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[51\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[51\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[57\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[57\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[10\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[10\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g2\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[40\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[40\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[59\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[59\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g3\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[1] gen_shunt_gy_g3\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[67\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[67\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g4\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[1]
+ gen_series_gy_g4\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[2\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[2\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g1\[3\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[3\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[50\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[50\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[56\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[56\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[69\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[69\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[58\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[58\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[66\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[66\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g2\[2\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[2\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g2\[55\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[55\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g5\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[68\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[68\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[9\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[9\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g2\[57\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[57\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[65\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[65\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[29\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[29\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[54\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[54\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[67\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[67\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[2\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[2\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[56\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[56\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[64\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[64\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[109\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[109\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g1\[16\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[16\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[53\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[53\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[66\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[66\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[9\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[9\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[2\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[2\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g3\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[55\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[55\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g5\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g11\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[63\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[63\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[15\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[15\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[4\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[9\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[9\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[108\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[108\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[24\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[24\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[52\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[52\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g5\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[65\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[65\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[29\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[29\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[54\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[54\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[62\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[62\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[107\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[107\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[4\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[51\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[51\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[64\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[64\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[11\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[11\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g2\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[109\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[109\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[16\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[16\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[53\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[53\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[61\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[61\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g4\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[1]
+ gen_series_gy_g4\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[10\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[10\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[9\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[9\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[106\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[106\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g3\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g11\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[50\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[50\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[63\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[63\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[15\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[15\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[4\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[108\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[108\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gygy_g1\[6\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[6\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[24\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[24\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[52\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[52\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[60\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[60\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[79\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[79\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[105\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[105\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[62\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[62\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[107\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[107\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[4\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[51\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[51\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[11\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[11\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[78\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[78\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g2\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[104\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[104\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[61\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[61\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g4\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[1]
+ gen_series_gy_g4\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[10\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[10\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[106\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[106\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[50\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[50\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[77\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[77\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[6\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[6\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g4\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[103\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[103\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[60\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[60\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[2\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[2\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[79\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[79\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[105\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[105\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[76\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[76\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[102\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[102\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g2\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[78\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[78\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[104\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[104\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g3\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[3]
+ gen_shunt_gygy_g3\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[75\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[75\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[101\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[101\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[77\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[77\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[103\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[103\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[17\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[17\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g2\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g1\[2\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[2\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[74\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[74\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[100\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[100\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[119\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[119\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[63\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[63\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[76\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[76\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g2\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[102\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[102\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[25\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[25\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[73\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[73\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[7\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[7\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g3\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[3]
+ gen_shunt_gygy_g3\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[118\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[118\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[62\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[62\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[75\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[75\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[101\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[101\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[12\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[12\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[72\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[72\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[17\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[17\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[117\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[117\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_gy_g1\[7\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[7\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[61\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[61\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g8\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[0] gen_shunt_g8\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[74\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[74\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g11\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[11\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[11\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[3\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[3\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[100\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[100\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[119\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[119\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[63\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[63\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[20\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[20\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[71\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[71\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[25\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[25\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[116\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[116\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[39\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[39\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[60\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[60\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[73\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[73\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[7\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[7\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[118\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[118\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[3\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[3\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[62\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[62\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[70\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[70\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[89\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[89\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[115\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[115\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[38\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[38\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

