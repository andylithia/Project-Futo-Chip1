magic
tech gf180mcuC
magscale 1 5
timestamp 1670013959
<< obsm1 >>
rect 672 1538 6408 6302
<< obsm2 >>
rect 910 1549 6394 6291
<< metal3 >>
rect 0 3976 400 4032
<< obsm3 >>
rect 400 4062 6399 6286
rect 430 3946 6399 4062
rect 400 1554 6399 3946
<< metal4 >>
rect 1299 1538 1459 6302
rect 2006 1538 2166 6302
rect 2713 1538 2873 6302
rect 3420 1538 3580 6302
rect 4127 1538 4287 6302
rect 4834 1538 4994 6302
rect 5541 1538 5701 6302
rect 6248 1538 6408 6302
<< labels >>
rlabel metal3 s 0 3976 400 4032 6 Y
port 1 nsew signal output
rlabel metal4 s 1299 1538 1459 6302 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 2713 1538 2873 6302 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 4127 1538 4287 6302 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 5541 1538 5701 6302 6 vdd
port 2 nsew power bidirectional
rlabel metal4 s 2006 1538 2166 6302 6 vss
port 3 nsew ground bidirectional
rlabel metal4 s 3420 1538 3580 6302 6 vss
port 3 nsew ground bidirectional
rlabel metal4 s 4834 1538 4994 6302 6 vss
port 3 nsew ground bidirectional
rlabel metal4 s 6248 1538 6408 6302 6 vss
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 186934
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/ringosc/runs/22_12_02_15_45/results/signoff/ringosc.magic.gds
string GDS_START 31626
<< end >>

