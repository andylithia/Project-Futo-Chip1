VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caparray_s2
  CLASS BLOCK ;
  FOREIGN caparray_s2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 200.000 ;
  PIN cap_series_gygyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 196.000 374.640 200.000 ;
    END
  END cap_series_gygyn
  PIN cap_series_gygyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.240 196.000 324.800 200.000 ;
    END
  END cap_series_gygyp
  PIN cap_series_gyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 196.000 274.960 200.000 ;
    END
  END cap_series_gyn
  PIN cap_series_gyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.560 196.000 225.120 200.000 ;
    END
  END cap_series_gyp
  PIN cap_shunt_gyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 196.000 175.280 200.000 ;
    END
  END cap_shunt_gyn
  PIN cap_shunt_gyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.880 196.000 125.440 200.000 ;
    END
  END cap_shunt_gyp
  PIN cap_shunt_n
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 196.000 75.600 200.000 ;
    END
  END cap_shunt_n
  PIN cap_shunt_p
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.200 196.000 25.760 200.000 ;
    END
  END cap_shunt_p
  PIN tune_series_gy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.920 0.000 144.480 4.000 ;
    END
  END tune_series_gy[0]
  PIN tune_series_gy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.240 0.000 156.800 4.000 ;
    END
  END tune_series_gy[1]
  PIN tune_series_gy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.560 0.000 169.120 4.000 ;
    END
  END tune_series_gy[2]
  PIN tune_series_gy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.880 0.000 181.440 4.000 ;
    END
  END tune_series_gy[3]
  PIN tune_series_gy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.200 0.000 193.760 4.000 ;
    END
  END tune_series_gy[4]
  PIN tune_series_gy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.520 0.000 206.080 4.000 ;
    END
  END tune_series_gy[5]
  PIN tune_series_gy[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.840 0.000 218.400 4.000 ;
    END
  END tune_series_gy[6]
  PIN tune_series_gy[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.160 0.000 230.720 4.000 ;
    END
  END tune_series_gy[7]
  PIN tune_series_gygy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 242.480 0.000 243.040 4.000 ;
    END
  END tune_series_gygy[0]
  PIN tune_series_gygy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 0.000 255.360 4.000 ;
    END
  END tune_series_gygy[1]
  PIN tune_series_gygy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.120 0.000 267.680 4.000 ;
    END
  END tune_series_gygy[2]
  PIN tune_series_gygy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 0.000 280.000 4.000 ;
    END
  END tune_series_gygy[3]
  PIN tune_series_gygy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 0.000 292.320 4.000 ;
    END
  END tune_series_gygy[4]
  PIN tune_series_gygy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.080 0.000 304.640 4.000 ;
    END
  END tune_series_gygy[5]
  PIN tune_series_gygy[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.400 0.000 316.960 4.000 ;
    END
  END tune_series_gygy[6]
  PIN tune_series_gygy[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 0.000 329.280 4.000 ;
    END
  END tune_series_gygy[7]
  PIN tune_shunt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.400 0.000 8.960 4.000 ;
    END
  END tune_shunt[0]
  PIN tune_shunt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 0.000 132.160 4.000 ;
    END
  END tune_shunt[10]
  PIN tune_shunt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.720 0.000 21.280 4.000 ;
    END
  END tune_shunt[1]
  PIN tune_shunt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.040 0.000 33.600 4.000 ;
    END
  END tune_shunt[2]
  PIN tune_shunt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 0.000 45.920 4.000 ;
    END
  END tune_shunt[3]
  PIN tune_shunt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 0.000 58.240 4.000 ;
    END
  END tune_shunt[4]
  PIN tune_shunt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 0.000 70.560 4.000 ;
    END
  END tune_shunt[5]
  PIN tune_shunt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.320 0.000 82.880 4.000 ;
    END
  END tune_shunt[6]
  PIN tune_shunt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.640 0.000 95.200 4.000 ;
    END
  END tune_shunt[7]
  PIN tune_shunt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.960 0.000 107.520 4.000 ;
    END
  END tune_shunt[8]
  PIN tune_shunt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.280 0.000 119.840 4.000 ;
    END
  END tune_shunt[9]
  PIN tune_shunt_gy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.040 0.000 341.600 4.000 ;
    END
  END tune_shunt_gy[0]
  PIN tune_shunt_gy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.360 0.000 353.920 4.000 ;
    END
  END tune_shunt_gy[1]
  PIN tune_shunt_gy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.680 0.000 366.240 4.000 ;
    END
  END tune_shunt_gy[2]
  PIN tune_shunt_gy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.000 0.000 378.560 4.000 ;
    END
  END tune_shunt_gy[3]
  PIN tune_shunt_gy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.320 0.000 390.880 4.000 ;
    END
  END tune_shunt_gy[4]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 20.540 15.380 25.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.540 15.380 75.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 120.540 15.380 125.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 170.540 15.380 175.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 220.540 15.380 225.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 270.540 15.380 275.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 320.540 15.380 325.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.540 15.380 375.540 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 45.540 15.380 50.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 95.540 15.380 100.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.540 15.380 150.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.540 15.380 200.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 245.540 15.380 250.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 295.540 15.380 300.540 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 345.540 15.380 350.540 184.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 393.120 184.540 ;
      LAYER Metal2 ;
        RECT 8.540 195.700 24.900 196.420 ;
        RECT 26.060 195.700 74.740 196.420 ;
        RECT 75.900 195.700 124.580 196.420 ;
        RECT 125.740 195.700 174.420 196.420 ;
        RECT 175.580 195.700 224.260 196.420 ;
        RECT 225.420 195.700 274.100 196.420 ;
        RECT 275.260 195.700 323.940 196.420 ;
        RECT 325.100 195.700 373.780 196.420 ;
        RECT 374.940 195.700 391.300 196.420 ;
        RECT 8.540 4.300 391.300 195.700 ;
        RECT 9.260 3.500 20.420 4.300 ;
        RECT 21.580 3.500 32.740 4.300 ;
        RECT 33.900 3.500 45.060 4.300 ;
        RECT 46.220 3.500 57.380 4.300 ;
        RECT 58.540 3.500 69.700 4.300 ;
        RECT 70.860 3.500 82.020 4.300 ;
        RECT 83.180 3.500 94.340 4.300 ;
        RECT 95.500 3.500 106.660 4.300 ;
        RECT 107.820 3.500 118.980 4.300 ;
        RECT 120.140 3.500 131.300 4.300 ;
        RECT 132.460 3.500 143.620 4.300 ;
        RECT 144.780 3.500 155.940 4.300 ;
        RECT 157.100 3.500 168.260 4.300 ;
        RECT 169.420 3.500 180.580 4.300 ;
        RECT 181.740 3.500 192.900 4.300 ;
        RECT 194.060 3.500 205.220 4.300 ;
        RECT 206.380 3.500 217.540 4.300 ;
        RECT 218.700 3.500 229.860 4.300 ;
        RECT 231.020 3.500 242.180 4.300 ;
        RECT 243.340 3.500 254.500 4.300 ;
        RECT 255.660 3.500 266.820 4.300 ;
        RECT 267.980 3.500 279.140 4.300 ;
        RECT 280.300 3.500 291.460 4.300 ;
        RECT 292.620 3.500 303.780 4.300 ;
        RECT 304.940 3.500 316.100 4.300 ;
        RECT 317.260 3.500 328.420 4.300 ;
        RECT 329.580 3.500 340.740 4.300 ;
        RECT 341.900 3.500 353.060 4.300 ;
        RECT 354.220 3.500 365.380 4.300 ;
        RECT 366.540 3.500 377.700 4.300 ;
        RECT 378.860 3.500 390.020 4.300 ;
        RECT 391.180 3.500 391.300 4.300 ;
      LAYER Metal3 ;
        RECT 11.850 15.540 391.350 184.380 ;
      LAYER Metal4 ;
        RECT 319.900 21.930 320.240 44.710 ;
        RECT 325.840 21.930 345.240 44.710 ;
        RECT 350.840 21.930 369.460 44.710 ;
  END
END caparray_s2
END LIBRARY

