module caparray_s1 (cap_series_gygyn,
    cap_series_gygyp,
    cap_series_gyn,
    cap_series_gyp,
    cap_shunt_gyn,
    cap_shunt_gyp,
    cap_shunt_n,
    cap_shunt_p,
    vdd,
    vss,
    tune_series_gy,
    tune_series_gygy,
    tune_shunt,
    tune_shunt_gy);
 inout cap_series_gygyn;
 inout cap_series_gygyp;
 inout cap_series_gyn;
 inout cap_series_gyp;
 inout cap_shunt_gyn;
 inout cap_shunt_gyp;
 inout cap_shunt_n;
 inout cap_shunt_p;
 input vdd;
 input vss;
 input [5:0] tune_series_gy;
 input [5:0] tune_series_gygy;
 input [7:0] tune_shunt;
 input [6:0] tune_shunt_gy;

 wire \gen_series_gy_g1[0].d1 ;
 wire \gen_series_gy_g1[0].d2 ;
 wire \gen_series_gy_g1[0].d3 ;
 wire \gen_series_gy_g1[0].d4 ;
 wire \gen_series_gy_g1[10].d1 ;
 wire \gen_series_gy_g1[10].d2 ;
 wire \gen_series_gy_g1[10].d3 ;
 wire \gen_series_gy_g1[10].d4 ;
 wire \gen_series_gy_g1[11].d1 ;
 wire \gen_series_gy_g1[11].d2 ;
 wire \gen_series_gy_g1[11].d3 ;
 wire \gen_series_gy_g1[11].d4 ;
 wire \gen_series_gy_g1[12].d1 ;
 wire \gen_series_gy_g1[12].d2 ;
 wire \gen_series_gy_g1[12].d3 ;
 wire \gen_series_gy_g1[12].d4 ;
 wire \gen_series_gy_g1[13].d1 ;
 wire \gen_series_gy_g1[13].d2 ;
 wire \gen_series_gy_g1[13].d3 ;
 wire \gen_series_gy_g1[13].d4 ;
 wire \gen_series_gy_g1[14].d1 ;
 wire \gen_series_gy_g1[14].d2 ;
 wire \gen_series_gy_g1[14].d3 ;
 wire \gen_series_gy_g1[14].d4 ;
 wire \gen_series_gy_g1[15].d1 ;
 wire \gen_series_gy_g1[15].d2 ;
 wire \gen_series_gy_g1[15].d3 ;
 wire \gen_series_gy_g1[15].d4 ;
 wire \gen_series_gy_g1[1].d1 ;
 wire \gen_series_gy_g1[1].d2 ;
 wire \gen_series_gy_g1[1].d3 ;
 wire \gen_series_gy_g1[1].d4 ;
 wire \gen_series_gy_g1[2].d1 ;
 wire \gen_series_gy_g1[2].d2 ;
 wire \gen_series_gy_g1[2].d3 ;
 wire \gen_series_gy_g1[2].d4 ;
 wire \gen_series_gy_g1[3].d1 ;
 wire \gen_series_gy_g1[3].d2 ;
 wire \gen_series_gy_g1[3].d3 ;
 wire \gen_series_gy_g1[3].d4 ;
 wire \gen_series_gy_g1[4].d1 ;
 wire \gen_series_gy_g1[4].d2 ;
 wire \gen_series_gy_g1[4].d3 ;
 wire \gen_series_gy_g1[4].d4 ;
 wire \gen_series_gy_g1[5].d1 ;
 wire \gen_series_gy_g1[5].d2 ;
 wire \gen_series_gy_g1[5].d3 ;
 wire \gen_series_gy_g1[5].d4 ;
 wire \gen_series_gy_g1[6].d1 ;
 wire \gen_series_gy_g1[6].d2 ;
 wire \gen_series_gy_g1[6].d3 ;
 wire \gen_series_gy_g1[6].d4 ;
 wire \gen_series_gy_g1[7].d1 ;
 wire \gen_series_gy_g1[7].d2 ;
 wire \gen_series_gy_g1[7].d3 ;
 wire \gen_series_gy_g1[7].d4 ;
 wire \gen_series_gy_g1[8].d1 ;
 wire \gen_series_gy_g1[8].d2 ;
 wire \gen_series_gy_g1[8].d3 ;
 wire \gen_series_gy_g1[8].d4 ;
 wire \gen_series_gy_g1[9].d1 ;
 wire \gen_series_gy_g1[9].d2 ;
 wire \gen_series_gy_g1[9].d3 ;
 wire \gen_series_gy_g1[9].d4 ;
 wire \gen_series_gy_g2[0].d1 ;
 wire \gen_series_gy_g2[0].d2 ;
 wire \gen_series_gy_g2[1].d1 ;
 wire \gen_series_gy_g2[1].d2 ;
 wire \gen_series_gy_g2[2].d1 ;
 wire \gen_series_gy_g2[2].d2 ;
 wire \gen_series_gy_g2[3].d1 ;
 wire \gen_series_gy_g2[3].d2 ;
 wire \gen_series_gy_g2[4].d1 ;
 wire \gen_series_gy_g2[4].d2 ;
 wire \gen_series_gy_g2[5].d1 ;
 wire \gen_series_gy_g2[5].d2 ;
 wire \gen_series_gy_g2[6].d1 ;
 wire \gen_series_gy_g2[6].d2 ;
 wire \gen_series_gy_g2[7].d1 ;
 wire \gen_series_gy_g2[7].d2 ;
 wire \gen_series_gy_g3[0].d1 ;
 wire \gen_series_gy_g3[0].d2 ;
 wire \gen_series_gy_g3[1].d1 ;
 wire \gen_series_gy_g3[1].d2 ;
 wire \gen_series_gy_g3[2].d1 ;
 wire \gen_series_gy_g3[2].d2 ;
 wire \gen_series_gy_g3[3].d1 ;
 wire \gen_series_gy_g3[3].d2 ;
 wire \gen_series_gy_g4[0].d1 ;
 wire \gen_series_gy_g4[0].d2 ;
 wire \gen_series_gy_g4[1].d1 ;
 wire \gen_series_gy_g4[1].d2 ;
 wire \gen_series_gy_g5[0].d1 ;
 wire \gen_series_gy_g5[0].d2 ;
 wire \gen_shunt_g1[0].d1 ;
 wire \gen_shunt_g1[0].d2 ;
 wire \gen_shunt_g1[10].d1 ;
 wire \gen_shunt_g1[10].d2 ;
 wire \gen_shunt_g1[11].d1 ;
 wire \gen_shunt_g1[11].d2 ;
 wire \gen_shunt_g1[12].d1 ;
 wire \gen_shunt_g1[12].d2 ;
 wire \gen_shunt_g1[13].d1 ;
 wire \gen_shunt_g1[13].d2 ;
 wire \gen_shunt_g1[14].d1 ;
 wire \gen_shunt_g1[14].d2 ;
 wire \gen_shunt_g1[15].d1 ;
 wire \gen_shunt_g1[15].d2 ;
 wire \gen_shunt_g1[16].d1 ;
 wire \gen_shunt_g1[16].d2 ;
 wire \gen_shunt_g1[17].d1 ;
 wire \gen_shunt_g1[17].d2 ;
 wire \gen_shunt_g1[18].d1 ;
 wire \gen_shunt_g1[18].d2 ;
 wire \gen_shunt_g1[19].d1 ;
 wire \gen_shunt_g1[19].d2 ;
 wire \gen_shunt_g1[1].d1 ;
 wire \gen_shunt_g1[1].d2 ;
 wire \gen_shunt_g1[20].d1 ;
 wire \gen_shunt_g1[20].d2 ;
 wire \gen_shunt_g1[21].d1 ;
 wire \gen_shunt_g1[21].d2 ;
 wire \gen_shunt_g1[22].d1 ;
 wire \gen_shunt_g1[22].d2 ;
 wire \gen_shunt_g1[23].d1 ;
 wire \gen_shunt_g1[23].d2 ;
 wire \gen_shunt_g1[24].d1 ;
 wire \gen_shunt_g1[24].d2 ;
 wire \gen_shunt_g1[25].d1 ;
 wire \gen_shunt_g1[25].d2 ;
 wire \gen_shunt_g1[26].d1 ;
 wire \gen_shunt_g1[26].d2 ;
 wire \gen_shunt_g1[27].d1 ;
 wire \gen_shunt_g1[27].d2 ;
 wire \gen_shunt_g1[28].d1 ;
 wire \gen_shunt_g1[28].d2 ;
 wire \gen_shunt_g1[29].d1 ;
 wire \gen_shunt_g1[29].d2 ;
 wire \gen_shunt_g1[2].d1 ;
 wire \gen_shunt_g1[2].d2 ;
 wire \gen_shunt_g1[30].d1 ;
 wire \gen_shunt_g1[30].d2 ;
 wire \gen_shunt_g1[31].d1 ;
 wire \gen_shunt_g1[31].d2 ;
 wire \gen_shunt_g1[32].d1 ;
 wire \gen_shunt_g1[32].d2 ;
 wire \gen_shunt_g1[33].d1 ;
 wire \gen_shunt_g1[33].d2 ;
 wire \gen_shunt_g1[34].d1 ;
 wire \gen_shunt_g1[34].d2 ;
 wire \gen_shunt_g1[35].d1 ;
 wire \gen_shunt_g1[35].d2 ;
 wire \gen_shunt_g1[36].d1 ;
 wire \gen_shunt_g1[36].d2 ;
 wire \gen_shunt_g1[37].d1 ;
 wire \gen_shunt_g1[37].d2 ;
 wire \gen_shunt_g1[38].d1 ;
 wire \gen_shunt_g1[38].d2 ;
 wire \gen_shunt_g1[39].d1 ;
 wire \gen_shunt_g1[39].d2 ;
 wire \gen_shunt_g1[3].d1 ;
 wire \gen_shunt_g1[3].d2 ;
 wire \gen_shunt_g1[40].d1 ;
 wire \gen_shunt_g1[40].d2 ;
 wire \gen_shunt_g1[41].d1 ;
 wire \gen_shunt_g1[41].d2 ;
 wire \gen_shunt_g1[42].d1 ;
 wire \gen_shunt_g1[42].d2 ;
 wire \gen_shunt_g1[43].d1 ;
 wire \gen_shunt_g1[43].d2 ;
 wire \gen_shunt_g1[44].d1 ;
 wire \gen_shunt_g1[44].d2 ;
 wire \gen_shunt_g1[45].d1 ;
 wire \gen_shunt_g1[45].d2 ;
 wire \gen_shunt_g1[46].d1 ;
 wire \gen_shunt_g1[46].d2 ;
 wire \gen_shunt_g1[47].d1 ;
 wire \gen_shunt_g1[47].d2 ;
 wire \gen_shunt_g1[48].d1 ;
 wire \gen_shunt_g1[48].d2 ;
 wire \gen_shunt_g1[49].d1 ;
 wire \gen_shunt_g1[49].d2 ;
 wire \gen_shunt_g1[4].d1 ;
 wire \gen_shunt_g1[4].d2 ;
 wire \gen_shunt_g1[50].d1 ;
 wire \gen_shunt_g1[50].d2 ;
 wire \gen_shunt_g1[51].d1 ;
 wire \gen_shunt_g1[51].d2 ;
 wire \gen_shunt_g1[52].d1 ;
 wire \gen_shunt_g1[52].d2 ;
 wire \gen_shunt_g1[53].d1 ;
 wire \gen_shunt_g1[53].d2 ;
 wire \gen_shunt_g1[54].d1 ;
 wire \gen_shunt_g1[54].d2 ;
 wire \gen_shunt_g1[55].d1 ;
 wire \gen_shunt_g1[55].d2 ;
 wire \gen_shunt_g1[56].d1 ;
 wire \gen_shunt_g1[56].d2 ;
 wire \gen_shunt_g1[57].d1 ;
 wire \gen_shunt_g1[57].d2 ;
 wire \gen_shunt_g1[58].d1 ;
 wire \gen_shunt_g1[58].d2 ;
 wire \gen_shunt_g1[59].d1 ;
 wire \gen_shunt_g1[59].d2 ;
 wire \gen_shunt_g1[5].d1 ;
 wire \gen_shunt_g1[5].d2 ;
 wire \gen_shunt_g1[60].d1 ;
 wire \gen_shunt_g1[60].d2 ;
 wire \gen_shunt_g1[61].d1 ;
 wire \gen_shunt_g1[61].d2 ;
 wire \gen_shunt_g1[62].d1 ;
 wire \gen_shunt_g1[62].d2 ;
 wire \gen_shunt_g1[63].d1 ;
 wire \gen_shunt_g1[63].d2 ;
 wire \gen_shunt_g1[64].d1 ;
 wire \gen_shunt_g1[64].d2 ;
 wire \gen_shunt_g1[65].d1 ;
 wire \gen_shunt_g1[65].d2 ;
 wire \gen_shunt_g1[66].d1 ;
 wire \gen_shunt_g1[66].d2 ;
 wire \gen_shunt_g1[67].d1 ;
 wire \gen_shunt_g1[67].d2 ;
 wire \gen_shunt_g1[68].d1 ;
 wire \gen_shunt_g1[68].d2 ;
 wire \gen_shunt_g1[69].d1 ;
 wire \gen_shunt_g1[69].d2 ;
 wire \gen_shunt_g1[6].d1 ;
 wire \gen_shunt_g1[6].d2 ;
 wire \gen_shunt_g1[70].d1 ;
 wire \gen_shunt_g1[70].d2 ;
 wire \gen_shunt_g1[71].d1 ;
 wire \gen_shunt_g1[71].d2 ;
 wire \gen_shunt_g1[72].d1 ;
 wire \gen_shunt_g1[72].d2 ;
 wire \gen_shunt_g1[73].d1 ;
 wire \gen_shunt_g1[73].d2 ;
 wire \gen_shunt_g1[74].d1 ;
 wire \gen_shunt_g1[74].d2 ;
 wire \gen_shunt_g1[75].d1 ;
 wire \gen_shunt_g1[75].d2 ;
 wire \gen_shunt_g1[76].d1 ;
 wire \gen_shunt_g1[76].d2 ;
 wire \gen_shunt_g1[77].d1 ;
 wire \gen_shunt_g1[77].d2 ;
 wire \gen_shunt_g1[78].d1 ;
 wire \gen_shunt_g1[78].d2 ;
 wire \gen_shunt_g1[79].d1 ;
 wire \gen_shunt_g1[79].d2 ;
 wire \gen_shunt_g1[7].d1 ;
 wire \gen_shunt_g1[7].d2 ;
 wire \gen_shunt_g1[80].d1 ;
 wire \gen_shunt_g1[80].d2 ;
 wire \gen_shunt_g1[81].d1 ;
 wire \gen_shunt_g1[81].d2 ;
 wire \gen_shunt_g1[82].d1 ;
 wire \gen_shunt_g1[82].d2 ;
 wire \gen_shunt_g1[83].d1 ;
 wire \gen_shunt_g1[83].d2 ;
 wire \gen_shunt_g1[84].d1 ;
 wire \gen_shunt_g1[84].d2 ;
 wire \gen_shunt_g1[85].d1 ;
 wire \gen_shunt_g1[85].d2 ;
 wire \gen_shunt_g1[86].d1 ;
 wire \gen_shunt_g1[86].d2 ;
 wire \gen_shunt_g1[87].d1 ;
 wire \gen_shunt_g1[87].d2 ;
 wire \gen_shunt_g1[88].d1 ;
 wire \gen_shunt_g1[88].d2 ;
 wire \gen_shunt_g1[89].d1 ;
 wire \gen_shunt_g1[89].d2 ;
 wire \gen_shunt_g1[8].d1 ;
 wire \gen_shunt_g1[8].d2 ;
 wire \gen_shunt_g1[90].d1 ;
 wire \gen_shunt_g1[90].d2 ;
 wire \gen_shunt_g1[91].d1 ;
 wire \gen_shunt_g1[91].d2 ;
 wire \gen_shunt_g1[92].d1 ;
 wire \gen_shunt_g1[92].d2 ;
 wire \gen_shunt_g1[93].d1 ;
 wire \gen_shunt_g1[93].d2 ;
 wire \gen_shunt_g1[94].d1 ;
 wire \gen_shunt_g1[94].d2 ;
 wire \gen_shunt_g1[95].d1 ;
 wire \gen_shunt_g1[95].d2 ;
 wire \gen_shunt_g1[9].d1 ;
 wire \gen_shunt_g1[9].d2 ;
 wire \gen_shunt_g2[0].d1 ;
 wire \gen_shunt_g2[0].d2 ;
 wire \gen_shunt_g2[10].d1 ;
 wire \gen_shunt_g2[10].d2 ;
 wire \gen_shunt_g2[11].d1 ;
 wire \gen_shunt_g2[11].d2 ;
 wire \gen_shunt_g2[12].d1 ;
 wire \gen_shunt_g2[12].d2 ;
 wire \gen_shunt_g2[13].d1 ;
 wire \gen_shunt_g2[13].d2 ;
 wire \gen_shunt_g2[14].d1 ;
 wire \gen_shunt_g2[14].d2 ;
 wire \gen_shunt_g2[15].d1 ;
 wire \gen_shunt_g2[15].d2 ;
 wire \gen_shunt_g2[16].d1 ;
 wire \gen_shunt_g2[16].d2 ;
 wire \gen_shunt_g2[17].d1 ;
 wire \gen_shunt_g2[17].d2 ;
 wire \gen_shunt_g2[18].d1 ;
 wire \gen_shunt_g2[18].d2 ;
 wire \gen_shunt_g2[19].d1 ;
 wire \gen_shunt_g2[19].d2 ;
 wire \gen_shunt_g2[1].d1 ;
 wire \gen_shunt_g2[1].d2 ;
 wire \gen_shunt_g2[20].d1 ;
 wire \gen_shunt_g2[20].d2 ;
 wire \gen_shunt_g2[21].d1 ;
 wire \gen_shunt_g2[21].d2 ;
 wire \gen_shunt_g2[22].d1 ;
 wire \gen_shunt_g2[22].d2 ;
 wire \gen_shunt_g2[23].d1 ;
 wire \gen_shunt_g2[23].d2 ;
 wire \gen_shunt_g2[24].d1 ;
 wire \gen_shunt_g2[24].d2 ;
 wire \gen_shunt_g2[25].d1 ;
 wire \gen_shunt_g2[25].d2 ;
 wire \gen_shunt_g2[26].d1 ;
 wire \gen_shunt_g2[26].d2 ;
 wire \gen_shunt_g2[27].d1 ;
 wire \gen_shunt_g2[27].d2 ;
 wire \gen_shunt_g2[28].d1 ;
 wire \gen_shunt_g2[28].d2 ;
 wire \gen_shunt_g2[29].d1 ;
 wire \gen_shunt_g2[29].d2 ;
 wire \gen_shunt_g2[2].d1 ;
 wire \gen_shunt_g2[2].d2 ;
 wire \gen_shunt_g2[30].d1 ;
 wire \gen_shunt_g2[30].d2 ;
 wire \gen_shunt_g2[31].d1 ;
 wire \gen_shunt_g2[31].d2 ;
 wire \gen_shunt_g2[32].d1 ;
 wire \gen_shunt_g2[32].d2 ;
 wire \gen_shunt_g2[33].d1 ;
 wire \gen_shunt_g2[33].d2 ;
 wire \gen_shunt_g2[34].d1 ;
 wire \gen_shunt_g2[34].d2 ;
 wire \gen_shunt_g2[35].d1 ;
 wire \gen_shunt_g2[35].d2 ;
 wire \gen_shunt_g2[36].d1 ;
 wire \gen_shunt_g2[36].d2 ;
 wire \gen_shunt_g2[37].d1 ;
 wire \gen_shunt_g2[37].d2 ;
 wire \gen_shunt_g2[38].d1 ;
 wire \gen_shunt_g2[38].d2 ;
 wire \gen_shunt_g2[39].d1 ;
 wire \gen_shunt_g2[39].d2 ;
 wire \gen_shunt_g2[3].d1 ;
 wire \gen_shunt_g2[3].d2 ;
 wire \gen_shunt_g2[40].d1 ;
 wire \gen_shunt_g2[40].d2 ;
 wire \gen_shunt_g2[41].d1 ;
 wire \gen_shunt_g2[41].d2 ;
 wire \gen_shunt_g2[42].d1 ;
 wire \gen_shunt_g2[42].d2 ;
 wire \gen_shunt_g2[43].d1 ;
 wire \gen_shunt_g2[43].d2 ;
 wire \gen_shunt_g2[44].d1 ;
 wire \gen_shunt_g2[44].d2 ;
 wire \gen_shunt_g2[45].d1 ;
 wire \gen_shunt_g2[45].d2 ;
 wire \gen_shunt_g2[46].d1 ;
 wire \gen_shunt_g2[46].d2 ;
 wire \gen_shunt_g2[47].d1 ;
 wire \gen_shunt_g2[47].d2 ;
 wire \gen_shunt_g2[4].d1 ;
 wire \gen_shunt_g2[4].d2 ;
 wire \gen_shunt_g2[5].d1 ;
 wire \gen_shunt_g2[5].d2 ;
 wire \gen_shunt_g2[6].d1 ;
 wire \gen_shunt_g2[6].d2 ;
 wire \gen_shunt_g2[7].d1 ;
 wire \gen_shunt_g2[7].d2 ;
 wire \gen_shunt_g2[8].d1 ;
 wire \gen_shunt_g2[8].d2 ;
 wire \gen_shunt_g2[9].d1 ;
 wire \gen_shunt_g2[9].d2 ;
 wire \gen_shunt_g3[0].d1 ;
 wire \gen_shunt_g3[0].d2 ;
 wire \gen_shunt_g3[10].d1 ;
 wire \gen_shunt_g3[10].d2 ;
 wire \gen_shunt_g3[11].d1 ;
 wire \gen_shunt_g3[11].d2 ;
 wire \gen_shunt_g3[12].d1 ;
 wire \gen_shunt_g3[12].d2 ;
 wire \gen_shunt_g3[13].d1 ;
 wire \gen_shunt_g3[13].d2 ;
 wire \gen_shunt_g3[14].d1 ;
 wire \gen_shunt_g3[14].d2 ;
 wire \gen_shunt_g3[15].d1 ;
 wire \gen_shunt_g3[15].d2 ;
 wire \gen_shunt_g3[16].d1 ;
 wire \gen_shunt_g3[16].d2 ;
 wire \gen_shunt_g3[17].d1 ;
 wire \gen_shunt_g3[17].d2 ;
 wire \gen_shunt_g3[18].d1 ;
 wire \gen_shunt_g3[18].d2 ;
 wire \gen_shunt_g3[19].d1 ;
 wire \gen_shunt_g3[19].d2 ;
 wire \gen_shunt_g3[1].d1 ;
 wire \gen_shunt_g3[1].d2 ;
 wire \gen_shunt_g3[20].d1 ;
 wire \gen_shunt_g3[20].d2 ;
 wire \gen_shunt_g3[21].d1 ;
 wire \gen_shunt_g3[21].d2 ;
 wire \gen_shunt_g3[22].d1 ;
 wire \gen_shunt_g3[22].d2 ;
 wire \gen_shunt_g3[23].d1 ;
 wire \gen_shunt_g3[23].d2 ;
 wire \gen_shunt_g3[2].d1 ;
 wire \gen_shunt_g3[2].d2 ;
 wire \gen_shunt_g3[3].d1 ;
 wire \gen_shunt_g3[3].d2 ;
 wire \gen_shunt_g3[4].d1 ;
 wire \gen_shunt_g3[4].d2 ;
 wire \gen_shunt_g3[5].d1 ;
 wire \gen_shunt_g3[5].d2 ;
 wire \gen_shunt_g3[6].d1 ;
 wire \gen_shunt_g3[6].d2 ;
 wire \gen_shunt_g3[7].d1 ;
 wire \gen_shunt_g3[7].d2 ;
 wire \gen_shunt_g3[8].d1 ;
 wire \gen_shunt_g3[8].d2 ;
 wire \gen_shunt_g3[9].d1 ;
 wire \gen_shunt_g3[9].d2 ;
 wire \gen_shunt_g4[0].d1 ;
 wire \gen_shunt_g4[0].d2 ;
 wire \gen_shunt_g4[10].d1 ;
 wire \gen_shunt_g4[10].d2 ;
 wire \gen_shunt_g4[11].d1 ;
 wire \gen_shunt_g4[11].d2 ;
 wire \gen_shunt_g4[1].d1 ;
 wire \gen_shunt_g4[1].d2 ;
 wire \gen_shunt_g4[2].d1 ;
 wire \gen_shunt_g4[2].d2 ;
 wire \gen_shunt_g4[3].d1 ;
 wire \gen_shunt_g4[3].d2 ;
 wire \gen_shunt_g4[4].d1 ;
 wire \gen_shunt_g4[4].d2 ;
 wire \gen_shunt_g4[5].d1 ;
 wire \gen_shunt_g4[5].d2 ;
 wire \gen_shunt_g4[6].d1 ;
 wire \gen_shunt_g4[6].d2 ;
 wire \gen_shunt_g4[7].d1 ;
 wire \gen_shunt_g4[7].d2 ;
 wire \gen_shunt_g4[8].d1 ;
 wire \gen_shunt_g4[8].d2 ;
 wire \gen_shunt_g4[9].d1 ;
 wire \gen_shunt_g4[9].d2 ;
 wire \gen_shunt_g5[0].d1 ;
 wire \gen_shunt_g5[0].d2 ;
 wire \gen_shunt_g5[1].d1 ;
 wire \gen_shunt_g5[1].d2 ;
 wire \gen_shunt_g5[2].d1 ;
 wire \gen_shunt_g5[2].d2 ;
 wire \gen_shunt_g5[3].d1 ;
 wire \gen_shunt_g5[3].d2 ;
 wire \gen_shunt_g5[4].d1 ;
 wire \gen_shunt_g5[4].d2 ;
 wire \gen_shunt_g5[5].d1 ;
 wire \gen_shunt_g5[5].d2 ;
 wire \gen_shunt_g6[0].d1 ;
 wire \gen_shunt_g6[0].d2 ;
 wire \gen_shunt_g6[1].d1 ;
 wire \gen_shunt_g6[1].d2 ;
 wire \gen_shunt_g6[2].d1 ;
 wire \gen_shunt_g6[2].d2 ;
 wire \gen_shunt_g7[0].d1 ;
 wire \gen_shunt_g7[0].d2 ;
 wire \gen_shunt_g7[1].d1 ;
 wire \gen_shunt_g7[1].d2 ;
 wire \gen_shunt_g8[0].d1 ;
 wire \gen_shunt_g8[0].d2 ;
 wire \gen_shunt_gy_g1[0].d1 ;
 wire \gen_shunt_gy_g1[0].d2 ;
 wire \gen_shunt_gy_g1[0].d3 ;
 wire \gen_shunt_gy_g1[0].d4 ;
 wire \gen_shunt_gy_g1[1].d1 ;
 wire \gen_shunt_gy_g1[1].d2 ;
 wire \gen_shunt_gy_g1[1].d3 ;
 wire \gen_shunt_gy_g1[1].d4 ;
 wire \gen_shunt_gy_g1[2].d1 ;
 wire \gen_shunt_gy_g1[2].d2 ;
 wire \gen_shunt_gy_g1[2].d3 ;
 wire \gen_shunt_gy_g1[2].d4 ;
 wire \gen_shunt_gy_g1[3].d1 ;
 wire \gen_shunt_gy_g1[3].d2 ;
 wire \gen_shunt_gy_g1[3].d3 ;
 wire \gen_shunt_gy_g1[3].d4 ;
 wire \gen_shunt_gy_g1[4].d1 ;
 wire \gen_shunt_gy_g1[4].d2 ;
 wire \gen_shunt_gy_g1[4].d3 ;
 wire \gen_shunt_gy_g1[4].d4 ;
 wire \gen_shunt_gy_g1[5].d1 ;
 wire \gen_shunt_gy_g1[5].d2 ;
 wire \gen_shunt_gy_g1[5].d3 ;
 wire \gen_shunt_gy_g1[5].d4 ;
 wire \gen_shunt_gy_g1[6].d1 ;
 wire \gen_shunt_gy_g1[6].d2 ;
 wire \gen_shunt_gy_g1[6].d3 ;
 wire \gen_shunt_gy_g1[6].d4 ;
 wire \gen_shunt_gy_g1[7].d1 ;
 wire \gen_shunt_gy_g1[7].d2 ;
 wire \gen_shunt_gy_g1[7].d3 ;
 wire \gen_shunt_gy_g1[7].d4 ;
 wire \gen_shunt_gy_g2[0].d1 ;
 wire \gen_shunt_gy_g2[0].d2 ;
 wire \gen_shunt_gy_g2[0].d3 ;
 wire \gen_shunt_gy_g2[0].d4 ;
 wire \gen_shunt_gy_g2[1].d1 ;
 wire \gen_shunt_gy_g2[1].d2 ;
 wire \gen_shunt_gy_g2[1].d3 ;
 wire \gen_shunt_gy_g2[1].d4 ;
 wire \gen_shunt_gy_g2[2].d1 ;
 wire \gen_shunt_gy_g2[2].d2 ;
 wire \gen_shunt_gy_g2[2].d3 ;
 wire \gen_shunt_gy_g2[2].d4 ;
 wire \gen_shunt_gy_g2[3].d1 ;
 wire \gen_shunt_gy_g2[3].d2 ;
 wire \gen_shunt_gy_g2[3].d3 ;
 wire \gen_shunt_gy_g2[3].d4 ;
 wire \gen_shunt_gy_g3[0].d1 ;
 wire \gen_shunt_gy_g3[0].d2 ;
 wire \gen_shunt_gy_g3[0].d3 ;
 wire \gen_shunt_gy_g3[0].d4 ;
 wire \gen_shunt_gy_g3[1].d1 ;
 wire \gen_shunt_gy_g3[1].d2 ;
 wire \gen_shunt_gy_g3[1].d3 ;
 wire \gen_shunt_gy_g3[1].d4 ;
 wire \gen_shunt_gy_g4[0].d1 ;
 wire \gen_shunt_gy_g4[0].d2 ;
 wire \gen_shunt_gygy_g1[0].d1 ;
 wire \gen_shunt_gygy_g1[0].d2 ;
 wire \gen_shunt_gygy_g1[1].d1 ;
 wire \gen_shunt_gygy_g1[1].d2 ;
 wire \gen_shunt_gygy_g1[2].d1 ;
 wire \gen_shunt_gygy_g1[2].d2 ;
 wire \gen_shunt_gygy_g1[3].d1 ;
 wire \gen_shunt_gygy_g1[3].d2 ;
 wire \gen_shunt_gygy_g1[4].d1 ;
 wire \gen_shunt_gygy_g1[4].d2 ;
 wire \gen_shunt_gygy_g1[5].d1 ;
 wire \gen_shunt_gygy_g1[5].d2 ;
 wire \gen_shunt_gygy_g1[6].d1 ;
 wire \gen_shunt_gygy_g1[6].d2 ;
 wire \gen_shunt_gygy_g1[7].d1 ;
 wire \gen_shunt_gygy_g1[7].d2 ;
 wire \gen_shunt_gygy_g2[0].d1 ;
 wire \gen_shunt_gygy_g2[0].d2 ;
 wire \gen_shunt_gygy_g2[1].d1 ;
 wire \gen_shunt_gygy_g2[1].d2 ;
 wire \gen_shunt_gygy_g2[2].d1 ;
 wire \gen_shunt_gygy_g2[2].d2 ;
 wire \gen_shunt_gygy_g2[3].d1 ;
 wire \gen_shunt_gygy_g2[3].d2 ;
 wire \gen_shunt_gygy_g3[0].d1 ;
 wire \gen_shunt_gygy_g3[0].d2 ;
 wire \gen_shunt_gygy_g3[1].d1 ;
 wire \gen_shunt_gygy_g3[1].d2 ;
 wire \gen_shunt_gygy_g6[0].d1 ;
 wire \gen_shunt_gygy_g6[0].d2 ;
 wire \gen_shunt_gygy_g6[0].d3 ;
 wire \gen_shunt_gygy_g6[0].d4 ;
 wire \gen_shunt_gygy_g6[0].d5 ;
 wire \gen_shunt_gygy_g6[0].d6 ;

 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[10].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[10].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[11].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[11].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[12].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[12].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[13].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[13].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[14].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[14].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[15].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[15].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[8].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[8].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[9].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g1[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g1[9].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g2[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g3[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g4[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g4[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[0]),
    .ZN(\gen_series_gy_g5[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[0]),
    .ZN(\gen_series_gy_g5[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[10].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[10].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[11].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[11].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[12].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[12].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[13].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[13].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[14].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[14].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[15].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[15].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[16].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[16].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[16].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[16].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[17].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[17].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[17].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[17].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[18].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[18].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[18].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[18].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[19].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[19].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[19].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[19].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[20].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[20].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[20].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[20].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[21].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[21].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[21].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[21].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[22].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[22].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[22].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[22].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[23].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[23].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[23].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[23].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[24].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[24].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[24].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[24].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[25].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[25].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[25].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[25].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[26].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[26].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[26].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[26].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[27].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[27].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[27].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[27].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[28].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[28].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[28].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[28].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[29].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[29].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[29].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[29].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[30].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[30].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[30].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[30].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[31].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[31].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[31].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[31].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[32].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[32].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[32].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[32].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[33].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[33].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[33].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[33].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[34].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[34].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[34].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[34].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[35].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[35].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[35].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[35].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[36].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[36].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[36].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[36].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[37].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[37].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[37].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[37].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[38].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[38].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[38].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[38].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[39].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[39].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[39].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[39].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[40].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[40].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[40].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[40].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[41].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[41].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[41].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[41].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[42].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[42].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[42].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[42].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[43].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[43].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[43].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[43].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[44].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[44].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[44].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[44].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[45].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[45].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[45].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[45].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[46].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[46].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[46].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[46].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[47].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[47].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[47].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[47].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[48].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[48].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[48].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[48].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[49].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[49].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[49].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[49].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[50].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[50].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[50].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[50].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[51].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[51].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[51].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[51].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[52].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[52].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[52].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[52].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[53].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[53].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[53].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[53].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[54].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[54].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[54].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[54].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[55].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[55].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[55].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[55].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[56].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[56].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[56].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[56].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[57].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[57].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[57].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[57].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[58].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[58].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[58].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[58].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[59].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[59].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[59].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[59].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[60].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[60].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[60].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[60].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[61].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[61].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[61].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[61].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[62].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[62].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[62].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[62].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[63].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[63].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[63].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[63].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[64].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[64].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[64].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[64].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[65].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[65].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[65].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[65].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[66].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[66].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[66].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[66].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[67].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[67].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[67].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[67].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[68].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[68].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[68].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[68].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[69].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[69].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[69].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[69].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[6].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[6].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[70].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[70].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[70].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[70].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[71].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[71].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[71].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[71].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[72].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[72].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[72].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[72].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[73].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[73].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[73].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[73].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[74].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[74].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[74].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[74].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[75].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[75].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[75].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[75].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[76].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[76].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[76].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[76].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[77].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[77].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[77].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[77].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[78].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[78].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[78].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[78].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[79].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[79].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[79].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[79].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[7].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[7].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[80].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[80].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[80].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[80].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[81].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[81].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[81].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[81].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[82].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[82].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[82].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[82].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[83].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[83].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[83].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[83].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[84].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[84].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[84].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[84].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[85].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[85].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[85].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[85].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[86].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[86].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[86].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[86].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[87].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[87].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[87].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[87].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[88].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[88].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[88].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[88].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[89].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[89].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[89].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[89].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[8].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[8].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[90].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[90].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[90].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[90].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[91].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[91].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[91].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[91].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[92].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[92].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[92].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[92].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[93].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[93].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[93].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[93].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[94].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[94].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[94].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[94].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[95].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[95].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[95].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[95].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[9].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[9].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g1[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[16].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[16].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[17].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[17].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[18].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[18].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[19].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[19].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[20].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[20].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[21].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[21].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[22].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[22].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[23].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[23].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[24].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[24].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[25].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[25].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[26].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[26].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[27].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[27].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[28].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[28].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[29].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[29].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[30].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[30].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[31].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[31].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[32].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[32].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[32].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[32].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[33].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[33].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[33].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[33].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[34].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[34].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[34].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[34].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[35].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[35].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[35].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[35].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[36].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[36].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[36].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[36].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[37].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[37].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[37].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[37].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[38].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[38].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[38].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[38].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[39].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[39].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[39].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[39].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[40].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[40].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[40].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[40].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[41].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[41].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[41].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[41].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[42].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[42].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[42].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[42].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[43].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[43].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[43].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[43].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[44].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[44].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[44].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[44].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[45].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[45].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[45].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[45].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[46].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[46].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[46].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[46].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[47].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[47].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[47].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[47].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g2[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[16].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[16].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[16].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[16].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[17].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[17].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[17].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[17].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[18].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[18].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[18].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[18].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[19].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[19].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[19].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[19].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[20].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[20].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[20].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[20].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[21].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[21].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[21].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[21].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[22].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[22].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[22].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[22].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[23].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[23].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[23].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[23].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g3[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[10].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[10].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[11].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[11].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[8].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[8].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[9].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[9].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g7[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g7[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g7[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g7[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g8[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[0]),
    .ZN(\gen_shunt_g8[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g8[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[0]),
    .ZN(\gen_shunt_g8[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[6]),
    .ZN(\gen_shunt_gy_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[5]),
    .ZN(\gen_shunt_gy_g1[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g2[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g4[0].u_shunt_n  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[0]),
    .ZN(\gen_shunt_gy_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g4[0].u_shunt_p  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[0]),
    .ZN(\gen_shunt_gy_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[0].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[0].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[1].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[1].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g6[0].u_shunt_gyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g6[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g6[0].u_shunt_gyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g6[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g6[0].u_shunt_gyn3  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[0]),
    .ZN(\gen_shunt_gygy_g6[0].d6 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g6[0].u_shunt_gyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g6[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g6[0].u_shunt_gyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g6[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g6[0].u_shunt_gyp3  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[0]),
    .ZN(\gen_shunt_gygy_g6[0].d5 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_329 (.VDD(vdd),
    .VSS(vss));
endmodule
