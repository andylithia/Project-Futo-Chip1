magic
tech gf180mcuC
magscale 1 5
timestamp 1669860616
<< metal1 >>
rect 672 4325 5320 4342
rect 672 4299 1188 4325
rect 1214 4299 1240 4325
rect 1266 4299 1292 4325
rect 1318 4299 2350 4325
rect 2376 4299 2402 4325
rect 2428 4299 2454 4325
rect 2480 4299 3512 4325
rect 3538 4299 3564 4325
rect 3590 4299 3616 4325
rect 3642 4299 4674 4325
rect 4700 4299 4726 4325
rect 4752 4299 4778 4325
rect 4804 4299 5320 4325
rect 672 4282 5320 4299
rect 1079 4073 1105 4079
rect 1079 4041 1105 4047
rect 1415 4073 1441 4079
rect 1415 4041 1441 4047
rect 1751 4073 1777 4079
rect 1751 4041 1777 4047
rect 1807 4073 1833 4079
rect 1807 4041 1833 4047
rect 2087 4073 2113 4079
rect 2087 4041 2113 4047
rect 2423 4073 2449 4079
rect 2423 4041 2449 4047
rect 1135 4017 1161 4023
rect 1135 3985 1161 3991
rect 1471 4017 1497 4023
rect 1471 3985 1497 3991
rect 2143 4017 2169 4023
rect 2143 3985 2169 3991
rect 2479 4017 2505 4023
rect 2479 3985 2505 3991
rect 672 3933 5400 3950
rect 672 3907 1769 3933
rect 1795 3907 1821 3933
rect 1847 3907 1873 3933
rect 1899 3907 2931 3933
rect 2957 3907 2983 3933
rect 3009 3907 3035 3933
rect 3061 3907 4093 3933
rect 4119 3907 4145 3933
rect 4171 3907 4197 3933
rect 4223 3907 5255 3933
rect 5281 3907 5307 3933
rect 5333 3907 5359 3933
rect 5385 3907 5400 3933
rect 672 3890 5400 3907
rect 1079 3737 1105 3743
rect 1079 3705 1105 3711
rect 1415 3737 1441 3743
rect 1415 3705 1441 3711
rect 1471 3737 1497 3743
rect 1471 3705 1497 3711
rect 1751 3737 1777 3743
rect 1751 3705 1777 3711
rect 2087 3737 2113 3743
rect 2087 3705 2113 3711
rect 2143 3737 2169 3743
rect 2143 3705 2169 3711
rect 2423 3737 2449 3743
rect 2423 3705 2449 3711
rect 2479 3737 2505 3743
rect 2479 3705 2505 3711
rect 2815 3737 2841 3743
rect 2815 3705 2841 3711
rect 3151 3737 3177 3743
rect 3151 3705 3177 3711
rect 5055 3737 5081 3743
rect 5055 3705 5081 3711
rect 1135 3625 1161 3631
rect 1135 3593 1161 3599
rect 1807 3625 1833 3631
rect 1807 3593 1833 3599
rect 2759 3625 2785 3631
rect 2759 3593 2785 3599
rect 3095 3625 3121 3631
rect 3095 3593 3121 3599
rect 4999 3625 5025 3631
rect 4999 3593 5025 3599
rect 672 3541 5320 3558
rect 672 3515 1188 3541
rect 1214 3515 1240 3541
rect 1266 3515 1292 3541
rect 1318 3515 2350 3541
rect 2376 3515 2402 3541
rect 2428 3515 2454 3541
rect 2480 3515 3512 3541
rect 3538 3515 3564 3541
rect 3590 3515 3616 3541
rect 3642 3515 4674 3541
rect 4700 3515 4726 3541
rect 4752 3515 4778 3541
rect 4804 3515 5320 3541
rect 672 3498 5320 3515
rect 5055 3401 5081 3407
rect 4881 3375 4887 3401
rect 4913 3375 4919 3401
rect 5055 3369 5081 3375
rect 4825 3319 4831 3345
rect 4857 3319 4863 3345
rect 967 3289 993 3295
rect 967 3257 993 3263
rect 1303 3289 1329 3295
rect 1303 3257 1329 3263
rect 1639 3289 1665 3295
rect 1639 3257 1665 3263
rect 1695 3289 1721 3295
rect 1695 3257 1721 3263
rect 1975 3289 2001 3295
rect 1975 3257 2001 3263
rect 2311 3289 2337 3295
rect 2311 3257 2337 3263
rect 2871 3289 2897 3295
rect 2871 3257 2897 3263
rect 3207 3289 3233 3295
rect 3207 3257 3233 3263
rect 3543 3289 3569 3295
rect 3543 3257 3569 3263
rect 3599 3289 3625 3295
rect 3599 3257 3625 3263
rect 4215 3289 4241 3295
rect 4215 3257 4241 3263
rect 1023 3233 1049 3239
rect 1023 3201 1049 3207
rect 1359 3233 1385 3239
rect 1359 3201 1385 3207
rect 2031 3233 2057 3239
rect 2031 3201 2057 3207
rect 2367 3233 2393 3239
rect 2367 3201 2393 3207
rect 2927 3233 2953 3239
rect 2927 3201 2953 3207
rect 3263 3233 3289 3239
rect 3263 3201 3289 3207
rect 4271 3233 4297 3239
rect 4271 3201 4297 3207
rect 672 3149 5400 3166
rect 672 3123 1769 3149
rect 1795 3123 1821 3149
rect 1847 3123 1873 3149
rect 1899 3123 2931 3149
rect 2957 3123 2983 3149
rect 3009 3123 3035 3149
rect 3061 3123 4093 3149
rect 4119 3123 4145 3149
rect 4171 3123 4197 3149
rect 4223 3123 5255 3149
rect 5281 3123 5307 3149
rect 5333 3123 5359 3149
rect 5385 3123 5400 3149
rect 672 3106 5400 3123
rect 4999 3065 5025 3071
rect 4999 3033 5025 3039
rect 911 3009 937 3015
rect 911 2977 937 2983
rect 967 3009 993 3015
rect 967 2977 993 2983
rect 1247 3009 1273 3015
rect 1247 2977 1273 2983
rect 1303 3009 1329 3015
rect 1303 2977 1329 2983
rect 1583 3009 1609 3015
rect 1583 2977 1609 2983
rect 1919 3009 1945 3015
rect 1919 2977 1945 2983
rect 2927 3009 2953 3015
rect 2927 2977 2953 2983
rect 3263 3009 3289 3015
rect 3263 2977 3289 2983
rect 3319 3009 3345 3015
rect 3319 2977 3345 2983
rect 3879 3009 3905 3015
rect 3879 2977 3905 2983
rect 4215 3009 4241 3015
rect 4215 2977 4241 2983
rect 2255 2953 2281 2959
rect 2255 2921 2281 2927
rect 2591 2953 2617 2959
rect 2591 2921 2617 2927
rect 5055 2953 5081 2959
rect 5055 2921 5081 2927
rect 1639 2841 1665 2847
rect 1639 2809 1665 2815
rect 1975 2841 2001 2847
rect 1975 2809 2001 2815
rect 2311 2841 2337 2847
rect 2311 2809 2337 2815
rect 2647 2841 2673 2847
rect 2647 2809 2673 2815
rect 2983 2841 3009 2847
rect 2983 2809 3009 2815
rect 3935 2841 3961 2847
rect 3935 2809 3961 2815
rect 4271 2841 4297 2847
rect 4271 2809 4297 2815
rect 672 2757 5320 2774
rect 672 2731 1188 2757
rect 1214 2731 1240 2757
rect 1266 2731 1292 2757
rect 1318 2731 2350 2757
rect 2376 2731 2402 2757
rect 2428 2731 2454 2757
rect 2480 2731 3512 2757
rect 3538 2731 3564 2757
rect 3590 2731 3616 2757
rect 3642 2731 4674 2757
rect 4700 2731 4726 2757
rect 4752 2731 4778 2757
rect 4804 2731 5320 2757
rect 672 2714 5320 2731
rect 1135 2673 1161 2679
rect 1135 2641 1161 2647
rect 1471 2673 1497 2679
rect 1471 2641 1497 2647
rect 2143 2673 2169 2679
rect 2143 2641 2169 2647
rect 3543 2673 3569 2679
rect 3543 2641 3569 2647
rect 3879 2673 3905 2679
rect 3879 2641 3905 2647
rect 4999 2673 5025 2679
rect 4999 2641 5025 2647
rect 1079 2561 1105 2567
rect 1079 2529 1105 2535
rect 1415 2561 1441 2567
rect 1415 2529 1441 2535
rect 1751 2561 1777 2567
rect 1751 2529 1777 2535
rect 1807 2561 1833 2567
rect 1807 2529 1833 2535
rect 3487 2561 3513 2567
rect 3487 2529 3513 2535
rect 4159 2561 4185 2567
rect 4159 2529 4185 2535
rect 4215 2561 4241 2567
rect 4215 2529 4241 2535
rect 5055 2561 5081 2567
rect 5055 2529 5081 2535
rect 2087 2505 2113 2511
rect 2087 2473 2113 2479
rect 2423 2505 2449 2511
rect 2423 2473 2449 2479
rect 2479 2505 2505 2511
rect 2479 2473 2505 2479
rect 2871 2505 2897 2511
rect 2871 2473 2897 2479
rect 2927 2505 2953 2511
rect 2927 2473 2953 2479
rect 3823 2505 3849 2511
rect 3823 2473 3849 2479
rect 4663 2505 4689 2511
rect 4663 2473 4689 2479
rect 4719 2449 4745 2455
rect 4719 2417 4745 2423
rect 672 2365 5400 2382
rect 672 2339 1769 2365
rect 1795 2339 1821 2365
rect 1847 2339 1873 2365
rect 1899 2339 2931 2365
rect 2957 2339 2983 2365
rect 3009 2339 3035 2365
rect 3061 2339 4093 2365
rect 4119 2339 4145 2365
rect 4171 2339 4197 2365
rect 4223 2339 5255 2365
rect 5281 2339 5307 2365
rect 5333 2339 5359 2365
rect 5385 2339 5400 2365
rect 672 2322 5400 2339
rect 1023 2281 1049 2287
rect 1023 2249 1049 2255
rect 1695 2281 1721 2287
rect 1695 2249 1721 2255
rect 3263 2281 3289 2287
rect 3263 2249 3289 2255
rect 3599 2281 3625 2287
rect 3599 2249 3625 2255
rect 967 2225 993 2231
rect 967 2193 993 2199
rect 1303 2225 1329 2231
rect 1303 2193 1329 2199
rect 1975 2225 2001 2231
rect 1975 2193 2001 2199
rect 3207 2225 3233 2231
rect 3207 2193 3233 2199
rect 3543 2225 3569 2231
rect 3543 2193 3569 2199
rect 3879 2225 3905 2231
rect 3879 2193 3905 2199
rect 1639 2169 1665 2175
rect 1639 2137 1665 2143
rect 2311 2169 2337 2175
rect 2311 2137 2337 2143
rect 2871 2169 2897 2175
rect 2871 2137 2897 2143
rect 4215 2169 4241 2175
rect 4215 2137 4241 2143
rect 4999 2169 5025 2175
rect 4999 2137 5025 2143
rect 1359 2057 1385 2063
rect 1359 2025 1385 2031
rect 2031 2057 2057 2063
rect 2031 2025 2057 2031
rect 2367 2057 2393 2063
rect 2367 2025 2393 2031
rect 2927 2057 2953 2063
rect 2927 2025 2953 2031
rect 3935 2057 3961 2063
rect 3935 2025 3961 2031
rect 4271 2057 4297 2063
rect 4271 2025 4297 2031
rect 5055 2057 5081 2063
rect 5055 2025 5081 2031
rect 672 1973 5320 1990
rect 672 1947 1188 1973
rect 1214 1947 1240 1973
rect 1266 1947 1292 1973
rect 1318 1947 2350 1973
rect 2376 1947 2402 1973
rect 2428 1947 2454 1973
rect 2480 1947 3512 1973
rect 3538 1947 3564 1973
rect 3590 1947 3616 1973
rect 3642 1947 4674 1973
rect 4700 1947 4726 1973
rect 4752 1947 4778 1973
rect 4804 1947 5320 1973
rect 672 1930 5320 1947
rect 2927 1889 2953 1895
rect 2927 1857 2953 1863
rect 3375 1889 3401 1895
rect 3375 1857 3401 1863
rect 3711 1889 3737 1895
rect 3711 1857 3737 1863
rect 3991 1889 4017 1895
rect 3991 1857 4017 1863
rect 4383 1833 4409 1839
rect 4383 1801 4409 1807
rect 5055 1833 5081 1839
rect 5055 1801 5081 1807
rect 1023 1777 1049 1783
rect 1023 1745 1049 1751
rect 1359 1777 1385 1783
rect 1359 1745 1385 1751
rect 3319 1777 3345 1783
rect 3319 1745 3345 1751
rect 3655 1777 3681 1783
rect 3655 1745 3681 1751
rect 4047 1777 4073 1783
rect 4047 1745 4073 1751
rect 4327 1777 4353 1783
rect 4327 1745 4353 1751
rect 967 1721 993 1727
rect 967 1689 993 1695
rect 1303 1721 1329 1727
rect 1303 1689 1329 1695
rect 1639 1721 1665 1727
rect 1639 1689 1665 1695
rect 1695 1721 1721 1727
rect 1695 1689 1721 1695
rect 1975 1721 2001 1727
rect 1975 1689 2001 1695
rect 2031 1721 2057 1727
rect 2031 1689 2057 1695
rect 2311 1721 2337 1727
rect 2311 1689 2337 1695
rect 2367 1721 2393 1727
rect 2367 1689 2393 1695
rect 2871 1721 2897 1727
rect 2871 1689 2897 1695
rect 4999 1721 5025 1727
rect 4999 1689 5025 1695
rect 672 1581 5400 1598
rect 672 1555 1769 1581
rect 1795 1555 1821 1581
rect 1847 1555 1873 1581
rect 1899 1555 2931 1581
rect 2957 1555 2983 1581
rect 3009 1555 3035 1581
rect 3061 1555 4093 1581
rect 4119 1555 4145 1581
rect 4171 1555 4197 1581
rect 4223 1555 5255 1581
rect 5281 1555 5307 1581
rect 5333 1555 5359 1581
rect 5385 1555 5400 1581
rect 672 1538 5400 1555
<< via1 >>
rect 1188 4299 1214 4325
rect 1240 4299 1266 4325
rect 1292 4299 1318 4325
rect 2350 4299 2376 4325
rect 2402 4299 2428 4325
rect 2454 4299 2480 4325
rect 3512 4299 3538 4325
rect 3564 4299 3590 4325
rect 3616 4299 3642 4325
rect 4674 4299 4700 4325
rect 4726 4299 4752 4325
rect 4778 4299 4804 4325
rect 1079 4047 1105 4073
rect 1415 4047 1441 4073
rect 1751 4047 1777 4073
rect 1807 4047 1833 4073
rect 2087 4047 2113 4073
rect 2423 4047 2449 4073
rect 1135 3991 1161 4017
rect 1471 3991 1497 4017
rect 2143 3991 2169 4017
rect 2479 3991 2505 4017
rect 1769 3907 1795 3933
rect 1821 3907 1847 3933
rect 1873 3907 1899 3933
rect 2931 3907 2957 3933
rect 2983 3907 3009 3933
rect 3035 3907 3061 3933
rect 4093 3907 4119 3933
rect 4145 3907 4171 3933
rect 4197 3907 4223 3933
rect 5255 3907 5281 3933
rect 5307 3907 5333 3933
rect 5359 3907 5385 3933
rect 1079 3711 1105 3737
rect 1415 3711 1441 3737
rect 1471 3711 1497 3737
rect 1751 3711 1777 3737
rect 2087 3711 2113 3737
rect 2143 3711 2169 3737
rect 2423 3711 2449 3737
rect 2479 3711 2505 3737
rect 2815 3711 2841 3737
rect 3151 3711 3177 3737
rect 5055 3711 5081 3737
rect 1135 3599 1161 3625
rect 1807 3599 1833 3625
rect 2759 3599 2785 3625
rect 3095 3599 3121 3625
rect 4999 3599 5025 3625
rect 1188 3515 1214 3541
rect 1240 3515 1266 3541
rect 1292 3515 1318 3541
rect 2350 3515 2376 3541
rect 2402 3515 2428 3541
rect 2454 3515 2480 3541
rect 3512 3515 3538 3541
rect 3564 3515 3590 3541
rect 3616 3515 3642 3541
rect 4674 3515 4700 3541
rect 4726 3515 4752 3541
rect 4778 3515 4804 3541
rect 4887 3375 4913 3401
rect 5055 3375 5081 3401
rect 4831 3319 4857 3345
rect 967 3263 993 3289
rect 1303 3263 1329 3289
rect 1639 3263 1665 3289
rect 1695 3263 1721 3289
rect 1975 3263 2001 3289
rect 2311 3263 2337 3289
rect 2871 3263 2897 3289
rect 3207 3263 3233 3289
rect 3543 3263 3569 3289
rect 3599 3263 3625 3289
rect 4215 3263 4241 3289
rect 1023 3207 1049 3233
rect 1359 3207 1385 3233
rect 2031 3207 2057 3233
rect 2367 3207 2393 3233
rect 2927 3207 2953 3233
rect 3263 3207 3289 3233
rect 4271 3207 4297 3233
rect 1769 3123 1795 3149
rect 1821 3123 1847 3149
rect 1873 3123 1899 3149
rect 2931 3123 2957 3149
rect 2983 3123 3009 3149
rect 3035 3123 3061 3149
rect 4093 3123 4119 3149
rect 4145 3123 4171 3149
rect 4197 3123 4223 3149
rect 5255 3123 5281 3149
rect 5307 3123 5333 3149
rect 5359 3123 5385 3149
rect 4999 3039 5025 3065
rect 911 2983 937 3009
rect 967 2983 993 3009
rect 1247 2983 1273 3009
rect 1303 2983 1329 3009
rect 1583 2983 1609 3009
rect 1919 2983 1945 3009
rect 2927 2983 2953 3009
rect 3263 2983 3289 3009
rect 3319 2983 3345 3009
rect 3879 2983 3905 3009
rect 4215 2983 4241 3009
rect 2255 2927 2281 2953
rect 2591 2927 2617 2953
rect 5055 2927 5081 2953
rect 1639 2815 1665 2841
rect 1975 2815 2001 2841
rect 2311 2815 2337 2841
rect 2647 2815 2673 2841
rect 2983 2815 3009 2841
rect 3935 2815 3961 2841
rect 4271 2815 4297 2841
rect 1188 2731 1214 2757
rect 1240 2731 1266 2757
rect 1292 2731 1318 2757
rect 2350 2731 2376 2757
rect 2402 2731 2428 2757
rect 2454 2731 2480 2757
rect 3512 2731 3538 2757
rect 3564 2731 3590 2757
rect 3616 2731 3642 2757
rect 4674 2731 4700 2757
rect 4726 2731 4752 2757
rect 4778 2731 4804 2757
rect 1135 2647 1161 2673
rect 1471 2647 1497 2673
rect 2143 2647 2169 2673
rect 3543 2647 3569 2673
rect 3879 2647 3905 2673
rect 4999 2647 5025 2673
rect 1079 2535 1105 2561
rect 1415 2535 1441 2561
rect 1751 2535 1777 2561
rect 1807 2535 1833 2561
rect 3487 2535 3513 2561
rect 4159 2535 4185 2561
rect 4215 2535 4241 2561
rect 5055 2535 5081 2561
rect 2087 2479 2113 2505
rect 2423 2479 2449 2505
rect 2479 2479 2505 2505
rect 2871 2479 2897 2505
rect 2927 2479 2953 2505
rect 3823 2479 3849 2505
rect 4663 2479 4689 2505
rect 4719 2423 4745 2449
rect 1769 2339 1795 2365
rect 1821 2339 1847 2365
rect 1873 2339 1899 2365
rect 2931 2339 2957 2365
rect 2983 2339 3009 2365
rect 3035 2339 3061 2365
rect 4093 2339 4119 2365
rect 4145 2339 4171 2365
rect 4197 2339 4223 2365
rect 5255 2339 5281 2365
rect 5307 2339 5333 2365
rect 5359 2339 5385 2365
rect 1023 2255 1049 2281
rect 1695 2255 1721 2281
rect 3263 2255 3289 2281
rect 3599 2255 3625 2281
rect 967 2199 993 2225
rect 1303 2199 1329 2225
rect 1975 2199 2001 2225
rect 3207 2199 3233 2225
rect 3543 2199 3569 2225
rect 3879 2199 3905 2225
rect 1639 2143 1665 2169
rect 2311 2143 2337 2169
rect 2871 2143 2897 2169
rect 4215 2143 4241 2169
rect 4999 2143 5025 2169
rect 1359 2031 1385 2057
rect 2031 2031 2057 2057
rect 2367 2031 2393 2057
rect 2927 2031 2953 2057
rect 3935 2031 3961 2057
rect 4271 2031 4297 2057
rect 5055 2031 5081 2057
rect 1188 1947 1214 1973
rect 1240 1947 1266 1973
rect 1292 1947 1318 1973
rect 2350 1947 2376 1973
rect 2402 1947 2428 1973
rect 2454 1947 2480 1973
rect 3512 1947 3538 1973
rect 3564 1947 3590 1973
rect 3616 1947 3642 1973
rect 4674 1947 4700 1973
rect 4726 1947 4752 1973
rect 4778 1947 4804 1973
rect 2927 1863 2953 1889
rect 3375 1863 3401 1889
rect 3711 1863 3737 1889
rect 3991 1863 4017 1889
rect 4383 1807 4409 1833
rect 5055 1807 5081 1833
rect 1023 1751 1049 1777
rect 1359 1751 1385 1777
rect 3319 1751 3345 1777
rect 3655 1751 3681 1777
rect 4047 1751 4073 1777
rect 4327 1751 4353 1777
rect 967 1695 993 1721
rect 1303 1695 1329 1721
rect 1639 1695 1665 1721
rect 1695 1695 1721 1721
rect 1975 1695 2001 1721
rect 2031 1695 2057 1721
rect 2311 1695 2337 1721
rect 2367 1695 2393 1721
rect 2871 1695 2897 1721
rect 4999 1695 5025 1721
rect 1769 1555 1795 1581
rect 1821 1555 1847 1581
rect 1873 1555 1899 1581
rect 2931 1555 2957 1581
rect 2983 1555 3009 1581
rect 3035 1555 3061 1581
rect 4093 1555 4119 1581
rect 4145 1555 4171 1581
rect 4197 1555 4223 1581
rect 5255 1555 5281 1581
rect 5307 1555 5333 1581
rect 5359 1555 5385 1581
<< metal2 >>
rect 4942 5362 4970 5367
rect 1187 4326 1319 4331
rect 1215 4298 1239 4326
rect 1267 4298 1291 4326
rect 1187 4293 1319 4298
rect 2349 4326 2481 4331
rect 2377 4298 2401 4326
rect 2429 4298 2453 4326
rect 2349 4293 2481 4298
rect 3511 4326 3643 4331
rect 3539 4298 3563 4326
rect 3591 4298 3615 4326
rect 3511 4293 3643 4298
rect 4673 4326 4805 4331
rect 4701 4298 4725 4326
rect 4753 4298 4777 4326
rect 4673 4293 4805 4298
rect 1134 4186 1162 4191
rect 1078 4074 1106 4079
rect 1134 4074 1162 4158
rect 4886 4186 4914 4191
rect 1078 4073 1162 4074
rect 1078 4047 1079 4073
rect 1105 4047 1162 4073
rect 1078 4046 1162 4047
rect 1078 4041 1106 4046
rect 1134 4017 1162 4046
rect 1414 4074 1442 4079
rect 1750 4074 1778 4079
rect 1806 4074 1834 4079
rect 1414 4073 1498 4074
rect 1414 4047 1415 4073
rect 1441 4047 1498 4073
rect 1414 4046 1498 4047
rect 1414 4041 1442 4046
rect 1134 3991 1135 4017
rect 1161 3991 1162 4017
rect 1078 3737 1106 3743
rect 1078 3711 1079 3737
rect 1105 3711 1106 3737
rect 1078 3626 1106 3711
rect 1134 3626 1162 3991
rect 1470 4017 1498 4046
rect 1470 3991 1471 4017
rect 1497 3991 1498 4017
rect 1414 3738 1442 3743
rect 1470 3738 1498 3991
rect 1078 3625 1162 3626
rect 1078 3599 1135 3625
rect 1161 3599 1162 3625
rect 1078 3598 1162 3599
rect 966 3289 994 3295
rect 966 3263 967 3289
rect 993 3263 994 3289
rect 966 3234 994 3263
rect 1022 3234 1050 3239
rect 1078 3234 1106 3598
rect 1134 3593 1162 3598
rect 1358 3737 1498 3738
rect 1358 3711 1415 3737
rect 1441 3711 1471 3737
rect 1497 3711 1498 3737
rect 1358 3710 1498 3711
rect 1694 4073 1834 4074
rect 1694 4047 1751 4073
rect 1777 4047 1807 4073
rect 1833 4047 1834 4073
rect 1694 4046 1834 4047
rect 1694 3738 1722 4046
rect 1750 4041 1778 4046
rect 1806 4041 1834 4046
rect 2086 4074 2114 4079
rect 2086 4073 2170 4074
rect 2086 4047 2087 4073
rect 2113 4047 2170 4073
rect 2086 4046 2170 4047
rect 2086 4041 2114 4046
rect 2142 4017 2170 4046
rect 2142 3991 2143 4017
rect 2169 3991 2170 4017
rect 1768 3934 1900 3939
rect 1796 3906 1820 3934
rect 1848 3906 1872 3934
rect 1768 3901 1900 3906
rect 1750 3738 1778 3743
rect 2086 3738 2114 3743
rect 2142 3738 2170 3991
rect 2422 4073 2450 4079
rect 2422 4047 2423 4073
rect 2449 4047 2450 4073
rect 2422 4018 2450 4047
rect 2478 4018 2506 4023
rect 2422 4017 2506 4018
rect 2422 3991 2479 4017
rect 2505 3991 2506 4017
rect 2422 3990 2506 3991
rect 2422 3738 2450 3990
rect 2478 3985 2506 3990
rect 2930 3934 3062 3939
rect 2958 3906 2982 3934
rect 3010 3906 3034 3934
rect 2930 3901 3062 3906
rect 4092 3934 4224 3939
rect 4120 3906 4144 3934
rect 4172 3906 4196 3934
rect 4092 3901 4224 3906
rect 2478 3738 2506 3743
rect 2814 3738 2842 3743
rect 3150 3738 3178 3743
rect 1694 3737 1778 3738
rect 1694 3711 1751 3737
rect 1777 3711 1778 3737
rect 1694 3710 1778 3711
rect 1187 3542 1319 3547
rect 1215 3514 1239 3542
rect 1267 3514 1291 3542
rect 1187 3509 1319 3514
rect 966 3233 1106 3234
rect 966 3207 1023 3233
rect 1049 3207 1106 3233
rect 966 3206 1106 3207
rect 1302 3289 1330 3295
rect 1302 3263 1303 3289
rect 1329 3263 1330 3289
rect 1302 3234 1330 3263
rect 1358 3234 1386 3710
rect 1414 3705 1442 3710
rect 1470 3705 1498 3710
rect 1750 3626 1778 3710
rect 2030 3737 2506 3738
rect 2030 3711 2087 3737
rect 2113 3711 2143 3737
rect 2169 3711 2423 3737
rect 2449 3711 2479 3737
rect 2505 3711 2506 3737
rect 2030 3710 2506 3711
rect 1806 3626 1834 3631
rect 1750 3625 1834 3626
rect 1750 3599 1807 3625
rect 1833 3599 1834 3625
rect 1750 3598 1834 3599
rect 1638 3290 1666 3295
rect 1694 3290 1722 3295
rect 1750 3290 1778 3598
rect 1806 3593 1834 3598
rect 1302 3233 1386 3234
rect 1302 3207 1359 3233
rect 1385 3207 1386 3233
rect 1302 3206 1386 3207
rect 910 3010 938 3015
rect 966 3010 994 3206
rect 1022 3201 1050 3206
rect 910 3009 966 3010
rect 910 2983 911 3009
rect 937 2983 966 3009
rect 910 2982 966 2983
rect 910 2977 938 2982
rect 966 2963 994 2982
rect 1246 3010 1274 3015
rect 1302 3010 1330 3206
rect 1358 3201 1386 3206
rect 1582 3289 1778 3290
rect 1582 3263 1639 3289
rect 1665 3263 1695 3289
rect 1721 3263 1778 3289
rect 1582 3262 1778 3263
rect 1974 3289 2002 3295
rect 1974 3263 1975 3289
rect 2001 3263 2002 3289
rect 1246 3009 1302 3010
rect 1246 2983 1247 3009
rect 1273 2983 1302 3009
rect 1246 2982 1302 2983
rect 1246 2977 1274 2982
rect 1302 2963 1330 2982
rect 1470 3010 1498 3015
rect 1187 2758 1319 2763
rect 1215 2730 1239 2758
rect 1267 2730 1291 2758
rect 1187 2725 1319 2730
rect 1134 2674 1162 2679
rect 1022 2646 1134 2674
rect 966 2562 994 2567
rect 966 2226 994 2534
rect 910 2225 994 2226
rect 910 2199 967 2225
rect 993 2199 994 2225
rect 910 2198 994 2199
rect 910 1722 938 2198
rect 966 2193 994 2198
rect 1022 2281 1050 2646
rect 1134 2627 1162 2646
rect 1302 2674 1330 2679
rect 1078 2562 1106 2567
rect 1078 2515 1106 2534
rect 1022 2255 1023 2281
rect 1049 2255 1050 2281
rect 1022 1777 1050 2255
rect 1302 2225 1330 2646
rect 1470 2674 1498 2982
rect 1582 3010 1610 3262
rect 1638 3257 1666 3262
rect 1694 3257 1722 3262
rect 1974 3234 2002 3263
rect 2030 3234 2058 3710
rect 2086 3705 2114 3710
rect 2142 3705 2170 3710
rect 2422 3705 2450 3710
rect 2478 3705 2506 3710
rect 2758 3737 2842 3738
rect 2758 3711 2815 3737
rect 2841 3711 2842 3737
rect 2758 3710 2842 3711
rect 2758 3625 2786 3710
rect 2814 3705 2842 3710
rect 3094 3737 3178 3738
rect 3094 3711 3151 3737
rect 3177 3711 3178 3737
rect 3094 3710 3178 3711
rect 2758 3599 2759 3625
rect 2785 3599 2786 3625
rect 2349 3542 2481 3547
rect 2377 3514 2401 3542
rect 2429 3514 2453 3542
rect 2349 3509 2481 3514
rect 1974 3233 2058 3234
rect 1974 3207 2031 3233
rect 2057 3207 2058 3233
rect 1974 3206 2058 3207
rect 1768 3150 1900 3155
rect 1796 3122 1820 3150
rect 1848 3122 1872 3150
rect 1768 3117 1900 3122
rect 1582 2963 1610 2982
rect 1750 3010 1778 3015
rect 1414 2562 1442 2567
rect 1414 2515 1442 2534
rect 1302 2199 1303 2225
rect 1329 2199 1330 2225
rect 1302 2193 1330 2199
rect 1470 2114 1498 2646
rect 1638 2841 1666 2847
rect 1638 2815 1639 2841
rect 1665 2815 1666 2841
rect 1638 2562 1666 2815
rect 1750 2562 1778 2982
rect 1918 3010 1946 3015
rect 1974 3010 2002 3206
rect 2030 3201 2058 3206
rect 2310 3289 2338 3295
rect 2310 3263 2311 3289
rect 2337 3263 2338 3289
rect 2310 3234 2338 3263
rect 2758 3290 2786 3599
rect 3094 3625 3122 3710
rect 3150 3705 3178 3710
rect 3094 3599 3095 3625
rect 3121 3599 3122 3625
rect 2870 3290 2898 3295
rect 2758 3262 2870 3290
rect 2366 3234 2394 3239
rect 2310 3233 2394 3234
rect 2310 3207 2367 3233
rect 2393 3207 2394 3233
rect 2310 3206 2394 3207
rect 1946 2982 2002 3010
rect 2142 3010 2170 3015
rect 1918 2963 1946 2982
rect 1974 2842 2002 2847
rect 2030 2842 2058 2847
rect 1974 2841 2030 2842
rect 1974 2815 1975 2841
rect 2001 2815 2030 2841
rect 1974 2814 2030 2815
rect 1974 2809 2002 2814
rect 1638 2529 1666 2534
rect 1694 2561 1778 2562
rect 1694 2535 1751 2561
rect 1777 2535 1778 2561
rect 1694 2534 1778 2535
rect 1694 2282 1722 2534
rect 1750 2529 1778 2534
rect 1806 2562 1834 2567
rect 1806 2515 1834 2534
rect 2030 2506 2058 2814
rect 2142 2673 2170 2982
rect 2254 2954 2282 2959
rect 2310 2954 2338 3206
rect 2366 3201 2394 3206
rect 2870 3234 2898 3262
rect 3094 3290 3122 3599
rect 4606 3626 4634 3631
rect 3511 3542 3643 3547
rect 3539 3514 3563 3542
rect 3591 3514 3615 3542
rect 3511 3509 3643 3514
rect 3094 3257 3122 3262
rect 3206 3290 3234 3295
rect 2926 3234 2954 3239
rect 2870 3233 2954 3234
rect 2870 3207 2927 3233
rect 2953 3207 2954 3233
rect 2870 3206 2954 3207
rect 2254 2953 2338 2954
rect 2254 2927 2255 2953
rect 2281 2927 2338 2953
rect 2254 2926 2338 2927
rect 2254 2921 2282 2926
rect 2310 2842 2338 2926
rect 2310 2809 2338 2814
rect 2590 2953 2618 2959
rect 2590 2927 2591 2953
rect 2617 2927 2618 2953
rect 2590 2842 2618 2927
rect 2646 2842 2674 2847
rect 2618 2841 2674 2842
rect 2618 2815 2647 2841
rect 2673 2815 2674 2841
rect 2618 2814 2674 2815
rect 2590 2809 2618 2814
rect 2646 2809 2674 2814
rect 2349 2758 2481 2763
rect 2377 2730 2401 2758
rect 2429 2730 2453 2758
rect 2349 2725 2481 2730
rect 2142 2647 2143 2673
rect 2169 2647 2170 2673
rect 2142 2641 2170 2647
rect 2086 2506 2114 2511
rect 2422 2506 2450 2511
rect 2478 2506 2506 2511
rect 2030 2505 2114 2506
rect 2030 2479 2087 2505
rect 2113 2479 2114 2505
rect 2030 2478 2114 2479
rect 1768 2366 1900 2371
rect 1796 2338 1820 2366
rect 1848 2338 1872 2366
rect 1768 2333 1900 2338
rect 1694 2281 2002 2282
rect 1694 2255 1695 2281
rect 1721 2255 2002 2281
rect 1694 2254 2002 2255
rect 1694 2249 1722 2254
rect 1974 2225 2002 2254
rect 1974 2199 1975 2225
rect 2001 2199 2002 2225
rect 1974 2193 2002 2199
rect 1414 2086 1498 2114
rect 1638 2169 1666 2175
rect 1638 2143 1639 2169
rect 1665 2143 1666 2169
rect 1358 2057 1386 2063
rect 1358 2031 1359 2057
rect 1385 2031 1386 2057
rect 1187 1974 1319 1979
rect 1215 1946 1239 1974
rect 1267 1946 1291 1974
rect 1187 1941 1319 1946
rect 1358 1890 1386 2031
rect 1022 1751 1023 1777
rect 1049 1751 1050 1777
rect 1022 1745 1050 1751
rect 1302 1862 1386 1890
rect 966 1722 994 1727
rect 910 1721 994 1722
rect 910 1695 967 1721
rect 993 1695 994 1721
rect 910 1694 994 1695
rect 966 1666 994 1694
rect 1302 1722 1330 1862
rect 1358 1778 1386 1783
rect 1414 1778 1442 2086
rect 1358 1777 1442 1778
rect 1358 1751 1359 1777
rect 1385 1751 1442 1777
rect 1358 1750 1442 1751
rect 1358 1745 1386 1750
rect 1302 1675 1330 1694
rect 1638 1722 1666 2143
rect 2030 2057 2058 2478
rect 2086 2473 2114 2478
rect 2366 2505 2506 2506
rect 2366 2479 2423 2505
rect 2449 2479 2479 2505
rect 2505 2479 2506 2505
rect 2366 2478 2506 2479
rect 2310 2169 2338 2175
rect 2310 2143 2311 2169
rect 2337 2143 2338 2169
rect 2310 2058 2338 2143
rect 2366 2058 2394 2478
rect 2422 2473 2450 2478
rect 2478 2473 2506 2478
rect 2870 2506 2898 3206
rect 2926 3201 2954 3206
rect 3206 3234 3234 3262
rect 3542 3290 3570 3295
rect 3598 3290 3626 3295
rect 3570 3289 3626 3290
rect 3570 3263 3599 3289
rect 3625 3263 3626 3289
rect 3570 3262 3626 3263
rect 3542 3243 3570 3262
rect 3598 3257 3626 3262
rect 4214 3290 4242 3295
rect 4214 3289 4298 3290
rect 4214 3263 4215 3289
rect 4241 3263 4298 3289
rect 4214 3262 4298 3263
rect 4214 3257 4242 3262
rect 3262 3234 3290 3239
rect 3206 3233 3290 3234
rect 3206 3207 3263 3233
rect 3289 3207 3290 3233
rect 3206 3206 3290 3207
rect 2930 3150 3062 3155
rect 2958 3122 2982 3150
rect 3010 3122 3034 3150
rect 2930 3117 3062 3122
rect 2926 3010 2954 3015
rect 3206 3010 3234 3206
rect 3262 3201 3290 3206
rect 4270 3234 4298 3262
rect 4270 3233 4354 3234
rect 4270 3207 4271 3233
rect 4297 3207 4354 3233
rect 4270 3206 4354 3207
rect 4270 3201 4298 3206
rect 4092 3150 4224 3155
rect 4120 3122 4144 3150
rect 4172 3122 4196 3150
rect 4092 3117 4224 3122
rect 3262 3010 3290 3015
rect 3318 3010 3346 3015
rect 3206 3009 3346 3010
rect 3206 2983 3263 3009
rect 3289 2983 3319 3009
rect 3345 2983 3346 3009
rect 3206 2982 3346 2983
rect 2926 2963 2954 2982
rect 3262 2977 3290 2982
rect 3318 2977 3346 2982
rect 3878 3010 3906 3015
rect 3878 2963 3906 2982
rect 4158 3010 4186 3015
rect 4214 3010 4242 3015
rect 4186 3009 4242 3010
rect 4186 2983 4215 3009
rect 4241 2983 4242 3009
rect 4186 2982 4242 2983
rect 2982 2841 3010 2847
rect 2982 2815 2983 2841
rect 3009 2815 3010 2841
rect 2982 2674 3010 2815
rect 3934 2842 3962 2847
rect 3511 2758 3643 2763
rect 3539 2730 3563 2758
rect 3591 2730 3615 2758
rect 3511 2725 3643 2730
rect 2982 2641 3010 2646
rect 3542 2674 3570 2679
rect 3486 2562 3514 2567
rect 3542 2562 3570 2646
rect 3878 2674 3906 2679
rect 3934 2674 3962 2814
rect 3906 2646 3962 2674
rect 3878 2608 3906 2646
rect 3486 2561 3570 2562
rect 3486 2535 3487 2561
rect 3513 2535 3570 2561
rect 3486 2534 3570 2535
rect 3486 2529 3514 2534
rect 2926 2506 2954 2511
rect 2870 2505 2954 2506
rect 2870 2479 2871 2505
rect 2897 2479 2927 2505
rect 2953 2479 2954 2505
rect 2870 2478 2954 2479
rect 2030 2031 2031 2057
rect 2057 2031 2058 2057
rect 1694 1722 1722 1727
rect 1638 1721 1722 1722
rect 1638 1695 1639 1721
rect 1665 1695 1695 1721
rect 1721 1695 1722 1721
rect 1638 1694 1722 1695
rect 1638 1689 1666 1694
rect 966 1498 994 1638
rect 1694 1666 1722 1694
rect 1694 1633 1722 1638
rect 1974 1722 2002 1727
rect 2030 1722 2058 2031
rect 1974 1721 2058 1722
rect 1974 1695 1975 1721
rect 2001 1695 2031 1721
rect 2057 1695 2058 1721
rect 1974 1694 2058 1695
rect 2254 2057 2394 2058
rect 2254 2031 2367 2057
rect 2393 2031 2394 2057
rect 2254 2030 2394 2031
rect 2254 1722 2282 2030
rect 2366 2025 2394 2030
rect 2870 2226 2898 2478
rect 2926 2473 2954 2478
rect 2930 2366 3062 2371
rect 2958 2338 2982 2366
rect 3010 2338 3034 2366
rect 2930 2333 3062 2338
rect 3262 2282 3290 2287
rect 3542 2282 3570 2534
rect 4158 2561 4186 2982
rect 4214 2977 4242 2982
rect 4270 2842 4298 2847
rect 4158 2535 4159 2561
rect 4185 2535 4186 2561
rect 4158 2529 4186 2535
rect 4214 2562 4242 2567
rect 4270 2562 4298 2814
rect 4242 2534 4298 2562
rect 4214 2515 4242 2534
rect 3822 2505 3850 2511
rect 3822 2479 3823 2505
rect 3849 2479 3850 2505
rect 3598 2282 3626 2287
rect 3262 2281 3626 2282
rect 3262 2255 3263 2281
rect 3289 2255 3599 2281
rect 3625 2255 3626 2281
rect 3262 2254 3626 2255
rect 2870 2169 2898 2198
rect 3206 2226 3234 2231
rect 3262 2226 3290 2254
rect 3206 2225 3290 2226
rect 3206 2199 3207 2225
rect 3233 2199 3290 2225
rect 3206 2198 3290 2199
rect 3206 2193 3234 2198
rect 2870 2143 2871 2169
rect 2897 2143 2898 2169
rect 2349 1974 2481 1979
rect 2377 1946 2401 1974
rect 2429 1946 2453 1974
rect 2349 1941 2481 1946
rect 2870 1890 2898 2143
rect 2926 2058 2954 2063
rect 2926 2011 2954 2030
rect 2926 1890 2954 1895
rect 3374 1890 3402 2254
rect 3542 2225 3570 2254
rect 3598 2249 3626 2254
rect 3542 2199 3543 2225
rect 3569 2199 3570 2225
rect 3542 2193 3570 2199
rect 3710 2058 3738 2063
rect 3511 1974 3643 1979
rect 3539 1946 3563 1974
rect 3591 1946 3615 1974
rect 3511 1941 3643 1946
rect 2870 1889 2954 1890
rect 2870 1863 2927 1889
rect 2953 1863 2954 1889
rect 2870 1862 2954 1863
rect 2310 1722 2338 1727
rect 2366 1722 2394 1727
rect 2254 1721 2394 1722
rect 2254 1695 2311 1721
rect 2337 1695 2367 1721
rect 2393 1695 2394 1721
rect 2254 1694 2394 1695
rect 1974 1666 2002 1694
rect 2030 1689 2058 1694
rect 1974 1633 2002 1638
rect 2310 1666 2338 1694
rect 2366 1689 2394 1694
rect 2870 1722 2898 1862
rect 2926 1857 2954 1862
rect 3318 1889 3682 1890
rect 3318 1863 3375 1889
rect 3401 1863 3682 1889
rect 3318 1862 3682 1863
rect 3318 1777 3346 1862
rect 3374 1857 3402 1862
rect 3318 1751 3319 1777
rect 3345 1751 3346 1777
rect 3318 1745 3346 1751
rect 3654 1777 3682 1862
rect 3710 1889 3738 2030
rect 3822 2058 3850 2479
rect 4326 2450 4354 3206
rect 4606 2562 4634 3598
rect 4673 3542 4805 3547
rect 4701 3514 4725 3542
rect 4753 3514 4777 3542
rect 4673 3509 4805 3514
rect 4886 3402 4914 4158
rect 4942 3514 4970 5334
rect 5254 3934 5386 3939
rect 5282 3906 5306 3934
rect 5334 3906 5358 3934
rect 5254 3901 5386 3906
rect 5054 3738 5082 3743
rect 5054 3737 5138 3738
rect 5054 3711 5055 3737
rect 5081 3711 5138 3737
rect 5054 3710 5138 3711
rect 5054 3705 5082 3710
rect 4998 3626 5026 3631
rect 4998 3579 5026 3598
rect 4942 3486 5026 3514
rect 4998 3402 5026 3486
rect 5054 3402 5082 3407
rect 4886 3401 4970 3402
rect 4886 3375 4887 3401
rect 4913 3375 4970 3401
rect 4886 3374 4970 3375
rect 4998 3401 5082 3402
rect 4998 3375 5055 3401
rect 5081 3375 5082 3401
rect 4998 3374 5082 3375
rect 4886 3369 4914 3374
rect 4830 3345 4858 3351
rect 4830 3319 4831 3345
rect 4857 3319 4858 3345
rect 4830 3010 4858 3319
rect 4942 3066 4970 3374
rect 5054 3369 5082 3374
rect 4998 3066 5026 3071
rect 4942 3065 5026 3066
rect 4942 3039 4999 3065
rect 5025 3039 5026 3065
rect 4942 3038 5026 3039
rect 4998 3033 5026 3038
rect 4830 2977 4858 2982
rect 4998 2954 5026 2959
rect 4673 2758 4805 2763
rect 4701 2730 4725 2758
rect 4753 2730 4777 2758
rect 4673 2725 4805 2730
rect 4998 2673 5026 2926
rect 5054 2954 5082 2959
rect 5110 2954 5138 3710
rect 5254 3150 5386 3155
rect 5282 3122 5306 3150
rect 5334 3122 5358 3150
rect 5254 3117 5386 3122
rect 5054 2953 5138 2954
rect 5054 2927 5055 2953
rect 5081 2927 5138 2953
rect 5054 2926 5138 2927
rect 5054 2921 5082 2926
rect 4998 2647 4999 2673
rect 5025 2647 5026 2673
rect 4998 2641 5026 2647
rect 4606 2529 4634 2534
rect 4942 2562 4970 2567
rect 5054 2562 5082 2567
rect 4970 2561 5082 2562
rect 4970 2535 5055 2561
rect 5081 2535 5082 2561
rect 4970 2534 5082 2535
rect 4662 2505 4690 2511
rect 4662 2479 4663 2505
rect 4689 2479 4690 2505
rect 4662 2450 4690 2479
rect 4718 2450 4746 2455
rect 4662 2422 4718 2450
rect 4326 2417 4354 2422
rect 4718 2403 4746 2422
rect 4092 2366 4224 2371
rect 4120 2338 4144 2366
rect 4172 2338 4196 2366
rect 4092 2333 4224 2338
rect 3878 2226 3906 2231
rect 3878 2179 3906 2198
rect 4214 2226 4242 2231
rect 4214 2170 4242 2198
rect 4214 2169 4354 2170
rect 4214 2143 4215 2169
rect 4241 2143 4354 2169
rect 4214 2142 4354 2143
rect 4214 2137 4242 2142
rect 3822 2025 3850 2030
rect 3934 2058 3962 2063
rect 3710 1863 3711 1889
rect 3737 1863 3738 1889
rect 3710 1857 3738 1863
rect 3934 1890 3962 2030
rect 4270 2057 4298 2063
rect 4270 2031 4271 2057
rect 4297 2031 4298 2057
rect 3990 1890 4018 1895
rect 3934 1889 4018 1890
rect 3934 1863 3991 1889
rect 4017 1863 4018 1889
rect 3934 1862 4018 1863
rect 3654 1751 3655 1777
rect 3681 1751 3682 1777
rect 3654 1745 3682 1751
rect 3990 1834 4018 1862
rect 3990 1778 4018 1806
rect 4270 1834 4298 2031
rect 4270 1801 4298 1806
rect 4046 1778 4074 1783
rect 3990 1777 4074 1778
rect 3990 1751 4047 1777
rect 4073 1751 4074 1777
rect 3990 1750 4074 1751
rect 4046 1745 4074 1750
rect 4326 1777 4354 2142
rect 4673 1974 4805 1979
rect 4701 1946 4725 1974
rect 4753 1946 4777 1974
rect 4673 1941 4805 1946
rect 4382 1834 4410 1839
rect 4382 1787 4410 1806
rect 4326 1751 4327 1777
rect 4353 1751 4354 1777
rect 4326 1745 4354 1751
rect 4942 1722 4970 2534
rect 5054 2529 5082 2534
rect 4998 2450 5026 2455
rect 4998 2170 5026 2422
rect 5110 2450 5138 2926
rect 5110 2417 5138 2422
rect 5254 2366 5386 2371
rect 5282 2338 5306 2366
rect 5334 2338 5358 2366
rect 5254 2333 5386 2338
rect 4998 2169 5082 2170
rect 4998 2143 4999 2169
rect 5025 2143 5082 2169
rect 4998 2142 5082 2143
rect 4998 2137 5026 2142
rect 5054 2057 5082 2142
rect 5054 2031 5055 2057
rect 5081 2031 5082 2057
rect 5054 1834 5082 2031
rect 5054 1787 5082 1806
rect 4998 1722 5026 1727
rect 4942 1721 5026 1722
rect 4942 1695 4999 1721
rect 5025 1695 5026 1721
rect 4942 1694 5026 1695
rect 2870 1675 2898 1694
rect 2310 1633 2338 1638
rect 1768 1582 1900 1587
rect 1796 1554 1820 1582
rect 1848 1554 1872 1582
rect 1768 1549 1900 1554
rect 2930 1582 3062 1587
rect 2958 1554 2982 1582
rect 3010 1554 3034 1582
rect 2930 1549 3062 1554
rect 4092 1582 4224 1587
rect 4120 1554 4144 1582
rect 4172 1554 4196 1582
rect 4092 1549 4224 1554
rect 966 1465 994 1470
rect 4998 658 5026 1694
rect 5254 1582 5386 1587
rect 5282 1554 5306 1582
rect 5334 1554 5358 1582
rect 5254 1549 5386 1554
rect 4998 625 5026 630
<< via2 >>
rect 4942 5334 4970 5362
rect 1187 4325 1215 4326
rect 1187 4299 1188 4325
rect 1188 4299 1214 4325
rect 1214 4299 1215 4325
rect 1187 4298 1215 4299
rect 1239 4325 1267 4326
rect 1239 4299 1240 4325
rect 1240 4299 1266 4325
rect 1266 4299 1267 4325
rect 1239 4298 1267 4299
rect 1291 4325 1319 4326
rect 1291 4299 1292 4325
rect 1292 4299 1318 4325
rect 1318 4299 1319 4325
rect 1291 4298 1319 4299
rect 2349 4325 2377 4326
rect 2349 4299 2350 4325
rect 2350 4299 2376 4325
rect 2376 4299 2377 4325
rect 2349 4298 2377 4299
rect 2401 4325 2429 4326
rect 2401 4299 2402 4325
rect 2402 4299 2428 4325
rect 2428 4299 2429 4325
rect 2401 4298 2429 4299
rect 2453 4325 2481 4326
rect 2453 4299 2454 4325
rect 2454 4299 2480 4325
rect 2480 4299 2481 4325
rect 2453 4298 2481 4299
rect 3511 4325 3539 4326
rect 3511 4299 3512 4325
rect 3512 4299 3538 4325
rect 3538 4299 3539 4325
rect 3511 4298 3539 4299
rect 3563 4325 3591 4326
rect 3563 4299 3564 4325
rect 3564 4299 3590 4325
rect 3590 4299 3591 4325
rect 3563 4298 3591 4299
rect 3615 4325 3643 4326
rect 3615 4299 3616 4325
rect 3616 4299 3642 4325
rect 3642 4299 3643 4325
rect 3615 4298 3643 4299
rect 4673 4325 4701 4326
rect 4673 4299 4674 4325
rect 4674 4299 4700 4325
rect 4700 4299 4701 4325
rect 4673 4298 4701 4299
rect 4725 4325 4753 4326
rect 4725 4299 4726 4325
rect 4726 4299 4752 4325
rect 4752 4299 4753 4325
rect 4725 4298 4753 4299
rect 4777 4325 4805 4326
rect 4777 4299 4778 4325
rect 4778 4299 4804 4325
rect 4804 4299 4805 4325
rect 4777 4298 4805 4299
rect 1134 4158 1162 4186
rect 4886 4158 4914 4186
rect 1768 3933 1796 3934
rect 1768 3907 1769 3933
rect 1769 3907 1795 3933
rect 1795 3907 1796 3933
rect 1768 3906 1796 3907
rect 1820 3933 1848 3934
rect 1820 3907 1821 3933
rect 1821 3907 1847 3933
rect 1847 3907 1848 3933
rect 1820 3906 1848 3907
rect 1872 3933 1900 3934
rect 1872 3907 1873 3933
rect 1873 3907 1899 3933
rect 1899 3907 1900 3933
rect 1872 3906 1900 3907
rect 2930 3933 2958 3934
rect 2930 3907 2931 3933
rect 2931 3907 2957 3933
rect 2957 3907 2958 3933
rect 2930 3906 2958 3907
rect 2982 3933 3010 3934
rect 2982 3907 2983 3933
rect 2983 3907 3009 3933
rect 3009 3907 3010 3933
rect 2982 3906 3010 3907
rect 3034 3933 3062 3934
rect 3034 3907 3035 3933
rect 3035 3907 3061 3933
rect 3061 3907 3062 3933
rect 3034 3906 3062 3907
rect 4092 3933 4120 3934
rect 4092 3907 4093 3933
rect 4093 3907 4119 3933
rect 4119 3907 4120 3933
rect 4092 3906 4120 3907
rect 4144 3933 4172 3934
rect 4144 3907 4145 3933
rect 4145 3907 4171 3933
rect 4171 3907 4172 3933
rect 4144 3906 4172 3907
rect 4196 3933 4224 3934
rect 4196 3907 4197 3933
rect 4197 3907 4223 3933
rect 4223 3907 4224 3933
rect 4196 3906 4224 3907
rect 1187 3541 1215 3542
rect 1187 3515 1188 3541
rect 1188 3515 1214 3541
rect 1214 3515 1215 3541
rect 1187 3514 1215 3515
rect 1239 3541 1267 3542
rect 1239 3515 1240 3541
rect 1240 3515 1266 3541
rect 1266 3515 1267 3541
rect 1239 3514 1267 3515
rect 1291 3541 1319 3542
rect 1291 3515 1292 3541
rect 1292 3515 1318 3541
rect 1318 3515 1319 3541
rect 1291 3514 1319 3515
rect 966 3009 994 3010
rect 966 2983 967 3009
rect 967 2983 993 3009
rect 993 2983 994 3009
rect 966 2982 994 2983
rect 1302 3009 1330 3010
rect 1302 2983 1303 3009
rect 1303 2983 1329 3009
rect 1329 2983 1330 3009
rect 1302 2982 1330 2983
rect 1470 2982 1498 3010
rect 1187 2757 1215 2758
rect 1187 2731 1188 2757
rect 1188 2731 1214 2757
rect 1214 2731 1215 2757
rect 1187 2730 1215 2731
rect 1239 2757 1267 2758
rect 1239 2731 1240 2757
rect 1240 2731 1266 2757
rect 1266 2731 1267 2757
rect 1239 2730 1267 2731
rect 1291 2757 1319 2758
rect 1291 2731 1292 2757
rect 1292 2731 1318 2757
rect 1318 2731 1319 2757
rect 1291 2730 1319 2731
rect 1134 2673 1162 2674
rect 1134 2647 1135 2673
rect 1135 2647 1161 2673
rect 1161 2647 1162 2673
rect 1134 2646 1162 2647
rect 966 2534 994 2562
rect 1302 2646 1330 2674
rect 1078 2561 1106 2562
rect 1078 2535 1079 2561
rect 1079 2535 1105 2561
rect 1105 2535 1106 2561
rect 1078 2534 1106 2535
rect 2349 3541 2377 3542
rect 2349 3515 2350 3541
rect 2350 3515 2376 3541
rect 2376 3515 2377 3541
rect 2349 3514 2377 3515
rect 2401 3541 2429 3542
rect 2401 3515 2402 3541
rect 2402 3515 2428 3541
rect 2428 3515 2429 3541
rect 2401 3514 2429 3515
rect 2453 3541 2481 3542
rect 2453 3515 2454 3541
rect 2454 3515 2480 3541
rect 2480 3515 2481 3541
rect 2453 3514 2481 3515
rect 1768 3149 1796 3150
rect 1768 3123 1769 3149
rect 1769 3123 1795 3149
rect 1795 3123 1796 3149
rect 1768 3122 1796 3123
rect 1820 3149 1848 3150
rect 1820 3123 1821 3149
rect 1821 3123 1847 3149
rect 1847 3123 1848 3149
rect 1820 3122 1848 3123
rect 1872 3149 1900 3150
rect 1872 3123 1873 3149
rect 1873 3123 1899 3149
rect 1899 3123 1900 3149
rect 1872 3122 1900 3123
rect 1582 3009 1610 3010
rect 1582 2983 1583 3009
rect 1583 2983 1609 3009
rect 1609 2983 1610 3009
rect 1582 2982 1610 2983
rect 1750 2982 1778 3010
rect 1470 2673 1498 2674
rect 1470 2647 1471 2673
rect 1471 2647 1497 2673
rect 1497 2647 1498 2673
rect 1470 2646 1498 2647
rect 1414 2561 1442 2562
rect 1414 2535 1415 2561
rect 1415 2535 1441 2561
rect 1441 2535 1442 2561
rect 1414 2534 1442 2535
rect 2870 3289 2898 3290
rect 2870 3263 2871 3289
rect 2871 3263 2897 3289
rect 2897 3263 2898 3289
rect 2870 3262 2898 3263
rect 1918 3009 1946 3010
rect 1918 2983 1919 3009
rect 1919 2983 1945 3009
rect 1945 2983 1946 3009
rect 1918 2982 1946 2983
rect 2142 2982 2170 3010
rect 2030 2814 2058 2842
rect 1638 2534 1666 2562
rect 1806 2561 1834 2562
rect 1806 2535 1807 2561
rect 1807 2535 1833 2561
rect 1833 2535 1834 2561
rect 1806 2534 1834 2535
rect 4606 3598 4634 3626
rect 3511 3541 3539 3542
rect 3511 3515 3512 3541
rect 3512 3515 3538 3541
rect 3538 3515 3539 3541
rect 3511 3514 3539 3515
rect 3563 3541 3591 3542
rect 3563 3515 3564 3541
rect 3564 3515 3590 3541
rect 3590 3515 3591 3541
rect 3563 3514 3591 3515
rect 3615 3541 3643 3542
rect 3615 3515 3616 3541
rect 3616 3515 3642 3541
rect 3642 3515 3643 3541
rect 3615 3514 3643 3515
rect 3094 3262 3122 3290
rect 3206 3289 3234 3290
rect 3206 3263 3207 3289
rect 3207 3263 3233 3289
rect 3233 3263 3234 3289
rect 3206 3262 3234 3263
rect 2310 2841 2338 2842
rect 2310 2815 2311 2841
rect 2311 2815 2337 2841
rect 2337 2815 2338 2841
rect 2310 2814 2338 2815
rect 2590 2814 2618 2842
rect 2349 2757 2377 2758
rect 2349 2731 2350 2757
rect 2350 2731 2376 2757
rect 2376 2731 2377 2757
rect 2349 2730 2377 2731
rect 2401 2757 2429 2758
rect 2401 2731 2402 2757
rect 2402 2731 2428 2757
rect 2428 2731 2429 2757
rect 2401 2730 2429 2731
rect 2453 2757 2481 2758
rect 2453 2731 2454 2757
rect 2454 2731 2480 2757
rect 2480 2731 2481 2757
rect 2453 2730 2481 2731
rect 1768 2365 1796 2366
rect 1768 2339 1769 2365
rect 1769 2339 1795 2365
rect 1795 2339 1796 2365
rect 1768 2338 1796 2339
rect 1820 2365 1848 2366
rect 1820 2339 1821 2365
rect 1821 2339 1847 2365
rect 1847 2339 1848 2365
rect 1820 2338 1848 2339
rect 1872 2365 1900 2366
rect 1872 2339 1873 2365
rect 1873 2339 1899 2365
rect 1899 2339 1900 2365
rect 1872 2338 1900 2339
rect 1187 1973 1215 1974
rect 1187 1947 1188 1973
rect 1188 1947 1214 1973
rect 1214 1947 1215 1973
rect 1187 1946 1215 1947
rect 1239 1973 1267 1974
rect 1239 1947 1240 1973
rect 1240 1947 1266 1973
rect 1266 1947 1267 1973
rect 1239 1946 1267 1947
rect 1291 1973 1319 1974
rect 1291 1947 1292 1973
rect 1292 1947 1318 1973
rect 1318 1947 1319 1973
rect 1291 1946 1319 1947
rect 1302 1721 1330 1722
rect 1302 1695 1303 1721
rect 1303 1695 1329 1721
rect 1329 1695 1330 1721
rect 1302 1694 1330 1695
rect 3542 3289 3570 3290
rect 3542 3263 3543 3289
rect 3543 3263 3569 3289
rect 3569 3263 3570 3289
rect 3542 3262 3570 3263
rect 2930 3149 2958 3150
rect 2930 3123 2931 3149
rect 2931 3123 2957 3149
rect 2957 3123 2958 3149
rect 2930 3122 2958 3123
rect 2982 3149 3010 3150
rect 2982 3123 2983 3149
rect 2983 3123 3009 3149
rect 3009 3123 3010 3149
rect 2982 3122 3010 3123
rect 3034 3149 3062 3150
rect 3034 3123 3035 3149
rect 3035 3123 3061 3149
rect 3061 3123 3062 3149
rect 3034 3122 3062 3123
rect 2926 3009 2954 3010
rect 2926 2983 2927 3009
rect 2927 2983 2953 3009
rect 2953 2983 2954 3009
rect 2926 2982 2954 2983
rect 4092 3149 4120 3150
rect 4092 3123 4093 3149
rect 4093 3123 4119 3149
rect 4119 3123 4120 3149
rect 4092 3122 4120 3123
rect 4144 3149 4172 3150
rect 4144 3123 4145 3149
rect 4145 3123 4171 3149
rect 4171 3123 4172 3149
rect 4144 3122 4172 3123
rect 4196 3149 4224 3150
rect 4196 3123 4197 3149
rect 4197 3123 4223 3149
rect 4223 3123 4224 3149
rect 4196 3122 4224 3123
rect 3878 3009 3906 3010
rect 3878 2983 3879 3009
rect 3879 2983 3905 3009
rect 3905 2983 3906 3009
rect 3878 2982 3906 2983
rect 4158 2982 4186 3010
rect 3934 2841 3962 2842
rect 3934 2815 3935 2841
rect 3935 2815 3961 2841
rect 3961 2815 3962 2841
rect 3934 2814 3962 2815
rect 3511 2757 3539 2758
rect 3511 2731 3512 2757
rect 3512 2731 3538 2757
rect 3538 2731 3539 2757
rect 3511 2730 3539 2731
rect 3563 2757 3591 2758
rect 3563 2731 3564 2757
rect 3564 2731 3590 2757
rect 3590 2731 3591 2757
rect 3563 2730 3591 2731
rect 3615 2757 3643 2758
rect 3615 2731 3616 2757
rect 3616 2731 3642 2757
rect 3642 2731 3643 2757
rect 3615 2730 3643 2731
rect 2982 2646 3010 2674
rect 3542 2673 3570 2674
rect 3542 2647 3543 2673
rect 3543 2647 3569 2673
rect 3569 2647 3570 2673
rect 3542 2646 3570 2647
rect 3878 2673 3906 2674
rect 3878 2647 3879 2673
rect 3879 2647 3905 2673
rect 3905 2647 3906 2673
rect 3878 2646 3906 2647
rect 966 1638 994 1666
rect 1694 1638 1722 1666
rect 2930 2365 2958 2366
rect 2930 2339 2931 2365
rect 2931 2339 2957 2365
rect 2957 2339 2958 2365
rect 2930 2338 2958 2339
rect 2982 2365 3010 2366
rect 2982 2339 2983 2365
rect 2983 2339 3009 2365
rect 3009 2339 3010 2365
rect 2982 2338 3010 2339
rect 3034 2365 3062 2366
rect 3034 2339 3035 2365
rect 3035 2339 3061 2365
rect 3061 2339 3062 2365
rect 3034 2338 3062 2339
rect 4270 2841 4298 2842
rect 4270 2815 4271 2841
rect 4271 2815 4297 2841
rect 4297 2815 4298 2841
rect 4270 2814 4298 2815
rect 4214 2561 4242 2562
rect 4214 2535 4215 2561
rect 4215 2535 4241 2561
rect 4241 2535 4242 2561
rect 4214 2534 4242 2535
rect 2870 2198 2898 2226
rect 2349 1973 2377 1974
rect 2349 1947 2350 1973
rect 2350 1947 2376 1973
rect 2376 1947 2377 1973
rect 2349 1946 2377 1947
rect 2401 1973 2429 1974
rect 2401 1947 2402 1973
rect 2402 1947 2428 1973
rect 2428 1947 2429 1973
rect 2401 1946 2429 1947
rect 2453 1973 2481 1974
rect 2453 1947 2454 1973
rect 2454 1947 2480 1973
rect 2480 1947 2481 1973
rect 2453 1946 2481 1947
rect 2926 2057 2954 2058
rect 2926 2031 2927 2057
rect 2927 2031 2953 2057
rect 2953 2031 2954 2057
rect 2926 2030 2954 2031
rect 3710 2030 3738 2058
rect 3511 1973 3539 1974
rect 3511 1947 3512 1973
rect 3512 1947 3538 1973
rect 3538 1947 3539 1973
rect 3511 1946 3539 1947
rect 3563 1973 3591 1974
rect 3563 1947 3564 1973
rect 3564 1947 3590 1973
rect 3590 1947 3591 1973
rect 3563 1946 3591 1947
rect 3615 1973 3643 1974
rect 3615 1947 3616 1973
rect 3616 1947 3642 1973
rect 3642 1947 3643 1973
rect 3615 1946 3643 1947
rect 1974 1638 2002 1666
rect 4673 3541 4701 3542
rect 4673 3515 4674 3541
rect 4674 3515 4700 3541
rect 4700 3515 4701 3541
rect 4673 3514 4701 3515
rect 4725 3541 4753 3542
rect 4725 3515 4726 3541
rect 4726 3515 4752 3541
rect 4752 3515 4753 3541
rect 4725 3514 4753 3515
rect 4777 3541 4805 3542
rect 4777 3515 4778 3541
rect 4778 3515 4804 3541
rect 4804 3515 4805 3541
rect 4777 3514 4805 3515
rect 5254 3933 5282 3934
rect 5254 3907 5255 3933
rect 5255 3907 5281 3933
rect 5281 3907 5282 3933
rect 5254 3906 5282 3907
rect 5306 3933 5334 3934
rect 5306 3907 5307 3933
rect 5307 3907 5333 3933
rect 5333 3907 5334 3933
rect 5306 3906 5334 3907
rect 5358 3933 5386 3934
rect 5358 3907 5359 3933
rect 5359 3907 5385 3933
rect 5385 3907 5386 3933
rect 5358 3906 5386 3907
rect 4998 3625 5026 3626
rect 4998 3599 4999 3625
rect 4999 3599 5025 3625
rect 5025 3599 5026 3625
rect 4998 3598 5026 3599
rect 4830 2982 4858 3010
rect 4998 2926 5026 2954
rect 4673 2757 4701 2758
rect 4673 2731 4674 2757
rect 4674 2731 4700 2757
rect 4700 2731 4701 2757
rect 4673 2730 4701 2731
rect 4725 2757 4753 2758
rect 4725 2731 4726 2757
rect 4726 2731 4752 2757
rect 4752 2731 4753 2757
rect 4725 2730 4753 2731
rect 4777 2757 4805 2758
rect 4777 2731 4778 2757
rect 4778 2731 4804 2757
rect 4804 2731 4805 2757
rect 4777 2730 4805 2731
rect 5254 3149 5282 3150
rect 5254 3123 5255 3149
rect 5255 3123 5281 3149
rect 5281 3123 5282 3149
rect 5254 3122 5282 3123
rect 5306 3149 5334 3150
rect 5306 3123 5307 3149
rect 5307 3123 5333 3149
rect 5333 3123 5334 3149
rect 5306 3122 5334 3123
rect 5358 3149 5386 3150
rect 5358 3123 5359 3149
rect 5359 3123 5385 3149
rect 5385 3123 5386 3149
rect 5358 3122 5386 3123
rect 4606 2534 4634 2562
rect 4942 2534 4970 2562
rect 4326 2422 4354 2450
rect 4718 2449 4746 2450
rect 4718 2423 4719 2449
rect 4719 2423 4745 2449
rect 4745 2423 4746 2449
rect 4718 2422 4746 2423
rect 4092 2365 4120 2366
rect 4092 2339 4093 2365
rect 4093 2339 4119 2365
rect 4119 2339 4120 2365
rect 4092 2338 4120 2339
rect 4144 2365 4172 2366
rect 4144 2339 4145 2365
rect 4145 2339 4171 2365
rect 4171 2339 4172 2365
rect 4144 2338 4172 2339
rect 4196 2365 4224 2366
rect 4196 2339 4197 2365
rect 4197 2339 4223 2365
rect 4223 2339 4224 2365
rect 4196 2338 4224 2339
rect 3878 2225 3906 2226
rect 3878 2199 3879 2225
rect 3879 2199 3905 2225
rect 3905 2199 3906 2225
rect 3878 2198 3906 2199
rect 4214 2198 4242 2226
rect 3822 2030 3850 2058
rect 3934 2057 3962 2058
rect 3934 2031 3935 2057
rect 3935 2031 3961 2057
rect 3961 2031 3962 2057
rect 3934 2030 3962 2031
rect 3990 1806 4018 1834
rect 4270 1806 4298 1834
rect 4673 1973 4701 1974
rect 4673 1947 4674 1973
rect 4674 1947 4700 1973
rect 4700 1947 4701 1973
rect 4673 1946 4701 1947
rect 4725 1973 4753 1974
rect 4725 1947 4726 1973
rect 4726 1947 4752 1973
rect 4752 1947 4753 1973
rect 4725 1946 4753 1947
rect 4777 1973 4805 1974
rect 4777 1947 4778 1973
rect 4778 1947 4804 1973
rect 4804 1947 4805 1973
rect 4777 1946 4805 1947
rect 4382 1833 4410 1834
rect 4382 1807 4383 1833
rect 4383 1807 4409 1833
rect 4409 1807 4410 1833
rect 4382 1806 4410 1807
rect 2870 1721 2898 1722
rect 2870 1695 2871 1721
rect 2871 1695 2897 1721
rect 2897 1695 2898 1721
rect 2870 1694 2898 1695
rect 4998 2422 5026 2450
rect 5110 2422 5138 2450
rect 5254 2365 5282 2366
rect 5254 2339 5255 2365
rect 5255 2339 5281 2365
rect 5281 2339 5282 2365
rect 5254 2338 5282 2339
rect 5306 2365 5334 2366
rect 5306 2339 5307 2365
rect 5307 2339 5333 2365
rect 5333 2339 5334 2365
rect 5306 2338 5334 2339
rect 5358 2365 5386 2366
rect 5358 2339 5359 2365
rect 5359 2339 5385 2365
rect 5385 2339 5386 2365
rect 5358 2338 5386 2339
rect 5054 1833 5082 1834
rect 5054 1807 5055 1833
rect 5055 1807 5081 1833
rect 5081 1807 5082 1833
rect 5054 1806 5082 1807
rect 2310 1638 2338 1666
rect 1768 1581 1796 1582
rect 1768 1555 1769 1581
rect 1769 1555 1795 1581
rect 1795 1555 1796 1581
rect 1768 1554 1796 1555
rect 1820 1581 1848 1582
rect 1820 1555 1821 1581
rect 1821 1555 1847 1581
rect 1847 1555 1848 1581
rect 1820 1554 1848 1555
rect 1872 1581 1900 1582
rect 1872 1555 1873 1581
rect 1873 1555 1899 1581
rect 1899 1555 1900 1581
rect 1872 1554 1900 1555
rect 2930 1581 2958 1582
rect 2930 1555 2931 1581
rect 2931 1555 2957 1581
rect 2957 1555 2958 1581
rect 2930 1554 2958 1555
rect 2982 1581 3010 1582
rect 2982 1555 2983 1581
rect 2983 1555 3009 1581
rect 3009 1555 3010 1581
rect 2982 1554 3010 1555
rect 3034 1581 3062 1582
rect 3034 1555 3035 1581
rect 3035 1555 3061 1581
rect 3061 1555 3062 1581
rect 3034 1554 3062 1555
rect 4092 1581 4120 1582
rect 4092 1555 4093 1581
rect 4093 1555 4119 1581
rect 4119 1555 4120 1581
rect 4092 1554 4120 1555
rect 4144 1581 4172 1582
rect 4144 1555 4145 1581
rect 4145 1555 4171 1581
rect 4171 1555 4172 1581
rect 4144 1554 4172 1555
rect 4196 1581 4224 1582
rect 4196 1555 4197 1581
rect 4197 1555 4223 1581
rect 4223 1555 4224 1581
rect 4196 1554 4224 1555
rect 966 1470 994 1498
rect 5254 1581 5282 1582
rect 5254 1555 5255 1581
rect 5255 1555 5281 1581
rect 5281 1555 5282 1581
rect 5254 1554 5282 1555
rect 5306 1581 5334 1582
rect 5306 1555 5307 1581
rect 5307 1555 5333 1581
rect 5333 1555 5334 1581
rect 5306 1554 5334 1555
rect 5358 1581 5386 1582
rect 5358 1555 5359 1581
rect 5359 1555 5385 1581
rect 5385 1555 5386 1581
rect 5358 1554 5386 1555
rect 4998 630 5026 658
<< metal3 >>
rect 5600 5362 6000 5376
rect 4937 5334 4942 5362
rect 4970 5334 6000 5362
rect 5600 5320 6000 5334
rect 0 4466 400 4480
rect 0 4438 658 4466
rect 0 4424 400 4438
rect 630 4242 658 4438
rect 1182 4298 1187 4326
rect 1215 4298 1239 4326
rect 1267 4298 1291 4326
rect 1319 4298 1324 4326
rect 2344 4298 2349 4326
rect 2377 4298 2401 4326
rect 2429 4298 2453 4326
rect 2481 4298 2486 4326
rect 3506 4298 3511 4326
rect 3539 4298 3563 4326
rect 3591 4298 3615 4326
rect 3643 4298 3648 4326
rect 4668 4298 4673 4326
rect 4701 4298 4725 4326
rect 4753 4298 4777 4326
rect 4805 4298 4810 4326
rect 630 4214 1162 4242
rect 1134 4186 1162 4214
rect 5600 4186 6000 4200
rect 1129 4158 1134 4186
rect 1162 4158 1167 4186
rect 4881 4158 4886 4186
rect 4914 4158 6000 4186
rect 5600 4144 6000 4158
rect 1763 3906 1768 3934
rect 1796 3906 1820 3934
rect 1848 3906 1872 3934
rect 1900 3906 1905 3934
rect 2925 3906 2930 3934
rect 2958 3906 2982 3934
rect 3010 3906 3034 3934
rect 3062 3906 3067 3934
rect 4087 3906 4092 3934
rect 4120 3906 4144 3934
rect 4172 3906 4196 3934
rect 4224 3906 4229 3934
rect 5249 3906 5254 3934
rect 5282 3906 5306 3934
rect 5334 3906 5358 3934
rect 5386 3906 5391 3934
rect 4601 3598 4606 3626
rect 4634 3598 4998 3626
rect 5026 3598 5031 3626
rect 1182 3514 1187 3542
rect 1215 3514 1239 3542
rect 1267 3514 1291 3542
rect 1319 3514 1324 3542
rect 2344 3514 2349 3542
rect 2377 3514 2401 3542
rect 2429 3514 2453 3542
rect 2481 3514 2486 3542
rect 3506 3514 3511 3542
rect 3539 3514 3563 3542
rect 3591 3514 3615 3542
rect 3643 3514 3648 3542
rect 4668 3514 4673 3542
rect 4701 3514 4725 3542
rect 4753 3514 4777 3542
rect 4805 3514 4810 3542
rect 2865 3262 2870 3290
rect 2898 3262 3094 3290
rect 3122 3262 3206 3290
rect 3234 3262 3542 3290
rect 3570 3262 3575 3290
rect 1763 3122 1768 3150
rect 1796 3122 1820 3150
rect 1848 3122 1872 3150
rect 1900 3122 1905 3150
rect 2925 3122 2930 3150
rect 2958 3122 2982 3150
rect 3010 3122 3034 3150
rect 3062 3122 3067 3150
rect 4087 3122 4092 3150
rect 4120 3122 4144 3150
rect 4172 3122 4196 3150
rect 4224 3122 4229 3150
rect 5249 3122 5254 3150
rect 5282 3122 5306 3150
rect 5334 3122 5358 3150
rect 5386 3122 5391 3150
rect 5600 3010 6000 3024
rect 961 2982 966 3010
rect 994 2982 1302 3010
rect 1330 2982 1470 3010
rect 1498 2982 1582 3010
rect 1610 2982 1750 3010
rect 1778 2982 1918 3010
rect 1946 2982 2142 3010
rect 2170 2982 2926 3010
rect 2954 2982 3878 3010
rect 3906 2982 4158 3010
rect 4186 2982 4191 3010
rect 4825 2982 4830 3010
rect 4858 2982 6000 3010
rect 4998 2954 5026 2982
rect 5600 2968 6000 2982
rect 4993 2926 4998 2954
rect 5026 2926 5031 2954
rect 2025 2814 2030 2842
rect 2058 2814 2310 2842
rect 2338 2814 2590 2842
rect 2618 2814 2623 2842
rect 3929 2814 3934 2842
rect 3962 2814 4270 2842
rect 4298 2814 4303 2842
rect 1182 2730 1187 2758
rect 1215 2730 1239 2758
rect 1267 2730 1291 2758
rect 1319 2730 1324 2758
rect 2344 2730 2349 2758
rect 2377 2730 2401 2758
rect 2429 2730 2453 2758
rect 2481 2730 2486 2758
rect 3506 2730 3511 2758
rect 3539 2730 3563 2758
rect 3591 2730 3615 2758
rect 3643 2730 3648 2758
rect 4668 2730 4673 2758
rect 4701 2730 4725 2758
rect 4753 2730 4777 2758
rect 4805 2730 4810 2758
rect 1129 2646 1134 2674
rect 1162 2646 1302 2674
rect 1330 2646 1470 2674
rect 1498 2646 1503 2674
rect 2977 2646 2982 2674
rect 3010 2646 3542 2674
rect 3570 2646 3878 2674
rect 3906 2646 3911 2674
rect 961 2534 966 2562
rect 994 2534 1078 2562
rect 1106 2534 1414 2562
rect 1442 2534 1638 2562
rect 1666 2534 1806 2562
rect 1834 2534 1839 2562
rect 4209 2534 4214 2562
rect 4242 2534 4606 2562
rect 4634 2534 4942 2562
rect 4970 2534 4975 2562
rect 4321 2422 4326 2450
rect 4354 2422 4718 2450
rect 4746 2422 4998 2450
rect 5026 2422 5110 2450
rect 5138 2422 5143 2450
rect 1763 2338 1768 2366
rect 1796 2338 1820 2366
rect 1848 2338 1872 2366
rect 1900 2338 1905 2366
rect 2925 2338 2930 2366
rect 2958 2338 2982 2366
rect 3010 2338 3034 2366
rect 3062 2338 3067 2366
rect 4087 2338 4092 2366
rect 4120 2338 4144 2366
rect 4172 2338 4196 2366
rect 4224 2338 4229 2366
rect 5249 2338 5254 2366
rect 5282 2338 5306 2366
rect 5334 2338 5358 2366
rect 5386 2338 5391 2366
rect 2865 2198 2870 2226
rect 2898 2198 3878 2226
rect 3906 2198 4214 2226
rect 4242 2198 4247 2226
rect 2921 2030 2926 2058
rect 2954 2030 3710 2058
rect 3738 2030 3822 2058
rect 3850 2030 3934 2058
rect 3962 2030 3967 2058
rect 1182 1946 1187 1974
rect 1215 1946 1239 1974
rect 1267 1946 1291 1974
rect 1319 1946 1324 1974
rect 2344 1946 2349 1974
rect 2377 1946 2401 1974
rect 2429 1946 2453 1974
rect 2481 1946 2486 1974
rect 3506 1946 3511 1974
rect 3539 1946 3563 1974
rect 3591 1946 3615 1974
rect 3643 1946 3648 1974
rect 4668 1946 4673 1974
rect 4701 1946 4725 1974
rect 4753 1946 4777 1974
rect 4805 1946 4810 1974
rect 5600 1834 6000 1848
rect 3985 1806 3990 1834
rect 4018 1806 4270 1834
rect 4298 1806 4382 1834
rect 4410 1806 5054 1834
rect 5082 1806 6000 1834
rect 5600 1792 6000 1806
rect 1297 1694 1302 1722
rect 1330 1694 1335 1722
rect 2478 1694 2870 1722
rect 2898 1694 2903 1722
rect 1302 1666 1330 1694
rect 2478 1666 2506 1694
rect 961 1638 966 1666
rect 994 1638 1694 1666
rect 1722 1638 1974 1666
rect 2002 1638 2310 1666
rect 2338 1638 2506 1666
rect 1763 1554 1768 1582
rect 1796 1554 1820 1582
rect 1848 1554 1872 1582
rect 1900 1554 1905 1582
rect 2925 1554 2930 1582
rect 2958 1554 2982 1582
rect 3010 1554 3034 1582
rect 3062 1554 3067 1582
rect 4087 1554 4092 1582
rect 4120 1554 4144 1582
rect 4172 1554 4196 1582
rect 4224 1554 4229 1582
rect 5249 1554 5254 1582
rect 5282 1554 5306 1582
rect 5334 1554 5358 1582
rect 5386 1554 5391 1582
rect 0 1498 400 1512
rect 0 1470 966 1498
rect 994 1470 999 1498
rect 0 1456 400 1470
rect 5600 658 6000 672
rect 4993 630 4998 658
rect 5026 630 6000 658
rect 5600 616 6000 630
<< via3 >>
rect 1187 4298 1215 4326
rect 1239 4298 1267 4326
rect 1291 4298 1319 4326
rect 2349 4298 2377 4326
rect 2401 4298 2429 4326
rect 2453 4298 2481 4326
rect 3511 4298 3539 4326
rect 3563 4298 3591 4326
rect 3615 4298 3643 4326
rect 4673 4298 4701 4326
rect 4725 4298 4753 4326
rect 4777 4298 4805 4326
rect 1768 3906 1796 3934
rect 1820 3906 1848 3934
rect 1872 3906 1900 3934
rect 2930 3906 2958 3934
rect 2982 3906 3010 3934
rect 3034 3906 3062 3934
rect 4092 3906 4120 3934
rect 4144 3906 4172 3934
rect 4196 3906 4224 3934
rect 5254 3906 5282 3934
rect 5306 3906 5334 3934
rect 5358 3906 5386 3934
rect 1187 3514 1215 3542
rect 1239 3514 1267 3542
rect 1291 3514 1319 3542
rect 2349 3514 2377 3542
rect 2401 3514 2429 3542
rect 2453 3514 2481 3542
rect 3511 3514 3539 3542
rect 3563 3514 3591 3542
rect 3615 3514 3643 3542
rect 4673 3514 4701 3542
rect 4725 3514 4753 3542
rect 4777 3514 4805 3542
rect 1768 3122 1796 3150
rect 1820 3122 1848 3150
rect 1872 3122 1900 3150
rect 2930 3122 2958 3150
rect 2982 3122 3010 3150
rect 3034 3122 3062 3150
rect 4092 3122 4120 3150
rect 4144 3122 4172 3150
rect 4196 3122 4224 3150
rect 5254 3122 5282 3150
rect 5306 3122 5334 3150
rect 5358 3122 5386 3150
rect 1187 2730 1215 2758
rect 1239 2730 1267 2758
rect 1291 2730 1319 2758
rect 2349 2730 2377 2758
rect 2401 2730 2429 2758
rect 2453 2730 2481 2758
rect 3511 2730 3539 2758
rect 3563 2730 3591 2758
rect 3615 2730 3643 2758
rect 4673 2730 4701 2758
rect 4725 2730 4753 2758
rect 4777 2730 4805 2758
rect 1768 2338 1796 2366
rect 1820 2338 1848 2366
rect 1872 2338 1900 2366
rect 2930 2338 2958 2366
rect 2982 2338 3010 2366
rect 3034 2338 3062 2366
rect 4092 2338 4120 2366
rect 4144 2338 4172 2366
rect 4196 2338 4224 2366
rect 5254 2338 5282 2366
rect 5306 2338 5334 2366
rect 5358 2338 5386 2366
rect 1187 1946 1215 1974
rect 1239 1946 1267 1974
rect 1291 1946 1319 1974
rect 2349 1946 2377 1974
rect 2401 1946 2429 1974
rect 2453 1946 2481 1974
rect 3511 1946 3539 1974
rect 3563 1946 3591 1974
rect 3615 1946 3643 1974
rect 4673 1946 4701 1974
rect 4725 1946 4753 1974
rect 4777 1946 4805 1974
rect 1768 1554 1796 1582
rect 1820 1554 1848 1582
rect 1872 1554 1900 1582
rect 2930 1554 2958 1582
rect 2982 1554 3010 1582
rect 3034 1554 3062 1582
rect 4092 1554 4120 1582
rect 4144 1554 4172 1582
rect 4196 1554 4224 1582
rect 5254 1554 5282 1582
rect 5306 1554 5334 1582
rect 5358 1554 5386 1582
<< metal4 >>
rect 1173 4326 1333 4342
rect 1173 4298 1187 4326
rect 1215 4298 1239 4326
rect 1267 4298 1291 4326
rect 1319 4298 1333 4326
rect 1173 3542 1333 4298
rect 1173 3514 1187 3542
rect 1215 3514 1239 3542
rect 1267 3514 1291 3542
rect 1319 3514 1333 3542
rect 1173 2758 1333 3514
rect 1173 2730 1187 2758
rect 1215 2730 1239 2758
rect 1267 2730 1291 2758
rect 1319 2730 1333 2758
rect 1173 1974 1333 2730
rect 1173 1946 1187 1974
rect 1215 1946 1239 1974
rect 1267 1946 1291 1974
rect 1319 1946 1333 1974
rect 1173 1538 1333 1946
rect 1754 3934 1914 4342
rect 1754 3906 1768 3934
rect 1796 3906 1820 3934
rect 1848 3906 1872 3934
rect 1900 3906 1914 3934
rect 1754 3150 1914 3906
rect 1754 3122 1768 3150
rect 1796 3122 1820 3150
rect 1848 3122 1872 3150
rect 1900 3122 1914 3150
rect 1754 2366 1914 3122
rect 1754 2338 1768 2366
rect 1796 2338 1820 2366
rect 1848 2338 1872 2366
rect 1900 2338 1914 2366
rect 1754 1582 1914 2338
rect 1754 1554 1768 1582
rect 1796 1554 1820 1582
rect 1848 1554 1872 1582
rect 1900 1554 1914 1582
rect 1754 1538 1914 1554
rect 2335 4326 2495 4342
rect 2335 4298 2349 4326
rect 2377 4298 2401 4326
rect 2429 4298 2453 4326
rect 2481 4298 2495 4326
rect 2335 3542 2495 4298
rect 2335 3514 2349 3542
rect 2377 3514 2401 3542
rect 2429 3514 2453 3542
rect 2481 3514 2495 3542
rect 2335 2758 2495 3514
rect 2335 2730 2349 2758
rect 2377 2730 2401 2758
rect 2429 2730 2453 2758
rect 2481 2730 2495 2758
rect 2335 1974 2495 2730
rect 2335 1946 2349 1974
rect 2377 1946 2401 1974
rect 2429 1946 2453 1974
rect 2481 1946 2495 1974
rect 2335 1538 2495 1946
rect 2916 3934 3076 4342
rect 2916 3906 2930 3934
rect 2958 3906 2982 3934
rect 3010 3906 3034 3934
rect 3062 3906 3076 3934
rect 2916 3150 3076 3906
rect 2916 3122 2930 3150
rect 2958 3122 2982 3150
rect 3010 3122 3034 3150
rect 3062 3122 3076 3150
rect 2916 2366 3076 3122
rect 2916 2338 2930 2366
rect 2958 2338 2982 2366
rect 3010 2338 3034 2366
rect 3062 2338 3076 2366
rect 2916 1582 3076 2338
rect 2916 1554 2930 1582
rect 2958 1554 2982 1582
rect 3010 1554 3034 1582
rect 3062 1554 3076 1582
rect 2916 1538 3076 1554
rect 3497 4326 3657 4342
rect 3497 4298 3511 4326
rect 3539 4298 3563 4326
rect 3591 4298 3615 4326
rect 3643 4298 3657 4326
rect 3497 3542 3657 4298
rect 3497 3514 3511 3542
rect 3539 3514 3563 3542
rect 3591 3514 3615 3542
rect 3643 3514 3657 3542
rect 3497 2758 3657 3514
rect 3497 2730 3511 2758
rect 3539 2730 3563 2758
rect 3591 2730 3615 2758
rect 3643 2730 3657 2758
rect 3497 1974 3657 2730
rect 3497 1946 3511 1974
rect 3539 1946 3563 1974
rect 3591 1946 3615 1974
rect 3643 1946 3657 1974
rect 3497 1538 3657 1946
rect 4078 3934 4238 4342
rect 4078 3906 4092 3934
rect 4120 3906 4144 3934
rect 4172 3906 4196 3934
rect 4224 3906 4238 3934
rect 4078 3150 4238 3906
rect 4078 3122 4092 3150
rect 4120 3122 4144 3150
rect 4172 3122 4196 3150
rect 4224 3122 4238 3150
rect 4078 2366 4238 3122
rect 4078 2338 4092 2366
rect 4120 2338 4144 2366
rect 4172 2338 4196 2366
rect 4224 2338 4238 2366
rect 4078 1582 4238 2338
rect 4078 1554 4092 1582
rect 4120 1554 4144 1582
rect 4172 1554 4196 1582
rect 4224 1554 4238 1582
rect 4078 1538 4238 1554
rect 4659 4326 4819 4342
rect 4659 4298 4673 4326
rect 4701 4298 4725 4326
rect 4753 4298 4777 4326
rect 4805 4298 4819 4326
rect 4659 3542 4819 4298
rect 4659 3514 4673 3542
rect 4701 3514 4725 3542
rect 4753 3514 4777 3542
rect 4805 3514 4819 3542
rect 4659 2758 4819 3514
rect 4659 2730 4673 2758
rect 4701 2730 4725 2758
rect 4753 2730 4777 2758
rect 4805 2730 4819 2758
rect 4659 1974 4819 2730
rect 4659 1946 4673 1974
rect 4701 1946 4725 1974
rect 4753 1946 4777 1974
rect 4805 1946 4819 1974
rect 4659 1538 4819 1946
rect 5240 3934 5400 4342
rect 5240 3906 5254 3934
rect 5282 3906 5306 3934
rect 5334 3906 5358 3934
rect 5386 3906 5400 3934
rect 5240 3150 5400 3906
rect 5240 3122 5254 3150
rect 5282 3122 5306 3150
rect 5334 3122 5358 3150
rect 5386 3122 5400 3150
rect 5240 2366 5400 3122
rect 5240 2338 5254 2366
rect 5282 2338 5306 2366
rect 5334 2338 5358 2366
rect 5386 2338 5400 2366
rect 5240 1582 5400 2338
rect 5240 1554 5254 1582
rect 5282 1554 5306 1582
rect 5334 1554 5358 1582
rect 5386 1554 5400 1582
rect 5240 1538 5400 1554
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8
timestamp 1667941163
transform 1 0 1120 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14
timestamp 1667941163
transform 1 0 1456 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20
timestamp 1667941163
transform 1 0 1792 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 2128 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32
timestamp 1667941163
transform 1 0 2464 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 3024 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50
timestamp 1667941163
transform 1 0 3472 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56
timestamp 1667941163
transform 1 0 3808 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62
timestamp 1667941163
transform 1 0 4144 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1667941163
transform 1 0 4480 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80
timestamp 1667941163
transform 1 0 5152 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_2
timestamp 1667941163
transform 1 0 784 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_8
timestamp 1667941163
transform 1 0 1120 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_14
timestamp 1667941163
transform 1 0 1456 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_20
timestamp 1667941163
transform 1 0 1792 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_26
timestamp 1667941163
transform 1 0 2128 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_32
timestamp 1667941163
transform 1 0 2464 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_36
timestamp 1667941163
transform 1 0 2688 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1667941163
transform 1 0 3024 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_48
timestamp 1667941163
transform 1 0 3360 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 3696 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_60
timestamp 1667941163
transform 1 0 4032 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_75
timestamp 1667941163
transform 1 0 4872 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_80
timestamp 1667941163
transform 1 0 5152 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_10
timestamp 1667941163
transform 1 0 1232 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_16
timestamp 1667941163
transform 1 0 1568 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_22
timestamp 1667941163
transform 1 0 1904 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_28
timestamp 1667941163
transform 1 0 2240 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_42
timestamp 1667941163
transform 1 0 3024 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_46
timestamp 1667941163
transform 1 0 3248 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_48
timestamp 1667941163
transform 1 0 3360 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_53
timestamp 1667941163
transform 1 0 3640 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_59
timestamp 1667941163
transform 1 0 3976 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_65
timestamp 1667941163
transform 1 0 4312 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_69
timestamp 1667941163
transform 1 0 4536 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_74
timestamp 1667941163
transform 1 0 4816 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_80
timestamp 1667941163
transform 1 0 5152 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_7
timestamp 1667941163
transform 1 0 1064 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_13
timestamp 1667941163
transform 1 0 1400 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_19
timestamp 1667941163
transform 1 0 1736 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_25
timestamp 1667941163
transform 1 0 2072 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_31
timestamp 1667941163
transform 1 0 2408 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_37
timestamp 1667941163
transform 1 0 2744 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_43
timestamp 1667941163
transform 1 0 3080 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_49
timestamp 1667941163
transform 1 0 3416 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_53
timestamp 1667941163
transform 1 0 3640 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 3752 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_60
timestamp 1667941163
transform 1 0 4032 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1667941163
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_75
timestamp 1667941163
transform 1 0 4872 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_80
timestamp 1667941163
transform 1 0 5152 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_8
timestamp 1667941163
transform 1 0 1120 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1667941163
transform 1 0 1456 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_20
timestamp 1667941163
transform 1 0 1792 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 2128 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_32
timestamp 1667941163
transform 1 0 2464 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_42
timestamp 1667941163
transform 1 0 3024 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_48
timestamp 1667941163
transform 1 0 3360 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_54 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 3696 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_66
timestamp 1667941163
transform 1 0 4368 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_80
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_10
timestamp 1667941163
transform 1 0 1232 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_16
timestamp 1667941163
transform 1 0 1568 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_22
timestamp 1667941163
transform 1 0 1904 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_28
timestamp 1667941163
transform 1 0 2240 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_34
timestamp 1667941163
transform 1 0 2576 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_40
timestamp 1667941163
transform 1 0 2912 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_46 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 3248 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_62
timestamp 1667941163
transform 1 0 4144 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_75
timestamp 1667941163
transform 1 0 4872 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_80
timestamp 1667941163
transform 1 0 5152 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_10
timestamp 1667941163
transform 1 0 1232 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_16
timestamp 1667941163
transform 1 0 1568 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_22
timestamp 1667941163
transform 1 0 1904 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_28
timestamp 1667941163
transform 1 0 2240 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_37 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_69
timestamp 1667941163
transform 1 0 4536 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_72
timestamp 1667941163
transform 1 0 4704 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_80
timestamp 1667941163
transform 1 0 5152 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 5320 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 5320 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 5320 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 5320 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 5320 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 5320 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 5320 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_14 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_15
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_16
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_17
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1667941163
transform 1 0 4592 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  oinvn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 5152 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  oinvp
timestamp 1667941163
transform -1 0 5152 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  oxor pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 4480 0 1 3136
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 4928 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 3416 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 4592 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 3472 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 4144 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 3136 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[3\].fbn
timestamp 1667941163
transform -1 0 4144 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 3248 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 4256 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 3808 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 4144 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 4088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 2800 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 2856 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 3808 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 4144 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 3584 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 3752 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 4928 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_amp.gen_X\[1\].crossp
timestamp 1667941163
transform -1 0 5152 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 3472 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 1680 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 3192 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 1568 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 2800 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 2016 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 2184 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 2352 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 1568 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 2352 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[1\].thrun
timestamp 1667941163
transform -1 0 2912 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 1176 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 1904 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 1344 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 2240 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 1344 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 2240 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 1008 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 2240 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 1232 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 2352 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 1680 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 3136 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 840 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[8\].thrun
timestamp 1667941163
transform -1 0 3248 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 2016 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 2800 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 1904 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[10\].thrun
timestamp 1667941163
transform 1 0 2800 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[10\].thrup
timestamp 1667941163
transform 1 0 1008 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[11\].thrun
timestamp 1667941163
transform 1 0 2520 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_T\[11\].thrup
timestamp 1667941163
transform 1 0 896 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 1848 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 1344 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 1232 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 1568 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 1680 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 896 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[3\].crossn
timestamp 1667941163
transform -1 0 1120 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 1232 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 1512 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 2016 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[5\].crossn
timestamp 1667941163
transform 1 0 1904 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_load.gen_X\[5\].crossp
timestamp 1667941163
transform 1 0 1008 0 1 2352
box -43 -43 267 435
<< labels >>
flabel metal3 s 0 4424 400 4480 0 FreeSans 224 0 0 0 nbus
port 0 nsew signal bidirectional
flabel metal3 s 5600 1792 6000 1848 0 FreeSans 224 0 0 0 outn
port 1 nsew signal bidirectional
flabel metal3 s 5600 4144 6000 4200 0 FreeSans 224 0 0 0 outnn
port 2 nsew signal tristate
flabel metal3 s 5600 616 6000 672 0 FreeSans 224 0 0 0 outp
port 3 nsew signal bidirectional
flabel metal3 s 5600 2968 6000 3024 0 FreeSans 224 0 0 0 outpn
port 4 nsew signal tristate
flabel metal3 s 5600 5320 6000 5376 0 FreeSans 224 0 0 0 outxor
port 5 nsew signal tristate
flabel metal3 s 0 1456 400 1512 0 FreeSans 224 0 0 0 pbus
port 6 nsew signal bidirectional
flabel metal4 s 1173 1538 1333 4342 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 2335 1538 2495 4342 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 3497 1538 3657 4342 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 4659 1538 4819 4342 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 1754 1538 1914 4342 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
flabel metal4 s 2916 1538 3076 4342 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
flabel metal4 s 4078 1538 4238 4342 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
flabel metal4 s 5240 1538 5400 4342 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
rlabel metal1 2996 4312 2996 4312 0 vdd
rlabel via1 3036 3920 3036 3920 0 vss
rlabel metal2 4172 2772 4172 2772 0 nbus
rlabel metal2 3724 1960 3724 1960 0 outn
rlabel metal2 4900 3780 4900 3780 0 outnn
rlabel metal2 3920 2660 3920 2660 0 outp
rlabel metal2 5012 2800 5012 2800 0 outpn
rlabel metal2 5040 3388 5040 3388 0 outxor
rlabel metal2 980 1596 980 1596 0 pbus
<< properties >>
string FIXED_BBOX 0 0 6000 6000
<< end >>
