// This is the unpowered netlist.
module injector (enable,
    outn,
    outp,
    signal,
    trim_n,
    trim_p);
 input enable;
 inout outn;
 inout outp;
 input signal;
 input [3:0] trim_n;
 input [3:0] trim_p;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire signal_n;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _29_ (.I(enable),
    .ZN(_00_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _30_ (.A1(signal_n),
    .A2(_00_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _31_ (.I(_04_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _32_ (.A1(enable),
    .A2(signal),
    .Z(_03_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _33_ (.I(_03_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _34_ (.Z(_05_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _35_ (.Z(_06_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _36_ (.Z(_07_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _37_ (.Z(_08_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _38_ (.Z(_09_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _39_ (.Z(_10_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _40_ (.Z(_11_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _41_ (.Z(_12_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _42_ (.Z(_13_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _43_ (.Z(_14_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _44_ (.Z(_15_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _45_ (.Z(_16_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _46_ (.Z(_17_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _47_ (.Z(_18_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _48_ (.Z(_19_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _49_ (.Z(_20_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _50_ (.Z(_21_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _51_ (.Z(_22_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _52_ (.Z(_23_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _53_ (.Z(_24_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _54_ (.Z(_25_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _55_ (.Z(_26_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _56_ (.Z(_27_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _57_ (.Z(_28_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[0].pdn  (.I(_05_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[0].pdp  (.I(_06_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[1].pdn  (.I(_07_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[1].pdp  (.I(_08_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[2].pdn  (.I(_09_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[2].pdp  (.I(_10_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[3].pdn  (.I(_11_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[3].pdp  (.I(_12_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[4].pdn  (.I(_13_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[4].pdp  (.I(_14_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[5].pdn  (.I(_15_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[5].pdp  (.I(_16_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[6].pdn  (.I(_17_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[6].pdp  (.I(_18_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[7].pdn  (.I(_19_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PD[7].pdp  (.I(_20_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[0].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[0].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[10].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[10].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[11].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[11].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[12].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[12].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[13].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[13].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[14].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[14].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[15].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[15].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[16].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[16].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[17].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[17].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[18].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[18].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[19].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[19].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[1].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[1].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[2].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[2].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[3].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[3].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[4].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[4].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[5].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[5].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[6].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[6].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[7].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[7].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[8].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[8].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[9].pun  (.I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_PU[9].pup  (.I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[0].ntrimn  (.EN(trim_n[0]),
    .I(_21_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[0].ntrimp  (.EN(trim_n[0]),
    .I(_22_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[0].ptrimn  (.EN(trim_p[0]),
    .I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[0].ptrimp  (.EN(trim_p[0]),
    .I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[1].ntrimn  (.EN(trim_n[1]),
    .I(_23_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[1].ntrimp  (.EN(trim_n[1]),
    .I(_24_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[1].ptrimn  (.EN(trim_p[1]),
    .I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[1].ptrimp  (.EN(trim_p[1]),
    .I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[2].ntrimn  (.EN(trim_n[2]),
    .I(_25_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[2].ntrimp  (.EN(trim_n[2]),
    .I(_26_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[2].ptrimn  (.EN(trim_p[2]),
    .I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[2].ptrimp  (.EN(trim_p[2]),
    .I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[3].ntrimn  (.EN(trim_n[3]),
    .I(_27_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[3].ntrimp  (.EN(trim_n[3]),
    .I(_28_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[3].ptrimn  (.EN(trim_p[3]),
    .I(_00_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \gen_TRIM[3].ptrimp  (.EN(trim_p[3]),
    .I(_00_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 nsijn (.I(_02_),
    .ZN(outn));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 psijp (.I(_01_),
    .ZN(outp));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 siginv (.I(signal),
    .ZN(signal_n));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_151 ();
endmodule

