magic
tech gf180mcuC
magscale 1 10
timestamp 1669830057
<< metal1 >>
rect 1344 8650 18592 8684
rect 1344 8598 3370 8650
rect 3422 8598 3474 8650
rect 3526 8598 3578 8650
rect 3630 8598 7682 8650
rect 7734 8598 7786 8650
rect 7838 8598 7890 8650
rect 7942 8598 11994 8650
rect 12046 8598 12098 8650
rect 12150 8598 12202 8650
rect 12254 8598 16306 8650
rect 16358 8598 16410 8650
rect 16462 8598 16514 8650
rect 16566 8598 18592 8650
rect 1344 8564 18592 8598
rect 10558 8370 10610 8382
rect 10558 8306 10610 8318
rect 16606 8370 16658 8382
rect 16606 8306 16658 8318
rect 4174 8258 4226 8270
rect 9886 8258 9938 8270
rect 2482 8206 2494 8258
rect 2546 8206 2558 8258
rect 7298 8206 7310 8258
rect 7362 8206 7374 8258
rect 8866 8206 8878 8258
rect 8930 8206 8942 8258
rect 11330 8206 11342 8258
rect 11394 8206 11406 8258
rect 12562 8206 12574 8258
rect 12626 8206 12638 8258
rect 14466 8206 14478 8258
rect 14530 8206 14542 8258
rect 15810 8206 15822 8258
rect 15874 8206 15886 8258
rect 4174 8194 4226 8206
rect 9886 8194 9938 8206
rect 1822 8146 1874 8158
rect 1822 8082 1874 8094
rect 3278 8146 3330 8158
rect 6750 8146 6802 8158
rect 4610 8094 4622 8146
rect 4674 8094 4686 8146
rect 3278 8082 3330 8094
rect 6750 8082 6802 8094
rect 8094 8146 8146 8158
rect 8094 8082 8146 8094
rect 10670 8146 10722 8158
rect 10670 8082 10722 8094
rect 12014 8146 12066 8158
rect 12014 8082 12066 8094
rect 13694 8146 13746 8158
rect 13694 8082 13746 8094
rect 15150 8146 15202 8158
rect 15150 8082 15202 8094
rect 16494 8146 16546 8158
rect 16494 8082 16546 8094
rect 17502 8146 17554 8158
rect 17502 8082 17554 8094
rect 1934 8034 1986 8046
rect 1934 7970 1986 7982
rect 4958 8034 5010 8046
rect 4958 7970 5010 7982
rect 6638 8034 6690 8046
rect 6638 7970 6690 7982
rect 9998 8034 10050 8046
rect 9998 7970 10050 7982
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 17614 8034 17666 8046
rect 17614 7970 17666 7982
rect 1344 7866 18752 7900
rect 1344 7814 5526 7866
rect 5578 7814 5630 7866
rect 5682 7814 5734 7866
rect 5786 7814 9838 7866
rect 9890 7814 9942 7866
rect 9994 7814 10046 7866
rect 10098 7814 14150 7866
rect 14202 7814 14254 7866
rect 14306 7814 14358 7866
rect 14410 7814 18462 7866
rect 18514 7814 18566 7866
rect 18618 7814 18670 7866
rect 18722 7814 18752 7866
rect 1344 7780 18752 7814
rect 1934 7698 1986 7710
rect 1934 7634 1986 7646
rect 16718 7698 16770 7710
rect 16718 7634 16770 7646
rect 17838 7698 17890 7710
rect 17838 7634 17890 7646
rect 1822 7474 1874 7486
rect 3278 7474 3330 7486
rect 2482 7422 2494 7474
rect 2546 7422 2558 7474
rect 1822 7410 1874 7422
rect 3278 7410 3330 7422
rect 4174 7474 4226 7486
rect 4174 7410 4226 7422
rect 4734 7474 4786 7486
rect 10110 7474 10162 7486
rect 7298 7422 7310 7474
rect 7362 7422 7374 7474
rect 8866 7422 8878 7474
rect 8930 7422 8942 7474
rect 4734 7410 4786 7422
rect 10110 7410 10162 7422
rect 10782 7474 10834 7486
rect 10782 7410 10834 7422
rect 11454 7474 11506 7486
rect 13806 7474 13858 7486
rect 16606 7474 16658 7486
rect 12338 7422 12350 7474
rect 12402 7422 12414 7474
rect 14578 7422 14590 7474
rect 14642 7422 14654 7474
rect 15810 7422 15822 7474
rect 15874 7422 15886 7474
rect 11454 7410 11506 7422
rect 13806 7410 13858 7422
rect 16606 7410 16658 7422
rect 17726 7474 17778 7486
rect 17726 7410 17778 7422
rect 8094 7362 8146 7374
rect 8094 7298 8146 7310
rect 12910 7362 12962 7374
rect 12910 7298 12962 7310
rect 15262 7362 15314 7374
rect 15262 7298 15314 7310
rect 4622 7250 4674 7262
rect 4622 7186 4674 7198
rect 10222 7250 10274 7262
rect 10222 7186 10274 7198
rect 10894 7250 10946 7262
rect 10894 7186 10946 7198
rect 11566 7250 11618 7262
rect 11566 7186 11618 7198
rect 1344 7082 18592 7116
rect 1344 7030 3370 7082
rect 3422 7030 3474 7082
rect 3526 7030 3578 7082
rect 3630 7030 7682 7082
rect 7734 7030 7786 7082
rect 7838 7030 7890 7082
rect 7942 7030 11994 7082
rect 12046 7030 12098 7082
rect 12150 7030 12202 7082
rect 12254 7030 16306 7082
rect 16358 7030 16410 7082
rect 16462 7030 16514 7082
rect 16566 7030 18592 7082
rect 1344 6996 18592 7030
rect 2158 6914 2210 6926
rect 2158 6850 2210 6862
rect 2494 6914 2546 6926
rect 2494 6850 2546 6862
rect 7646 6914 7698 6926
rect 7646 6850 7698 6862
rect 8318 6914 8370 6926
rect 8318 6850 8370 6862
rect 15822 6914 15874 6926
rect 15822 6850 15874 6862
rect 6862 6802 6914 6814
rect 6862 6738 6914 6750
rect 2718 6690 2770 6702
rect 2718 6626 2770 6638
rect 13694 6690 13746 6702
rect 13694 6626 13746 6638
rect 14366 6690 14418 6702
rect 14366 6626 14418 6638
rect 15038 6690 15090 6702
rect 15038 6626 15090 6638
rect 15710 6690 15762 6702
rect 15710 6626 15762 6638
rect 7534 6578 7586 6590
rect 3266 6526 3278 6578
rect 3330 6526 3342 6578
rect 7534 6514 7586 6526
rect 8206 6578 8258 6590
rect 8206 6514 8258 6526
rect 8878 6578 8930 6590
rect 8878 6514 8930 6526
rect 9550 6578 9602 6590
rect 9550 6514 9602 6526
rect 10222 6578 10274 6590
rect 10222 6514 10274 6526
rect 10894 6578 10946 6590
rect 10894 6514 10946 6526
rect 11566 6578 11618 6590
rect 11566 6514 11618 6526
rect 12238 6578 12290 6590
rect 12238 6514 12290 6526
rect 16382 6578 16434 6590
rect 16382 6514 16434 6526
rect 17054 6578 17106 6590
rect 17054 6514 17106 6526
rect 17726 6578 17778 6590
rect 17726 6514 17778 6526
rect 3614 6466 3666 6478
rect 3614 6402 3666 6414
rect 8990 6466 9042 6478
rect 8990 6402 9042 6414
rect 9662 6466 9714 6478
rect 9662 6402 9714 6414
rect 10334 6466 10386 6478
rect 10334 6402 10386 6414
rect 11006 6466 11058 6478
rect 11006 6402 11058 6414
rect 11678 6466 11730 6478
rect 11678 6402 11730 6414
rect 12350 6466 12402 6478
rect 12350 6402 12402 6414
rect 13806 6466 13858 6478
rect 13806 6402 13858 6414
rect 14478 6466 14530 6478
rect 14478 6402 14530 6414
rect 15150 6466 15202 6478
rect 15150 6402 15202 6414
rect 16494 6466 16546 6478
rect 16494 6402 16546 6414
rect 17166 6466 17218 6478
rect 17166 6402 17218 6414
rect 17838 6466 17890 6478
rect 17838 6402 17890 6414
rect 1344 6298 18752 6332
rect 1344 6246 5526 6298
rect 5578 6246 5630 6298
rect 5682 6246 5734 6298
rect 5786 6246 9838 6298
rect 9890 6246 9942 6298
rect 9994 6246 10046 6298
rect 10098 6246 14150 6298
rect 14202 6246 14254 6298
rect 14306 6246 14358 6298
rect 14410 6246 18462 6298
rect 18514 6246 18566 6298
rect 18618 6246 18670 6298
rect 18722 6246 18752 6298
rect 1344 6212 18752 6246
rect 3054 6130 3106 6142
rect 2370 6078 2382 6130
rect 2434 6078 2446 6130
rect 3054 6066 3106 6078
rect 8990 6130 9042 6142
rect 8990 6066 9042 6078
rect 11118 6130 11170 6142
rect 11118 6066 11170 6078
rect 14478 6130 14530 6142
rect 14478 6066 14530 6078
rect 15822 6130 15874 6142
rect 15822 6066 15874 6078
rect 6302 6018 6354 6030
rect 6302 5954 6354 5966
rect 8878 6018 8930 6030
rect 8878 5954 8930 5966
rect 13694 6018 13746 6030
rect 13694 5954 13746 5966
rect 15038 6018 15090 6030
rect 15038 5954 15090 5966
rect 2046 5906 2098 5918
rect 2046 5842 2098 5854
rect 2942 5906 2994 5918
rect 2942 5842 2994 5854
rect 6190 5906 6242 5918
rect 6190 5842 6242 5854
rect 6862 5906 6914 5918
rect 6862 5842 6914 5854
rect 6974 5906 7026 5918
rect 6974 5842 7026 5854
rect 7534 5906 7586 5918
rect 7534 5842 7586 5854
rect 7646 5906 7698 5918
rect 7646 5842 7698 5854
rect 10334 5906 10386 5918
rect 10334 5842 10386 5854
rect 11006 5906 11058 5918
rect 11006 5842 11058 5854
rect 11678 5906 11730 5918
rect 11678 5842 11730 5854
rect 12350 5906 12402 5918
rect 12350 5842 12402 5854
rect 13022 5906 13074 5918
rect 13022 5842 13074 5854
rect 14366 5906 14418 5918
rect 14366 5842 14418 5854
rect 15710 5906 15762 5918
rect 15710 5842 15762 5854
rect 1822 5794 1874 5806
rect 1822 5730 1874 5742
rect 5630 5794 5682 5806
rect 5630 5730 5682 5742
rect 16494 5794 16546 5806
rect 16494 5730 16546 5742
rect 8318 5682 8370 5694
rect 8318 5618 8370 5630
rect 10446 5682 10498 5694
rect 10446 5618 10498 5630
rect 11790 5682 11842 5694
rect 11790 5618 11842 5630
rect 12462 5682 12514 5694
rect 12462 5618 12514 5630
rect 13134 5682 13186 5694
rect 13134 5618 13186 5630
rect 13806 5682 13858 5694
rect 13806 5618 13858 5630
rect 15150 5682 15202 5694
rect 15150 5618 15202 5630
rect 17726 5682 17778 5694
rect 17726 5618 17778 5630
rect 1344 5514 18592 5548
rect 1344 5462 3370 5514
rect 3422 5462 3474 5514
rect 3526 5462 3578 5514
rect 3630 5462 7682 5514
rect 7734 5462 7786 5514
rect 7838 5462 7890 5514
rect 7942 5462 11994 5514
rect 12046 5462 12098 5514
rect 12150 5462 12202 5514
rect 12254 5462 16306 5514
rect 16358 5462 16410 5514
rect 16462 5462 16514 5514
rect 16566 5462 18592 5514
rect 1344 5428 18592 5462
rect 4958 5346 5010 5358
rect 4958 5282 5010 5294
rect 6414 5346 6466 5358
rect 6414 5282 6466 5294
rect 6974 5346 7026 5358
rect 6974 5282 7026 5294
rect 4286 5234 4338 5246
rect 4286 5170 4338 5182
rect 8430 5234 8482 5246
rect 8430 5170 8482 5182
rect 9102 5234 9154 5246
rect 9102 5170 9154 5182
rect 9774 5234 9826 5246
rect 9774 5170 9826 5182
rect 10446 5234 10498 5246
rect 10446 5170 10498 5182
rect 11118 5234 11170 5246
rect 11118 5170 11170 5182
rect 14478 5234 14530 5246
rect 14478 5170 14530 5182
rect 15710 5234 15762 5246
rect 15710 5170 15762 5182
rect 7646 5122 7698 5134
rect 7646 5058 7698 5070
rect 8990 5122 9042 5134
rect 8990 5058 9042 5070
rect 9662 5122 9714 5134
rect 9662 5058 9714 5070
rect 10334 5122 10386 5134
rect 10334 5058 10386 5070
rect 11006 5122 11058 5134
rect 11006 5058 11058 5070
rect 11678 5122 11730 5134
rect 11678 5058 11730 5070
rect 12350 5122 12402 5134
rect 12350 5058 12402 5070
rect 12462 5122 12514 5134
rect 12462 5058 12514 5070
rect 13694 5122 13746 5134
rect 13694 5058 13746 5070
rect 13806 5122 13858 5134
rect 13806 5058 13858 5070
rect 14366 5122 14418 5134
rect 14366 5058 14418 5070
rect 15150 5122 15202 5134
rect 15150 5058 15202 5070
rect 16382 5122 16434 5134
rect 16382 5058 16434 5070
rect 17278 5122 17330 5134
rect 17826 5070 17838 5122
rect 17890 5070 17902 5122
rect 17278 5058 17330 5070
rect 7758 5010 7810 5022
rect 7758 4946 7810 4958
rect 11790 4898 11842 4910
rect 11790 4834 11842 4846
rect 15038 4898 15090 4910
rect 15038 4834 15090 4846
rect 1344 4730 18752 4764
rect 1344 4678 5526 4730
rect 5578 4678 5630 4730
rect 5682 4678 5734 4730
rect 5786 4678 9838 4730
rect 9890 4678 9942 4730
rect 9994 4678 10046 4730
rect 10098 4678 14150 4730
rect 14202 4678 14254 4730
rect 14306 4678 14358 4730
rect 14410 4678 18462 4730
rect 18514 4678 18566 4730
rect 18618 4678 18670 4730
rect 18722 4678 18752 4730
rect 1344 4644 18752 4678
rect 10782 4562 10834 4574
rect 10782 4498 10834 4510
rect 11454 4562 11506 4574
rect 11454 4498 11506 4510
rect 15038 4562 15090 4574
rect 15038 4498 15090 4510
rect 15710 4562 15762 4574
rect 15710 4498 15762 4510
rect 16382 4562 16434 4574
rect 16382 4498 16434 4510
rect 17838 4562 17890 4574
rect 17838 4498 17890 4510
rect 3502 4450 3554 4462
rect 3502 4386 3554 4398
rect 7982 4450 8034 4462
rect 7982 4386 8034 4398
rect 10894 4450 10946 4462
rect 10894 4386 10946 4398
rect 11566 4450 11618 4462
rect 11566 4386 11618 4398
rect 12910 4450 12962 4462
rect 12910 4386 12962 4398
rect 14926 4450 14978 4462
rect 14926 4386 14978 4398
rect 16270 4450 16322 4462
rect 16270 4386 16322 4398
rect 7086 4338 7138 4350
rect 12014 4338 12066 4350
rect 15598 4338 15650 4350
rect 2706 4286 2718 4338
rect 2770 4286 2782 4338
rect 4274 4286 4286 4338
rect 4338 4286 4350 4338
rect 8642 4286 8654 4338
rect 8706 4286 8718 4338
rect 13458 4286 13470 4338
rect 13522 4286 13534 4338
rect 14466 4286 14478 4338
rect 14530 4335 14542 4338
rect 14802 4335 14814 4338
rect 14530 4289 14814 4335
rect 14530 4286 14542 4289
rect 14802 4286 14814 4289
rect 14866 4286 14878 4338
rect 7086 4274 7138 4286
rect 12014 4274 12066 4286
rect 15598 4274 15650 4286
rect 17726 4338 17778 4350
rect 17726 4274 17778 4286
rect 5966 4226 6018 4238
rect 5966 4162 6018 4174
rect 6638 4226 6690 4238
rect 6638 4162 6690 4174
rect 14366 4226 14418 4238
rect 14366 4162 14418 4174
rect 5294 4114 5346 4126
rect 5294 4050 5346 4062
rect 10222 4114 10274 4126
rect 10222 4050 10274 4062
rect 1344 3946 18592 3980
rect 1344 3894 3370 3946
rect 3422 3894 3474 3946
rect 3526 3894 3578 3946
rect 3630 3894 7682 3946
rect 7734 3894 7786 3946
rect 7838 3894 7890 3946
rect 7942 3894 11994 3946
rect 12046 3894 12098 3946
rect 12150 3894 12202 3946
rect 12254 3894 16306 3946
rect 16358 3894 16410 3946
rect 16462 3894 16514 3946
rect 16566 3894 18592 3946
rect 1344 3860 18592 3894
rect 6078 3778 6130 3790
rect 6078 3714 6130 3726
rect 9998 3778 10050 3790
rect 9998 3714 10050 3726
rect 10670 3778 10722 3790
rect 10670 3714 10722 3726
rect 14366 3778 14418 3790
rect 14366 3714 14418 3726
rect 17502 3778 17554 3790
rect 17502 3714 17554 3726
rect 2158 3666 2210 3678
rect 2158 3602 2210 3614
rect 3502 3666 3554 3678
rect 3502 3602 3554 3614
rect 4958 3666 5010 3678
rect 4958 3602 5010 3614
rect 6750 3666 6802 3678
rect 6750 3602 6802 3614
rect 8094 3666 8146 3678
rect 8094 3602 8146 3614
rect 12014 3666 12066 3678
rect 12014 3602 12066 3614
rect 15934 3666 15986 3678
rect 15934 3602 15986 3614
rect 2606 3554 2658 3566
rect 7198 3554 7250 3566
rect 11118 3554 11170 3566
rect 13694 3554 13746 3566
rect 4050 3502 4062 3554
rect 4114 3502 4126 3554
rect 8642 3502 8654 3554
rect 8706 3502 8718 3554
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 15138 3502 15150 3554
rect 15202 3502 15214 3554
rect 16706 3502 16718 3554
rect 16770 3502 16782 3554
rect 2606 3490 2658 3502
rect 7198 3490 7250 3502
rect 11118 3490 11170 3502
rect 13694 3490 13746 3502
rect 13582 3330 13634 3342
rect 13582 3266 13634 3278
rect 1344 3162 18752 3196
rect 1344 3110 5526 3162
rect 5578 3110 5630 3162
rect 5682 3110 5734 3162
rect 5786 3110 9838 3162
rect 9890 3110 9942 3162
rect 9994 3110 10046 3162
rect 10098 3110 14150 3162
rect 14202 3110 14254 3162
rect 14306 3110 14358 3162
rect 14410 3110 18462 3162
rect 18514 3110 18566 3162
rect 18618 3110 18670 3162
rect 18722 3110 18752 3162
rect 1344 3076 18752 3110
<< via1 >>
rect 3370 8598 3422 8650
rect 3474 8598 3526 8650
rect 3578 8598 3630 8650
rect 7682 8598 7734 8650
rect 7786 8598 7838 8650
rect 7890 8598 7942 8650
rect 11994 8598 12046 8650
rect 12098 8598 12150 8650
rect 12202 8598 12254 8650
rect 16306 8598 16358 8650
rect 16410 8598 16462 8650
rect 16514 8598 16566 8650
rect 10558 8318 10610 8370
rect 16606 8318 16658 8370
rect 2494 8206 2546 8258
rect 4174 8206 4226 8258
rect 7310 8206 7362 8258
rect 8878 8206 8930 8258
rect 9886 8206 9938 8258
rect 11342 8206 11394 8258
rect 12574 8206 12626 8258
rect 14478 8206 14530 8258
rect 15822 8206 15874 8258
rect 1822 8094 1874 8146
rect 3278 8094 3330 8146
rect 4622 8094 4674 8146
rect 6750 8094 6802 8146
rect 8094 8094 8146 8146
rect 10670 8094 10722 8146
rect 12014 8094 12066 8146
rect 13694 8094 13746 8146
rect 15150 8094 15202 8146
rect 16494 8094 16546 8146
rect 17502 8094 17554 8146
rect 1934 7982 1986 8034
rect 4958 7982 5010 8034
rect 6638 7982 6690 8034
rect 9998 7982 10050 8034
rect 13582 7982 13634 8034
rect 17614 7982 17666 8034
rect 5526 7814 5578 7866
rect 5630 7814 5682 7866
rect 5734 7814 5786 7866
rect 9838 7814 9890 7866
rect 9942 7814 9994 7866
rect 10046 7814 10098 7866
rect 14150 7814 14202 7866
rect 14254 7814 14306 7866
rect 14358 7814 14410 7866
rect 18462 7814 18514 7866
rect 18566 7814 18618 7866
rect 18670 7814 18722 7866
rect 1934 7646 1986 7698
rect 16718 7646 16770 7698
rect 17838 7646 17890 7698
rect 1822 7422 1874 7474
rect 2494 7422 2546 7474
rect 3278 7422 3330 7474
rect 4174 7422 4226 7474
rect 4734 7422 4786 7474
rect 7310 7422 7362 7474
rect 8878 7422 8930 7474
rect 10110 7422 10162 7474
rect 10782 7422 10834 7474
rect 11454 7422 11506 7474
rect 12350 7422 12402 7474
rect 13806 7422 13858 7474
rect 14590 7422 14642 7474
rect 15822 7422 15874 7474
rect 16606 7422 16658 7474
rect 17726 7422 17778 7474
rect 8094 7310 8146 7362
rect 12910 7310 12962 7362
rect 15262 7310 15314 7362
rect 4622 7198 4674 7250
rect 10222 7198 10274 7250
rect 10894 7198 10946 7250
rect 11566 7198 11618 7250
rect 3370 7030 3422 7082
rect 3474 7030 3526 7082
rect 3578 7030 3630 7082
rect 7682 7030 7734 7082
rect 7786 7030 7838 7082
rect 7890 7030 7942 7082
rect 11994 7030 12046 7082
rect 12098 7030 12150 7082
rect 12202 7030 12254 7082
rect 16306 7030 16358 7082
rect 16410 7030 16462 7082
rect 16514 7030 16566 7082
rect 2158 6862 2210 6914
rect 2494 6862 2546 6914
rect 7646 6862 7698 6914
rect 8318 6862 8370 6914
rect 15822 6862 15874 6914
rect 6862 6750 6914 6802
rect 2718 6638 2770 6690
rect 13694 6638 13746 6690
rect 14366 6638 14418 6690
rect 15038 6638 15090 6690
rect 15710 6638 15762 6690
rect 3278 6526 3330 6578
rect 7534 6526 7586 6578
rect 8206 6526 8258 6578
rect 8878 6526 8930 6578
rect 9550 6526 9602 6578
rect 10222 6526 10274 6578
rect 10894 6526 10946 6578
rect 11566 6526 11618 6578
rect 12238 6526 12290 6578
rect 16382 6526 16434 6578
rect 17054 6526 17106 6578
rect 17726 6526 17778 6578
rect 3614 6414 3666 6466
rect 8990 6414 9042 6466
rect 9662 6414 9714 6466
rect 10334 6414 10386 6466
rect 11006 6414 11058 6466
rect 11678 6414 11730 6466
rect 12350 6414 12402 6466
rect 13806 6414 13858 6466
rect 14478 6414 14530 6466
rect 15150 6414 15202 6466
rect 16494 6414 16546 6466
rect 17166 6414 17218 6466
rect 17838 6414 17890 6466
rect 5526 6246 5578 6298
rect 5630 6246 5682 6298
rect 5734 6246 5786 6298
rect 9838 6246 9890 6298
rect 9942 6246 9994 6298
rect 10046 6246 10098 6298
rect 14150 6246 14202 6298
rect 14254 6246 14306 6298
rect 14358 6246 14410 6298
rect 18462 6246 18514 6298
rect 18566 6246 18618 6298
rect 18670 6246 18722 6298
rect 2382 6078 2434 6130
rect 3054 6078 3106 6130
rect 8990 6078 9042 6130
rect 11118 6078 11170 6130
rect 14478 6078 14530 6130
rect 15822 6078 15874 6130
rect 6302 5966 6354 6018
rect 8878 5966 8930 6018
rect 13694 5966 13746 6018
rect 15038 5966 15090 6018
rect 2046 5854 2098 5906
rect 2942 5854 2994 5906
rect 6190 5854 6242 5906
rect 6862 5854 6914 5906
rect 6974 5854 7026 5906
rect 7534 5854 7586 5906
rect 7646 5854 7698 5906
rect 10334 5854 10386 5906
rect 11006 5854 11058 5906
rect 11678 5854 11730 5906
rect 12350 5854 12402 5906
rect 13022 5854 13074 5906
rect 14366 5854 14418 5906
rect 15710 5854 15762 5906
rect 1822 5742 1874 5794
rect 5630 5742 5682 5794
rect 16494 5742 16546 5794
rect 8318 5630 8370 5682
rect 10446 5630 10498 5682
rect 11790 5630 11842 5682
rect 12462 5630 12514 5682
rect 13134 5630 13186 5682
rect 13806 5630 13858 5682
rect 15150 5630 15202 5682
rect 17726 5630 17778 5682
rect 3370 5462 3422 5514
rect 3474 5462 3526 5514
rect 3578 5462 3630 5514
rect 7682 5462 7734 5514
rect 7786 5462 7838 5514
rect 7890 5462 7942 5514
rect 11994 5462 12046 5514
rect 12098 5462 12150 5514
rect 12202 5462 12254 5514
rect 16306 5462 16358 5514
rect 16410 5462 16462 5514
rect 16514 5462 16566 5514
rect 4958 5294 5010 5346
rect 6414 5294 6466 5346
rect 6974 5294 7026 5346
rect 4286 5182 4338 5234
rect 8430 5182 8482 5234
rect 9102 5182 9154 5234
rect 9774 5182 9826 5234
rect 10446 5182 10498 5234
rect 11118 5182 11170 5234
rect 14478 5182 14530 5234
rect 15710 5182 15762 5234
rect 7646 5070 7698 5122
rect 8990 5070 9042 5122
rect 9662 5070 9714 5122
rect 10334 5070 10386 5122
rect 11006 5070 11058 5122
rect 11678 5070 11730 5122
rect 12350 5070 12402 5122
rect 12462 5070 12514 5122
rect 13694 5070 13746 5122
rect 13806 5070 13858 5122
rect 14366 5070 14418 5122
rect 15150 5070 15202 5122
rect 16382 5070 16434 5122
rect 17278 5070 17330 5122
rect 17838 5070 17890 5122
rect 7758 4958 7810 5010
rect 11790 4846 11842 4898
rect 15038 4846 15090 4898
rect 5526 4678 5578 4730
rect 5630 4678 5682 4730
rect 5734 4678 5786 4730
rect 9838 4678 9890 4730
rect 9942 4678 9994 4730
rect 10046 4678 10098 4730
rect 14150 4678 14202 4730
rect 14254 4678 14306 4730
rect 14358 4678 14410 4730
rect 18462 4678 18514 4730
rect 18566 4678 18618 4730
rect 18670 4678 18722 4730
rect 10782 4510 10834 4562
rect 11454 4510 11506 4562
rect 15038 4510 15090 4562
rect 15710 4510 15762 4562
rect 16382 4510 16434 4562
rect 17838 4510 17890 4562
rect 3502 4398 3554 4450
rect 7982 4398 8034 4450
rect 10894 4398 10946 4450
rect 11566 4398 11618 4450
rect 12910 4398 12962 4450
rect 14926 4398 14978 4450
rect 16270 4398 16322 4450
rect 2718 4286 2770 4338
rect 4286 4286 4338 4338
rect 7086 4286 7138 4338
rect 8654 4286 8706 4338
rect 12014 4286 12066 4338
rect 13470 4286 13522 4338
rect 14478 4286 14530 4338
rect 14814 4286 14866 4338
rect 15598 4286 15650 4338
rect 17726 4286 17778 4338
rect 5966 4174 6018 4226
rect 6638 4174 6690 4226
rect 14366 4174 14418 4226
rect 5294 4062 5346 4114
rect 10222 4062 10274 4114
rect 3370 3894 3422 3946
rect 3474 3894 3526 3946
rect 3578 3894 3630 3946
rect 7682 3894 7734 3946
rect 7786 3894 7838 3946
rect 7890 3894 7942 3946
rect 11994 3894 12046 3946
rect 12098 3894 12150 3946
rect 12202 3894 12254 3946
rect 16306 3894 16358 3946
rect 16410 3894 16462 3946
rect 16514 3894 16566 3946
rect 6078 3726 6130 3778
rect 9998 3726 10050 3778
rect 10670 3726 10722 3778
rect 14366 3726 14418 3778
rect 17502 3726 17554 3778
rect 2158 3614 2210 3666
rect 3502 3614 3554 3666
rect 4958 3614 5010 3666
rect 6750 3614 6802 3666
rect 8094 3614 8146 3666
rect 12014 3614 12066 3666
rect 15934 3614 15986 3666
rect 2606 3502 2658 3554
rect 4062 3502 4114 3554
rect 7198 3502 7250 3554
rect 8654 3502 8706 3554
rect 11118 3502 11170 3554
rect 12574 3502 12626 3554
rect 13694 3502 13746 3554
rect 15150 3502 15202 3554
rect 16718 3502 16770 3554
rect 13582 3278 13634 3330
rect 5526 3110 5578 3162
rect 5630 3110 5682 3162
rect 5734 3110 5786 3162
rect 9838 3110 9890 3162
rect 9942 3110 9994 3162
rect 10046 3110 10098 3162
rect 14150 3110 14202 3162
rect 14254 3110 14306 3162
rect 14358 3110 14410 3162
rect 18462 3110 18514 3162
rect 18566 3110 18618 3162
rect 18670 3110 18722 3162
<< metal2 >>
rect 2464 11200 2576 12000
rect 7392 11200 7504 12000
rect 12320 11200 12432 12000
rect 17248 11200 17360 12000
rect 2044 8372 2100 8382
rect 1820 8148 1876 8158
rect 1820 8054 1876 8092
rect 1932 8034 1988 8046
rect 1932 7982 1934 8034
rect 1986 7982 1988 8034
rect 1932 7924 1988 7982
rect 1932 7858 1988 7868
rect 1932 7700 1988 7710
rect 1932 7606 1988 7644
rect 1820 7474 1876 7486
rect 1820 7422 1822 7474
rect 1874 7422 1876 7474
rect 1820 6580 1876 7422
rect 1820 6514 1876 6524
rect 2044 7476 2100 8316
rect 2492 8258 2548 11200
rect 3368 8652 3632 8662
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3368 8586 3632 8596
rect 7420 8428 7476 11200
rect 7680 8652 7944 8662
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7680 8586 7944 8596
rect 11992 8652 12256 8662
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 11992 8586 12256 8596
rect 7308 8372 7476 8428
rect 10556 8372 10612 8382
rect 2492 8206 2494 8258
rect 2546 8206 2548 8258
rect 2044 5906 2100 7420
rect 2156 8036 2212 8046
rect 2156 6914 2212 7980
rect 2492 7474 2548 8206
rect 4172 8258 4228 8270
rect 4172 8206 4174 8258
rect 4226 8206 4228 8258
rect 3276 8146 3332 8158
rect 3276 8094 3278 8146
rect 3330 8094 3332 8146
rect 3276 7700 3332 8094
rect 2492 7422 2494 7474
rect 2546 7422 2548 7474
rect 2492 7410 2548 7422
rect 3164 7644 3276 7700
rect 3052 7364 3108 7374
rect 2716 7252 2772 7262
rect 2156 6862 2158 6914
rect 2210 6862 2212 6914
rect 2156 6850 2212 6862
rect 2492 6916 2548 6926
rect 2492 6822 2548 6860
rect 2716 6690 2772 7196
rect 2716 6638 2718 6690
rect 2770 6638 2772 6690
rect 2716 6626 2772 6638
rect 3052 6916 3108 7308
rect 2380 6132 2436 6142
rect 2380 6038 2436 6076
rect 3052 6130 3108 6860
rect 3052 6078 3054 6130
rect 3106 6078 3108 6130
rect 3052 6066 3108 6078
rect 2044 5854 2046 5906
rect 2098 5854 2100 5906
rect 2044 5842 2100 5854
rect 2940 5906 2996 5918
rect 2940 5854 2942 5906
rect 2994 5854 2996 5906
rect 1820 5794 1876 5806
rect 1820 5742 1822 5794
rect 1874 5742 1876 5794
rect 1820 5012 1876 5742
rect 1820 2996 1876 4956
rect 2940 5012 2996 5854
rect 3164 5908 3220 7644
rect 3276 7634 3332 7644
rect 3388 7924 3444 7934
rect 3276 7476 3332 7486
rect 3388 7476 3444 7868
rect 3276 7474 3444 7476
rect 3276 7422 3278 7474
rect 3330 7422 3444 7474
rect 3276 7420 3444 7422
rect 3724 7924 3780 7934
rect 3276 7410 3332 7420
rect 3368 7084 3632 7094
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3368 7018 3632 7028
rect 3276 6580 3332 6590
rect 3276 6486 3332 6524
rect 3612 6466 3668 6478
rect 3612 6414 3614 6466
rect 3666 6414 3668 6466
rect 3612 6132 3668 6414
rect 3612 6066 3668 6076
rect 3164 5348 3220 5852
rect 3368 5516 3632 5526
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3368 5450 3632 5460
rect 3164 5292 3556 5348
rect 2940 4946 2996 4956
rect 3500 4450 3556 5292
rect 3500 4398 3502 4450
rect 3554 4398 3556 4450
rect 3500 4386 3556 4398
rect 2716 4338 2772 4350
rect 2716 4286 2718 4338
rect 2770 4286 2772 4338
rect 2156 3666 2212 3678
rect 2156 3614 2158 3666
rect 2210 3614 2212 3666
rect 2156 3556 2212 3614
rect 2604 3556 2660 3566
rect 2156 3554 2660 3556
rect 2156 3502 2606 3554
rect 2658 3502 2660 3554
rect 2156 3500 2660 3502
rect 2604 3490 2660 3500
rect 2716 3556 2772 4286
rect 3368 3948 3632 3958
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3368 3882 3632 3892
rect 3500 3668 3556 3678
rect 3724 3668 3780 7868
rect 4172 7474 4228 8206
rect 7308 8258 7364 8372
rect 10556 8370 10948 8372
rect 10556 8318 10558 8370
rect 10610 8318 10948 8370
rect 10556 8316 10948 8318
rect 10556 8306 10612 8316
rect 7308 8206 7310 8258
rect 7362 8206 7364 8258
rect 4620 8148 4676 8158
rect 4620 8054 4676 8092
rect 6748 8146 6804 8158
rect 6748 8094 6750 8146
rect 6802 8094 6804 8146
rect 4956 8036 5012 8046
rect 4956 7942 5012 7980
rect 6636 8036 6692 8046
rect 6636 7942 6692 7980
rect 5524 7868 5788 7878
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5524 7802 5788 7812
rect 4172 7422 4174 7474
rect 4226 7422 4228 7474
rect 4172 7364 4228 7422
rect 4732 7476 4788 7486
rect 4732 7382 4788 7420
rect 4172 7298 4228 7308
rect 6748 7364 6804 8094
rect 7308 7474 7364 8206
rect 8876 8258 8932 8270
rect 8876 8206 8878 8258
rect 8930 8206 8932 8258
rect 8092 8146 8148 8158
rect 8092 8094 8094 8146
rect 8146 8094 8148 8146
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 7308 7410 7364 7422
rect 7532 8036 7588 8046
rect 4620 7252 4676 7262
rect 4620 7158 4676 7196
rect 6300 6804 6356 6814
rect 4956 6692 5012 6702
rect 4956 5346 5012 6636
rect 5524 6300 5788 6310
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5524 6234 5788 6244
rect 6300 6018 6356 6748
rect 6748 6580 6804 7308
rect 7532 6916 7588 7980
rect 8092 8036 8148 8094
rect 8092 7970 8148 7980
rect 8876 7474 8932 8206
rect 9884 8260 9940 8270
rect 9884 8258 10388 8260
rect 9884 8206 9886 8258
rect 9938 8206 10388 8258
rect 9884 8204 10388 8206
rect 9884 8194 9940 8204
rect 10332 8148 10388 8204
rect 10668 8148 10724 8158
rect 10332 8146 10836 8148
rect 10332 8094 10670 8146
rect 10722 8094 10836 8146
rect 10332 8092 10836 8094
rect 10668 8082 10724 8092
rect 9996 8036 10052 8046
rect 9996 8034 10388 8036
rect 9996 7982 9998 8034
rect 10050 7982 10388 8034
rect 9996 7980 10388 7982
rect 9996 7970 10052 7980
rect 9836 7868 10100 7878
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 9836 7802 10100 7812
rect 8876 7422 8878 7474
rect 8930 7422 8932 7474
rect 8092 7362 8148 7374
rect 8092 7310 8094 7362
rect 8146 7310 8148 7362
rect 7680 7084 7944 7094
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7680 7018 7944 7028
rect 7644 6916 7700 6926
rect 7532 6860 7644 6916
rect 6860 6804 6916 6814
rect 7644 6784 7700 6860
rect 6860 6710 6916 6748
rect 6748 6514 6804 6524
rect 7532 6580 7588 6590
rect 7532 6486 7588 6524
rect 6300 5966 6302 6018
rect 6354 5966 6356 6018
rect 6300 5954 6356 5966
rect 6188 5908 6244 5918
rect 6188 5814 6244 5852
rect 6860 5908 6916 5918
rect 6860 5814 6916 5852
rect 6972 5906 7028 5918
rect 6972 5854 6974 5906
rect 7026 5854 7028 5906
rect 5628 5796 5684 5806
rect 5628 5702 5684 5740
rect 4956 5294 4958 5346
rect 5010 5294 5012 5346
rect 4956 5282 5012 5294
rect 6412 5348 6468 5358
rect 6412 5254 6468 5292
rect 6972 5346 7028 5854
rect 6972 5294 6974 5346
rect 7026 5294 7028 5346
rect 6972 5282 7028 5294
rect 7420 5908 7476 5918
rect 4284 5234 4340 5246
rect 4284 5182 4286 5234
rect 4338 5182 4340 5234
rect 4284 4338 4340 5182
rect 7420 5124 7476 5852
rect 7532 5906 7588 5918
rect 7532 5854 7534 5906
rect 7586 5854 7588 5906
rect 7532 5348 7588 5854
rect 7644 5908 7700 5918
rect 7644 5814 7700 5852
rect 8092 5908 8148 7310
rect 8316 6916 8372 6926
rect 8204 6580 8260 6590
rect 8204 6486 8260 6524
rect 8316 6468 8372 6860
rect 8316 5908 8372 6412
rect 8876 6580 8932 7422
rect 10108 7474 10164 7486
rect 10108 7422 10110 7474
rect 10162 7422 10164 7474
rect 8876 6018 8932 6524
rect 9548 6580 9604 6590
rect 9548 6486 9604 6524
rect 10108 6580 10164 7422
rect 10220 7252 10276 7262
rect 10332 7252 10388 7980
rect 10220 7250 10388 7252
rect 10220 7198 10222 7250
rect 10274 7198 10388 7250
rect 10220 7196 10388 7198
rect 10220 7186 10276 7196
rect 10220 6580 10276 6590
rect 10164 6578 10276 6580
rect 10164 6526 10222 6578
rect 10274 6526 10276 6578
rect 10164 6524 10276 6526
rect 8988 6468 9044 6478
rect 8988 6132 9044 6412
rect 8988 6038 9044 6076
rect 9660 6466 9716 6478
rect 9660 6414 9662 6466
rect 9714 6414 9716 6466
rect 10108 6448 10164 6524
rect 9660 6132 9716 6414
rect 9836 6300 10100 6310
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 9836 6234 10100 6244
rect 9660 6066 9716 6076
rect 8876 5966 8878 6018
rect 8930 5966 8932 6018
rect 8876 5954 8932 5966
rect 8092 5684 8148 5852
rect 8092 5618 8148 5628
rect 8204 5852 8372 5908
rect 10220 5908 10276 6524
rect 10332 6468 10388 7196
rect 10780 7474 10836 8092
rect 10780 7422 10782 7474
rect 10834 7422 10836 7474
rect 10780 6580 10836 7422
rect 10892 7252 10948 8316
rect 11340 8260 11396 8270
rect 12348 8260 12404 11200
rect 16304 8652 16568 8662
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16304 8586 16568 8596
rect 15260 8372 15316 8382
rect 12572 8260 12628 8270
rect 11340 8258 11508 8260
rect 11340 8206 11342 8258
rect 11394 8206 11508 8258
rect 11340 8204 11508 8206
rect 11340 8194 11396 8204
rect 11452 7474 11508 8204
rect 12348 8258 12628 8260
rect 12348 8206 12574 8258
rect 12626 8206 12628 8258
rect 12348 8204 12628 8206
rect 11452 7422 11454 7474
rect 11506 7422 11508 7474
rect 10892 7250 11172 7252
rect 10892 7198 10894 7250
rect 10946 7198 11172 7250
rect 10892 7196 11172 7198
rect 10892 7186 10948 7196
rect 10892 6580 10948 6590
rect 10780 6578 10948 6580
rect 10780 6526 10894 6578
rect 10946 6526 10948 6578
rect 10780 6524 10948 6526
rect 10332 6374 10388 6412
rect 10668 6020 10724 6030
rect 10332 5908 10388 5918
rect 10220 5852 10332 5908
rect 7680 5516 7944 5526
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7680 5450 7944 5460
rect 7532 5282 7588 5292
rect 7644 5124 7700 5134
rect 7420 5122 7700 5124
rect 7420 5070 7646 5122
rect 7698 5070 7700 5122
rect 7420 5068 7700 5070
rect 7644 4788 7700 5068
rect 7756 5012 7812 5022
rect 7756 5010 8148 5012
rect 7756 4958 7758 5010
rect 7810 4958 8148 5010
rect 7756 4956 8148 4958
rect 7756 4946 7812 4956
rect 5524 4732 5788 4742
rect 7644 4732 8036 4788
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5524 4666 5788 4676
rect 7980 4450 8036 4732
rect 7980 4398 7982 4450
rect 8034 4398 8036 4450
rect 7980 4386 8036 4398
rect 4284 4286 4286 4338
rect 4338 4286 4340 4338
rect 4284 4274 4340 4286
rect 5964 4340 6020 4350
rect 5964 4226 6020 4284
rect 7084 4340 7140 4350
rect 7084 4246 7140 4284
rect 5964 4174 5966 4226
rect 6018 4174 6020 4226
rect 5964 4162 6020 4174
rect 6636 4228 6692 4238
rect 6636 4134 6692 4172
rect 5292 4116 5348 4126
rect 5292 4022 5348 4060
rect 7680 3948 7944 3958
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7680 3882 7944 3892
rect 8092 3892 8148 4956
rect 8092 3826 8148 3836
rect 6076 3780 6132 3790
rect 6076 3686 6132 3724
rect 3500 3666 3780 3668
rect 3500 3614 3502 3666
rect 3554 3614 3780 3666
rect 3500 3612 3780 3614
rect 4956 3668 5012 3678
rect 3500 3602 3556 3612
rect 4956 3574 5012 3612
rect 6748 3666 6804 3678
rect 6748 3614 6750 3666
rect 6802 3614 6804 3666
rect 1820 2930 1876 2940
rect 2716 2660 2772 3500
rect 4060 3556 4116 3566
rect 4060 3462 4116 3500
rect 6748 3444 6804 3614
rect 7196 3668 7252 3678
rect 7196 3554 7252 3612
rect 8092 3668 8148 3678
rect 8204 3668 8260 5852
rect 8316 5682 8372 5694
rect 8316 5630 8318 5682
rect 8370 5630 8372 5682
rect 8316 5348 8372 5630
rect 8316 5282 8372 5292
rect 9100 5684 9156 5694
rect 8428 5236 8484 5246
rect 9100 5236 9156 5628
rect 8428 5234 9044 5236
rect 8428 5182 8430 5234
rect 8482 5182 9044 5234
rect 8428 5180 9044 5182
rect 8428 5170 8484 5180
rect 8988 5122 9044 5180
rect 9100 5142 9156 5180
rect 9772 5236 9828 5246
rect 9772 5142 9828 5180
rect 8988 5070 8990 5122
rect 9042 5070 9044 5122
rect 8988 5058 9044 5070
rect 9660 5124 9716 5134
rect 9660 5030 9716 5068
rect 10332 5124 10388 5852
rect 10444 5682 10500 5694
rect 10444 5630 10446 5682
rect 10498 5630 10500 5682
rect 10444 5236 10500 5630
rect 10444 5142 10500 5180
rect 10332 4992 10388 5068
rect 9836 4732 10100 4742
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 9836 4666 10100 4676
rect 9996 4452 10052 4462
rect 8092 3666 8260 3668
rect 8092 3614 8094 3666
rect 8146 3614 8260 3666
rect 8092 3612 8260 3614
rect 8652 4338 8708 4350
rect 8652 4286 8654 4338
rect 8706 4286 8708 4338
rect 8092 3602 8148 3612
rect 7196 3502 7198 3554
rect 7250 3502 7252 3554
rect 7196 3490 7252 3502
rect 7420 3556 7476 3566
rect 6748 3378 6804 3388
rect 5524 3164 5788 3174
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5524 3098 5788 3108
rect 2492 2604 2772 2660
rect 2492 800 2548 2604
rect 7420 800 7476 3500
rect 8652 3556 8708 4286
rect 9884 4116 9940 4126
rect 9884 3668 9940 4060
rect 9996 3778 10052 4396
rect 10220 4116 10276 4126
rect 10220 4022 10276 4060
rect 9996 3726 9998 3778
rect 10050 3726 10052 3778
rect 9996 3714 10052 3726
rect 10668 3778 10724 5964
rect 10892 5908 10948 6524
rect 11004 6468 11060 6478
rect 11004 6374 11060 6412
rect 11116 6132 11172 7196
rect 11452 6580 11508 7422
rect 12012 8146 12068 8158
rect 12012 8094 12014 8146
rect 12066 8094 12068 8146
rect 11564 7252 11620 7262
rect 12012 7252 12068 8094
rect 12348 7474 12404 8204
rect 12572 8194 12628 8204
rect 14476 8258 14532 8270
rect 14476 8206 14478 8258
rect 14530 8206 14532 8258
rect 13692 8146 13748 8158
rect 13692 8094 13694 8146
rect 13746 8094 13748 8146
rect 12348 7422 12350 7474
rect 12402 7422 12404 7474
rect 12348 7410 12404 7422
rect 13580 8034 13636 8046
rect 13580 7982 13582 8034
rect 13634 7982 13636 8034
rect 12908 7364 12964 7374
rect 13580 7364 13636 7982
rect 13692 7476 13748 8094
rect 14148 7868 14412 7878
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14148 7802 14412 7812
rect 13804 7476 13860 7486
rect 13692 7420 13804 7476
rect 12908 7362 13636 7364
rect 12908 7310 12910 7362
rect 12962 7310 13636 7362
rect 12908 7308 13636 7310
rect 11564 7250 11732 7252
rect 11564 7198 11566 7250
rect 11618 7198 11732 7250
rect 11564 7196 11732 7198
rect 12012 7196 12404 7252
rect 11564 7186 11620 7196
rect 11564 6580 11620 6590
rect 11452 6578 11620 6580
rect 11452 6526 11566 6578
rect 11618 6526 11620 6578
rect 11452 6524 11620 6526
rect 11116 6038 11172 6076
rect 11004 5908 11060 5918
rect 10892 5852 11004 5908
rect 11564 5908 11620 6524
rect 11676 6468 11732 7196
rect 11992 7084 12256 7094
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 11992 7018 12256 7028
rect 12236 6578 12292 6590
rect 12236 6526 12238 6578
rect 12290 6526 12292 6578
rect 11676 6466 11844 6468
rect 11676 6414 11678 6466
rect 11730 6414 11844 6466
rect 11676 6412 11844 6414
rect 11676 6402 11732 6412
rect 11788 6132 11844 6412
rect 11676 5908 11732 5918
rect 11564 5852 11676 5908
rect 10780 5236 10836 5246
rect 10780 4562 10836 5180
rect 10780 4510 10782 4562
rect 10834 4510 10836 4562
rect 10780 4498 10836 4510
rect 11004 5122 11060 5852
rect 11116 5236 11172 5246
rect 11116 5142 11172 5180
rect 11452 5236 11508 5246
rect 11004 5070 11006 5122
rect 11058 5070 11060 5122
rect 10892 4452 10948 4462
rect 11004 4452 11060 5070
rect 11452 4562 11508 5180
rect 11452 4510 11454 4562
rect 11506 4510 11508 4562
rect 11452 4498 11508 4510
rect 11676 5122 11732 5852
rect 11676 5070 11678 5122
rect 11730 5070 11732 5122
rect 10892 4450 11060 4452
rect 10892 4398 10894 4450
rect 10946 4398 11060 4450
rect 10892 4396 11060 4398
rect 11564 4452 11620 4462
rect 11676 4452 11732 5070
rect 11788 5682 11844 6076
rect 12236 5908 12292 6526
rect 12348 6468 12404 7196
rect 12404 6412 12516 6468
rect 12348 6336 12404 6412
rect 12348 5908 12404 5918
rect 12236 5852 12348 5908
rect 11788 5630 11790 5682
rect 11842 5630 11844 5682
rect 11788 5124 11844 5630
rect 11992 5516 12256 5526
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 11992 5450 12256 5460
rect 11788 5058 11844 5068
rect 11900 5236 11956 5246
rect 11788 4900 11844 4910
rect 11900 4900 11956 5180
rect 12348 5122 12404 5852
rect 12460 5684 12516 6412
rect 12908 5684 12964 7308
rect 13692 6692 13748 6702
rect 13804 6692 13860 7420
rect 14476 7476 14532 8206
rect 15148 8146 15204 8158
rect 15148 8094 15150 8146
rect 15202 8094 15204 8146
rect 14588 7476 14644 7486
rect 14476 7420 14588 7476
rect 13692 6690 13860 6692
rect 13692 6638 13694 6690
rect 13746 6638 13860 6690
rect 13692 6636 13860 6638
rect 14364 6692 14420 6702
rect 14476 6692 14532 7420
rect 14588 7382 14644 7420
rect 14364 6690 14532 6692
rect 14364 6638 14366 6690
rect 14418 6638 14532 6690
rect 14364 6636 14532 6638
rect 15036 6804 15092 6814
rect 15036 6690 15092 6748
rect 15036 6638 15038 6690
rect 15090 6638 15092 6690
rect 13692 6018 13748 6636
rect 14364 6626 14420 6636
rect 14812 6580 14868 6590
rect 13692 5966 13694 6018
rect 13746 5966 13748 6018
rect 13020 5908 13076 5918
rect 13020 5814 13076 5852
rect 13692 5908 13748 5966
rect 13132 5684 13188 5694
rect 12460 5682 12628 5684
rect 12460 5630 12462 5682
rect 12514 5630 12628 5682
rect 12460 5628 12628 5630
rect 12908 5682 13188 5684
rect 12908 5630 13134 5682
rect 13186 5630 13188 5682
rect 12908 5628 13188 5630
rect 12460 5618 12516 5628
rect 12572 5236 12628 5628
rect 12572 5170 12628 5180
rect 12908 5236 12964 5246
rect 12348 5070 12350 5122
rect 12402 5070 12404 5122
rect 12348 5058 12404 5070
rect 12460 5124 12516 5134
rect 11788 4898 11956 4900
rect 11788 4846 11790 4898
rect 11842 4846 11956 4898
rect 11788 4844 11956 4846
rect 11788 4834 11844 4844
rect 11564 4450 11732 4452
rect 11564 4398 11566 4450
rect 11618 4398 11732 4450
rect 11564 4396 11732 4398
rect 10892 4386 10948 4396
rect 11564 4386 11620 4396
rect 12012 4340 12068 4350
rect 11788 4338 12068 4340
rect 11788 4286 12014 4338
rect 12066 4286 12068 4338
rect 11788 4284 12068 4286
rect 10668 3726 10670 3778
rect 10722 3726 10724 3778
rect 10668 3714 10724 3726
rect 11116 3780 11172 3790
rect 9884 3602 9940 3612
rect 8652 3424 8708 3500
rect 11116 3554 11172 3724
rect 11116 3502 11118 3554
rect 11170 3502 11172 3554
rect 11116 3490 11172 3502
rect 11788 3444 11844 4284
rect 12012 4274 12068 4284
rect 11992 3948 12256 3958
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 11992 3882 12256 3892
rect 12460 3780 12516 5068
rect 12908 4450 12964 5180
rect 13132 5124 13188 5628
rect 13132 5058 13188 5068
rect 13580 5684 13636 5694
rect 12908 4398 12910 4450
rect 12962 4398 12964 4450
rect 12908 4386 12964 4398
rect 12012 3724 12516 3780
rect 12572 4340 12628 4350
rect 12012 3666 12068 3724
rect 12012 3614 12014 3666
rect 12066 3614 12068 3666
rect 12012 3602 12068 3614
rect 12572 3556 12628 4284
rect 13468 4340 13524 4350
rect 13468 4246 13524 4284
rect 11788 3378 11844 3388
rect 12348 3554 12628 3556
rect 12348 3502 12574 3554
rect 12626 3502 12628 3554
rect 12348 3500 12628 3502
rect 13580 3556 13636 5628
rect 13692 5122 13748 5852
rect 13804 6466 13860 6478
rect 13804 6414 13806 6466
rect 13858 6414 13860 6466
rect 13804 5684 13860 6414
rect 14476 6468 14532 6478
rect 14148 6300 14412 6310
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14148 6234 14412 6244
rect 14476 6130 14532 6412
rect 14476 6078 14478 6130
rect 14530 6078 14532 6130
rect 14476 6066 14532 6078
rect 14364 5908 14420 5918
rect 13804 5682 13972 5684
rect 13804 5630 13806 5682
rect 13858 5630 13972 5682
rect 13804 5628 13972 5630
rect 13804 5618 13860 5628
rect 13916 5236 13972 5628
rect 13916 5170 13972 5180
rect 13692 5070 13694 5122
rect 13746 5070 13748 5122
rect 13692 5058 13748 5070
rect 13804 5124 13860 5134
rect 13692 3556 13748 3566
rect 13580 3554 13748 3556
rect 13580 3502 13694 3554
rect 13746 3502 13748 3554
rect 13580 3500 13748 3502
rect 9836 3164 10100 3174
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 9836 3098 10100 3108
rect 12348 800 12404 3500
rect 12572 3490 12628 3500
rect 13692 3490 13748 3500
rect 13580 3332 13636 3342
rect 13804 3332 13860 5068
rect 14364 5122 14420 5852
rect 14588 5908 14644 5918
rect 14476 5236 14532 5246
rect 14476 5142 14532 5180
rect 14364 5070 14366 5122
rect 14418 5070 14420 5122
rect 14364 5058 14420 5070
rect 14148 4732 14412 4742
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14148 4666 14412 4676
rect 14476 4338 14532 4350
rect 14476 4286 14478 4338
rect 14530 4286 14532 4338
rect 14364 4228 14420 4238
rect 14476 4228 14532 4286
rect 14364 4226 14532 4228
rect 14364 4174 14366 4226
rect 14418 4174 14532 4226
rect 14364 4172 14532 4174
rect 14364 4162 14420 4172
rect 14588 3892 14644 5852
rect 14812 4338 14868 6524
rect 15036 6018 15092 6638
rect 15148 6468 15204 8094
rect 15148 6374 15204 6412
rect 15260 7362 15316 8316
rect 15932 8372 15988 8382
rect 15820 8260 15876 8270
rect 15260 7310 15262 7362
rect 15314 7310 15316 7362
rect 15036 5966 15038 6018
rect 15090 5966 15092 6018
rect 15036 5954 15092 5966
rect 15148 5684 15204 5694
rect 15260 5684 15316 7310
rect 15708 7476 15764 7486
rect 15708 6804 15764 7420
rect 15820 7474 15876 8204
rect 15820 7422 15822 7474
rect 15874 7422 15876 7474
rect 15820 7410 15876 7422
rect 15820 6916 15876 6926
rect 15932 6916 15988 8316
rect 16604 8372 16660 8382
rect 16492 8148 16548 8158
rect 16492 7476 16548 8092
rect 16604 7700 16660 8316
rect 17276 8260 17332 11200
rect 17276 8194 17332 8204
rect 17836 8932 17892 8942
rect 17836 8484 17892 8876
rect 17500 8148 17556 8158
rect 17500 8054 17556 8092
rect 17612 8034 17668 8046
rect 17612 7982 17614 8034
rect 17666 7982 17668 8034
rect 16716 7700 16772 7710
rect 16604 7698 16772 7700
rect 16604 7646 16718 7698
rect 16770 7646 16772 7698
rect 16604 7644 16772 7646
rect 16716 7634 16772 7644
rect 17612 7588 17668 7982
rect 17836 7698 17892 8428
rect 18460 7868 18724 7878
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18460 7802 18724 7812
rect 17836 7646 17838 7698
rect 17890 7646 17892 7698
rect 17836 7634 17892 7646
rect 17500 7532 17668 7588
rect 16604 7476 16660 7486
rect 16548 7474 16660 7476
rect 16548 7422 16606 7474
rect 16658 7422 16660 7474
rect 16548 7420 16660 7422
rect 16492 7344 16548 7420
rect 16604 7410 16660 7420
rect 16304 7084 16568 7094
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16304 7018 16568 7028
rect 15820 6914 15988 6916
rect 15820 6862 15822 6914
rect 15874 6862 15988 6914
rect 15820 6860 15988 6862
rect 15820 6850 15876 6860
rect 15708 6690 15764 6748
rect 15708 6638 15710 6690
rect 15762 6638 15764 6690
rect 15708 6626 15764 6638
rect 16380 6580 16436 6590
rect 16380 6486 16436 6524
rect 17052 6578 17108 6590
rect 17052 6526 17054 6578
rect 17106 6526 17108 6578
rect 15820 6468 15876 6478
rect 15820 6130 15876 6412
rect 16492 6468 16548 6478
rect 16492 6374 16548 6412
rect 15820 6078 15822 6130
rect 15874 6078 15876 6130
rect 15708 5908 15764 5918
rect 15708 5814 15764 5852
rect 15148 5682 15316 5684
rect 15148 5630 15150 5682
rect 15202 5630 15316 5682
rect 15148 5628 15316 5630
rect 15148 5460 15204 5628
rect 15148 5394 15204 5404
rect 14924 5348 14980 5358
rect 14924 4450 14980 5292
rect 15708 5236 15764 5246
rect 15148 5234 15764 5236
rect 15148 5182 15710 5234
rect 15762 5182 15764 5234
rect 15148 5180 15764 5182
rect 15036 5124 15092 5134
rect 15036 4898 15092 5068
rect 15148 5122 15204 5180
rect 15708 5170 15764 5180
rect 15148 5070 15150 5122
rect 15202 5070 15204 5122
rect 15148 5058 15204 5070
rect 15036 4846 15038 4898
rect 15090 4846 15092 4898
rect 15036 4564 15092 4846
rect 15708 4564 15764 4574
rect 15820 4564 15876 6078
rect 16156 5796 16212 5806
rect 16156 5124 16212 5740
rect 16492 5796 16548 5806
rect 16492 5702 16548 5740
rect 17052 5796 17108 6526
rect 17164 6468 17220 6478
rect 17276 6468 17332 6478
rect 17164 6466 17276 6468
rect 17164 6414 17166 6466
rect 17218 6414 17276 6466
rect 17164 6412 17276 6414
rect 17164 6402 17220 6412
rect 17052 5730 17108 5740
rect 16304 5516 16568 5526
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16304 5450 16568 5460
rect 16380 5124 16436 5134
rect 16156 5122 16436 5124
rect 16156 5070 16382 5122
rect 16434 5070 16436 5122
rect 16156 5068 16436 5070
rect 16380 5058 16436 5068
rect 16492 5124 16548 5134
rect 15036 4562 15876 4564
rect 15036 4510 15038 4562
rect 15090 4510 15710 4562
rect 15762 4510 15876 4562
rect 15036 4508 15876 4510
rect 16380 4564 16436 4574
rect 16492 4564 16548 5068
rect 17276 5122 17332 6412
rect 17500 6468 17556 7532
rect 17724 7476 17780 7486
rect 17612 7474 17780 7476
rect 17612 7422 17726 7474
rect 17778 7422 17780 7474
rect 17612 7420 17780 7422
rect 17612 6692 17668 7420
rect 17724 7410 17780 7420
rect 17612 6626 17668 6636
rect 17500 6402 17556 6412
rect 17724 6578 17780 6590
rect 17724 6526 17726 6578
rect 17778 6526 17780 6578
rect 17724 6020 17780 6526
rect 17836 6468 17892 6478
rect 17836 6374 17892 6412
rect 18460 6300 18724 6310
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18460 6234 18724 6244
rect 17724 5954 17780 5964
rect 17724 5684 17780 5694
rect 17724 5590 17780 5628
rect 17276 5070 17278 5122
rect 17330 5070 17332 5122
rect 16380 4562 16548 4564
rect 16380 4510 16382 4562
rect 16434 4510 16548 4562
rect 16380 4508 16548 4510
rect 16828 5012 16884 5022
rect 15036 4498 15092 4508
rect 15708 4498 15764 4508
rect 14924 4398 14926 4450
rect 14978 4398 14980 4450
rect 14924 4386 14980 4398
rect 16268 4452 16324 4462
rect 16268 4358 16324 4396
rect 14812 4286 14814 4338
rect 14866 4286 14868 4338
rect 14812 4274 14868 4286
rect 15596 4338 15652 4350
rect 15596 4286 15598 4338
rect 15650 4286 15652 4338
rect 15596 4116 15652 4286
rect 16380 4116 16436 4508
rect 15596 4050 15652 4060
rect 15932 4060 16436 4116
rect 14364 3836 14644 3892
rect 14364 3778 14420 3836
rect 14364 3726 14366 3778
rect 14418 3726 14420 3778
rect 14364 3714 14420 3726
rect 15148 3668 15204 3678
rect 15148 3554 15204 3612
rect 15932 3666 15988 4060
rect 16304 3948 16568 3958
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16304 3882 16568 3892
rect 15932 3614 15934 3666
rect 15986 3614 15988 3666
rect 15932 3602 15988 3614
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3490 15204 3502
rect 16716 3556 16772 3566
rect 16828 3556 16884 4956
rect 16716 3554 16884 3556
rect 16716 3502 16718 3554
rect 16770 3502 16884 3554
rect 16716 3500 16884 3502
rect 16716 3490 16772 3500
rect 13580 3330 13860 3332
rect 13580 3278 13582 3330
rect 13634 3278 13860 3330
rect 13580 3276 13860 3278
rect 13580 3266 13636 3276
rect 14148 3164 14412 3174
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14148 3098 14412 3108
rect 16828 2772 16884 3500
rect 17276 2996 17332 5070
rect 17724 5124 17780 5134
rect 17724 4788 17780 5068
rect 17836 5122 17892 5134
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5012 17892 5070
rect 17836 4946 17892 4956
rect 17724 4732 17892 4788
rect 17836 4562 17892 4732
rect 18460 4732 18724 4742
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18460 4666 18724 4676
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 17724 4338 17780 4350
rect 17724 4286 17726 4338
rect 17778 4286 17780 4338
rect 17724 4228 17780 4286
rect 17724 4162 17780 4172
rect 17500 3780 17556 3790
rect 17500 3686 17556 3724
rect 18460 3164 18724 3174
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18460 3098 18724 3108
rect 17276 2930 17332 2940
rect 16828 2716 17332 2772
rect 17276 800 17332 2716
rect 2464 0 2576 800
rect 7392 0 7504 800
rect 12320 0 12432 800
rect 17248 0 17360 800
<< via2 >>
rect 2044 8316 2100 8372
rect 1820 8146 1876 8148
rect 1820 8094 1822 8146
rect 1822 8094 1874 8146
rect 1874 8094 1876 8146
rect 1820 8092 1876 8094
rect 1932 7868 1988 7924
rect 1932 7698 1988 7700
rect 1932 7646 1934 7698
rect 1934 7646 1986 7698
rect 1986 7646 1988 7698
rect 1932 7644 1988 7646
rect 1820 6524 1876 6580
rect 3368 8650 3424 8652
rect 3368 8598 3370 8650
rect 3370 8598 3422 8650
rect 3422 8598 3424 8650
rect 3368 8596 3424 8598
rect 3472 8650 3528 8652
rect 3472 8598 3474 8650
rect 3474 8598 3526 8650
rect 3526 8598 3528 8650
rect 3472 8596 3528 8598
rect 3576 8650 3632 8652
rect 3576 8598 3578 8650
rect 3578 8598 3630 8650
rect 3630 8598 3632 8650
rect 3576 8596 3632 8598
rect 7680 8650 7736 8652
rect 7680 8598 7682 8650
rect 7682 8598 7734 8650
rect 7734 8598 7736 8650
rect 7680 8596 7736 8598
rect 7784 8650 7840 8652
rect 7784 8598 7786 8650
rect 7786 8598 7838 8650
rect 7838 8598 7840 8650
rect 7784 8596 7840 8598
rect 7888 8650 7944 8652
rect 7888 8598 7890 8650
rect 7890 8598 7942 8650
rect 7942 8598 7944 8650
rect 7888 8596 7944 8598
rect 11992 8650 12048 8652
rect 11992 8598 11994 8650
rect 11994 8598 12046 8650
rect 12046 8598 12048 8650
rect 11992 8596 12048 8598
rect 12096 8650 12152 8652
rect 12096 8598 12098 8650
rect 12098 8598 12150 8650
rect 12150 8598 12152 8650
rect 12096 8596 12152 8598
rect 12200 8650 12256 8652
rect 12200 8598 12202 8650
rect 12202 8598 12254 8650
rect 12254 8598 12256 8650
rect 12200 8596 12256 8598
rect 2044 7420 2100 7476
rect 2156 7980 2212 8036
rect 3276 7644 3332 7700
rect 3052 7308 3108 7364
rect 2716 7196 2772 7252
rect 2492 6914 2548 6916
rect 2492 6862 2494 6914
rect 2494 6862 2546 6914
rect 2546 6862 2548 6914
rect 2492 6860 2548 6862
rect 3052 6860 3108 6916
rect 2380 6130 2436 6132
rect 2380 6078 2382 6130
rect 2382 6078 2434 6130
rect 2434 6078 2436 6130
rect 2380 6076 2436 6078
rect 1820 4956 1876 5012
rect 3388 7868 3444 7924
rect 3724 7868 3780 7924
rect 3368 7082 3424 7084
rect 3368 7030 3370 7082
rect 3370 7030 3422 7082
rect 3422 7030 3424 7082
rect 3368 7028 3424 7030
rect 3472 7082 3528 7084
rect 3472 7030 3474 7082
rect 3474 7030 3526 7082
rect 3526 7030 3528 7082
rect 3472 7028 3528 7030
rect 3576 7082 3632 7084
rect 3576 7030 3578 7082
rect 3578 7030 3630 7082
rect 3630 7030 3632 7082
rect 3576 7028 3632 7030
rect 3276 6578 3332 6580
rect 3276 6526 3278 6578
rect 3278 6526 3330 6578
rect 3330 6526 3332 6578
rect 3276 6524 3332 6526
rect 3612 6076 3668 6132
rect 3164 5852 3220 5908
rect 3368 5514 3424 5516
rect 3368 5462 3370 5514
rect 3370 5462 3422 5514
rect 3422 5462 3424 5514
rect 3368 5460 3424 5462
rect 3472 5514 3528 5516
rect 3472 5462 3474 5514
rect 3474 5462 3526 5514
rect 3526 5462 3528 5514
rect 3472 5460 3528 5462
rect 3576 5514 3632 5516
rect 3576 5462 3578 5514
rect 3578 5462 3630 5514
rect 3630 5462 3632 5514
rect 3576 5460 3632 5462
rect 2940 4956 2996 5012
rect 3368 3946 3424 3948
rect 3368 3894 3370 3946
rect 3370 3894 3422 3946
rect 3422 3894 3424 3946
rect 3368 3892 3424 3894
rect 3472 3946 3528 3948
rect 3472 3894 3474 3946
rect 3474 3894 3526 3946
rect 3526 3894 3528 3946
rect 3472 3892 3528 3894
rect 3576 3946 3632 3948
rect 3576 3894 3578 3946
rect 3578 3894 3630 3946
rect 3630 3894 3632 3946
rect 3576 3892 3632 3894
rect 4620 8146 4676 8148
rect 4620 8094 4622 8146
rect 4622 8094 4674 8146
rect 4674 8094 4676 8146
rect 4620 8092 4676 8094
rect 4956 8034 5012 8036
rect 4956 7982 4958 8034
rect 4958 7982 5010 8034
rect 5010 7982 5012 8034
rect 4956 7980 5012 7982
rect 6636 8034 6692 8036
rect 6636 7982 6638 8034
rect 6638 7982 6690 8034
rect 6690 7982 6692 8034
rect 6636 7980 6692 7982
rect 5524 7866 5580 7868
rect 5524 7814 5526 7866
rect 5526 7814 5578 7866
rect 5578 7814 5580 7866
rect 5524 7812 5580 7814
rect 5628 7866 5684 7868
rect 5628 7814 5630 7866
rect 5630 7814 5682 7866
rect 5682 7814 5684 7866
rect 5628 7812 5684 7814
rect 5732 7866 5788 7868
rect 5732 7814 5734 7866
rect 5734 7814 5786 7866
rect 5786 7814 5788 7866
rect 5732 7812 5788 7814
rect 4732 7474 4788 7476
rect 4732 7422 4734 7474
rect 4734 7422 4786 7474
rect 4786 7422 4788 7474
rect 4732 7420 4788 7422
rect 4172 7308 4228 7364
rect 7532 7980 7588 8036
rect 6748 7308 6804 7364
rect 4620 7250 4676 7252
rect 4620 7198 4622 7250
rect 4622 7198 4674 7250
rect 4674 7198 4676 7250
rect 4620 7196 4676 7198
rect 6300 6748 6356 6804
rect 4956 6636 5012 6692
rect 5524 6298 5580 6300
rect 5524 6246 5526 6298
rect 5526 6246 5578 6298
rect 5578 6246 5580 6298
rect 5524 6244 5580 6246
rect 5628 6298 5684 6300
rect 5628 6246 5630 6298
rect 5630 6246 5682 6298
rect 5682 6246 5684 6298
rect 5628 6244 5684 6246
rect 5732 6298 5788 6300
rect 5732 6246 5734 6298
rect 5734 6246 5786 6298
rect 5786 6246 5788 6298
rect 5732 6244 5788 6246
rect 8092 7980 8148 8036
rect 9836 7866 9892 7868
rect 9836 7814 9838 7866
rect 9838 7814 9890 7866
rect 9890 7814 9892 7866
rect 9836 7812 9892 7814
rect 9940 7866 9996 7868
rect 9940 7814 9942 7866
rect 9942 7814 9994 7866
rect 9994 7814 9996 7866
rect 9940 7812 9996 7814
rect 10044 7866 10100 7868
rect 10044 7814 10046 7866
rect 10046 7814 10098 7866
rect 10098 7814 10100 7866
rect 10044 7812 10100 7814
rect 7680 7082 7736 7084
rect 7680 7030 7682 7082
rect 7682 7030 7734 7082
rect 7734 7030 7736 7082
rect 7680 7028 7736 7030
rect 7784 7082 7840 7084
rect 7784 7030 7786 7082
rect 7786 7030 7838 7082
rect 7838 7030 7840 7082
rect 7784 7028 7840 7030
rect 7888 7082 7944 7084
rect 7888 7030 7890 7082
rect 7890 7030 7942 7082
rect 7942 7030 7944 7082
rect 7888 7028 7944 7030
rect 7644 6914 7700 6916
rect 7644 6862 7646 6914
rect 7646 6862 7698 6914
rect 7698 6862 7700 6914
rect 7644 6860 7700 6862
rect 6860 6802 6916 6804
rect 6860 6750 6862 6802
rect 6862 6750 6914 6802
rect 6914 6750 6916 6802
rect 6860 6748 6916 6750
rect 6748 6524 6804 6580
rect 7532 6578 7588 6580
rect 7532 6526 7534 6578
rect 7534 6526 7586 6578
rect 7586 6526 7588 6578
rect 7532 6524 7588 6526
rect 6188 5906 6244 5908
rect 6188 5854 6190 5906
rect 6190 5854 6242 5906
rect 6242 5854 6244 5906
rect 6188 5852 6244 5854
rect 6860 5906 6916 5908
rect 6860 5854 6862 5906
rect 6862 5854 6914 5906
rect 6914 5854 6916 5906
rect 6860 5852 6916 5854
rect 5628 5794 5684 5796
rect 5628 5742 5630 5794
rect 5630 5742 5682 5794
rect 5682 5742 5684 5794
rect 5628 5740 5684 5742
rect 6412 5346 6468 5348
rect 6412 5294 6414 5346
rect 6414 5294 6466 5346
rect 6466 5294 6468 5346
rect 6412 5292 6468 5294
rect 7420 5852 7476 5908
rect 7644 5906 7700 5908
rect 7644 5854 7646 5906
rect 7646 5854 7698 5906
rect 7698 5854 7700 5906
rect 7644 5852 7700 5854
rect 8316 6914 8372 6916
rect 8316 6862 8318 6914
rect 8318 6862 8370 6914
rect 8370 6862 8372 6914
rect 8316 6860 8372 6862
rect 8204 6578 8260 6580
rect 8204 6526 8206 6578
rect 8206 6526 8258 6578
rect 8258 6526 8260 6578
rect 8204 6524 8260 6526
rect 8316 6412 8372 6468
rect 8876 6578 8932 6580
rect 8876 6526 8878 6578
rect 8878 6526 8930 6578
rect 8930 6526 8932 6578
rect 8876 6524 8932 6526
rect 9548 6578 9604 6580
rect 9548 6526 9550 6578
rect 9550 6526 9602 6578
rect 9602 6526 9604 6578
rect 9548 6524 9604 6526
rect 10108 6524 10164 6580
rect 8988 6466 9044 6468
rect 8988 6414 8990 6466
rect 8990 6414 9042 6466
rect 9042 6414 9044 6466
rect 8988 6412 9044 6414
rect 8988 6130 9044 6132
rect 8988 6078 8990 6130
rect 8990 6078 9042 6130
rect 9042 6078 9044 6130
rect 8988 6076 9044 6078
rect 9836 6298 9892 6300
rect 9836 6246 9838 6298
rect 9838 6246 9890 6298
rect 9890 6246 9892 6298
rect 9836 6244 9892 6246
rect 9940 6298 9996 6300
rect 9940 6246 9942 6298
rect 9942 6246 9994 6298
rect 9994 6246 9996 6298
rect 9940 6244 9996 6246
rect 10044 6298 10100 6300
rect 10044 6246 10046 6298
rect 10046 6246 10098 6298
rect 10098 6246 10100 6298
rect 10044 6244 10100 6246
rect 9660 6076 9716 6132
rect 8092 5852 8148 5908
rect 8092 5628 8148 5684
rect 16304 8650 16360 8652
rect 16304 8598 16306 8650
rect 16306 8598 16358 8650
rect 16358 8598 16360 8650
rect 16304 8596 16360 8598
rect 16408 8650 16464 8652
rect 16408 8598 16410 8650
rect 16410 8598 16462 8650
rect 16462 8598 16464 8650
rect 16408 8596 16464 8598
rect 16512 8650 16568 8652
rect 16512 8598 16514 8650
rect 16514 8598 16566 8650
rect 16566 8598 16568 8650
rect 16512 8596 16568 8598
rect 15260 8316 15316 8372
rect 10332 6466 10388 6468
rect 10332 6414 10334 6466
rect 10334 6414 10386 6466
rect 10386 6414 10388 6466
rect 10332 6412 10388 6414
rect 10668 5964 10724 6020
rect 10332 5906 10388 5908
rect 10332 5854 10334 5906
rect 10334 5854 10386 5906
rect 10386 5854 10388 5906
rect 10332 5852 10388 5854
rect 7680 5514 7736 5516
rect 7680 5462 7682 5514
rect 7682 5462 7734 5514
rect 7734 5462 7736 5514
rect 7680 5460 7736 5462
rect 7784 5514 7840 5516
rect 7784 5462 7786 5514
rect 7786 5462 7838 5514
rect 7838 5462 7840 5514
rect 7784 5460 7840 5462
rect 7888 5514 7944 5516
rect 7888 5462 7890 5514
rect 7890 5462 7942 5514
rect 7942 5462 7944 5514
rect 7888 5460 7944 5462
rect 7532 5292 7588 5348
rect 5524 4730 5580 4732
rect 5524 4678 5526 4730
rect 5526 4678 5578 4730
rect 5578 4678 5580 4730
rect 5524 4676 5580 4678
rect 5628 4730 5684 4732
rect 5628 4678 5630 4730
rect 5630 4678 5682 4730
rect 5682 4678 5684 4730
rect 5628 4676 5684 4678
rect 5732 4730 5788 4732
rect 5732 4678 5734 4730
rect 5734 4678 5786 4730
rect 5786 4678 5788 4730
rect 5732 4676 5788 4678
rect 5964 4284 6020 4340
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 6636 4226 6692 4228
rect 6636 4174 6638 4226
rect 6638 4174 6690 4226
rect 6690 4174 6692 4226
rect 6636 4172 6692 4174
rect 5292 4114 5348 4116
rect 5292 4062 5294 4114
rect 5294 4062 5346 4114
rect 5346 4062 5348 4114
rect 5292 4060 5348 4062
rect 7680 3946 7736 3948
rect 7680 3894 7682 3946
rect 7682 3894 7734 3946
rect 7734 3894 7736 3946
rect 7680 3892 7736 3894
rect 7784 3946 7840 3948
rect 7784 3894 7786 3946
rect 7786 3894 7838 3946
rect 7838 3894 7840 3946
rect 7784 3892 7840 3894
rect 7888 3946 7944 3948
rect 7888 3894 7890 3946
rect 7890 3894 7942 3946
rect 7942 3894 7944 3946
rect 7888 3892 7944 3894
rect 8092 3836 8148 3892
rect 6076 3778 6132 3780
rect 6076 3726 6078 3778
rect 6078 3726 6130 3778
rect 6130 3726 6132 3778
rect 6076 3724 6132 3726
rect 4956 3666 5012 3668
rect 4956 3614 4958 3666
rect 4958 3614 5010 3666
rect 5010 3614 5012 3666
rect 4956 3612 5012 3614
rect 2716 3500 2772 3556
rect 1820 2940 1876 2996
rect 4060 3554 4116 3556
rect 4060 3502 4062 3554
rect 4062 3502 4114 3554
rect 4114 3502 4116 3554
rect 4060 3500 4116 3502
rect 7196 3612 7252 3668
rect 8316 5292 8372 5348
rect 9100 5628 9156 5684
rect 9100 5234 9156 5236
rect 9100 5182 9102 5234
rect 9102 5182 9154 5234
rect 9154 5182 9156 5234
rect 9100 5180 9156 5182
rect 9772 5234 9828 5236
rect 9772 5182 9774 5234
rect 9774 5182 9826 5234
rect 9826 5182 9828 5234
rect 9772 5180 9828 5182
rect 9660 5122 9716 5124
rect 9660 5070 9662 5122
rect 9662 5070 9714 5122
rect 9714 5070 9716 5122
rect 9660 5068 9716 5070
rect 10444 5234 10500 5236
rect 10444 5182 10446 5234
rect 10446 5182 10498 5234
rect 10498 5182 10500 5234
rect 10444 5180 10500 5182
rect 10332 5122 10388 5124
rect 10332 5070 10334 5122
rect 10334 5070 10386 5122
rect 10386 5070 10388 5122
rect 10332 5068 10388 5070
rect 9836 4730 9892 4732
rect 9836 4678 9838 4730
rect 9838 4678 9890 4730
rect 9890 4678 9892 4730
rect 9836 4676 9892 4678
rect 9940 4730 9996 4732
rect 9940 4678 9942 4730
rect 9942 4678 9994 4730
rect 9994 4678 9996 4730
rect 9940 4676 9996 4678
rect 10044 4730 10100 4732
rect 10044 4678 10046 4730
rect 10046 4678 10098 4730
rect 10098 4678 10100 4730
rect 10044 4676 10100 4678
rect 9996 4396 10052 4452
rect 7420 3500 7476 3556
rect 6748 3388 6804 3444
rect 5524 3162 5580 3164
rect 5524 3110 5526 3162
rect 5526 3110 5578 3162
rect 5578 3110 5580 3162
rect 5524 3108 5580 3110
rect 5628 3162 5684 3164
rect 5628 3110 5630 3162
rect 5630 3110 5682 3162
rect 5682 3110 5684 3162
rect 5628 3108 5684 3110
rect 5732 3162 5788 3164
rect 5732 3110 5734 3162
rect 5734 3110 5786 3162
rect 5786 3110 5788 3162
rect 5732 3108 5788 3110
rect 9884 4060 9940 4116
rect 10220 4114 10276 4116
rect 10220 4062 10222 4114
rect 10222 4062 10274 4114
rect 10274 4062 10276 4114
rect 10220 4060 10276 4062
rect 11004 6466 11060 6468
rect 11004 6414 11006 6466
rect 11006 6414 11058 6466
rect 11058 6414 11060 6466
rect 11004 6412 11060 6414
rect 14148 7866 14204 7868
rect 14148 7814 14150 7866
rect 14150 7814 14202 7866
rect 14202 7814 14204 7866
rect 14148 7812 14204 7814
rect 14252 7866 14308 7868
rect 14252 7814 14254 7866
rect 14254 7814 14306 7866
rect 14306 7814 14308 7866
rect 14252 7812 14308 7814
rect 14356 7866 14412 7868
rect 14356 7814 14358 7866
rect 14358 7814 14410 7866
rect 14410 7814 14412 7866
rect 14356 7812 14412 7814
rect 13804 7474 13860 7476
rect 13804 7422 13806 7474
rect 13806 7422 13858 7474
rect 13858 7422 13860 7474
rect 13804 7420 13860 7422
rect 11116 6130 11172 6132
rect 11116 6078 11118 6130
rect 11118 6078 11170 6130
rect 11170 6078 11172 6130
rect 11116 6076 11172 6078
rect 11004 5906 11060 5908
rect 11004 5854 11006 5906
rect 11006 5854 11058 5906
rect 11058 5854 11060 5906
rect 11004 5852 11060 5854
rect 11992 7082 12048 7084
rect 11992 7030 11994 7082
rect 11994 7030 12046 7082
rect 12046 7030 12048 7082
rect 11992 7028 12048 7030
rect 12096 7082 12152 7084
rect 12096 7030 12098 7082
rect 12098 7030 12150 7082
rect 12150 7030 12152 7082
rect 12096 7028 12152 7030
rect 12200 7082 12256 7084
rect 12200 7030 12202 7082
rect 12202 7030 12254 7082
rect 12254 7030 12256 7082
rect 12200 7028 12256 7030
rect 11788 6076 11844 6132
rect 11676 5906 11732 5908
rect 11676 5854 11678 5906
rect 11678 5854 11730 5906
rect 11730 5854 11732 5906
rect 11676 5852 11732 5854
rect 10780 5180 10836 5236
rect 11116 5234 11172 5236
rect 11116 5182 11118 5234
rect 11118 5182 11170 5234
rect 11170 5182 11172 5234
rect 11116 5180 11172 5182
rect 11452 5180 11508 5236
rect 12348 6466 12404 6468
rect 12348 6414 12350 6466
rect 12350 6414 12402 6466
rect 12402 6414 12404 6466
rect 12348 6412 12404 6414
rect 12348 5906 12404 5908
rect 12348 5854 12350 5906
rect 12350 5854 12402 5906
rect 12402 5854 12404 5906
rect 12348 5852 12404 5854
rect 11992 5514 12048 5516
rect 11992 5462 11994 5514
rect 11994 5462 12046 5514
rect 12046 5462 12048 5514
rect 11992 5460 12048 5462
rect 12096 5514 12152 5516
rect 12096 5462 12098 5514
rect 12098 5462 12150 5514
rect 12150 5462 12152 5514
rect 12096 5460 12152 5462
rect 12200 5514 12256 5516
rect 12200 5462 12202 5514
rect 12202 5462 12254 5514
rect 12254 5462 12256 5514
rect 12200 5460 12256 5462
rect 11788 5068 11844 5124
rect 11900 5180 11956 5236
rect 14588 7474 14644 7476
rect 14588 7422 14590 7474
rect 14590 7422 14642 7474
rect 14642 7422 14644 7474
rect 14588 7420 14644 7422
rect 15036 6748 15092 6804
rect 14812 6524 14868 6580
rect 13020 5906 13076 5908
rect 13020 5854 13022 5906
rect 13022 5854 13074 5906
rect 13074 5854 13076 5906
rect 13020 5852 13076 5854
rect 13692 5852 13748 5908
rect 12572 5180 12628 5236
rect 12908 5180 12964 5236
rect 12460 5122 12516 5124
rect 12460 5070 12462 5122
rect 12462 5070 12514 5122
rect 12514 5070 12516 5122
rect 12460 5068 12516 5070
rect 11116 3724 11172 3780
rect 9884 3612 9940 3668
rect 8652 3554 8708 3556
rect 8652 3502 8654 3554
rect 8654 3502 8706 3554
rect 8706 3502 8708 3554
rect 8652 3500 8708 3502
rect 11992 3946 12048 3948
rect 11992 3894 11994 3946
rect 11994 3894 12046 3946
rect 12046 3894 12048 3946
rect 11992 3892 12048 3894
rect 12096 3946 12152 3948
rect 12096 3894 12098 3946
rect 12098 3894 12150 3946
rect 12150 3894 12152 3946
rect 12096 3892 12152 3894
rect 12200 3946 12256 3948
rect 12200 3894 12202 3946
rect 12202 3894 12254 3946
rect 12254 3894 12256 3946
rect 12200 3892 12256 3894
rect 13132 5068 13188 5124
rect 13580 5628 13636 5684
rect 12572 4284 12628 4340
rect 13468 4338 13524 4340
rect 13468 4286 13470 4338
rect 13470 4286 13522 4338
rect 13522 4286 13524 4338
rect 13468 4284 13524 4286
rect 11788 3388 11844 3444
rect 14476 6466 14532 6468
rect 14476 6414 14478 6466
rect 14478 6414 14530 6466
rect 14530 6414 14532 6466
rect 14476 6412 14532 6414
rect 14148 6298 14204 6300
rect 14148 6246 14150 6298
rect 14150 6246 14202 6298
rect 14202 6246 14204 6298
rect 14148 6244 14204 6246
rect 14252 6298 14308 6300
rect 14252 6246 14254 6298
rect 14254 6246 14306 6298
rect 14306 6246 14308 6298
rect 14252 6244 14308 6246
rect 14356 6298 14412 6300
rect 14356 6246 14358 6298
rect 14358 6246 14410 6298
rect 14410 6246 14412 6298
rect 14356 6244 14412 6246
rect 14364 5906 14420 5908
rect 14364 5854 14366 5906
rect 14366 5854 14418 5906
rect 14418 5854 14420 5906
rect 14364 5852 14420 5854
rect 13916 5180 13972 5236
rect 13804 5122 13860 5124
rect 13804 5070 13806 5122
rect 13806 5070 13858 5122
rect 13858 5070 13860 5122
rect 13804 5068 13860 5070
rect 9836 3162 9892 3164
rect 9836 3110 9838 3162
rect 9838 3110 9890 3162
rect 9890 3110 9892 3162
rect 9836 3108 9892 3110
rect 9940 3162 9996 3164
rect 9940 3110 9942 3162
rect 9942 3110 9994 3162
rect 9994 3110 9996 3162
rect 9940 3108 9996 3110
rect 10044 3162 10100 3164
rect 10044 3110 10046 3162
rect 10046 3110 10098 3162
rect 10098 3110 10100 3162
rect 10044 3108 10100 3110
rect 14588 5852 14644 5908
rect 14476 5234 14532 5236
rect 14476 5182 14478 5234
rect 14478 5182 14530 5234
rect 14530 5182 14532 5234
rect 14476 5180 14532 5182
rect 14148 4730 14204 4732
rect 14148 4678 14150 4730
rect 14150 4678 14202 4730
rect 14202 4678 14204 4730
rect 14148 4676 14204 4678
rect 14252 4730 14308 4732
rect 14252 4678 14254 4730
rect 14254 4678 14306 4730
rect 14306 4678 14308 4730
rect 14252 4676 14308 4678
rect 14356 4730 14412 4732
rect 14356 4678 14358 4730
rect 14358 4678 14410 4730
rect 14410 4678 14412 4730
rect 14356 4676 14412 4678
rect 15148 6466 15204 6468
rect 15148 6414 15150 6466
rect 15150 6414 15202 6466
rect 15202 6414 15204 6466
rect 15148 6412 15204 6414
rect 15932 8316 15988 8372
rect 15820 8258 15876 8260
rect 15820 8206 15822 8258
rect 15822 8206 15874 8258
rect 15874 8206 15876 8258
rect 15820 8204 15876 8206
rect 15708 7420 15764 7476
rect 16604 8370 16660 8372
rect 16604 8318 16606 8370
rect 16606 8318 16658 8370
rect 16658 8318 16660 8370
rect 16604 8316 16660 8318
rect 16492 8146 16548 8148
rect 16492 8094 16494 8146
rect 16494 8094 16546 8146
rect 16546 8094 16548 8146
rect 16492 8092 16548 8094
rect 17276 8204 17332 8260
rect 17836 8876 17892 8932
rect 17836 8428 17892 8484
rect 17500 8146 17556 8148
rect 17500 8094 17502 8146
rect 17502 8094 17554 8146
rect 17554 8094 17556 8146
rect 17500 8092 17556 8094
rect 18460 7866 18516 7868
rect 18460 7814 18462 7866
rect 18462 7814 18514 7866
rect 18514 7814 18516 7866
rect 18460 7812 18516 7814
rect 18564 7866 18620 7868
rect 18564 7814 18566 7866
rect 18566 7814 18618 7866
rect 18618 7814 18620 7866
rect 18564 7812 18620 7814
rect 18668 7866 18724 7868
rect 18668 7814 18670 7866
rect 18670 7814 18722 7866
rect 18722 7814 18724 7866
rect 18668 7812 18724 7814
rect 16492 7420 16548 7476
rect 16304 7082 16360 7084
rect 16304 7030 16306 7082
rect 16306 7030 16358 7082
rect 16358 7030 16360 7082
rect 16304 7028 16360 7030
rect 16408 7082 16464 7084
rect 16408 7030 16410 7082
rect 16410 7030 16462 7082
rect 16462 7030 16464 7082
rect 16408 7028 16464 7030
rect 16512 7082 16568 7084
rect 16512 7030 16514 7082
rect 16514 7030 16566 7082
rect 16566 7030 16568 7082
rect 16512 7028 16568 7030
rect 15708 6748 15764 6804
rect 16380 6578 16436 6580
rect 16380 6526 16382 6578
rect 16382 6526 16434 6578
rect 16434 6526 16436 6578
rect 16380 6524 16436 6526
rect 15820 6412 15876 6468
rect 16492 6466 16548 6468
rect 16492 6414 16494 6466
rect 16494 6414 16546 6466
rect 16546 6414 16548 6466
rect 16492 6412 16548 6414
rect 15708 5906 15764 5908
rect 15708 5854 15710 5906
rect 15710 5854 15762 5906
rect 15762 5854 15764 5906
rect 15708 5852 15764 5854
rect 15148 5404 15204 5460
rect 14924 5292 14980 5348
rect 15036 5068 15092 5124
rect 16156 5740 16212 5796
rect 16492 5794 16548 5796
rect 16492 5742 16494 5794
rect 16494 5742 16546 5794
rect 16546 5742 16548 5794
rect 16492 5740 16548 5742
rect 17276 6412 17332 6468
rect 17052 5740 17108 5796
rect 16304 5514 16360 5516
rect 16304 5462 16306 5514
rect 16306 5462 16358 5514
rect 16358 5462 16360 5514
rect 16304 5460 16360 5462
rect 16408 5514 16464 5516
rect 16408 5462 16410 5514
rect 16410 5462 16462 5514
rect 16462 5462 16464 5514
rect 16408 5460 16464 5462
rect 16512 5514 16568 5516
rect 16512 5462 16514 5514
rect 16514 5462 16566 5514
rect 16566 5462 16568 5514
rect 16512 5460 16568 5462
rect 16492 5068 16548 5124
rect 17612 6636 17668 6692
rect 17500 6412 17556 6468
rect 17836 6466 17892 6468
rect 17836 6414 17838 6466
rect 17838 6414 17890 6466
rect 17890 6414 17892 6466
rect 17836 6412 17892 6414
rect 18460 6298 18516 6300
rect 18460 6246 18462 6298
rect 18462 6246 18514 6298
rect 18514 6246 18516 6298
rect 18460 6244 18516 6246
rect 18564 6298 18620 6300
rect 18564 6246 18566 6298
rect 18566 6246 18618 6298
rect 18618 6246 18620 6298
rect 18564 6244 18620 6246
rect 18668 6298 18724 6300
rect 18668 6246 18670 6298
rect 18670 6246 18722 6298
rect 18722 6246 18724 6298
rect 18668 6244 18724 6246
rect 17724 5964 17780 6020
rect 17724 5682 17780 5684
rect 17724 5630 17726 5682
rect 17726 5630 17778 5682
rect 17778 5630 17780 5682
rect 17724 5628 17780 5630
rect 16828 4956 16884 5012
rect 16268 4450 16324 4452
rect 16268 4398 16270 4450
rect 16270 4398 16322 4450
rect 16322 4398 16324 4450
rect 16268 4396 16324 4398
rect 15596 4060 15652 4116
rect 15148 3612 15204 3668
rect 16304 3946 16360 3948
rect 16304 3894 16306 3946
rect 16306 3894 16358 3946
rect 16358 3894 16360 3946
rect 16304 3892 16360 3894
rect 16408 3946 16464 3948
rect 16408 3894 16410 3946
rect 16410 3894 16462 3946
rect 16462 3894 16464 3946
rect 16408 3892 16464 3894
rect 16512 3946 16568 3948
rect 16512 3894 16514 3946
rect 16514 3894 16566 3946
rect 16566 3894 16568 3946
rect 16512 3892 16568 3894
rect 14148 3162 14204 3164
rect 14148 3110 14150 3162
rect 14150 3110 14202 3162
rect 14202 3110 14204 3162
rect 14148 3108 14204 3110
rect 14252 3162 14308 3164
rect 14252 3110 14254 3162
rect 14254 3110 14306 3162
rect 14306 3110 14308 3162
rect 14252 3108 14308 3110
rect 14356 3162 14412 3164
rect 14356 3110 14358 3162
rect 14358 3110 14410 3162
rect 14410 3110 14412 3162
rect 14356 3108 14412 3110
rect 17724 5068 17780 5124
rect 17836 4956 17892 5012
rect 18460 4730 18516 4732
rect 18460 4678 18462 4730
rect 18462 4678 18514 4730
rect 18514 4678 18516 4730
rect 18460 4676 18516 4678
rect 18564 4730 18620 4732
rect 18564 4678 18566 4730
rect 18566 4678 18618 4730
rect 18618 4678 18620 4730
rect 18564 4676 18620 4678
rect 18668 4730 18724 4732
rect 18668 4678 18670 4730
rect 18670 4678 18722 4730
rect 18722 4678 18724 4730
rect 18668 4676 18724 4678
rect 17724 4172 17780 4228
rect 17500 3778 17556 3780
rect 17500 3726 17502 3778
rect 17502 3726 17554 3778
rect 17554 3726 17556 3778
rect 17500 3724 17556 3726
rect 18460 3162 18516 3164
rect 18460 3110 18462 3162
rect 18462 3110 18514 3162
rect 18514 3110 18516 3162
rect 18460 3108 18516 3110
rect 18564 3162 18620 3164
rect 18564 3110 18566 3162
rect 18566 3110 18618 3162
rect 18618 3110 18620 3162
rect 18564 3108 18620 3110
rect 18668 3162 18724 3164
rect 18668 3110 18670 3162
rect 18670 3110 18722 3162
rect 18722 3110 18724 3162
rect 18668 3108 18724 3110
rect 17276 2940 17332 2996
<< metal3 >>
rect 0 8932 800 8960
rect 19200 8932 20000 8960
rect 0 8876 2100 8932
rect 17826 8876 17836 8932
rect 17892 8876 20000 8932
rect 0 8848 800 8876
rect 2044 8372 2100 8876
rect 19200 8848 20000 8876
rect 3358 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3642 8652
rect 7670 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7954 8652
rect 11982 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12266 8652
rect 16294 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16578 8652
rect 15260 8428 17836 8484
rect 17892 8428 17902 8484
rect 15260 8372 15316 8428
rect 15820 8372 15876 8428
rect 16716 8372 16772 8428
rect 2034 8316 2044 8372
rect 2100 8316 2110 8372
rect 15250 8316 15260 8372
rect 15316 8316 15326 8372
rect 15820 8316 15932 8372
rect 15988 8316 15998 8372
rect 16594 8316 16604 8372
rect 16660 8316 16772 8372
rect 15810 8204 15820 8260
rect 15876 8204 17276 8260
rect 17332 8204 17342 8260
rect 1810 8092 1820 8148
rect 1876 8092 4620 8148
rect 4676 8092 4686 8148
rect 16482 8092 16492 8148
rect 16548 8092 17500 8148
rect 17556 8092 17566 8148
rect 2146 7980 2156 8036
rect 2212 7980 4956 8036
rect 5012 7980 5022 8036
rect 5292 7980 6636 8036
rect 6692 7980 7532 8036
rect 7588 7980 8092 8036
rect 8148 7980 8158 8036
rect 5292 7924 5348 7980
rect 1922 7868 1932 7924
rect 1988 7868 3388 7924
rect 3444 7868 3724 7924
rect 3780 7868 5348 7924
rect 5514 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5798 7868
rect 9826 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10110 7868
rect 14138 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14422 7868
rect 18450 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18734 7868
rect 1922 7644 1932 7700
rect 1988 7644 3276 7700
rect 3332 7644 3342 7700
rect 2034 7420 2044 7476
rect 2100 7420 4732 7476
rect 4788 7420 4798 7476
rect 13794 7420 13804 7476
rect 13860 7420 14588 7476
rect 14644 7420 15708 7476
rect 15764 7420 16492 7476
rect 16548 7420 16558 7476
rect 3042 7308 3052 7364
rect 3108 7308 4172 7364
rect 4228 7308 6748 7364
rect 6804 7308 6814 7364
rect 2706 7196 2716 7252
rect 2772 7196 4620 7252
rect 4676 7196 4686 7252
rect 3358 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3642 7084
rect 7670 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7954 7084
rect 11982 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12266 7084
rect 16294 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16578 7084
rect 2482 6860 2492 6916
rect 2548 6860 3052 6916
rect 3108 6860 3118 6916
rect 7634 6860 7644 6916
rect 7700 6860 8316 6916
rect 8372 6860 8382 6916
rect 6290 6748 6300 6804
rect 6356 6748 6860 6804
rect 6916 6748 6926 6804
rect 15026 6748 15036 6804
rect 15092 6748 15708 6804
rect 15764 6748 15774 6804
rect 4946 6636 4956 6692
rect 5012 6636 17612 6692
rect 17668 6636 17678 6692
rect 1810 6524 1820 6580
rect 1876 6524 3276 6580
rect 3332 6524 3342 6580
rect 6738 6524 6748 6580
rect 6804 6524 7532 6580
rect 7588 6524 8204 6580
rect 8260 6524 8876 6580
rect 8932 6524 9548 6580
rect 9604 6524 10108 6580
rect 10164 6524 10174 6580
rect 14802 6524 14812 6580
rect 14868 6524 16380 6580
rect 16436 6524 16446 6580
rect 8306 6412 8316 6468
rect 8372 6412 8988 6468
rect 9044 6412 9054 6468
rect 10322 6412 10332 6468
rect 10388 6412 11004 6468
rect 11060 6412 12348 6468
rect 12404 6412 12414 6468
rect 14466 6412 14476 6468
rect 14532 6412 15148 6468
rect 15204 6412 15820 6468
rect 15876 6412 16492 6468
rect 16548 6412 17276 6468
rect 17332 6412 17500 6468
rect 17556 6412 17836 6468
rect 17892 6412 17902 6468
rect 5514 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5798 6300
rect 9826 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10110 6300
rect 14138 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14422 6300
rect 18450 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18734 6300
rect 2370 6076 2380 6132
rect 2436 6076 3612 6132
rect 3668 6076 3678 6132
rect 8978 6076 8988 6132
rect 9044 6076 9660 6132
rect 9716 6076 11116 6132
rect 11172 6076 11788 6132
rect 11844 6076 11854 6132
rect 10658 5964 10668 6020
rect 10724 5964 17724 6020
rect 17780 5964 17790 6020
rect 3154 5852 3164 5908
rect 3220 5852 6188 5908
rect 6244 5852 6860 5908
rect 6916 5852 7420 5908
rect 7476 5852 7644 5908
rect 7700 5852 8092 5908
rect 8148 5852 8158 5908
rect 10322 5852 10332 5908
rect 10388 5852 11004 5908
rect 11060 5852 11676 5908
rect 11732 5852 12348 5908
rect 12404 5852 13020 5908
rect 13076 5852 13692 5908
rect 13748 5852 14364 5908
rect 14420 5852 14430 5908
rect 14578 5852 14588 5908
rect 14644 5852 15708 5908
rect 15764 5852 15774 5908
rect 5618 5740 5628 5796
rect 5684 5740 16156 5796
rect 16212 5740 16222 5796
rect 16482 5740 16492 5796
rect 16548 5740 17052 5796
rect 17108 5740 17118 5796
rect 8082 5628 8092 5684
rect 8148 5628 9100 5684
rect 9156 5628 9166 5684
rect 13570 5628 13580 5684
rect 13636 5628 17724 5684
rect 17780 5628 17790 5684
rect 3358 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3642 5516
rect 7670 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7954 5516
rect 11982 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12266 5516
rect 16294 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16578 5516
rect 15138 5404 15148 5460
rect 15204 5404 15214 5460
rect 6402 5292 6412 5348
rect 6468 5292 7532 5348
rect 7588 5292 7598 5348
rect 8306 5292 8316 5348
rect 8372 5292 14924 5348
rect 14980 5292 14990 5348
rect 15148 5236 15204 5404
rect 9090 5180 9100 5236
rect 9156 5180 9772 5236
rect 9828 5180 10444 5236
rect 10500 5180 10780 5236
rect 10836 5180 11116 5236
rect 11172 5180 11452 5236
rect 11508 5180 11900 5236
rect 11956 5180 12572 5236
rect 12628 5180 12908 5236
rect 12964 5180 13916 5236
rect 13972 5180 14476 5236
rect 14532 5180 16548 5236
rect 16492 5124 16548 5180
rect 9650 5068 9660 5124
rect 9716 5068 10332 5124
rect 10388 5068 10398 5124
rect 11778 5068 11788 5124
rect 11844 5068 12460 5124
rect 12516 5068 13132 5124
rect 13188 5068 13804 5124
rect 13860 5068 15036 5124
rect 15092 5068 15102 5124
rect 16482 5068 16492 5124
rect 16548 5068 17724 5124
rect 17780 5068 17790 5124
rect 1810 4956 1820 5012
rect 1876 4956 2940 5012
rect 2996 4956 3006 5012
rect 16818 4956 16828 5012
rect 16884 4956 17836 5012
rect 17892 4956 17902 5012
rect 5514 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5798 4732
rect 9826 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10110 4732
rect 14138 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14422 4732
rect 18450 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18734 4732
rect 9986 4396 9996 4452
rect 10052 4396 16268 4452
rect 16324 4396 16334 4452
rect 5954 4284 5964 4340
rect 6020 4284 7084 4340
rect 7140 4284 7150 4340
rect 12562 4284 12572 4340
rect 12628 4284 13468 4340
rect 13524 4284 13534 4340
rect 6626 4172 6636 4228
rect 6692 4172 17724 4228
rect 17780 4172 17790 4228
rect 5282 4060 5292 4116
rect 5348 4060 9884 4116
rect 9940 4060 9950 4116
rect 10210 4060 10220 4116
rect 10276 4060 15596 4116
rect 15652 4060 15662 4116
rect 8372 3948 11844 4004
rect 3358 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3642 3948
rect 7670 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7954 3948
rect 8372 3892 8428 3948
rect 8082 3836 8092 3892
rect 8148 3836 8428 3892
rect 11788 3780 11844 3948
rect 11982 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12266 3948
rect 16294 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16578 3948
rect 6066 3724 6076 3780
rect 6132 3724 11116 3780
rect 11172 3724 11182 3780
rect 11788 3724 17500 3780
rect 17556 3724 17566 3780
rect 4946 3612 4956 3668
rect 5012 3612 7196 3668
rect 7252 3612 7262 3668
rect 9874 3612 9884 3668
rect 9940 3612 15148 3668
rect 15204 3612 15214 3668
rect 2706 3500 2716 3556
rect 2772 3500 4060 3556
rect 4116 3500 4126 3556
rect 7410 3500 7420 3556
rect 7476 3500 8652 3556
rect 8708 3500 8718 3556
rect 6738 3388 6748 3444
rect 6804 3388 11788 3444
rect 11844 3388 11854 3444
rect 5514 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5798 3164
rect 9826 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10110 3164
rect 14138 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14422 3164
rect 18450 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18734 3164
rect 0 2996 800 3024
rect 19200 2996 20000 3024
rect 0 2940 1820 2996
rect 1876 2940 1886 2996
rect 17266 2940 17276 2996
rect 17332 2940 20000 2996
rect 0 2912 800 2940
rect 19200 2912 20000 2940
<< via3 >>
rect 3368 8596 3424 8652
rect 3472 8596 3528 8652
rect 3576 8596 3632 8652
rect 7680 8596 7736 8652
rect 7784 8596 7840 8652
rect 7888 8596 7944 8652
rect 11992 8596 12048 8652
rect 12096 8596 12152 8652
rect 12200 8596 12256 8652
rect 16304 8596 16360 8652
rect 16408 8596 16464 8652
rect 16512 8596 16568 8652
rect 5524 7812 5580 7868
rect 5628 7812 5684 7868
rect 5732 7812 5788 7868
rect 9836 7812 9892 7868
rect 9940 7812 9996 7868
rect 10044 7812 10100 7868
rect 14148 7812 14204 7868
rect 14252 7812 14308 7868
rect 14356 7812 14412 7868
rect 18460 7812 18516 7868
rect 18564 7812 18620 7868
rect 18668 7812 18724 7868
rect 3368 7028 3424 7084
rect 3472 7028 3528 7084
rect 3576 7028 3632 7084
rect 7680 7028 7736 7084
rect 7784 7028 7840 7084
rect 7888 7028 7944 7084
rect 11992 7028 12048 7084
rect 12096 7028 12152 7084
rect 12200 7028 12256 7084
rect 16304 7028 16360 7084
rect 16408 7028 16464 7084
rect 16512 7028 16568 7084
rect 5524 6244 5580 6300
rect 5628 6244 5684 6300
rect 5732 6244 5788 6300
rect 9836 6244 9892 6300
rect 9940 6244 9996 6300
rect 10044 6244 10100 6300
rect 14148 6244 14204 6300
rect 14252 6244 14308 6300
rect 14356 6244 14412 6300
rect 18460 6244 18516 6300
rect 18564 6244 18620 6300
rect 18668 6244 18724 6300
rect 3368 5460 3424 5516
rect 3472 5460 3528 5516
rect 3576 5460 3632 5516
rect 7680 5460 7736 5516
rect 7784 5460 7840 5516
rect 7888 5460 7944 5516
rect 11992 5460 12048 5516
rect 12096 5460 12152 5516
rect 12200 5460 12256 5516
rect 16304 5460 16360 5516
rect 16408 5460 16464 5516
rect 16512 5460 16568 5516
rect 5524 4676 5580 4732
rect 5628 4676 5684 4732
rect 5732 4676 5788 4732
rect 9836 4676 9892 4732
rect 9940 4676 9996 4732
rect 10044 4676 10100 4732
rect 14148 4676 14204 4732
rect 14252 4676 14308 4732
rect 14356 4676 14412 4732
rect 18460 4676 18516 4732
rect 18564 4676 18620 4732
rect 18668 4676 18724 4732
rect 3368 3892 3424 3948
rect 3472 3892 3528 3948
rect 3576 3892 3632 3948
rect 7680 3892 7736 3948
rect 7784 3892 7840 3948
rect 7888 3892 7944 3948
rect 11992 3892 12048 3948
rect 12096 3892 12152 3948
rect 12200 3892 12256 3948
rect 16304 3892 16360 3948
rect 16408 3892 16464 3948
rect 16512 3892 16568 3948
rect 5524 3108 5580 3164
rect 5628 3108 5684 3164
rect 5732 3108 5788 3164
rect 9836 3108 9892 3164
rect 9940 3108 9996 3164
rect 10044 3108 10100 3164
rect 14148 3108 14204 3164
rect 14252 3108 14308 3164
rect 14356 3108 14412 3164
rect 18460 3108 18516 3164
rect 18564 3108 18620 3164
rect 18668 3108 18724 3164
<< metal4 >>
rect 3340 8652 3660 8684
rect 3340 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3660 8652
rect 3340 7084 3660 8596
rect 3340 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3660 7084
rect 3340 5516 3660 7028
rect 3340 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3660 5516
rect 3340 3948 3660 5460
rect 3340 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3660 3948
rect 3340 3076 3660 3892
rect 5496 7868 5816 8684
rect 5496 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5816 7868
rect 5496 6300 5816 7812
rect 5496 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5816 6300
rect 5496 4732 5816 6244
rect 5496 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5816 4732
rect 5496 3164 5816 4676
rect 5496 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5816 3164
rect 5496 3076 5816 3108
rect 7652 8652 7972 8684
rect 7652 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7972 8652
rect 7652 7084 7972 8596
rect 7652 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7972 7084
rect 7652 5516 7972 7028
rect 7652 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7972 5516
rect 7652 3948 7972 5460
rect 7652 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7972 3948
rect 7652 3076 7972 3892
rect 9808 7868 10128 8684
rect 9808 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10128 7868
rect 9808 6300 10128 7812
rect 9808 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10128 6300
rect 9808 4732 10128 6244
rect 9808 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10128 4732
rect 9808 3164 10128 4676
rect 9808 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10128 3164
rect 9808 3076 10128 3108
rect 11964 8652 12284 8684
rect 11964 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12284 8652
rect 11964 7084 12284 8596
rect 11964 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12284 7084
rect 11964 5516 12284 7028
rect 11964 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12284 5516
rect 11964 3948 12284 5460
rect 11964 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12284 3948
rect 11964 3076 12284 3892
rect 14120 7868 14440 8684
rect 14120 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14440 7868
rect 14120 6300 14440 7812
rect 14120 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14440 6300
rect 14120 4732 14440 6244
rect 14120 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14440 4732
rect 14120 3164 14440 4676
rect 14120 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14440 3164
rect 14120 3076 14440 3108
rect 16276 8652 16596 8684
rect 16276 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16596 8652
rect 16276 7084 16596 8596
rect 16276 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16596 7084
rect 16276 5516 16596 7028
rect 16276 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16596 5516
rect 16276 3948 16596 5460
rect 16276 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16596 3948
rect 16276 3076 16596 3892
rect 18432 7868 18752 8684
rect 18432 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18752 7868
rect 18432 6300 18752 7812
rect 18432 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18752 6300
rect 18432 4732 18752 6244
rect 18432 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18752 4732
rect 18432 3164 18752 4676
rect 18432 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18752 3164
rect 18432 3076 18752 3108
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9
timestamp 1667941163
transform 1 0 2352 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28
timestamp 1667941163
transform 1 0 4480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1667941163
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39
timestamp 1667941163
transform 1 0 5712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44
timestamp 1667941163
transform 1 0 6272 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50
timestamp 1667941163
transform 1 0 6944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1667941163
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74
timestamp 1667941163
transform 1 0 9632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79
timestamp 1667941163
transform 1 0 10192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 10864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1667941163
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112
timestamp 1667941163
transform 1 0 13888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 14560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1667941163
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147
timestamp 1667941163
transform 1 0 17808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_151
timestamp 1667941163
transform 1 0 18256 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_10
timestamp 1667941163
transform 1 0 2464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_28
timestamp 1667941163
transform 1 0 4480 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_32
timestamp 1667941163
transform 1 0 4928 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_37
timestamp 1667941163
transform 1 0 5488 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_43
timestamp 1667941163
transform 1 0 6160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_49
timestamp 1667941163
transform 1 0 6832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1667941163
transform 1 0 8960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_73
timestamp 1667941163
transform 1 0 9520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_81
timestamp 1667941163
transform 1 0 10416 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_87
timestamp 1667941163
transform 1 0 11088 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_93
timestamp 1667941163
transform 1 0 11760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1667941163
transform 1 0 13888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_118
timestamp 1667941163
transform 1 0 14560 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_124
timestamp 1667941163
transform 1 0 15232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_130
timestamp 1667941163
transform 1 0 15904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_136
timestamp 1667941163
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_140
timestamp 1667941163
transform 1 0 17024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1667941163
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_149
timestamp 1667941163
transform 1 0 18032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_151
timestamp 1667941163
transform 1 0 18256 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_18
timestamp 1667941163
transform 1 0 3360 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_22
timestamp 1667941163
transform 1 0 3808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_28
timestamp 1667941163
transform 1 0 4480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1667941163
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_41
timestamp 1667941163
transform 1 0 5936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_47
timestamp 1667941163
transform 1 0 6608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_53
timestamp 1667941163
transform 1 0 7280 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_59
timestamp 1667941163
transform 1 0 7952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_65
timestamp 1667941163
transform 1 0 8624 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_71
timestamp 1667941163
transform 1 0 9296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_77
timestamp 1667941163
transform 1 0 9968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_83
timestamp 1667941163
transform 1 0 10640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_89
timestamp 1667941163
transform 1 0 11312 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_95
timestamp 1667941163
transform 1 0 11984 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1667941163
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1667941163
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_113
timestamp 1667941163
transform 1 0 14000 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_119
timestamp 1667941163
transform 1 0 14672 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_125
timestamp 1667941163
transform 1 0 15344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_131
timestamp 1667941163
transform 1 0 16016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_133
timestamp 1667941163
transform 1 0 16240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_151
timestamp 1667941163
transform 1 0 18256 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_11
timestamp 1667941163
transform 1 0 2576 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_17
timestamp 1667941163
transform 1 0 3248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_33
timestamp 1667941163
transform 1 0 5040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_35
timestamp 1667941163
transform 1 0 5264 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_40
timestamp 1667941163
transform 1 0 5824 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_46
timestamp 1667941163
transform 1 0 6496 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_52
timestamp 1667941163
transform 1 0 7168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_58
timestamp 1667941163
transform 1 0 7840 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_64
timestamp 1667941163
transform 1 0 8512 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_73
timestamp 1667941163
transform 1 0 9520 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_77
timestamp 1667941163
transform 1 0 9968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_83
timestamp 1667941163
transform 1 0 10640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_89
timestamp 1667941163
transform 1 0 11312 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_95
timestamp 1667941163
transform 1 0 11984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_101
timestamp 1667941163
transform 1 0 12656 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_107
timestamp 1667941163
transform 1 0 13328 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 14000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_119
timestamp 1667941163
transform 1 0 14672 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_125
timestamp 1667941163
transform 1 0 15344 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_131
timestamp 1667941163
transform 1 0 16016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1667941163
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_149
timestamp 1667941163
transform 1 0 18032 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_151
timestamp 1667941163
transform 1 0 18256 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1667941163
transform 1 0 1568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1667941163
transform 1 0 2912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_22
timestamp 1667941163
transform 1 0 3808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_30
timestamp 1667941163
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_37
timestamp 1667941163
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_45
timestamp 1667941163
transform 1 0 6384 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_47
timestamp 1667941163
transform 1 0 6608 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_52
timestamp 1667941163
transform 1 0 7168 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_58
timestamp 1667941163
transform 1 0 7840 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_64
timestamp 1667941163
transform 1 0 8512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_70
timestamp 1667941163
transform 1 0 9184 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_76
timestamp 1667941163
transform 1 0 9856 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 10528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_88
timestamp 1667941163
transform 1 0 11200 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_94
timestamp 1667941163
transform 1 0 11872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_100
timestamp 1667941163
transform 1 0 12544 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_104
timestamp 1667941163
transform 1 0 12992 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1667941163
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_113
timestamp 1667941163
transform 1 0 14000 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_119
timestamp 1667941163
transform 1 0 14672 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_125
timestamp 1667941163
transform 1 0 15344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_131
timestamp 1667941163
transform 1 0 16016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_137
timestamp 1667941163
transform 1 0 16688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_143
timestamp 1667941163
transform 1 0 17360 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_149
timestamp 1667941163
transform 1 0 18032 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_151
timestamp 1667941163
transform 1 0 18256 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1667941163
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_7
timestamp 1667941163
transform 1 0 2128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_26
timestamp 1667941163
transform 1 0 4256 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_32
timestamp 1667941163
transform 1 0 4928 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_48
timestamp 1667941163
transform 1 0 6720 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_69
timestamp 1667941163
transform 1 0 9072 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_73
timestamp 1667941163
transform 1 0 9520 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_81
timestamp 1667941163
transform 1 0 10416 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_87
timestamp 1667941163
transform 1 0 11088 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_93
timestamp 1667941163
transform 1 0 11760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_112
timestamp 1667941163
transform 1 0 13888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_133
timestamp 1667941163
transform 1 0 16240 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_139
timestamp 1667941163
transform 1 0 16912 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1667941163
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_149
timestamp 1667941163
transform 1 0 18032 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_151
timestamp 1667941163
transform 1 0 18256 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1667941163
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_7
timestamp 1667941163
transform 1 0 2128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 4256 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_37
timestamp 1667941163
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_45
timestamp 1667941163
transform 1 0 6384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_50
timestamp 1667941163
transform 1 0 6944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_69
timestamp 1667941163
transform 1 0 9072 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_72
timestamp 1667941163
transform 1 0 9408 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_74
timestamp 1667941163
transform 1 0 9632 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_79
timestamp 1667941163
transform 1 0 10192 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 10864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1667941163
transform 1 0 12992 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_107
timestamp 1667941163
transform 1 0 13328 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_112
timestamp 1667941163
transform 1 0 13888 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_114
timestamp 1667941163
transform 1 0 14112 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_132
timestamp 1667941163
transform 1 0 16128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 16800 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_142
timestamp 1667941163
transform 1 0 17248 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_147
timestamp 1667941163
transform 1 0 17808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_151
timestamp 1667941163
transform 1 0 18256 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 18592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 18592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 18592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 18592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_14 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_15
timestamp 1667941163
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_16
timestamp 1667941163
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_17
timestamp 1667941163
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18
timestamp 1667941163
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1667941163
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1667941163
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1667941163
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_23
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24
timestamp 1667941163
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1667941163
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1667941163
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1667941163
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1667941163
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1667941163
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1667941163
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1667941163
transform 1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _29_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2800 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _30_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 2912 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _31_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 5152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _32_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1680 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _33_
timestamp 1667941163
transform -1 0 3808 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _34_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 9744 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _35_
timestamp 1667941163
transform 1 0 14112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _36_
timestamp 1667941163
transform -1 0 17808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _37_
timestamp 1667941163
transform 1 0 8064 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _38_
timestamp 1667941163
transform 1 0 6160 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _39_
timestamp 1667941163
transform 1 0 9968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _40_
timestamp 1667941163
transform -1 0 7280 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _41_
timestamp 1667941163
transform 1 0 16240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _42_
timestamp 1667941163
transform 1 0 8176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _43_
timestamp 1667941163
transform -1 0 16016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _44_
timestamp 1667941163
transform -1 0 7168 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _45_
timestamp 1667941163
transform 1 0 10416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _46_
timestamp 1667941163
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _47_
timestamp 1667941163
transform 1 0 14112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _48_
timestamp 1667941163
transform 1 0 6384 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _49_
timestamp 1667941163
transform -1 0 18032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _50_
timestamp 1667941163
transform 1 0 4032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _51_
timestamp 1667941163
transform 1 0 1904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _52_
timestamp 1667941163
transform 1 0 5712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _53_
timestamp 1667941163
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _54_
timestamp 1667941163
transform 1 0 6496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _55_
timestamp 1667941163
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _56_
timestamp 1667941163
transform 1 0 5040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _57_
timestamp 1667941163
transform 1 0 5376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[0\].pdn
timestamp 1667941163
transform 1 0 16128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[0\].pdp
timestamp 1667941163
transform 1 0 16240 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[1\].pdn
timestamp 1667941163
transform -1 0 7952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[1\].pdp
timestamp 1667941163
transform 1 0 14784 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[2\].pdn
timestamp 1667941163
transform 1 0 7392 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[2\].pdp
timestamp 1667941163
transform 1 0 15456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[3\].pdn
timestamp 1667941163
transform -1 0 7168 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[3\].pdp
timestamp 1667941163
transform 1 0 16912 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[4\].pdn
timestamp 1667941163
transform 1 0 8848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[4\].pdp
timestamp 1667941163
transform -1 0 15344 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[5\].pdn
timestamp 1667941163
transform -1 0 6496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[5\].pdp
timestamp 1667941163
transform 1 0 17584 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[6\].pdn
timestamp 1667941163
transform 1 0 17584 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[6\].pdp
timestamp 1667941163
transform 1 0 15568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[7\].pdn
timestamp 1667941163
transform 1 0 17584 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PD\[7\].pdp
timestamp 1667941163
transform -1 0 13888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[0\].pun
timestamp 1667941163
transform 1 0 11536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[0\].pup
timestamp 1667941163
transform 1 0 8736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[1\].pun
timestamp 1667941163
transform 1 0 9744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[1\].pup
timestamp 1667941163
transform 1 0 14224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[2\].pun
timestamp 1667941163
transform 1 0 10192 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[2\].pup
timestamp 1667941163
transform 1 0 11536 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[3\].pun
timestamp 1667941163
transform 1 0 15568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[3\].pup
timestamp 1667941163
transform 1 0 9408 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[4\].pun
timestamp 1667941163
transform 1 0 9520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[4\].pup
timestamp 1667941163
transform 1 0 10640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[5\].pun
timestamp 1667941163
transform 1 0 10864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[5\].pup
timestamp 1667941163
transform -1 0 13888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[6\].pun
timestamp 1667941163
transform 1 0 13552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[6\].pup
timestamp 1667941163
transform 1 0 17360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[7\].pun
timestamp 1667941163
transform 1 0 16464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[7\].pup
timestamp 1667941163
transform 1 0 12880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[8\].pun
timestamp 1667941163
transform 1 0 14224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[8\].pup
timestamp 1667941163
transform 1 0 14224 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[9\].pun
timestamp 1667941163
transform 1 0 12208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[9\].pup
timestamp 1667941163
transform 1 0 8064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[10\].pun
timestamp 1667941163
transform -1 0 11760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[10\].pup
timestamp 1667941163
transform -1 0 6944 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[11\].pun
timestamp 1667941163
transform 1 0 9968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[11\].pup
timestamp 1667941163
transform 1 0 11312 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[12\].pun
timestamp 1667941163
transform 1 0 12096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[12\].pup
timestamp 1667941163
transform 1 0 13552 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[13\].pun
timestamp 1667941163
transform 1 0 16352 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[13\].pup
timestamp 1667941163
transform 1 0 11424 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[14\].pun
timestamp 1667941163
transform 1 0 10080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[14\].pup
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[15\].pun
timestamp 1667941163
transform 1 0 10192 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[15\].pup
timestamp 1667941163
transform -1 0 10864 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[16\].pun
timestamp 1667941163
transform 1 0 13552 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[16\].pup
timestamp 1667941163
transform 1 0 10864 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[17\].pun
timestamp 1667941163
transform 1 0 10752 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[17\].pup
timestamp 1667941163
transform 1 0 12208 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[18\].pun
timestamp 1667941163
transform -1 0 11088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[18\].pup
timestamp 1667941163
transform 1 0 14896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[19\].pun
timestamp 1667941163
transform 1 0 14896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_PU\[19\].pup
timestamp 1667941163
transform 1 0 7392 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[0\].ntrimn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2576 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[0\].ntrimp
timestamp 1667941163
transform -1 0 4480 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[0\].ptrimn
timestamp 1667941163
transform 1 0 2352 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[0\].ptrimp
timestamp 1667941163
transform 1 0 2352 0 -1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[1\].ntrimn
timestamp 1667941163
transform -1 0 8960 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[1\].ntrimp
timestamp 1667941163
transform -1 0 9072 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[1\].ptrimn
timestamp 1667941163
transform 1 0 7168 0 -1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[1\].ptrimp
timestamp 1667941163
transform 1 0 7168 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[2\].ntrimn
timestamp 1667941163
transform -1 0 13888 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[2\].ntrimp
timestamp 1667941163
transform -1 0 12992 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[2\].ptrimn
timestamp 1667941163
transform -1 0 12992 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[2\].ptrimp
timestamp 1667941163
transform 1 0 11984 0 -1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[3\].ntrimn
timestamp 1667941163
transform -1 0 16912 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[3\].ntrimp
timestamp 1667941163
transform -1 0 18256 0 1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[3\].ptrimn
timestamp 1667941163
transform -1 0 16240 0 -1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  gen_TRIM\[3\].ptrimp
timestamp 1667941163
transform -1 0 16128 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  nsijn
timestamp 1667941163
transform 1 0 1680 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  psijp
timestamp 1667941163
transform 1 0 1680 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  siginv
timestamp 1667941163
transform -1 0 4928 0 -1 7840
box -86 -86 534 870
<< labels >>
flabel metal3 s 0 2912 800 3024 0 FreeSans 448 0 0 0 enable
port 0 nsew signal input
flabel metal3 s 19200 8848 20000 8960 0 FreeSans 448 0 0 0 outn
port 1 nsew signal bidirectional
flabel metal3 s 19200 2912 20000 3024 0 FreeSans 448 0 0 0 outp
port 2 nsew signal bidirectional
flabel metal3 s 0 8848 800 8960 0 FreeSans 448 0 0 0 signal
port 3 nsew signal input
flabel metal2 s 2464 0 2576 800 0 FreeSans 448 90 0 0 trim_n[0]
port 4 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 trim_n[1]
port 5 nsew signal input
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 trim_n[2]
port 6 nsew signal input
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 trim_n[3]
port 7 nsew signal input
flabel metal2 s 2464 11200 2576 12000 0 FreeSans 448 90 0 0 trim_p[0]
port 8 nsew signal input
flabel metal2 s 7392 11200 7504 12000 0 FreeSans 448 90 0 0 trim_p[1]
port 9 nsew signal input
flabel metal2 s 12320 11200 12432 12000 0 FreeSans 448 90 0 0 trim_p[2]
port 10 nsew signal input
flabel metal2 s 17248 11200 17360 12000 0 FreeSans 448 90 0 0 trim_p[3]
port 11 nsew signal input
flabel metal4 s 3340 3076 3660 8684 0 FreeSans 1280 90 0 0 vdd
port 12 nsew power bidirectional
flabel metal4 s 7652 3076 7972 8684 0 FreeSans 1280 90 0 0 vdd
port 12 nsew power bidirectional
flabel metal4 s 11964 3076 12284 8684 0 FreeSans 1280 90 0 0 vdd
port 12 nsew power bidirectional
flabel metal4 s 16276 3076 16596 8684 0 FreeSans 1280 90 0 0 vdd
port 12 nsew power bidirectional
flabel metal4 s 5496 3076 5816 8684 0 FreeSans 1280 90 0 0 vss
port 13 nsew ground bidirectional
flabel metal4 s 9808 3076 10128 8684 0 FreeSans 1280 90 0 0 vss
port 13 nsew ground bidirectional
flabel metal4 s 14120 3076 14440 8684 0 FreeSans 1280 90 0 0 vss
port 13 nsew ground bidirectional
flabel metal4 s 18432 3076 18752 8684 0 FreeSans 1280 90 0 0 vss
port 13 nsew ground bidirectional
rlabel metal1 9968 8624 9968 8624 0 vdd
rlabel via1 10048 7840 10048 7840 0 vss
rlabel metal3 7896 6552 7896 6552 0 _00_
rlabel metal3 3248 8120 3248 8120 0 _01_
rlabel metal3 2576 6552 2576 6552 0 _02_
rlabel metal3 3024 6104 3024 6104 0 _03_
rlabel metal2 2184 7448 2184 7448 0 _04_
rlabel metal2 10024 4088 10024 4088 0 _05_
rlabel metal2 14448 4200 14448 4200 0 _06_
rlabel metal2 8120 4424 8120 4424 0 _07_
rlabel metal2 8344 5488 8344 5488 0 _08_
rlabel metal3 7000 5320 7000 5320 0 _09_
rlabel metal3 12936 4088 12936 4088 0 _10_
rlabel metal2 7000 5600 7000 5600 0 _11_
rlabel metal3 16800 5768 16800 5768 0 _12_
rlabel metal2 9016 5152 9016 5152 0 _13_
rlabel metal2 15176 5152 15176 5152 0 _14_
rlabel metal2 6328 6384 6328 6384 0 _15_
rlabel metal2 10696 4872 10696 4872 0 _16_
rlabel metal2 4984 5992 4984 5992 0 _17_
rlabel metal2 14392 3808 14392 3808 0 _18_
rlabel metal2 17752 4256 17752 4256 0 _19_
rlabel metal2 13664 3528 13664 3528 0 _20_
rlabel metal2 4312 4760 4312 4760 0 _21_
rlabel metal2 2184 3584 2184 3584 0 _22_
rlabel metal2 5992 4256 5992 4256 0 _23_
rlabel metal3 6104 3640 6104 3640 0 _24_
rlabel metal2 6776 3528 6776 3528 0 _25_
rlabel metal2 11144 3640 11144 3640 0 _26_
rlabel metal2 9912 3864 9912 3864 0 _27_
rlabel metal2 16184 5432 16184 5432 0 _28_
rlabel metal2 1848 4368 1848 4368 0 enable
rlabel metal2 3304 7896 3304 7896 0 outn
rlabel metal2 3360 7448 3360 7448 0 outp
rlabel metal2 2072 7112 2072 7112 0 signal
rlabel metal2 2744 6944 2744 6944 0 signal_n
rlabel metal2 2744 3472 2744 3472 0 trim_n[0]
rlabel metal2 7448 2142 7448 2142 0 trim_n[1]
rlabel metal2 12488 3528 12488 3528 0 trim_n[2]
rlabel metal2 16800 3528 16800 3528 0 trim_n[3]
rlabel metal2 2520 7840 2520 7840 0 trim_p[0]
rlabel metal2 7336 7840 7336 7840 0 trim_p[1]
rlabel metal2 12488 8232 12488 8232 0 trim_p[2]
rlabel metal3 16576 8232 16576 8232 0 trim_p[3]
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
