module captune_1p (cap,
    vdd,
    vss,
    tune);
 inout cap;
 input vdd;
 input vss;
 input [63:0] tune;

 wire \gen_cap[0].loose_end ;
 wire \gen_cap[10].loose_end ;
 wire \gen_cap[11].loose_end ;
 wire \gen_cap[12].loose_end ;
 wire \gen_cap[13].loose_end ;
 wire \gen_cap[14].loose_end ;
 wire \gen_cap[15].loose_end ;
 wire \gen_cap[16].loose_end ;
 wire \gen_cap[17].loose_end ;
 wire \gen_cap[18].loose_end ;
 wire \gen_cap[19].loose_end ;
 wire \gen_cap[1].loose_end ;
 wire \gen_cap[20].loose_end ;
 wire \gen_cap[21].loose_end ;
 wire \gen_cap[22].loose_end ;
 wire \gen_cap[23].loose_end ;
 wire \gen_cap[24].loose_end ;
 wire \gen_cap[25].loose_end ;
 wire \gen_cap[26].loose_end ;
 wire \gen_cap[27].loose_end ;
 wire \gen_cap[28].loose_end ;
 wire \gen_cap[29].loose_end ;
 wire \gen_cap[2].loose_end ;
 wire \gen_cap[30].loose_end ;
 wire \gen_cap[31].loose_end ;
 wire \gen_cap[32].loose_end ;
 wire \gen_cap[33].loose_end ;
 wire \gen_cap[34].loose_end ;
 wire \gen_cap[35].loose_end ;
 wire \gen_cap[36].loose_end ;
 wire \gen_cap[37].loose_end ;
 wire \gen_cap[38].loose_end ;
 wire \gen_cap[39].loose_end ;
 wire \gen_cap[3].loose_end ;
 wire \gen_cap[40].loose_end ;
 wire \gen_cap[41].loose_end ;
 wire \gen_cap[42].loose_end ;
 wire \gen_cap[43].loose_end ;
 wire \gen_cap[44].loose_end ;
 wire \gen_cap[45].loose_end ;
 wire \gen_cap[46].loose_end ;
 wire \gen_cap[47].loose_end ;
 wire \gen_cap[48].loose_end ;
 wire \gen_cap[49].loose_end ;
 wire \gen_cap[4].loose_end ;
 wire \gen_cap[50].loose_end ;
 wire \gen_cap[51].loose_end ;
 wire \gen_cap[52].loose_end ;
 wire \gen_cap[53].loose_end ;
 wire \gen_cap[54].loose_end ;
 wire \gen_cap[55].loose_end ;
 wire \gen_cap[56].loose_end ;
 wire \gen_cap[57].loose_end ;
 wire \gen_cap[58].loose_end ;
 wire \gen_cap[59].loose_end ;
 wire \gen_cap[5].loose_end ;
 wire \gen_cap[60].loose_end ;
 wire \gen_cap[61].loose_end ;
 wire \gen_cap[62].loose_end ;
 wire \gen_cap[63].loose_end ;
 wire \gen_cap[6].loose_end ;
 wire \gen_cap[7].loose_end ;
 wire \gen_cap[8].loose_end ;
 wire \gen_cap[9].loose_end ;

 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[0].u_cap  (.A1(tune[0]),
    .A2(tune[0]),
    .B(cap),
    .ZN(\gen_cap[0].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[10].u_cap  (.A1(tune[10]),
    .A2(tune[10]),
    .B(cap),
    .ZN(\gen_cap[10].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[11].u_cap  (.A1(tune[11]),
    .A2(tune[11]),
    .B(cap),
    .ZN(\gen_cap[11].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[12].u_cap  (.A1(tune[12]),
    .A2(tune[12]),
    .B(cap),
    .ZN(\gen_cap[12].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[13].u_cap  (.A1(tune[13]),
    .A2(tune[13]),
    .B(cap),
    .ZN(\gen_cap[13].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[14].u_cap  (.A1(tune[14]),
    .A2(tune[14]),
    .B(cap),
    .ZN(\gen_cap[14].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[15].u_cap  (.A1(tune[15]),
    .A2(tune[15]),
    .B(cap),
    .ZN(\gen_cap[15].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[16].u_cap  (.A1(tune[16]),
    .A2(tune[16]),
    .B(cap),
    .ZN(\gen_cap[16].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[17].u_cap  (.A1(tune[17]),
    .A2(tune[17]),
    .B(cap),
    .ZN(\gen_cap[17].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[18].u_cap  (.A1(tune[18]),
    .A2(tune[18]),
    .B(cap),
    .ZN(\gen_cap[18].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[19].u_cap  (.A1(tune[19]),
    .A2(tune[19]),
    .B(cap),
    .ZN(\gen_cap[19].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[1].u_cap  (.A1(tune[1]),
    .A2(tune[1]),
    .B(cap),
    .ZN(\gen_cap[1].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[20].u_cap  (.A1(tune[20]),
    .A2(tune[20]),
    .B(cap),
    .ZN(\gen_cap[20].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[21].u_cap  (.A1(tune[21]),
    .A2(tune[21]),
    .B(cap),
    .ZN(\gen_cap[21].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[22].u_cap  (.A1(tune[22]),
    .A2(tune[22]),
    .B(cap),
    .ZN(\gen_cap[22].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[23].u_cap  (.A1(tune[23]),
    .A2(tune[23]),
    .B(cap),
    .ZN(\gen_cap[23].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[24].u_cap  (.A1(tune[24]),
    .A2(tune[24]),
    .B(cap),
    .ZN(\gen_cap[24].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[25].u_cap  (.A1(tune[25]),
    .A2(tune[25]),
    .B(cap),
    .ZN(\gen_cap[25].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[26].u_cap  (.A1(tune[26]),
    .A2(tune[26]),
    .B(cap),
    .ZN(\gen_cap[26].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[27].u_cap  (.A1(tune[27]),
    .A2(tune[27]),
    .B(cap),
    .ZN(\gen_cap[27].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[28].u_cap  (.A1(tune[28]),
    .A2(tune[28]),
    .B(cap),
    .ZN(\gen_cap[28].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[29].u_cap  (.A1(tune[29]),
    .A2(tune[29]),
    .B(cap),
    .ZN(\gen_cap[29].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[2].u_cap  (.A1(tune[2]),
    .A2(tune[2]),
    .B(cap),
    .ZN(\gen_cap[2].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[30].u_cap  (.A1(tune[30]),
    .A2(tune[30]),
    .B(cap),
    .ZN(\gen_cap[30].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[31].u_cap  (.A1(tune[31]),
    .A2(tune[31]),
    .B(cap),
    .ZN(\gen_cap[31].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[32].u_cap  (.A1(tune[32]),
    .A2(tune[32]),
    .B(cap),
    .ZN(\gen_cap[32].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[33].u_cap  (.A1(tune[33]),
    .A2(tune[33]),
    .B(cap),
    .ZN(\gen_cap[33].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[34].u_cap  (.A1(tune[34]),
    .A2(tune[34]),
    .B(cap),
    .ZN(\gen_cap[34].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[35].u_cap  (.A1(tune[35]),
    .A2(tune[35]),
    .B(cap),
    .ZN(\gen_cap[35].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[36].u_cap  (.A1(tune[36]),
    .A2(tune[36]),
    .B(cap),
    .ZN(\gen_cap[36].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[37].u_cap  (.A1(tune[37]),
    .A2(tune[37]),
    .B(cap),
    .ZN(\gen_cap[37].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[38].u_cap  (.A1(tune[38]),
    .A2(tune[38]),
    .B(cap),
    .ZN(\gen_cap[38].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[39].u_cap  (.A1(tune[39]),
    .A2(tune[39]),
    .B(cap),
    .ZN(\gen_cap[39].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[3].u_cap  (.A1(tune[3]),
    .A2(tune[3]),
    .B(cap),
    .ZN(\gen_cap[3].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[40].u_cap  (.A1(tune[40]),
    .A2(tune[40]),
    .B(cap),
    .ZN(\gen_cap[40].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[41].u_cap  (.A1(tune[41]),
    .A2(tune[41]),
    .B(cap),
    .ZN(\gen_cap[41].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[42].u_cap  (.A1(tune[42]),
    .A2(tune[42]),
    .B(cap),
    .ZN(\gen_cap[42].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[43].u_cap  (.A1(tune[43]),
    .A2(tune[43]),
    .B(cap),
    .ZN(\gen_cap[43].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[44].u_cap  (.A1(tune[44]),
    .A2(tune[44]),
    .B(cap),
    .ZN(\gen_cap[44].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[45].u_cap  (.A1(tune[45]),
    .A2(tune[45]),
    .B(cap),
    .ZN(\gen_cap[45].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[46].u_cap  (.A1(tune[46]),
    .A2(tune[46]),
    .B(cap),
    .ZN(\gen_cap[46].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[47].u_cap  (.A1(tune[47]),
    .A2(tune[47]),
    .B(cap),
    .ZN(\gen_cap[47].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[48].u_cap  (.A1(tune[48]),
    .A2(tune[48]),
    .B(cap),
    .ZN(\gen_cap[48].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[49].u_cap  (.A1(tune[49]),
    .A2(tune[49]),
    .B(cap),
    .ZN(\gen_cap[49].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[4].u_cap  (.A1(tune[4]),
    .A2(tune[4]),
    .B(cap),
    .ZN(\gen_cap[4].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[50].u_cap  (.A1(tune[50]),
    .A2(tune[50]),
    .B(cap),
    .ZN(\gen_cap[50].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[51].u_cap  (.A1(tune[51]),
    .A2(tune[51]),
    .B(cap),
    .ZN(\gen_cap[51].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[52].u_cap  (.A1(tune[52]),
    .A2(tune[52]),
    .B(cap),
    .ZN(\gen_cap[52].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[53].u_cap  (.A1(tune[53]),
    .A2(tune[53]),
    .B(cap),
    .ZN(\gen_cap[53].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[54].u_cap  (.A1(tune[54]),
    .A2(tune[54]),
    .B(cap),
    .ZN(\gen_cap[54].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[55].u_cap  (.A1(tune[55]),
    .A2(tune[55]),
    .B(cap),
    .ZN(\gen_cap[55].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[56].u_cap  (.A1(tune[56]),
    .A2(tune[56]),
    .B(cap),
    .ZN(\gen_cap[56].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[57].u_cap  (.A1(tune[57]),
    .A2(tune[57]),
    .B(cap),
    .ZN(\gen_cap[57].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[58].u_cap  (.A1(tune[58]),
    .A2(tune[58]),
    .B(cap),
    .ZN(\gen_cap[58].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[59].u_cap  (.A1(tune[59]),
    .A2(tune[59]),
    .B(cap),
    .ZN(\gen_cap[59].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[5].u_cap  (.A1(tune[5]),
    .A2(tune[5]),
    .B(cap),
    .ZN(\gen_cap[5].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[60].u_cap  (.A1(tune[60]),
    .A2(tune[60]),
    .B(cap),
    .ZN(\gen_cap[60].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[61].u_cap  (.A1(tune[61]),
    .A2(tune[61]),
    .B(cap),
    .ZN(\gen_cap[61].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[62].u_cap  (.A1(tune[62]),
    .A2(tune[62]),
    .B(cap),
    .ZN(\gen_cap[62].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[63].u_cap  (.A1(tune[63]),
    .A2(tune[63]),
    .B(cap),
    .ZN(\gen_cap[63].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[6].u_cap  (.A1(tune[6]),
    .A2(tune[6]),
    .B(cap),
    .ZN(\gen_cap[6].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[7].u_cap  (.A1(tune[7]),
    .A2(tune[7]),
    .B(cap),
    .ZN(\gen_cap[7].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[8].u_cap  (.A1(tune[8]),
    .A2(tune[8]),
    .B(cap),
    .ZN(\gen_cap[8].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_cap[9].u_cap  (.A1(tune[9]),
    .A2(tune[9]),
    .B(cap),
    .ZN(\gen_cap[9].loose_end ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_151 (.VDD(vdd),
    .VSS(vss));
endmodule
