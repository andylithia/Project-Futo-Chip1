VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caparray_s1
  CLASS BLOCK ;
  FOREIGN caparray_s1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 300.000 ;
  PIN cap_series_gygyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 296.000 186.480 300.000 ;
    END
  END cap_series_gygyn
  PIN cap_series_gygyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 296.000 161.840 300.000 ;
    END
  END cap_series_gygyp
  PIN cap_series_gyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 296.000 137.200 300.000 ;
    END
  END cap_series_gyn
  PIN cap_series_gyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 296.000 112.560 300.000 ;
    END
  END cap_series_gyp
  PIN cap_shunt_gyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 296.000 87.920 300.000 ;
    END
  END cap_shunt_gyn
  PIN cap_shunt_gyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 296.000 63.280 300.000 ;
    END
  END cap_shunt_gyp
  PIN cap_shunt_n
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 296.000 38.640 300.000 ;
    END
  END cap_shunt_n
  PIN cap_shunt_p
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 296.000 14.000 300.000 ;
    END
  END cap_shunt_p
  PIN tune_series_gy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END tune_series_gy[0]
  PIN tune_series_gy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 0.000 50.400 4.000 ;
    END
  END tune_series_gy[1]
  PIN tune_series_gy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END tune_series_gy[2]
  PIN tune_series_gy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.920 0.000 116.480 4.000 ;
    END
  END tune_series_gy[3]
  PIN tune_series_gy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END tune_series_gy[4]
  PIN tune_series_gy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.000 0.000 182.560 4.000 ;
    END
  END tune_series_gy[5]
  PIN tune_series_gygy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 11.760 200.000 12.320 ;
    END
  END tune_series_gygy[0]
  PIN tune_series_gygy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 34.720 200.000 35.280 ;
    END
  END tune_series_gygy[1]
  PIN tune_series_gygy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 57.680 200.000 58.240 ;
    END
  END tune_series_gygy[2]
  PIN tune_series_gygy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 80.640 200.000 81.200 ;
    END
  END tune_series_gygy[3]
  PIN tune_series_gygy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 103.600 200.000 104.160 ;
    END
  END tune_series_gygy[4]
  PIN tune_series_gygy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 126.560 200.000 127.120 ;
    END
  END tune_series_gygy[5]
  PIN tune_shunt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END tune_shunt[0]
  PIN tune_shunt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END tune_shunt[1]
  PIN tune_shunt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END tune_shunt[2]
  PIN tune_shunt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END tune_shunt[3]
  PIN tune_shunt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END tune_shunt[4]
  PIN tune_shunt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END tune_shunt[5]
  PIN tune_shunt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END tune_shunt[6]
  PIN tune_shunt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END tune_shunt[7]
  PIN tune_shunt_gy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 149.520 200.000 150.080 ;
    END
  END tune_shunt_gy[0]
  PIN tune_shunt_gy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 172.480 200.000 173.040 ;
    END
  END tune_shunt_gy[1]
  PIN tune_shunt_gy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 195.440 200.000 196.000 ;
    END
  END tune_shunt_gy[2]
  PIN tune_shunt_gy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 218.400 200.000 218.960 ;
    END
  END tune_shunt_gy[3]
  PIN tune_shunt_gy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 241.360 200.000 241.920 ;
    END
  END tune_shunt_gy[4]
  PIN tune_shunt_gy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 264.320 200.000 264.880 ;
    END
  END tune_shunt_gy[5]
  PIN tune_shunt_gy[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 287.280 200.000 287.840 ;
    END
  END tune_shunt_gy[6]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 193.200 282.540 ;
      LAYER Metal2 ;
        RECT 9.100 295.700 13.140 296.000 ;
        RECT 14.300 295.700 37.780 296.000 ;
        RECT 38.940 295.700 62.420 296.000 ;
        RECT 63.580 295.700 87.060 296.000 ;
        RECT 88.220 295.700 111.700 296.000 ;
        RECT 112.860 295.700 136.340 296.000 ;
        RECT 137.500 295.700 160.980 296.000 ;
        RECT 162.140 295.700 185.620 296.000 ;
        RECT 186.780 295.700 190.820 296.000 ;
        RECT 9.100 4.300 190.820 295.700 ;
        RECT 9.100 3.500 16.500 4.300 ;
        RECT 17.660 3.500 49.540 4.300 ;
        RECT 50.700 3.500 82.580 4.300 ;
        RECT 83.740 3.500 115.620 4.300 ;
        RECT 116.780 3.500 148.660 4.300 ;
        RECT 149.820 3.500 181.700 4.300 ;
        RECT 182.860 3.500 190.820 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 286.980 195.700 287.700 ;
        RECT 4.000 279.740 196.000 286.980 ;
        RECT 4.300 278.580 196.000 279.740 ;
        RECT 4.000 265.180 196.000 278.580 ;
        RECT 4.000 264.020 195.700 265.180 ;
        RECT 4.000 242.780 196.000 264.020 ;
        RECT 4.300 242.220 196.000 242.780 ;
        RECT 4.300 241.620 195.700 242.220 ;
        RECT 4.000 241.060 195.700 241.620 ;
        RECT 4.000 219.260 196.000 241.060 ;
        RECT 4.000 218.100 195.700 219.260 ;
        RECT 4.000 205.820 196.000 218.100 ;
        RECT 4.300 204.660 196.000 205.820 ;
        RECT 4.000 196.300 196.000 204.660 ;
        RECT 4.000 195.140 195.700 196.300 ;
        RECT 4.000 173.340 196.000 195.140 ;
        RECT 4.000 172.180 195.700 173.340 ;
        RECT 4.000 168.860 196.000 172.180 ;
        RECT 4.300 167.700 196.000 168.860 ;
        RECT 4.000 150.380 196.000 167.700 ;
        RECT 4.000 149.220 195.700 150.380 ;
        RECT 4.000 131.900 196.000 149.220 ;
        RECT 4.300 130.740 196.000 131.900 ;
        RECT 4.000 127.420 196.000 130.740 ;
        RECT 4.000 126.260 195.700 127.420 ;
        RECT 4.000 104.460 196.000 126.260 ;
        RECT 4.000 103.300 195.700 104.460 ;
        RECT 4.000 94.940 196.000 103.300 ;
        RECT 4.300 93.780 196.000 94.940 ;
        RECT 4.000 81.500 196.000 93.780 ;
        RECT 4.000 80.340 195.700 81.500 ;
        RECT 4.000 58.540 196.000 80.340 ;
        RECT 4.000 57.980 195.700 58.540 ;
        RECT 4.300 57.380 195.700 57.980 ;
        RECT 4.300 56.820 196.000 57.380 ;
        RECT 4.000 35.580 196.000 56.820 ;
        RECT 4.000 34.420 195.700 35.580 ;
        RECT 4.000 21.020 196.000 34.420 ;
        RECT 4.300 19.860 196.000 21.020 ;
        RECT 4.000 12.620 196.000 19.860 ;
        RECT 4.000 11.900 195.700 12.620 ;
      LAYER Metal4 ;
        RECT 178.220 33.130 178.500 58.150 ;
  END
END caparray_s1
END LIBRARY

