// This is the unpowered netlist.
module filterstage (nbusin_nshunt,
    nbusout,
    nseries_gy,
    nseries_gygy,
    nshunt_gy,
    pbusin_pshunt,
    pbusout,
    pseries_gy,
    pseries_gygy,
    pshunt_gy);
 inout nbusin_nshunt;
 inout nbusout;
 inout nseries_gy;
 inout nseries_gygy;
 inout nshunt_gy;
 inout pbusin_pshunt;
 inout pbusout;
 inout pseries_gy;
 inout pseries_gygy;
 inout pshunt_gy;


 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[0].fbn  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[0].fbp  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[1].fbn  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[1].fbp  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[2].fbn  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[2].fbp  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[3].fbn  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_FB[3].fbp  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[0].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[0].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[1].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[1].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[2].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[2].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[3].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[3].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[4].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[4].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[5].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[5].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[6].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[6].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[7].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[7].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[8].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[8].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[9].thrun  (.I(pbusout),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_T[9].thrup  (.I(pbusin_pshunt),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[0].crossn  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[0].crossp  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[1].crossn  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[1].crossp  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[2].crossn  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[2].crossp  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[3].crossn  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[3].crossp  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[4].crossn  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f1.gen_X[4].crossp  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[0].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[0].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[1].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[1].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[2].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[2].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[3].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_FB[3].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[0].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[0].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[1].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[1].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[2].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[2].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[3].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[3].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[4].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[4].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[5].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[5].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[6].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[6].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[7].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[7].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[8].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[8].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[9].thrun  (.I(nbusout),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_T[9].thrup  (.I(nbusin_nshunt),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[0].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[0].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[1].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[1].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[2].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[2].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[3].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[3].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[4].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_f2.gen_X[4].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[0].fbn  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[0].fbp  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[1].fbn  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[1].fbp  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[2].fbn  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[2].fbp  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[3].fbn  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_FB[3].fbp  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[0].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[0].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[1].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[1].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[2].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[2].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[3].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[3].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[4].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[4].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[5].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[5].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[6].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[6].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[7].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[7].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[8].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[8].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[9].thrun  (.I(pseries_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_T[9].thrup  (.I(nseries_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[0].crossn  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[0].crossp  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[1].crossn  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[1].crossp  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[2].crossn  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[2].crossp  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[3].crossn  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[3].crossp  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[4].crossn  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r1.gen_X[4].crossp  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[0].fbn  (.I(pbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[0].fbp  (.I(nbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[1].fbn  (.I(pbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[1].fbp  (.I(nbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[2].fbn  (.I(pbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[2].fbp  (.I(nbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[3].fbn  (.I(pbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_FB[3].fbp  (.I(nbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[0].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[0].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[1].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[1].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[2].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[2].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[3].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[3].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[4].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[4].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[5].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[5].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[6].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[6].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[7].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[7].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[8].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[8].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[9].thrun  (.I(nseries_gy),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_T[9].thrup  (.I(pseries_gy),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[0].crossn  (.I(nbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[0].crossp  (.I(pbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[1].crossn  (.I(nbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[1].crossp  (.I(pbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[2].crossn  (.I(nbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[2].crossp  (.I(pbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[3].crossn  (.I(nbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[3].crossp  (.I(pbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[4].crossn  (.I(nbusout),
    .ZN(pbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_series_r2.gen_X[4].crossp  (.I(pbusout),
    .ZN(nbusout));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[0].fbn  (.I(nseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[0].fbp  (.I(pseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[1].fbn  (.I(nseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[1].fbp  (.I(pseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[2].fbn  (.I(nseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[2].fbp  (.I(pseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[3].fbn  (.I(nseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_FB[3].fbp  (.I(pseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[0].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[0].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[1].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[1].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[2].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[2].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[3].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[3].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[4].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[4].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[5].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[5].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[6].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[6].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[7].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[7].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[8].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[8].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[9].thrun  (.I(pseries_gy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_T[9].thrup  (.I(nseries_gy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[0].crossn  (.I(pseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[0].crossp  (.I(nseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[1].crossn  (.I(pseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[1].crossp  (.I(nseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[2].crossn  (.I(pseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[2].crossp  (.I(nseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[3].crossn  (.I(pseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[3].crossp  (.I(nseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[4].crossn  (.I(pseries_gygy),
    .ZN(nseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_f.gen_X[4].crossp  (.I(nseries_gygy),
    .ZN(pseries_gygy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[0].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[0].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[1].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[1].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[2].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[2].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[3].fbn  (.I(nseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_FB[3].fbp  (.I(pseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[0].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[0].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[1].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[1].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[2].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[2].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[3].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[3].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[4].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[4].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[5].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[5].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[6].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[6].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[7].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[7].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[8].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[8].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[9].thrun  (.I(nseries_gygy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_T[9].thrup  (.I(pseries_gygy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[0].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[0].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[1].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[1].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[2].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[2].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[3].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[3].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[4].crossn  (.I(pseries_gy),
    .ZN(nseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_seriesgy.u_nauta_r.gen_X[4].crossp  (.I(nseries_gy),
    .ZN(pseries_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[0].fbn  (.I(nshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[0].fbp  (.I(pshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[1].fbn  (.I(nshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[1].fbp  (.I(pshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[2].fbn  (.I(nshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[2].fbp  (.I(pshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[3].fbn  (.I(nshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_FB[3].fbp  (.I(pshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[0].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[0].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[1].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[1].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[2].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[2].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[3].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[3].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[4].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[4].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[5].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[5].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[6].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[6].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[7].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[7].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[8].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[8].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[9].thrun  (.I(pbusin_pshunt),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_T[9].thrup  (.I(nbusin_nshunt),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[0].crossn  (.I(pshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[0].crossp  (.I(nshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[1].crossn  (.I(pshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[1].crossp  (.I(nshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[2].crossn  (.I(pshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[2].crossp  (.I(nshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[3].crossn  (.I(pshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[3].crossp  (.I(nshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[4].crossn  (.I(pshunt_gy),
    .ZN(nshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_f.gen_X[4].crossp  (.I(nshunt_gy),
    .ZN(pshunt_gy));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[0].fbn  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[0].fbp  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[1].fbn  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[1].fbp  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[2].fbn  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[2].fbp  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[3].fbn  (.I(nbusin_nshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_FB[3].fbp  (.I(pbusin_pshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[0].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[0].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[1].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[1].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[2].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[2].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[3].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[3].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[4].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[4].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[5].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[5].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[6].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[6].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[7].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[7].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[8].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[8].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[9].thrun  (.I(nshunt_gy),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_T[9].thrup  (.I(pshunt_gy),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[0].crossn  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[0].crossp  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[1].crossn  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[1].crossp  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[2].crossn  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[2].crossp  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[3].crossn  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[3].crossp  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[4].crossn  (.I(pbusin_pshunt),
    .ZN(nbusin_nshunt));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_shuntgy.u_nauta_r.gen_X[4].crossp  (.I(nbusin_nshunt),
    .ZN(pbusin_pshunt));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_187 ();
endmodule

