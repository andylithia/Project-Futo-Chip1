* NGSPICE file created from injector_flat.ext - technology: gf180mcuC

.subckt injector_flat enable outn outp signal trim_n[0] trim_n[1] trim_n[2] trim_n[3]
+ trim_p[0] trim_p[1] trim_p[2] trim_p[3] vss vdd
X0 _13_ a_8301_4728# vdd vdd pmos_6p0 w=1.22u l=0.5u
X1 vdd a_9644_7080# a_9556_7124# vdd pmos_6p0 w=1.22u l=1u
X2 a_3055_3728# a_2612_3229# vdd vdd pmos_6p0 w=0.62u l=0.5u
X3 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X4 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X5 vdd trim_p[0] a_2388_7933# vdd pmos_6p0 w=0.62u l=0.5u
X6 _09_ a_6285_4728# vdd vdd pmos_6p0 w=1.22u l=0.5u
X7 vdd a_3036_5079# a_2948_5176# vdd pmos_6p0 w=1.22u l=1u
X8 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X9 a_5948_7080# a_5860_7124# vss vss nmos_6p0 w=0.82u l=1u
X10 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X11 vdd _20_ outp vdd pmos_6p0 w=1.22u l=0.5u
X12 vss trim_p[1] a_7204_7933# vss nmos_6p0 w=0.36u l=0.6u
X13 a_15496_8308# trim_p[3] vdd vdd pmos_6p0 w=0.62u l=0.5u
X14 outp _18_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X15 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X16 a_3820_5512# a_3732_5556# vss vss nmos_6p0 w=0.82u l=1u
X17 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X18 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X19 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X20 vdd a_5052_7080# a_4964_7124# vdd pmos_6p0 w=1.22u l=1u
X21 a_8573_7889# _00_ vss vss nmos_6p0 w=0.36u l=0.6u
X22 a_14703_8432# a_15496_8308# a_14723_7933# vdd pmos_6p0 w=0.62u l=0.5u
X23 a_3932_6647# a_3844_6744# vss vss nmos_6p0 w=0.82u l=1u
X24 a_7636_7675# a_7204_7156# vss vss nmos_6p0 w=0.36u l=0.6u
X25 _06_ a_14237_3944# vdd vdd pmos_6p0 w=1.22u l=0.5u
X26 vdd a_3484_5079# a_3396_5176# vdd pmos_6p0 w=1.22u l=1u
X27 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X28 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X29 vdd _15_ outn vdd pmos_6p0 w=1.22u l=0.5u
X30 a_9869_3160# a_9869_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X31 a_16280_3604# trim_n[3] vss vss nmos_6p0 w=0.36u l=0.6u
X32 a_6621_3160# a_6621_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X33 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X34 vdd _26_ a_11124_3229# vdd pmos_6p0 w=0.62u l=0.5u
X35 vdd a_2140_3944# a_2052_3988# vdd pmos_6p0 w=1.22u l=1u
X36 vdd a_3981_4417# a_3004_4020# vdd pmos_6p0 w=0.62u l=0.5u
X37 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X38 vss signal_n a_2161_6296# vss nmos_6p0 w=0.36u l=0.6u
X39 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X40 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X41 outp a_14703_8432# vdd vdd pmos_6p0 w=1.095u l=0.5u
X42 a_16280_3604# trim_n[3] vdd vdd pmos_6p0 w=0.62u l=0.5u
X43 outn a_7555_4539# vss vss nmos_6p0 w=0.82u l=0.6u
X44 a_16700_3944# a_16612_3988# vss vss nmos_6p0 w=0.82u l=1u
X45 vdd a_2140_5079# a_2052_5176# vdd pmos_6p0 w=1.22u l=1u
X46 vss a_3757_7889# a_2820_7933# vss nmos_6p0 w=0.36u l=0.6u
X47 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X48 vdd a_8573_7553# a_7596_7156# vdd pmos_6p0 w=0.62u l=0.5u
X49 a_16851_4797# a_16388_4797# vss vss nmos_6p0 w=0.36u l=0.6u
X50 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X51 a_15487_3728# a_16280_3604# a_15507_3229# vdd pmos_6p0 w=0.62u l=0.5u
X52 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X53 vdd a_3004_4020# outn vdd pmos_6p0 w=1.095u l=0.5u
X54 a_12463_3988# a_12020_4539# vdd vdd pmos_6p0 w=0.62u l=0.5u
X55 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X56 vdd a_4828_6647# a_4740_6744# vdd pmos_6p0 w=1.22u l=1u
X57 vss _22_ a_2612_3229# vss nmos_6p0 w=0.36u l=0.6u
X58 vss signal a_1924_6040# vss nmos_6p0 w=0.365u l=0.6u
X59 vss _07_ outn vss nmos_6p0 w=0.82u l=0.6u
X60 a_12360_8308# trim_p[2] vss vss nmos_6p0 w=0.36u l=0.6u
X61 _10_ a_10093_3944# vdd vdd pmos_6p0 w=1.22u l=0.5u
X62 vdd a_6060_8215# a_5972_8312# vdd pmos_6p0 w=1.22u l=1u
X63 _03_ a_1716_6040# vdd vdd pmos_6p0 w=1.215u l=0.5u
X64 a_12780_5079# a_12692_5176# vss vss nmos_6p0 w=0.82u l=1u
X65 vdd a_17932_8215# a_17844_8312# vdd pmos_6p0 w=1.22u l=1u
X66 _03_ a_1716_6040# vss vss nmos_6p0 w=0.815u l=0.6u
X67 vdd a_8573_7889# a_7596_8400# vdd pmos_6p0 w=0.62u l=0.5u
X68 a_7667_3229# trim_n[1] a_7647_3728# vss nmos_6p0 w=0.36u l=0.6u
X69 a_10541_3160# a_10541_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X70 a_4268_5512# a_4180_5556# vss vss nmos_6p0 w=0.82u l=1u
X71 outn _09_ vss vss nmos_6p0 w=0.82u l=0.6u
X72 a_12483_4539# a_12020_4539# vss vss nmos_6p0 w=0.36u l=0.6u
X73 a_7667_3229# a_7204_3229# vss vss nmos_6p0 w=0.36u l=0.6u
X74 vss _25_ a_12020_4539# vss nmos_6p0 w=0.36u l=0.6u
X75 a_3004_4020# trim_n[0] vdd vdd pmos_6p0 w=0.62u l=0.5u
X76 a_1692_6647# a_1604_6744# vss vss nmos_6p0 w=0.82u l=1u
X77 vss trim_p[2] a_12020_7156# vss nmos_6p0 w=0.36u l=0.6u
X78 vss a_16280_3604# a_15507_3229# vss nmos_6p0 w=0.36u l=0.6u
X79 a_3055_3728# a_3848_3604# a_3075_3229# vdd pmos_6p0 w=0.62u l=0.5u
X80 _28_ a_5501_5512# vdd vdd pmos_6p0 w=1.22u l=0.5u
X81 vss _00_ outn vss nmos_6p0 w=0.82u l=0.6u
X82 a_8189_5512# a_8189_5512# vss vss nmos_6p0 w=0.82u l=0.6u
X83 a_3757_7889# _00_ vss vss nmos_6p0 w=0.36u l=0.6u
X84 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X85 a_8573_7553# _00_ vdd vdd pmos_6p0 w=0.62u l=0.5u
X86 a_2161_6296# _00_ vss vss nmos_6p0 w=0.36u l=0.6u
X87 outn a_14835_7675# vss vss nmos_6p0 w=0.82u l=0.6u
X88 a_6844_7080# a_6756_7124# vss vss nmos_6p0 w=0.82u l=1u
X89 vdd a_9644_3944# a_9556_3988# vdd pmos_6p0 w=1.22u l=1u
X90 vdd a_4716_5512# a_4628_5556# vdd pmos_6p0 w=1.22u l=1u
X91 a_5612_6647# a_5524_6744# vss vss nmos_6p0 w=0.82u l=1u
X92 a_14815_7124# a_15608_7112# a_14835_7675# vdd pmos_6p0 w=0.62u l=0.5u
X93 a_7596_7156# trim_p[1] a_7636_7675# vss nmos_6p0 w=0.36u l=0.6u
X94 vss _00_ outn vss nmos_6p0 w=0.82u l=0.6u
X95 vdd a_3932_6647# a_3844_6744# vdd pmos_6p0 w=1.22u l=1u
X96 vss a_2820_7675# outp vss nmos_6p0 w=0.82u l=0.6u
X97 vdd trim_n[1] a_7535_3988# vdd pmos_6p0 w=0.62u l=0.5u
X98 vdd signal a_1716_6040# vdd pmos_6p0 w=0.6u l=0.5u
X99 a_12412_7156# trim_p[2] a_12452_7675# vss nmos_6p0 w=0.36u l=0.6u
X100 _05_ a_9869_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X101 _25_ a_6621_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X102 a_16831_5296# a_17624_5172# a_16851_4797# vdd pmos_6p0 w=0.62u l=0.5u
X103 vdd a_7596_7156# outn vdd pmos_6p0 w=1.095u l=0.5u
X104 vss a_17699_6040# a_17699_6040# vss nmos_6p0 w=0.82u l=0.6u
X105 vdd trim_n[1] a_7647_3728# vdd pmos_6p0 w=0.62u l=0.5u
X106 a_2780_7156# trim_p[0] vdd vdd pmos_6p0 w=0.62u l=0.5u
X107 vdd _00_ outp vdd pmos_6p0 w=1.22u l=0.5u
X108 vdd a_14012_7080# a_13924_7124# vdd pmos_6p0 w=1.22u l=1u
X109 a_5500_7080# a_5412_7124# vss vss nmos_6p0 w=0.82u l=1u
X110 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X111 a_8573_7889# _00_ vdd vdd pmos_6p0 w=0.62u l=0.5u
X112 vdd a_3296_6296# _02_ vdd pmos_6p0 w=1.22u l=0.5u
X113 a_3372_5512# a_3284_5556# vss vss nmos_6p0 w=0.82u l=1u
X114 vss a_12360_8308# a_11587_7933# vss nmos_6p0 w=0.36u l=0.6u
X115 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X116 a_2820_7933# a_2388_7933# a_2780_8400# vdd pmos_6p0 w=0.62u l=0.5u
X117 a_5612_8215# a_5524_8312# vss vss nmos_6p0 w=0.82u l=1u
X118 a_2161_6296# signal_n a_2553_6875# vdd pmos_6p0 w=0.565u l=0.5u
X119 a_11587_3229# a_11124_3229# vss vss nmos_6p0 w=0.36u l=0.6u
X120 vdd trim_n[0] a_3055_3728# vdd pmos_6p0 w=0.62u l=0.5u
X121 vdd signal signal_n vdd pmos_6p0 w=1.22u l=0.5u
X122 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X123 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X124 a_15507_3229# trim_n[3] a_15487_3728# vss nmos_6p0 w=0.36u l=0.6u
X125 vss a_2820_7933# outn vss nmos_6p0 w=0.82u l=0.6u
X126 outp _10_ vss vss nmos_6p0 w=0.82u l=0.6u
X127 vdd a_3820_5512# a_3732_5556# vdd pmos_6p0 w=1.22u l=1u
X128 outp _06_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X129 vdd a_7596_8400# outp vdd pmos_6p0 w=1.095u l=0.5u
X130 a_14237_3160# a_14237_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X131 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X132 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X133 a_3296_6296# _03_ vss vss nmos_6p0 w=0.36u l=0.6u
X134 a_16831_5296# a_16388_4797# vdd vdd pmos_6p0 w=0.62u l=0.5u
X135 outn _05_ vss vss nmos_6p0 w=0.82u l=0.6u
X136 vdd a_6947_4772# _11_ vdd pmos_6p0 w=1.22u l=0.5u
X137 outp _12_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X138 outn a_12483_4539# vss vss nmos_6p0 w=0.82u l=0.6u
X139 _16_ a_10541_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X140 a_4829_4728# a_4829_4728# vss vss nmos_6p0 w=0.82u l=0.6u
X141 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X142 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X143 a_7647_3728# a_7204_3229# vdd vdd pmos_6p0 w=0.62u l=0.5u
X144 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X145 a_12452_7675# a_12020_7156# vss vss nmos_6p0 w=0.36u l=0.6u
X146 vdd trim_n[2] a_11567_3728# vdd pmos_6p0 w=0.62u l=0.5u
X147 vdd a_1692_6647# a_1604_6744# vdd pmos_6p0 w=1.22u l=1u
X148 vdd _00_ outp vdd pmos_6p0 w=1.22u l=0.5u
X149 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X150 a_3757_7553# _00_ vdd vdd pmos_6p0 w=0.62u l=0.5u
X151 vdd _07_ outn vdd pmos_6p0 w=1.22u l=0.5u
X152 a_12668_6647# a_12580_6744# vss vss nmos_6p0 w=0.82u l=1u
X153 vdd a_12780_5079# a_12692_5176# vdd pmos_6p0 w=1.22u l=1u
X154 vdd _27_ a_15044_3229# vdd pmos_6p0 w=0.62u l=0.5u
X155 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X156 vdd a_16700_3944# a_16612_3988# vdd pmos_6p0 w=1.22u l=1u
X157 vdd a_5612_6647# a_5524_6744# vdd pmos_6p0 w=1.22u l=1u
X158 a_11587_7933# trim_p[2] a_11567_8432# vss nmos_6p0 w=0.36u l=0.6u
X159 a_9644_5512# a_9556_5556# vss vss nmos_6p0 w=0.82u l=1u
X160 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X161 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X162 a_5837_3944# a_5837_3944# vss vss nmos_6p0 w=0.82u l=0.6u
X163 vss _28_ a_16388_4797# vss nmos_6p0 w=0.36u l=0.6u
X164 a_2780_8400# trim_p[0] a_2820_7933# vss nmos_6p0 w=0.36u l=0.6u
X165 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X166 vdd a_6835_6340# _15_ vdd pmos_6p0 w=1.22u l=0.5u
X167 a_6509_3944# a_6509_3944# vss vss nmos_6p0 w=0.82u l=0.6u
X168 a_3757_7889# _00_ vdd vdd pmos_6p0 w=0.62u l=0.5u
X169 a_1716_6040# enable vdd vdd pmos_6p0 w=0.6u l=0.5u
X170 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X171 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X172 outp _08_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X173 a_16365_5512# a_16365_5512# vss vss nmos_6p0 w=0.82u l=0.6u
X174 a_14723_7933# trim_p[3] a_14703_8432# vss nmos_6p0 w=0.36u l=0.6u
X175 a_6396_7080# a_6308_7124# vss vss nmos_6p0 w=0.82u l=1u
X176 a_11567_3728# a_11124_3229# vdd vdd pmos_6p0 w=0.62u l=0.5u
X177 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X178 a_4640_7864# _04_ vss vss nmos_6p0 w=0.36u l=0.6u
X179 vdd a_4268_5512# a_4180_5556# vdd pmos_6p0 w=1.22u l=1u
X180 a_9644_7080# a_9556_7124# vss vss nmos_6p0 w=0.82u l=1u
X181 vss a_17475_3204# a_17475_3204# vss nmos_6p0 w=0.82u l=0.6u
X182 vss trim_p[1] a_7204_7156# vss nmos_6p0 w=0.36u l=0.6u
X183 a_3981_4417# _21_ vdd vdd pmos_6p0 w=0.62u l=0.5u
X184 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X185 vss a_7636_7675# outn vss nmos_6p0 w=0.82u l=0.6u
X186 vdd trim_n[2] a_12463_3988# vdd pmos_6p0 w=0.62u l=0.5u
X187 outn _17_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X188 outn _17_ vss vss nmos_6p0 w=0.82u l=0.6u
X189 a_8573_7553# _00_ vss vss nmos_6p0 w=0.36u l=0.6u
X190 a_7596_7156# trim_p[1] vdd vdd pmos_6p0 w=0.62u l=0.5u
X191 vdd _00_ outp vdd pmos_6p0 w=1.22u l=0.5u
X192 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X193 vdd _00_ outn vdd pmos_6p0 w=1.22u l=0.5u
X194 _08_ a_8189_5512# vdd vdd pmos_6p0 w=1.22u l=0.5u
X195 a_4380_6647# a_4292_6744# vss vss nmos_6p0 w=0.82u l=1u
X196 _18_ a_14237_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X197 outp _16_ vss vss nmos_6p0 w=0.82u l=0.6u
X198 a_12412_7156# trim_p[2] vdd vdd pmos_6p0 w=0.62u l=0.5u
X199 a_5052_7080# a_4964_7124# vss vss nmos_6p0 w=0.82u l=1u
X200 a_15496_8308# trim_p[3] vss vss nmos_6p0 w=0.36u l=0.6u
X201 vss a_2161_6296# _04_ vss nmos_6p0 w=0.82u l=0.6u
X202 a_16812_5512# a_16724_5556# vss vss nmos_6p0 w=0.82u l=1u
X203 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X204 a_13389_7553# _00_ vdd vdd pmos_6p0 w=0.62u l=0.5u
X205 vdd _00_ outn vdd pmos_6p0 w=1.22u l=0.5u
X206 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X207 a_3981_4417# _21_ vss vss nmos_6p0 w=0.36u l=0.6u
X208 a_7636_7933# a_7204_7933# a_7596_8400# vdd pmos_6p0 w=0.62u l=0.5u
X209 a_7535_3988# a_8328_3976# a_7555_4539# vdd pmos_6p0 w=0.62u l=0.5u
X210 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X211 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X212 vss _23_ a_7092_4539# vss nmos_6p0 w=0.36u l=0.6u
X213 vdd trim_p[1] a_7204_7933# vdd pmos_6p0 w=0.62u l=0.5u
X214 vdd _00_ a_11124_7933# vdd pmos_6p0 w=0.62u l=0.5u
X215 a_8328_3976# trim_n[1] vss vss nmos_6p0 w=0.36u l=0.6u
X216 vss a_3757_7553# a_2820_7675# vss nmos_6p0 w=0.36u l=0.6u
X217 a_2820_7933# a_2388_7933# vss vss nmos_6p0 w=0.36u l=0.6u
X218 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X219 vdd trim_p[0] a_2388_7156# vdd pmos_6p0 w=0.62u l=0.5u
X220 vdd trim_p[2] a_11567_8432# vdd pmos_6p0 w=0.62u l=0.5u
X221 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X222 vss a_7636_7933# outp vss nmos_6p0 w=0.82u l=0.6u
X223 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X224 vdd a_3372_5512# a_3284_5556# vdd pmos_6p0 w=1.22u l=1u
X225 outp a_7647_3728# vdd vdd pmos_6p0 w=1.095u l=0.5u
X226 vss _11_ outn vss nmos_6p0 w=0.82u l=0.6u
X227 vdd a_12668_6647# a_12580_6744# vdd pmos_6p0 w=1.22u l=1u
X228 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X229 vss _00_ a_14372_7675# vss nmos_6p0 w=0.36u l=0.6u
X230 _17_ a_4829_4728# vdd vdd pmos_6p0 w=1.22u l=0.5u
X231 _00_ enable vdd vdd pmos_6p0 w=1.22u l=0.5u
X232 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X233 vdd a_15683_4772# _14_ vdd pmos_6p0 w=1.22u l=0.5u
X234 vss _26_ a_11124_3229# vss nmos_6p0 w=0.36u l=0.6u
X235 outp a_7667_3229# vss vss nmos_6p0 w=0.82u l=0.6u
X236 vdd _00_ a_14260_7933# vdd pmos_6p0 w=0.62u l=0.5u
X237 vdd _25_ a_12020_4539# vdd pmos_6p0 w=0.62u l=0.5u
X238 outp a_3055_3728# vdd vdd pmos_6p0 w=1.095u l=0.5u
X239 a_15507_3229# a_15044_3229# vss vss nmos_6p0 w=0.36u l=0.6u
X240 vdd trim_p[3] a_14703_8432# vdd pmos_6p0 w=0.62u l=0.5u
X241 vss a_15496_8308# a_14723_7933# vss nmos_6p0 w=0.36u l=0.6u
X242 outp a_3075_3229# vss vss nmos_6p0 w=0.82u l=0.6u
X243 vss a_8573_7889# a_7636_7933# vss nmos_6p0 w=0.36u l=0.6u
X244 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X245 a_3757_7553# _00_ vss vss nmos_6p0 w=0.36u l=0.6u
X246 vdd _23_ a_7092_4539# vdd pmos_6p0 w=0.62u l=0.5u
X247 outp a_16831_5296# vdd vdd pmos_6p0 w=1.095u l=0.5u
X248 vss trim_p[0] a_2388_7933# vss nmos_6p0 w=0.36u l=0.6u
X249 a_6060_6647# a_5972_6744# vss vss nmos_6p0 w=0.82u l=1u
X250 outp a_11567_3728# vdd vdd pmos_6p0 w=1.095u l=0.5u
X251 a_14684_3511# a_14596_3608# vss vss nmos_6p0 w=0.82u l=1u
X252 vdd a_4380_6647# a_4292_6744# vdd pmos_6p0 w=1.22u l=1u
X253 a_3075_3229# trim_n[0] a_3055_3728# vss nmos_6p0 w=0.36u l=0.6u
X254 a_17932_3511# a_17844_3608# vss vss nmos_6p0 w=0.82u l=1u
X255 a_4604_3944# a_4516_3988# vss vss nmos_6p0 w=0.82u l=1u
X256 vdd trim_n[3] a_15487_3728# vdd pmos_6p0 w=0.62u l=0.5u
X257 outn _13_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X258 vdd a_9644_5512# a_9556_5556# vdd pmos_6p0 w=1.22u l=1u
X259 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X260 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X261 _23_ a_5837_3944# vdd vdd pmos_6p0 w=1.22u l=0.5u
X262 a_11587_7933# a_11124_7933# vss vss nmos_6p0 w=0.36u l=0.6u
X263 outn _19_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X264 outp a_11587_3229# vss vss nmos_6p0 w=0.82u l=0.6u
X265 outn a_15487_3728# vdd vdd pmos_6p0 w=1.095u l=0.5u
X266 vdd a_5948_7080# a_5860_7124# vdd pmos_6p0 w=1.22u l=1u
X267 a_4157_4728# a_4157_4728# vss vss nmos_6p0 w=0.82u l=0.6u
X268 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X269 vss a_3981_4417# a_3044_4539# vss nmos_6p0 w=0.36u l=0.6u
X270 vdd a_17699_6040# _20_ vdd pmos_6p0 w=1.22u l=0.5u
X271 _19_ a_6509_3944# vdd vdd pmos_6p0 w=1.22u l=0.5u
X272 outp _18_ vss vss nmos_6p0 w=0.82u l=0.6u
X273 a_14012_7080# a_13924_7124# vss vss nmos_6p0 w=0.82u l=1u
X274 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X275 a_6060_8215# a_5972_8312# vss vss nmos_6p0 w=0.82u l=1u
X276 vdd a_3757_7553# a_2780_7156# vdd pmos_6p0 w=0.62u l=0.5u
X277 vss a_3044_4539# outn vss nmos_6p0 w=0.82u l=0.6u
X278 a_17932_8215# a_17844_8312# vss vss nmos_6p0 w=0.82u l=1u
X279 _12_ a_16365_5512# vdd vdd pmos_6p0 w=1.22u l=0.5u
X280 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X281 vss signal signal_n vss nmos_6p0 w=0.82u l=0.6u
X282 outn a_11587_7933# vss vss nmos_6p0 w=0.82u l=0.6u
X283 a_14723_7933# a_14260_7933# vss vss nmos_6p0 w=0.36u l=0.6u
X284 a_12463_3988# a_13256_3976# a_12483_4539# vdd pmos_6p0 w=0.62u l=0.5u
X285 vdd _22_ a_2612_3229# vdd pmos_6p0 w=0.62u l=0.5u
X286 a_5165_3944# a_5165_3944# vss vss nmos_6p0 w=0.82u l=0.6u
X287 a_7636_7933# a_7204_7933# vss vss nmos_6p0 w=0.36u l=0.6u
X288 vdd _00_ a_14372_7675# vdd pmos_6p0 w=0.62u l=0.5u
X289 vdd trim_n[0] a_2612_4020# vdd pmos_6p0 w=0.62u l=0.5u
X290 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X291 vss a_12452_7675# outp vss nmos_6p0 w=0.82u l=0.6u
X292 vss _24_ a_7204_3229# vss nmos_6p0 w=0.36u l=0.6u
X293 a_2588_5079# a_2500_5176# vss vss nmos_6p0 w=0.82u l=1u
X294 outp _10_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X295 a_7555_4539# trim_n[1] a_7535_3988# vss nmos_6p0 w=0.36u l=0.6u
X296 a_15487_3728# a_15044_3229# vdd vdd pmos_6p0 w=0.62u l=0.5u
X297 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X298 a_13389_7553# _00_ vss vss nmos_6p0 w=0.36u l=0.6u
X299 outn a_11567_8432# vdd vdd pmos_6p0 w=1.095u l=0.5u
X300 a_13256_3976# trim_n[2] vss vss nmos_6p0 w=0.36u l=0.6u
X301 a_8440_3604# trim_n[1] vss vss nmos_6p0 w=0.36u l=0.6u
X302 a_1692_3944# a_1604_3988# vss vss nmos_6p0 w=0.82u l=1u
X303 vdd trim_p[2] a_12020_7156# vdd pmos_6p0 w=0.62u l=0.5u
X304 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X305 vdd a_3757_7889# a_2780_8400# vdd pmos_6p0 w=0.62u l=0.5u
X306 a_8328_3976# trim_n[1] vdd vdd pmos_6p0 w=0.62u l=0.5u
X307 vdd a_16812_5512# a_16724_5556# vdd pmos_6p0 w=1.22u l=1u
X308 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X309 vss a_6947_4772# a_6947_4772# vss nmos_6p0 w=0.82u l=0.6u
X310 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X311 a_4829_3160# a_4829_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X312 vdd trim_n[3] a_16831_5296# vdd pmos_6p0 w=0.62u l=0.5u
X313 a_8440_3604# trim_n[1] vdd vdd pmos_6p0 w=0.62u l=0.5u
X314 a_2820_7675# a_2388_7156# a_2780_7156# vdd pmos_6p0 w=0.62u l=0.5u
X315 vss _14_ outp vss nmos_6p0 w=0.82u l=0.6u
X316 a_3848_3604# trim_n[0] vss vss nmos_6p0 w=0.36u l=0.6u
X317 vss a_17624_5172# a_16851_4797# vss nmos_6p0 w=0.36u l=0.6u
X318 a_14835_7675# trim_p[3] a_14815_7124# vss nmos_6p0 w=0.36u l=0.6u
X319 outp _06_ vss vss nmos_6p0 w=0.82u l=0.6u
X320 vss _00_ outp vss nmos_6p0 w=0.82u l=0.6u
X321 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X322 vdd a_6060_6647# a_5972_6744# vdd pmos_6p0 w=1.22u l=1u
X323 vdd a_14684_3511# a_14596_3608# vdd pmos_6p0 w=1.22u l=1u
X324 a_7647_3728# a_8440_3604# a_7667_3229# vdd pmos_6p0 w=0.62u l=0.5u
X325 vdd a_17932_3511# a_17844_3608# vdd pmos_6p0 w=1.22u l=1u
X326 vdd _11_ outn vdd pmos_6p0 w=1.22u l=0.5u
X327 outp _08_ vss vss nmos_6p0 w=0.82u l=0.6u
X328 a_3044_4539# a_2612_4020# vss vss nmos_6p0 w=0.36u l=0.6u
X329 a_2780_7156# trim_p[0] a_2820_7675# vss nmos_6p0 w=0.36u l=0.6u
X330 vdd a_5612_8215# a_5524_8312# vdd pmos_6p0 w=1.22u l=1u
X331 a_3848_3604# trim_n[0] vdd vdd pmos_6p0 w=0.62u l=0.5u
X332 outp _12_ vss vss nmos_6p0 w=0.82u l=0.6u
X333 a_14815_7124# a_14372_7675# vdd vdd pmos_6p0 w=0.62u l=0.5u
X334 a_2780_8400# trim_p[0] vdd vdd pmos_6p0 w=0.62u l=0.5u
X335 a_1692_5079# a_1604_5176# vss vss nmos_6p0 w=0.82u l=1u
X336 a_2553_6875# _00_ vdd vdd pmos_6p0 w=0.565u l=0.5u
X337 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X338 a_15608_7112# trim_p[3] vss vss nmos_6p0 w=0.36u l=0.6u
X339 vdd a_2780_7156# outp vdd pmos_6p0 w=1.095u l=0.5u
X340 a_5949_3160# a_5949_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X341 a_12360_3604# trim_n[2] vss vss nmos_6p0 w=0.36u l=0.6u
X342 outn a_7535_3988# vdd vdd pmos_6p0 w=1.095u l=0.5u
X343 a_15608_7112# trim_p[3] vdd vdd pmos_6p0 w=0.62u l=0.5u
X344 outp a_16851_4797# vss vss nmos_6p0 w=0.82u l=0.6u
X345 a_1924_6040# enable a_1716_6040# vss nmos_6p0 w=0.365u l=0.6u
X346 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X347 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X348 a_5612_5079# a_5524_5176# vss vss nmos_6p0 w=0.82u l=1u
X349 vdd a_6844_7080# a_6756_7124# vdd pmos_6p0 w=1.22u l=1u
X350 vss a_13256_3976# a_12483_4539# vss nmos_6p0 w=0.36u l=0.6u
X351 vss a_8440_3604# a_7667_3229# vss nmos_6p0 w=0.36u l=0.6u
X352 vss _27_ a_15044_3229# vss nmos_6p0 w=0.36u l=0.6u
X353 a_17624_5172# trim_n[3] vdd vdd pmos_6p0 w=0.62u l=0.5u
X354 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X355 a_8301_4728# a_8301_4728# vss vss nmos_6p0 w=0.82u l=0.6u
X356 a_14237_3944# a_14237_3944# vss vss nmos_6p0 w=0.82u l=0.6u
X357 a_11567_8432# a_11124_7933# vdd vdd pmos_6p0 w=0.62u l=0.5u
X358 vss _15_ outn vss nmos_6p0 w=0.82u l=0.6u
X359 a_12360_3604# trim_n[2] vdd vdd pmos_6p0 w=0.62u l=0.5u
X360 a_6285_4728# a_6285_4728# vss vss nmos_6p0 w=0.82u l=0.6u
X361 a_3036_5079# a_2948_5176# vss vss nmos_6p0 w=0.82u l=1u
X362 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X363 outn _09_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X364 outp _01_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X365 a_2140_3944# a_2052_3988# vss vss nmos_6p0 w=0.82u l=1u
X366 vss _00_ outp vss nmos_6p0 w=0.82u l=0.6u
X367 vss a_6835_6340# a_6835_6340# vss nmos_6p0 w=0.82u l=0.6u
X368 a_7596_8400# trim_p[1] a_7636_7933# vss nmos_6p0 w=0.36u l=0.6u
X369 _21_ a_4157_4728# vdd vdd pmos_6p0 w=1.22u l=0.5u
X370 vdd a_2780_8400# outn vdd pmos_6p0 w=1.095u l=0.5u
X371 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X372 a_11567_3728# a_12360_3604# a_11587_3229# vdd pmos_6p0 w=0.62u l=0.5u
X373 vss a_3848_3604# a_3075_3229# vss nmos_6p0 w=0.36u l=0.6u
X374 a_16851_4797# trim_n[3] a_16831_5296# vss nmos_6p0 w=0.36u l=0.6u
X375 vss a_8328_3976# a_7555_4539# vss nmos_6p0 w=0.36u l=0.6u
X376 vdd a_5500_7080# a_5412_7124# vdd pmos_6p0 w=1.22u l=1u
X377 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X378 a_2029_3160# a_2029_3160# vss vss nmos_6p0 w=0.82u l=0.6u
X379 outn _02_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X380 outn _02_ vss vss nmos_6p0 w=0.82u l=0.6u
X381 vdd a_4604_3944# a_4516_3988# vdd pmos_6p0 w=1.22u l=1u
X382 outp _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X383 vss trim_n[0] a_2612_4020# vss nmos_6p0 w=0.36u l=0.6u
X384 outn _00_ vss vss nmos_6p0 w=0.82u l=0.6u
X385 a_3484_5079# a_3396_5176# vss vss nmos_6p0 w=0.82u l=1u
X386 a_2820_7675# a_2388_7156# vss vss nmos_6p0 w=0.36u l=0.6u
X387 _00_ enable vss vss nmos_6p0 w=0.82u l=0.6u
X388 vdd a_13389_7553# a_12412_7156# vdd pmos_6p0 w=0.62u l=0.5u
X389 vdd a_4640_7864# _01_ vdd pmos_6p0 w=1.22u l=0.5u
X390 outp _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X391 a_3075_3229# a_2612_3229# vss vss nmos_6p0 w=0.36u l=0.6u
X392 _24_ a_4829_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X393 a_14703_8432# a_14260_7933# vdd vdd pmos_6p0 w=0.62u l=0.5u
X394 outn _00_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X395 vss _20_ outp vss nmos_6p0 w=0.82u l=0.6u
X396 vss _00_ a_11124_7933# vss nmos_6p0 w=0.36u l=0.6u
X397 a_3296_6296# _03_ vdd vdd pmos_6p0 w=0.565u l=0.5u
X398 vss a_15608_7112# a_14835_7675# vss nmos_6p0 w=0.36u l=0.6u
X399 vdd a_2588_5079# a_2500_5176# vdd pmos_6p0 w=1.22u l=1u
X400 a_10093_3944# a_10093_3944# vss vss nmos_6p0 w=0.82u l=0.6u
X401 vss a_12360_3604# a_11587_3229# vss nmos_6p0 w=0.36u l=0.6u
X402 outn a_15507_3229# vss vss nmos_6p0 w=0.82u l=0.6u
X403 vdd a_12412_7156# outp vdd pmos_6p0 w=1.095u l=0.5u
X404 a_12483_4539# trim_n[2] a_12463_3988# vss nmos_6p0 w=0.36u l=0.6u
X405 a_2140_5079# a_2052_5176# vss vss nmos_6p0 w=0.82u l=1u
X406 a_7535_3988# a_7092_4539# vdd vdd pmos_6p0 w=0.62u l=0.5u
X407 a_13256_3976# trim_n[2] vdd vdd pmos_6p0 w=0.62u l=0.5u
X408 vss a_15683_4772# a_15683_4772# vss nmos_6p0 w=0.82u l=0.6u
X409 outp _01_ vss vss nmos_6p0 w=0.82u l=0.6u
X410 _27_ a_5165_3944# vdd vdd pmos_6p0 w=1.22u l=0.5u
X411 vdd _14_ outp vdd pmos_6p0 w=1.22u l=0.5u
X412 a_5501_5512# a_5501_5512# vss vss nmos_6p0 w=0.82u l=0.6u
X413 a_7636_7675# a_7204_7156# a_7596_7156# vdd pmos_6p0 w=0.62u l=0.5u
X414 vss _00_ a_14260_7933# vss nmos_6p0 w=0.36u l=0.6u
X415 vss _00_ outp vss nmos_6p0 w=0.82u l=0.6u
X416 a_12452_7675# a_12020_7156# a_12412_7156# vdd pmos_6p0 w=0.62u l=0.5u
X417 _26_ a_5949_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X418 vdd trim_p[1] a_7204_7156# vdd pmos_6p0 w=0.62u l=0.5u
X419 vss a_8573_7553# a_7636_7675# vss nmos_6p0 w=0.36u l=0.6u
X420 vss a_3296_6296# _02_ vss nmos_6p0 w=0.82u l=0.6u
X421 vdd a_1692_3944# a_1604_3988# vdd pmos_6p0 w=1.22u l=1u
X422 vss a_13389_7553# a_12452_7675# vss nmos_6p0 w=0.36u l=0.6u
X423 a_9644_3944# a_9556_3988# vss vss nmos_6p0 w=0.82u l=1u
X424 a_4716_5512# a_4628_5556# vss vss nmos_6p0 w=0.82u l=1u
X425 a_7555_4539# a_7092_4539# vss vss nmos_6p0 w=0.36u l=0.6u
X426 vdd _28_ a_16388_4797# vdd pmos_6p0 w=0.62u l=0.5u
X427 vdd trim_p[3] a_14815_7124# vdd pmos_6p0 w=0.62u l=0.5u
X428 vss trim_p[0] a_2388_7156# vss nmos_6p0 w=0.36u l=0.6u
X429 outn _05_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X430 a_7596_8400# trim_p[1] vdd vdd pmos_6p0 w=0.62u l=0.5u
X431 vss a_4640_7864# _01_ vss nmos_6p0 w=0.82u l=0.6u
X432 outn _19_ vss vss nmos_6p0 w=0.82u l=0.6u
X433 vdd a_17475_3204# _07_ vdd pmos_6p0 w=1.22u l=0.5u
X434 a_17624_5172# trim_n[3] vss vss nmos_6p0 w=0.36u l=0.6u
X435 vdd a_1692_5079# a_1604_5176# vdd pmos_6p0 w=1.22u l=1u
X436 a_4828_6647# a_4740_6744# vss vss nmos_6p0 w=0.82u l=1u
X437 a_12360_8308# trim_p[2] vdd vdd pmos_6p0 w=0.62u l=0.5u
X438 outn a_14815_7124# vdd vdd pmos_6p0 w=1.095u l=0.5u
X439 vdd _24_ a_7204_3229# vdd pmos_6p0 w=0.62u l=0.5u
X440 outp a_14723_7933# vss vss nmos_6p0 w=0.82u l=0.6u
X441 a_3004_4020# trim_n[0] a_3044_4539# vss nmos_6p0 w=0.36u l=0.6u
X442 a_4640_7864# _04_ vdd vdd pmos_6p0 w=0.565u l=0.5u
X443 a_11567_8432# a_12360_8308# a_11587_7933# vdd pmos_6p0 w=0.62u l=0.5u
X444 _22_ a_2029_3160# vdd vdd pmos_6p0 w=1.22u l=0.5u
X445 outp _16_ vdd vdd pmos_6p0 w=1.22u l=0.5u
X446 outn a_12463_3988# vdd vdd pmos_6p0 w=1.095u l=0.5u
X447 outn _13_ vss vss nmos_6p0 w=0.82u l=0.6u
X448 vdd a_5612_5079# a_5524_5176# vdd pmos_6p0 w=1.22u l=1u
X449 a_14835_7675# a_14372_7675# vss vss nmos_6p0 w=0.36u l=0.6u
X450 a_11587_3229# trim_n[2] a_11567_3728# vss nmos_6p0 w=0.36u l=0.6u
X451 a_3044_4539# a_2612_4020# a_3004_4020# vdd pmos_6p0 w=0.62u l=0.5u
X452 vdd a_2161_6296# _04_ vdd pmos_6p0 w=1.22u l=0.5u
X453 vdd a_6396_7080# a_6308_7124# vdd pmos_6p0 w=1.22u l=1u
C0 _27_ _07_ 2.90fF
C1 outp vdd 5.81fF
C2 _10_ _19_ 3.02fF
C3 outn vdd 5.93fF
C4 _00_ vdd 3.45fF
C5 _00_ _17_ 2.81fF
C6 _08_ outn 3.45fF
C7 outp outn 5.06fF
C8 _00_ outp 6.12fF
C9 _28_ outn 2.17fF
C10 _00_ _28_ 2.35fF
C11 _16_ _00_ 2.42fF
C12 _00_ outn 6.24fF
C13 trim_n[2] vss 2.73fF
C14 trim_n[1] vss 2.75fF
C15 trim_n[0] vss 2.69fF
C16 trim_n[3] vss 2.90fF
C17 trim_p[3] vss 2.63fF
C18 trim_p[2] vss 2.71fF
C19 trim_p[1] vss 2.58fF
C20 outn vss 7.10fF
C21 trim_p[0] vss 2.57fF
C22 outp vss 7.76fF
C23 vdd vss 178.33fF
C24 _00_ vss 22.42fF $ **FLOATING
.ends
