VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caparray_s1
  CLASS BLOCK ;
  FOREIGN caparray_s1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 350.000 ;
  PIN cap_series_gygyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.400 346.000 232.960 350.000 ;
    END
  END cap_series_gygyn
  PIN cap_series_gygyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 346.000 202.160 350.000 ;
    END
  END cap_series_gygyp
  PIN cap_series_gyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 346.000 171.360 350.000 ;
    END
  END cap_series_gyn
  PIN cap_series_gyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 346.000 140.560 350.000 ;
    END
  END cap_series_gyp
  PIN cap_shunt_gyn
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.200 346.000 109.760 350.000 ;
    END
  END cap_shunt_gyn
  PIN cap_shunt_gyp
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 346.000 78.960 350.000 ;
    END
  END cap_shunt_gyp
  PIN cap_shunt_n
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.600 346.000 48.160 350.000 ;
    END
  END cap_shunt_n
  PIN cap_shunt_p
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 346.000 17.360 350.000 ;
    END
  END cap_shunt_p
  PIN tune_series_gy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.720 0.000 21.280 4.000 ;
    END
  END tune_series_gy[0]
  PIN tune_series_gy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.160 0.000 62.720 4.000 ;
    END
  END tune_series_gy[1]
  PIN tune_series_gy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.600 0.000 104.160 4.000 ;
    END
  END tune_series_gy[2]
  PIN tune_series_gy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.040 0.000 145.600 4.000 ;
    END
  END tune_series_gy[3]
  PIN tune_series_gy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.480 0.000 187.040 4.000 ;
    END
  END tune_series_gy[4]
  PIN tune_series_gy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.920 0.000 228.480 4.000 ;
    END
  END tune_series_gy[5]
  PIN tune_series_gygy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 13.440 250.000 14.000 ;
    END
  END tune_series_gygy[0]
  PIN tune_series_gygy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 40.320 250.000 40.880 ;
    END
  END tune_series_gygy[1]
  PIN tune_series_gygy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 67.200 250.000 67.760 ;
    END
  END tune_series_gygy[2]
  PIN tune_series_gygy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 94.080 250.000 94.640 ;
    END
  END tune_series_gygy[3]
  PIN tune_series_gygy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 120.960 250.000 121.520 ;
    END
  END tune_series_gygy[4]
  PIN tune_series_gygy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 147.840 250.000 148.400 ;
    END
  END tune_series_gygy[5]
  PIN tune_shunt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.840 4.000 22.400 ;
    END
  END tune_shunt[0]
  PIN tune_shunt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 65.520 4.000 66.080 ;
    END
  END tune_shunt[1]
  PIN tune_shunt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.200 4.000 109.760 ;
    END
  END tune_shunt[2]
  PIN tune_shunt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.880 4.000 153.440 ;
    END
  END tune_shunt[3]
  PIN tune_shunt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.560 4.000 197.120 ;
    END
  END tune_shunt[4]
  PIN tune_shunt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.240 4.000 240.800 ;
    END
  END tune_shunt[5]
  PIN tune_shunt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.920 4.000 284.480 ;
    END
  END tune_shunt[6]
  PIN tune_shunt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 327.600 4.000 328.160 ;
    END
  END tune_shunt[7]
  PIN tune_shunt_gy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 174.720 250.000 175.280 ;
    END
  END tune_shunt_gy[0]
  PIN tune_shunt_gy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 201.600 250.000 202.160 ;
    END
  END tune_shunt_gy[1]
  PIN tune_shunt_gy[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 228.480 250.000 229.040 ;
    END
  END tune_shunt_gy[2]
  PIN tune_shunt_gy[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 255.360 250.000 255.920 ;
    END
  END tune_shunt_gy[3]
  PIN tune_shunt_gy[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 282.240 250.000 282.800 ;
    END
  END tune_shunt_gy[4]
  PIN tune_shunt_gy[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 309.120 250.000 309.680 ;
    END
  END tune_shunt_gy[5]
  PIN tune_shunt_gy[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 336.000 250.000 336.560 ;
    END
  END tune_shunt_gy[6]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 333.500 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 333.500 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 243.040 333.500 ;
      LAYER Metal2 ;
        RECT 9.100 345.700 16.500 346.500 ;
        RECT 17.660 345.700 47.300 346.500 ;
        RECT 48.460 345.700 78.100 346.500 ;
        RECT 79.260 345.700 108.900 346.500 ;
        RECT 110.060 345.700 139.700 346.500 ;
        RECT 140.860 345.700 170.500 346.500 ;
        RECT 171.660 345.700 201.300 346.500 ;
        RECT 202.460 345.700 232.100 346.500 ;
        RECT 233.260 345.700 240.660 346.500 ;
        RECT 9.100 4.300 240.660 345.700 ;
        RECT 9.100 4.000 20.420 4.300 ;
        RECT 21.580 4.000 61.860 4.300 ;
        RECT 63.020 4.000 103.300 4.300 ;
        RECT 104.460 4.000 144.740 4.300 ;
        RECT 145.900 4.000 186.180 4.300 ;
        RECT 187.340 4.000 227.620 4.300 ;
        RECT 228.780 4.000 240.660 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 335.700 245.700 336.420 ;
        RECT 4.000 328.460 246.820 335.700 ;
        RECT 4.300 327.300 246.820 328.460 ;
        RECT 4.000 309.980 246.820 327.300 ;
        RECT 4.000 308.820 245.700 309.980 ;
        RECT 4.000 284.780 246.820 308.820 ;
        RECT 4.300 283.620 246.820 284.780 ;
        RECT 4.000 283.100 246.820 283.620 ;
        RECT 4.000 281.940 245.700 283.100 ;
        RECT 4.000 256.220 246.820 281.940 ;
        RECT 4.000 255.060 245.700 256.220 ;
        RECT 4.000 241.100 246.820 255.060 ;
        RECT 4.300 239.940 246.820 241.100 ;
        RECT 4.000 229.340 246.820 239.940 ;
        RECT 4.000 228.180 245.700 229.340 ;
        RECT 4.000 202.460 246.820 228.180 ;
        RECT 4.000 201.300 245.700 202.460 ;
        RECT 4.000 197.420 246.820 201.300 ;
        RECT 4.300 196.260 246.820 197.420 ;
        RECT 4.000 175.580 246.820 196.260 ;
        RECT 4.000 174.420 245.700 175.580 ;
        RECT 4.000 153.740 246.820 174.420 ;
        RECT 4.300 152.580 246.820 153.740 ;
        RECT 4.000 148.700 246.820 152.580 ;
        RECT 4.000 147.540 245.700 148.700 ;
        RECT 4.000 121.820 246.820 147.540 ;
        RECT 4.000 120.660 245.700 121.820 ;
        RECT 4.000 110.060 246.820 120.660 ;
        RECT 4.300 108.900 246.820 110.060 ;
        RECT 4.000 94.940 246.820 108.900 ;
        RECT 4.000 93.780 245.700 94.940 ;
        RECT 4.000 68.060 246.820 93.780 ;
        RECT 4.000 66.900 245.700 68.060 ;
        RECT 4.000 66.380 246.820 66.900 ;
        RECT 4.300 65.220 246.820 66.380 ;
        RECT 4.000 41.180 246.820 65.220 ;
        RECT 4.000 40.020 245.700 41.180 ;
        RECT 4.000 22.700 246.820 40.020 ;
        RECT 4.300 21.540 246.820 22.700 ;
        RECT 4.000 14.300 246.820 21.540 ;
        RECT 4.000 13.580 245.700 14.300 ;
      LAYER Metal4 ;
        RECT 42.140 229.130 42.420 236.230 ;
  END
END caparray_s1
END LIBRARY

