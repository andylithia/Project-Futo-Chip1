* NGSPICE file created from user_proj_example.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_1 EN I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18]
+ la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29]
+ la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45]
+ la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50]
+ la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56]
+ la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__036__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_206 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[6\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PD\[3\].pdp_22 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[2\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_207 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_inj.gen_TRIM\[2\].ptrimn_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_inj.psijn_215 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_TRIM\[1\].ptrimp_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_inj.gen_PU\[17\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input3_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[0\].pdp_16 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_208 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_inj.gen_PU\[13\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PD\[4\].pdn_23 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_TRIM\[0\].ntrimn u_inj.trim_n_r\[0\] net31 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA__039__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_209 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[6\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__037__D net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[1\].pdn_17 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[2\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_TRIM\[1\].ptrimn_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_TRIM\[0\].ptrimp_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_TRIM\[0\].ntrimp u_inj.trim_n_r\[0\] net32 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_190 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_040_ net9 net10 u_inj.trim_n_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_TRIM\[1\].ptrimn u_inj.trim_p_r\[1\] net14 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_180 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_191 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_TRIM\[3\].ntrimn u_inj.trim_n_r\[3\] net37 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_170 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_181 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_192 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[7\].pdn net29 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_90 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_inj.nsijn _001_ u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[16\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_TRIM\[1\].ptrimp u_inj.trim_p_r\[1\] net14 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_171 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_160 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_182 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_193 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_u_inj.gen_TRIM\[0\].ptrimn_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_80 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_91 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PD\[6\].pdn net27 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[12\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_TRIM\[3\].ntrimp u_inj.trim_n_r\[3\] net38 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.siginv_39 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_172 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_161 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_150 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_183 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_194 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[7\].pdp net30 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_16_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__031__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_70 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_proj_example_81 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_92 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.nsijp net214 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[5\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[5\].pdn net25 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_inj.gen_PD\[2\].pdp_20 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout13_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_140 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_173 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_151 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_162 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_184 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_195 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_TRIM\[0\].ntrimp_32 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_71 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_60 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_82 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_93 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PD\[6\].pdp net28 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[1\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[6\].pdp_28 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[16\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_130 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_141 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_174 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_163 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_152 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_185 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_196 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xu_inj.gen_PD\[4\].pdn net23 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_inj.gen_TRIM\[1\].ntrimp_34 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_72 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_61 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_50 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_83 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_94 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__035__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[3\].pdn_21 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[5\].pdp net26 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_u_inj.gen_PU\[12\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_131 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_120 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_142 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_153 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_175 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_164 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input8_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_197 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_186 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[3\].pdn net21 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_16_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.siginv net39 u_inj.signal_n vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_73 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_62 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_51 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_40 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_84 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_95 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout11 net13 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_inj.gen_PD\[7\].pdn_29 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_inj.gen_TRIM\[2\].ntrimp_36 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_inj.gen_PU\[5\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_inj.gen_PD\[0\].pdn_15 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_176 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_132 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_165 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_121 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_154 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_110 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_143 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_187 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xu_inj.gen_PD\[4\].pdp net24 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xuser_proj_example_198 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_52 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_41 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_74 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_63 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_85 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_96 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout12 net13 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[2\].pdn net19 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_TRIM\[3\].ntrimp_38 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_u_inj.gen_PU\[1\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 io_in[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_177 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_133 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_166 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_122 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_155 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_111 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_144 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_199 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_188 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_100 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[18\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__038__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[3\].pdp net22 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_16_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_75 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_64 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_53 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_42 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_86 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_97 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout13 net14 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_10_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 io_in[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PD\[1\].pdn net17 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_112 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_101 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_178 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_134 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_167 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_123 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_156 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_145 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_189 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[17\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__040__D net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_76 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_65 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_54 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_43 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_87 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_98 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout14 _000_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__035__D net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[2\].pdp net20 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput4 io_in[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_135 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_113 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_124 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_102 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_179 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_168 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_157 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_146 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[18\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_16_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PD\[0\].pdn net15 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_039_ net8 net10 u_inj.trim_n_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__038__D net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_77 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_66 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_55 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_44 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_88 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_99 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[16\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 io_in[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_TRIM\[0\].ptrimn u_inj.trim_p_r\[0\] net14 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_0_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[1\].pdp net18 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[15\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_136 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_169 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_125 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_158 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_114 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_147 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_103 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_038_ net7 net10 u_inj.trim_n_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[17\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_78 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_67 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_56 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_45 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_89 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_TRIM\[2\].ntrimn u_inj.trim_n_r\[2\] net35 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput6 io_in[5] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PU\[15\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_137 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_126 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_159 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_148 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_115 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_104 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[8\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PD\[0\].pdp net16 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_16_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_037_ net6 net10 u_inj.trim_n_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_68 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_57 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_46 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_79 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[16\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 io_in[6] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_TRIM\[0\].ptrimp u_inj.trim_p_r\[0\] net14 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_inj.gen_PU\[4\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_138 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_127 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_116 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_105 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_149 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 io_in[9] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_036_ net5 net10 u_inj.trim_p_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PU\[14\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_69 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_58 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_47 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_inj.gen_TRIM\[2\].ntrimp u_inj.trim_n_r\[2\] net36 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
Xu_inj.gen_PD\[5\].pdp_26 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 io_in[7] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_inj.gen_PU\[0\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[15\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_106 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_117 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_139 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_128 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[15\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_035_ net4 net10 u_inj.trim_p_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_59 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_48 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_TRIM\[3\].ptrimn u_inj.trim_p_r\[3\] net14 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PU\[13\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_inj.gen_PU\[9\].pun net13 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_10_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_TRIM\[0\].ntrimn_31 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput9 io_in[8] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[11\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_129 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_118 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_107 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_034_ net3 net10 u_inj.trim_p_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_inj.gen_PU\[14\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PD\[6\].pdn_27 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_49 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.psijn net215 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_input10_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PU\[12\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[8\].pun net13 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_15_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_TRIM\[1\].ntrimn_33 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_119 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_108 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_inj.gen_PU\[4\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_033_ net2 net10 u_inj.trim_p_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_TRIM\[3\].ptrimp u_inj.trim_p_r\[3\] net14 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
Xu_inj.gen_PU\[13\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__034__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[9\].pup net13 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__242__I u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[0\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_109 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PU\[11\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_inj.gen_TRIM\[2\].ntrimn_35 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[7\].pun net13 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_032_ _002_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.psijp _001_ u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[12\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_inj.gen_PU\[8\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_031_ net14 u_inj.signal_n _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_TRIM\[3\].ntrimn_37 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_inj.gen_PU\[10\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[6\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[11\].pup net13 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[7\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_030_ net1 _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__037__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[18\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_inj.gen_PU\[5\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_inj.gen_PU\[14\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PU\[10\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PU\[6\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PD\[7\].pdp_30 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xu_inj.gen_PU\[4\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_u_inj.gen_PU\[10\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_243_ u_inj.outn la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[7\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PU\[5\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__036__D net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_242_ u_inj.outp la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_inj.gen_TRIM\[1\].ntrimn u_inj.trim_n_r\[1\] net33 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_15_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PD\[4\].pdp_24 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[3\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__039__D net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_PU\[18\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[4\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[14\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_210 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_inj.gen_PD\[1\].pdp_18 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xu_inj.gen_PU\[2\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__040__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PD\[5\].pdn_25 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_inj.gen_PU\[10\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_TRIM\[1\].ntrimp u_inj.trim_n_r\[1\] net34 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_PU\[3\].pup net13 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_211 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_200 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PU\[1\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_inj.gen_TRIM\[3\].ptrimp_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_TRIM\[2\].ptrimn u_inj.trim_p_r\[2\] net14 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[3\].pun_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_inj.gen_PD\[2\].pdn_19 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_212 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_201 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__030__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_inj.gen_PU\[2\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input7_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_inj.gen_PU\[0\].pun net12 u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_6_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_213 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_202 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_inj.gen_PU\[1\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_inj.nsijp_214 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_10_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_inj.gen_TRIM\[2\].ptrimp u_inj.trim_p_r\[2\] net14 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_203 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__033__CLK net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_inj.gen_PU\[0\].pup net11 u_inj.outp vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_TRIM\[3\].ptrimn_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_inj.gen_TRIM\[2\].ptrimp_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_204 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_inj.gen_PU\[17\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__243__I u_inj.outn vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_inj.gen_PU\[13\].pup_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_205 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

