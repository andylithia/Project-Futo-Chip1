magic
tech gf180mcuC
magscale 1 10
timestamp 1669957629
<< nwell >>
rect 1000 1317 1300 2905
rect 1000 486 1300 954
<< pwell >>
rect 1000 2905 1300 3259
rect 1000 954 1300 1317
rect 1000 0 1300 486
<< psubdiff >>
rect 1100 3210 1200 3230
rect 1100 2960 1120 3210
rect 1180 2960 1200 3210
rect 1100 2940 1200 2960
rect 1100 1260 1200 1280
rect 1100 1010 1120 1260
rect 1180 1010 1200 1260
rect 1100 990 1200 1010
rect 1100 430 1200 450
rect 1100 50 1120 430
rect 1180 50 1200 430
rect 1100 30 1200 50
<< nsubdiff >>
rect 1100 2850 1200 2870
rect 1100 1370 1120 2850
rect 1180 1370 1200 2850
rect 1100 1350 1200 1370
rect 1100 900 1200 920
rect 1100 540 1120 900
rect 1180 540 1200 900
rect 1100 520 1200 540
<< psubdiffcont >>
rect 1120 2960 1180 3210
rect 1120 1010 1180 1260
rect 1120 50 1180 430
<< nsubdiffcont >>
rect 1120 1370 1180 2850
rect 1120 540 1180 900
<< metal1 >>
rect 1110 3210 1190 3230
rect 1110 2960 1120 3210
rect 1180 2960 1190 3210
rect 1110 2940 1190 2960
rect 1110 2850 1190 2870
rect 1110 1370 1120 2850
rect 1180 1370 1190 2850
rect 1110 1350 1190 1370
rect 1110 1260 1190 1280
rect 1110 1010 1120 1260
rect 1180 1010 1190 1260
rect 1110 990 1190 1010
rect 1110 900 1190 920
rect 1110 540 1120 900
rect 1180 540 1190 900
rect 1110 520 1190 540
rect 1110 430 1190 450
rect 1110 50 1120 430
rect 1180 50 1190 430
rect 1110 30 1190 50
<< via1 >>
rect 1120 2960 1180 3210
rect 1120 1370 1180 2850
rect 1120 1010 1180 1260
rect 1120 540 1180 900
rect 1120 50 1180 430
<< metal2 >>
rect 1100 3210 1200 3230
rect 1100 3030 1120 3210
rect 1180 3030 1200 3210
rect 1100 2950 1110 3030
rect 1190 2950 1200 3030
rect 1100 2940 1200 2950
rect 1100 2850 1200 2870
rect 1100 1440 1120 2850
rect 1180 1440 1200 2850
rect 1100 1360 1110 1440
rect 1190 1360 1200 1440
rect 1100 1350 1200 1360
rect 1100 1260 1200 1280
rect 1100 1080 1120 1260
rect 1180 1080 1200 1260
rect 1100 1000 1110 1080
rect 1190 1000 1200 1080
rect 1100 990 1200 1000
rect 1100 910 1200 920
rect 1100 830 1110 910
rect 1190 830 1200 910
rect 1100 540 1120 830
rect 1180 540 1200 830
rect 1100 520 1200 540
rect 1100 430 1200 450
rect 1100 130 1120 430
rect 1180 130 1200 430
rect 1100 40 1110 130
rect 1190 40 1200 130
rect 1100 30 1200 40
<< via2 >>
rect 1110 2960 1120 3030
rect 1120 2960 1180 3030
rect 1180 2960 1190 3030
rect 1110 2950 1190 2960
rect 1110 1370 1120 1440
rect 1120 1370 1180 1440
rect 1180 1370 1190 1440
rect 1110 1360 1190 1370
rect 1110 1010 1120 1080
rect 1120 1010 1180 1080
rect 1180 1010 1190 1080
rect 1110 1000 1190 1010
rect 1110 900 1190 910
rect 1110 830 1120 900
rect 1120 830 1180 900
rect 1180 830 1190 900
rect 1110 50 1120 130
rect 1120 50 1180 130
rect 1180 50 1190 130
rect 1110 40 1190 50
<< metal3 >>
rect 1100 3030 1200 3040
rect 1100 2950 1110 3030
rect 1190 2950 1200 3030
rect 1100 2940 1200 2950
rect 1100 1440 1200 1450
rect 1100 1360 1110 1440
rect 1190 1360 1200 1440
rect 1100 1350 1200 1360
rect 1100 1080 1200 1090
rect 1100 1000 1110 1080
rect 1190 1000 1200 1080
rect 1100 990 1200 1000
rect 1100 910 1200 920
rect 1100 830 1110 910
rect 1190 830 1200 910
rect 1100 820 1200 830
rect 1100 130 1200 140
rect 1100 40 1110 130
rect 1190 40 1200 130
rect 1100 30 1200 40
<< via3 >>
rect 1110 2950 1190 3030
rect 1110 1360 1190 1440
rect 1110 1000 1190 1080
rect 1110 830 1190 910
rect 1110 40 1190 130
<< metal4 >>
rect 1100 3030 1200 3040
rect 1100 2950 1110 3030
rect 1190 2950 1200 3030
rect 1100 2940 1200 2950
rect 920 1440 1200 1450
rect 920 1360 930 1440
rect 1010 1360 1110 1440
rect 1190 1360 1200 1440
rect 920 1350 1200 1360
rect 740 1080 1200 1090
rect 740 1000 750 1080
rect 830 1000 1110 1080
rect 1190 1000 1200 1080
rect 740 990 1200 1000
rect 560 910 1190 920
rect 560 830 570 910
rect 650 830 1110 910
rect 560 820 1190 830
rect 380 130 1200 140
rect 380 120 1110 130
rect 380 40 390 120
rect 470 40 1110 120
rect 1190 40 1200 130
rect 380 30 1200 40
<< via4 >>
rect 1110 2950 1190 3030
rect 930 1360 1010 1440
rect 750 1000 830 1080
rect 570 830 650 910
rect 390 40 470 120
<< metal5 >>
rect 380 120 480 3350
rect 380 40 390 120
rect 470 40 480 120
rect 380 0 480 40
rect 560 910 660 3350
rect 560 830 570 910
rect 650 830 660 910
rect 560 -30 660 830
rect 740 1080 840 3350
rect 740 1000 750 1080
rect 830 1000 840 1080
rect 740 -30 840 1000
rect 920 1440 1020 3350
rect 920 1360 930 1440
rect 1010 1360 1020 1440
rect 920 -30 1020 1360
rect 1100 3030 1200 3350
rect 1100 2950 1110 3030
rect 1190 2950 1200 3030
rect 1100 -30 1200 2950
<< comment >>
rect 594 2905 597 2915
rect 597 2895 600 2905
rect 594 1317 597 1327
rect 597 1307 600 1317
rect 594 954 597 964
rect 597 944 600 954
rect 594 486 597 496
rect 597 476 600 486
rect 597 0 600 10
rect 594 -10 597 0
<< end >>
