magic
tech gf180mcuC
magscale 1 10
timestamp 1669496281
<< nwell >>
rect 132 1758 648 3714
rect 132 710 648 1268
<< pwell >>
rect 132 3714 648 4240
rect 132 1268 648 1758
rect 132 184 648 710
<< metal1 >>
rect 296 4154 484 4156
rect 296 4098 308 4154
rect 364 4098 416 4154
rect 472 4098 484 4154
rect 296 4096 484 4098
rect 154 4064 214 4076
rect 154 4008 156 4064
rect 212 4040 214 4064
rect 566 4064 626 4076
rect 566 4040 568 4064
rect 212 4008 237 4040
rect 154 3956 237 4008
rect 154 3900 156 3956
rect 212 3924 237 3956
rect 543 4008 568 4040
rect 624 4008 626 4064
rect 543 3956 626 4008
rect 543 3924 568 3956
rect 212 3900 214 3924
rect 154 3888 214 3900
rect 566 3900 568 3924
rect 624 3900 626 3956
rect 566 3888 626 3900
rect 305 3868 490 3869
rect 296 3847 490 3868
rect 296 3808 508 3847
rect 296 3748 673 3808
rect 296 3650 484 3652
rect 296 3594 308 3650
rect 364 3594 416 3650
rect 472 3594 484 3650
rect 296 3592 484 3594
rect 342 3569 438 3592
rect 226 3466 286 3478
rect 226 3410 228 3466
rect 284 3410 286 3466
rect 226 3358 286 3410
rect 226 3302 228 3358
rect 284 3302 286 3358
rect 226 3250 286 3302
rect 226 3194 228 3250
rect 284 3194 286 3250
rect 226 3142 286 3194
rect 226 3086 228 3142
rect 284 3086 286 3142
rect 226 3034 286 3086
rect 226 2978 228 3034
rect 284 2978 286 3034
rect 226 2926 286 2978
rect 226 2870 228 2926
rect 284 2870 286 2926
rect 226 2818 286 2870
rect 226 2762 228 2818
rect 284 2762 286 2818
rect 226 2710 286 2762
rect 226 2654 228 2710
rect 284 2654 286 2710
rect 226 2602 286 2654
rect 226 2546 228 2602
rect 284 2546 286 2602
rect 226 2494 286 2546
rect 226 2438 228 2494
rect 284 2438 286 2494
rect 226 2386 286 2438
rect 226 2330 228 2386
rect 284 2330 286 2386
rect 226 2278 286 2330
rect 226 2222 228 2278
rect 284 2222 286 2278
rect 226 2170 286 2222
rect 226 2114 228 2170
rect 284 2114 286 2170
rect 226 2062 286 2114
rect 226 2006 228 2062
rect 284 2006 286 2062
rect 226 1994 286 2006
rect 494 3466 554 3478
rect 494 3410 496 3466
rect 552 3410 554 3466
rect 494 3358 554 3410
rect 494 3302 496 3358
rect 552 3302 554 3358
rect 494 3250 554 3302
rect 494 3194 496 3250
rect 552 3194 554 3250
rect 494 3142 554 3194
rect 494 3086 496 3142
rect 552 3086 554 3142
rect 494 3034 554 3086
rect 494 2978 496 3034
rect 552 2978 554 3034
rect 494 2926 554 2978
rect 494 2870 496 2926
rect 552 2870 554 2926
rect 494 2818 554 2870
rect 494 2762 496 2818
rect 552 2762 554 2818
rect 494 2710 554 2762
rect 494 2654 496 2710
rect 552 2654 554 2710
rect 494 2602 554 2654
rect 494 2546 496 2602
rect 552 2546 554 2602
rect 494 2494 554 2546
rect 494 2438 496 2494
rect 552 2438 554 2494
rect 494 2386 554 2438
rect 494 2330 496 2386
rect 552 2330 554 2386
rect 494 2278 554 2330
rect 494 2222 496 2278
rect 552 2222 554 2278
rect 494 2170 554 2222
rect 494 2114 496 2170
rect 552 2114 554 2170
rect 494 2062 554 2114
rect 494 2006 496 2062
rect 552 2006 554 2062
rect 494 1994 554 2006
rect 342 1880 438 1903
rect 296 1878 484 1880
rect 296 1822 308 1878
rect 364 1822 416 1878
rect 472 1822 484 1878
rect 296 1820 484 1822
rect 296 1747 484 1749
rect 296 1691 308 1747
rect 364 1691 416 1747
rect 472 1691 484 1747
rect 296 1689 484 1691
rect 332 1666 448 1689
rect 613 1631 673 3748
rect 512 1609 673 1631
rect 107 1419 276 1607
rect 107 1395 266 1419
rect 496 1416 673 1609
rect 107 676 167 1395
rect 332 1337 448 1360
rect 296 1335 484 1337
rect 296 1279 308 1335
rect 364 1279 416 1335
rect 472 1279 484 1335
rect 296 1277 484 1279
rect 296 1202 484 1204
rect 296 1146 308 1202
rect 364 1146 416 1202
rect 472 1146 484 1202
rect 296 1144 484 1146
rect 342 1121 438 1144
rect 226 1070 286 1082
rect 226 1014 228 1070
rect 284 1014 286 1070
rect 226 962 286 1014
rect 226 906 228 962
rect 284 906 286 962
rect 226 894 286 906
rect 494 1070 554 1082
rect 494 1014 496 1070
rect 552 1014 554 1070
rect 494 962 554 1014
rect 494 906 496 962
rect 552 906 554 962
rect 494 894 554 906
rect 342 832 438 855
rect 296 830 484 832
rect 296 774 308 830
rect 364 774 416 830
rect 472 774 484 830
rect 296 772 484 774
rect 107 616 484 676
rect 272 577 484 616
rect 290 556 484 577
rect 290 555 475 556
rect 154 524 214 536
rect 154 468 156 524
rect 212 500 214 524
rect 566 524 626 536
rect 566 500 568 524
rect 212 468 237 500
rect 154 416 237 468
rect 154 360 156 416
rect 212 384 237 416
rect 543 468 568 500
rect 624 468 626 524
rect 543 416 626 468
rect 543 384 568 416
rect 212 360 214 384
rect 154 348 214 360
rect 566 360 568 384
rect 624 360 626 416
rect 566 348 626 360
rect 296 326 484 328
rect 296 270 308 326
rect 364 270 416 326
rect 472 270 484 326
rect 296 268 484 270
<< via1 >>
rect 308 4098 364 4154
rect 416 4098 472 4154
rect 156 4008 212 4064
rect 156 3900 212 3956
rect 568 4008 624 4064
rect 568 3900 624 3956
rect 308 3594 364 3650
rect 416 3594 472 3650
rect 228 3410 284 3466
rect 228 3302 284 3358
rect 228 3194 284 3250
rect 228 3086 284 3142
rect 228 2978 284 3034
rect 228 2870 284 2926
rect 228 2762 284 2818
rect 228 2654 284 2710
rect 228 2546 284 2602
rect 228 2438 284 2494
rect 228 2330 284 2386
rect 228 2222 284 2278
rect 228 2114 284 2170
rect 228 2006 284 2062
rect 496 3410 552 3466
rect 496 3302 552 3358
rect 496 3194 552 3250
rect 496 3086 552 3142
rect 496 2978 552 3034
rect 496 2870 552 2926
rect 496 2762 552 2818
rect 496 2654 552 2710
rect 496 2546 552 2602
rect 496 2438 552 2494
rect 496 2330 552 2386
rect 496 2222 552 2278
rect 496 2114 552 2170
rect 496 2006 552 2062
rect 308 1822 364 1878
rect 416 1822 472 1878
rect 308 1691 364 1747
rect 416 1691 472 1747
rect 308 1279 364 1335
rect 416 1279 472 1335
rect 308 1146 364 1202
rect 416 1146 472 1202
rect 228 1014 284 1070
rect 228 906 284 962
rect 496 1014 552 1070
rect 496 906 552 962
rect 308 774 364 830
rect 416 774 472 830
rect 156 468 212 524
rect 156 360 212 416
rect 568 468 624 524
rect 568 360 624 416
rect 308 270 364 326
rect 416 270 472 326
<< metal2 >>
rect 296 4154 484 4156
rect 296 4098 308 4154
rect 364 4098 416 4154
rect 472 4098 484 4154
rect 296 4096 484 4098
rect 132 4064 214 4076
rect 132 4008 156 4064
rect 212 4040 214 4064
rect 566 4064 673 4076
rect 566 4040 568 4064
rect 212 4008 568 4040
rect 624 4008 673 4064
rect 132 3956 673 4008
rect 132 3900 156 3956
rect 212 3924 568 3956
rect 212 3900 214 3924
rect 132 3888 214 3900
rect 566 3900 568 3924
rect 624 3900 673 3956
rect 566 3888 673 3900
rect 296 3650 484 3652
rect 296 3594 308 3650
rect 364 3594 416 3650
rect 472 3594 484 3650
rect 296 3592 484 3594
rect 226 3466 286 3478
rect 226 3408 228 3466
rect 284 3408 286 3466
rect 226 3360 286 3408
rect 226 3302 228 3360
rect 284 3302 286 3360
rect 226 3250 286 3302
rect 226 3192 228 3250
rect 284 3192 286 3250
rect 226 3144 286 3192
rect 226 3086 228 3144
rect 284 3086 286 3144
rect 226 3034 286 3086
rect 226 2976 228 3034
rect 284 2976 286 3034
rect 226 2928 286 2976
rect 226 2870 228 2928
rect 284 2870 286 2928
rect 226 2818 286 2870
rect 226 2760 228 2818
rect 284 2760 286 2818
rect 226 2712 286 2760
rect 226 2654 228 2712
rect 284 2654 286 2712
rect 226 2602 286 2654
rect 226 2544 228 2602
rect 284 2544 286 2602
rect 226 2496 286 2544
rect 226 2438 228 2496
rect 284 2438 286 2496
rect 226 2386 286 2438
rect 226 2328 228 2386
rect 284 2328 286 2386
rect 226 2280 286 2328
rect 226 2222 228 2280
rect 284 2222 286 2280
rect 226 2170 286 2222
rect 226 2112 228 2170
rect 284 2112 286 2170
rect 226 2064 286 2112
rect 226 2006 228 2064
rect 284 2006 286 2064
rect 226 1994 286 2006
rect 342 1880 438 3592
rect 494 3466 554 3478
rect 494 3408 496 3466
rect 552 3408 554 3466
rect 494 3360 554 3408
rect 494 3302 496 3360
rect 552 3302 554 3360
rect 494 3250 554 3302
rect 494 3192 496 3250
rect 552 3192 554 3250
rect 494 3144 554 3192
rect 494 3086 496 3144
rect 552 3086 554 3144
rect 494 3034 554 3086
rect 494 2976 496 3034
rect 552 2976 554 3034
rect 494 2928 554 2976
rect 494 2870 496 2928
rect 552 2870 554 2928
rect 494 2818 554 2870
rect 494 2760 496 2818
rect 552 2760 554 2818
rect 494 2712 554 2760
rect 494 2654 496 2712
rect 552 2654 554 2712
rect 494 2602 554 2654
rect 494 2544 496 2602
rect 552 2544 554 2602
rect 494 2496 554 2544
rect 494 2438 496 2496
rect 552 2438 554 2496
rect 494 2386 554 2438
rect 494 2328 496 2386
rect 552 2328 554 2386
rect 494 2280 554 2328
rect 494 2222 496 2280
rect 552 2222 554 2280
rect 494 2170 554 2222
rect 494 2112 496 2170
rect 552 2112 554 2170
rect 494 2064 554 2112
rect 494 2006 496 2064
rect 552 2006 554 2064
rect 494 1994 554 2006
rect 296 1878 484 1880
rect 296 1822 308 1878
rect 364 1822 416 1878
rect 472 1822 484 1878
rect 296 1747 484 1822
rect 296 1691 308 1747
rect 364 1691 416 1747
rect 472 1691 484 1747
rect 296 1689 484 1691
rect 332 1337 448 1689
rect 296 1335 484 1337
rect 296 1279 308 1335
rect 364 1279 416 1335
rect 472 1279 484 1335
rect 296 1202 484 1279
rect 296 1146 308 1202
rect 364 1146 416 1202
rect 472 1146 484 1202
rect 296 1144 484 1146
rect 226 1070 286 1082
rect 226 1012 228 1070
rect 284 1012 286 1070
rect 226 964 286 1012
rect 226 906 228 964
rect 284 906 286 964
rect 226 894 286 906
rect 342 832 438 1144
rect 494 1070 554 1082
rect 494 1012 496 1070
rect 552 1012 554 1070
rect 494 964 554 1012
rect 494 906 496 964
rect 552 906 554 964
rect 494 894 554 906
rect 296 830 484 832
rect 296 774 308 830
rect 364 774 416 830
rect 472 774 484 830
rect 296 772 484 774
rect 333 764 449 772
rect 107 524 214 536
rect 107 468 156 524
rect 212 500 214 524
rect 566 524 648 536
rect 566 500 568 524
rect 212 468 568 500
rect 624 468 648 524
rect 107 416 648 468
rect 107 360 156 416
rect 212 384 568 416
rect 212 360 214 384
rect 107 348 214 360
rect 566 360 568 384
rect 624 360 648 416
rect 566 348 648 360
rect 296 326 484 328
rect 296 270 308 326
rect 364 270 416 326
rect 472 270 484 326
rect 296 268 484 270
<< via2 >>
rect 228 3410 284 3464
rect 228 3408 284 3410
rect 228 3358 284 3360
rect 228 3304 284 3358
rect 228 3194 284 3248
rect 228 3192 284 3194
rect 228 3142 284 3144
rect 228 3088 284 3142
rect 228 2978 284 3032
rect 228 2976 284 2978
rect 228 2926 284 2928
rect 228 2872 284 2926
rect 228 2762 284 2816
rect 228 2760 284 2762
rect 228 2710 284 2712
rect 228 2656 284 2710
rect 228 2546 284 2600
rect 228 2544 284 2546
rect 228 2494 284 2496
rect 228 2440 284 2494
rect 228 2330 284 2384
rect 228 2328 284 2330
rect 228 2278 284 2280
rect 228 2224 284 2278
rect 228 2114 284 2168
rect 228 2112 284 2114
rect 228 2062 284 2064
rect 228 2008 284 2062
rect 496 3410 552 3464
rect 496 3408 552 3410
rect 496 3358 552 3360
rect 496 3304 552 3358
rect 496 3194 552 3248
rect 496 3192 552 3194
rect 496 3142 552 3144
rect 496 3088 552 3142
rect 496 2978 552 3032
rect 496 2976 552 2978
rect 496 2926 552 2928
rect 496 2872 552 2926
rect 496 2762 552 2816
rect 496 2760 552 2762
rect 496 2710 552 2712
rect 496 2656 552 2710
rect 496 2546 552 2600
rect 496 2544 552 2546
rect 496 2494 552 2496
rect 496 2440 552 2494
rect 496 2330 552 2384
rect 496 2328 552 2330
rect 496 2278 552 2280
rect 496 2224 552 2278
rect 496 2114 552 2168
rect 496 2112 552 2114
rect 496 2062 552 2064
rect 496 2008 552 2062
rect 228 1014 284 1068
rect 228 1012 284 1014
rect 228 962 284 964
rect 228 908 284 962
rect 496 1014 552 1068
rect 496 1012 552 1014
rect 496 962 552 964
rect 496 908 552 962
<< metal3 >>
rect 226 3464 286 3478
rect 226 3408 228 3464
rect 284 3408 286 3464
rect 226 3360 286 3408
rect 226 3304 228 3360
rect 284 3304 286 3360
rect 226 3248 286 3304
rect 226 3192 228 3248
rect 284 3192 286 3248
rect 226 3144 286 3192
rect 226 3088 228 3144
rect 284 3088 286 3144
rect 226 3032 286 3088
rect 226 2976 228 3032
rect 284 2976 286 3032
rect 226 2928 286 2976
rect 226 2872 228 2928
rect 284 2872 286 2928
rect 226 2819 286 2872
rect 494 3464 554 3478
rect 494 3408 496 3464
rect 552 3408 554 3464
rect 494 3360 554 3408
rect 494 3304 496 3360
rect 552 3304 554 3360
rect 494 3248 554 3304
rect 494 3192 496 3248
rect 552 3192 554 3248
rect 494 3144 554 3192
rect 494 3088 496 3144
rect 552 3088 554 3144
rect 494 3032 554 3088
rect 494 2976 496 3032
rect 552 2976 554 3032
rect 494 2928 554 2976
rect 494 2872 496 2928
rect 552 2872 554 2928
rect 494 2819 554 2872
rect 132 2816 673 2819
rect 132 2760 228 2816
rect 284 2760 496 2816
rect 552 2760 673 2816
rect 132 2712 673 2760
rect 132 2656 228 2712
rect 284 2656 496 2712
rect 552 2656 673 2712
rect 132 2654 673 2656
rect 226 2600 286 2654
rect 226 2544 228 2600
rect 284 2544 286 2600
rect 226 2496 286 2544
rect 226 2440 228 2496
rect 284 2440 286 2496
rect 226 2384 286 2440
rect 226 2328 228 2384
rect 284 2328 286 2384
rect 226 2280 286 2328
rect 226 2224 228 2280
rect 284 2224 286 2280
rect 226 2168 286 2224
rect 226 2112 228 2168
rect 284 2112 286 2168
rect 226 2064 286 2112
rect 226 2008 228 2064
rect 284 2008 286 2064
rect 226 1994 286 2008
rect 494 2600 554 2654
rect 494 2544 496 2600
rect 552 2544 554 2600
rect 494 2496 554 2544
rect 494 2440 496 2496
rect 552 2440 554 2496
rect 494 2384 554 2440
rect 494 2328 496 2384
rect 552 2328 554 2384
rect 494 2280 554 2328
rect 494 2224 496 2280
rect 552 2224 554 2280
rect 494 2168 554 2224
rect 494 2112 496 2168
rect 552 2112 554 2168
rect 494 2064 554 2112
rect 494 2008 496 2064
rect 552 2008 554 2064
rect 494 1994 554 2008
rect 132 1068 648 1082
rect 132 1012 228 1068
rect 284 1012 496 1068
rect 552 1012 648 1068
rect 132 964 648 1012
rect 132 908 228 964
rect 284 908 496 964
rect 552 908 648 964
rect 132 894 648 908
use nmos_6p0_ZS2JNU  nmos_6p0_ZS2JNU_0
timestamp 1669491903
transform 0 1 390 1 0 3982
box -180 -244 180 244
use nmos_6p0_ZS2JNU  nmos_6p0_ZS2JNU_1
timestamp 1669491903
transform 1 0 390 0 -1 1513
box -180 -244 180 244
use nmos_6p0_ZS2JNU  nmos_6p0_ZS2JNU_2
timestamp 1669491903
transform 0 -1 390 -1 0 442
box -180 -244 180 244
use pmos_6p0_SPFY8K  pmos_6p0_SPFY8K_0
timestamp 1669496281
transform 1 0 390 0 -1 988
box -258 -278 258 278
use pmos_6p0_SPFYFH  pmos_6p0_SPFYFH_0
timestamp 1669496281
transform 1 0 390 0 1 2736
box -258 -978 258 978
<< end >>
