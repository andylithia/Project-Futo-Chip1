magic
tech gf180mcuC
magscale 1 5
timestamp 1669696112
<< obsm1 >>
rect 672 1538 6408 5126
<< metal2 >>
rect 840 0 896 400
rect 2576 0 2632 400
rect 4312 0 4368 400
rect 6048 0 6104 400
<< obsm2 >>
rect 854 430 6394 5115
rect 926 350 2546 430
rect 2662 350 4282 430
rect 4398 350 6018 430
rect 6134 350 6394 430
<< obsm3 >>
rect 1129 1554 6399 5110
<< metal4 >>
rect 1299 1538 1459 5126
rect 2006 1538 2166 5126
rect 2713 1538 2873 5126
rect 3420 1538 3580 5126
rect 4127 1538 4287 5126
rect 4834 1538 4994 5126
rect 5541 1538 5701 5126
rect 6248 1538 6408 5126
<< labels >>
rlabel metal2 s 2576 0 2632 400 6 nbus
port 1 nsew signal bidirectional
rlabel metal2 s 6048 0 6104 400 6 nload
port 2 nsew signal bidirectional
rlabel metal2 s 840 0 896 400 6 pbus
port 3 nsew signal bidirectional
rlabel metal2 s 4312 0 4368 400 6 pload
port 4 nsew signal bidirectional
rlabel metal4 s 1299 1538 1459 5126 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 2713 1538 2873 5126 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 4127 1538 4287 5126 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 5541 1538 5701 5126 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 2006 1538 2166 5126 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 3420 1538 3580 5126 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 4834 1538 4994 5126 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 6248 1538 6408 5126 6 vss
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7000 7000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 125154
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/dlc/runs/22_11_28_23_28/results/signoff/gyrator.magic.gds
string GDS_START 29176
<< end >>

