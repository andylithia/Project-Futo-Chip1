magic
tech gf180mcuC
magscale 1 10
timestamp 1670875428
<< error_s >>
rect 148 963 159 1009
rect 64 871 75 917
rect 232 871 243 917
rect 148 779 159 825
<< metal1 >>
rect -460 1050 -230 1090
rect -460 60 -420 1050
rect -270 60 -230 1050
rect -460 30 -230 60
<< via1 >>
rect -420 60 -270 1050
<< metal2 >>
rect -460 1050 -230 1090
rect -460 60 -420 1050
rect -270 60 -230 1050
rect -460 30 -230 60
use nmos_3p3_BD67EX  nmos_3p3_BD67EX_0
timestamp 1670875428
transform 1 0 182 0 1 894
box -282 -244 282 244
use ppolyf_s_EWZ6SG  ppolyf_s_EWZ6SG_0
timestamp 1670875428
transform 1 0 198 0 1 264
box -258 -324 258 324
<< end >>
