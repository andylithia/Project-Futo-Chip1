* NGSPICE file created from hold_flat.ext - technology: gf180mcuC

.subckt hold_flat Z VDD VSS
X0 a_168_69# Z VSS VSS nmos_6p0 w=0.82u l=0.6u
X1 VDD a_168_69# Z VDD pmos_6p0 w=0.32u l=2u
X2 a_168_69# Z VDD VDD pmos_6p0 w=1.22u l=0.5u
X3 VSS a_168_69# Z VSS nmos_6p0 w=0.32u l=2u
.ends
