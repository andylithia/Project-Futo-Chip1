magic
tech gf180mcuC
magscale 1 5
timestamp 1669696111
<< metal1 >>
rect 672 5109 6328 5126
rect 672 5083 1314 5109
rect 1340 5083 1366 5109
rect 1392 5083 1418 5109
rect 1444 5083 2728 5109
rect 2754 5083 2780 5109
rect 2806 5083 2832 5109
rect 2858 5083 4142 5109
rect 4168 5083 4194 5109
rect 4220 5083 4246 5109
rect 4272 5083 5556 5109
rect 5582 5083 5608 5109
rect 5634 5083 5660 5109
rect 5686 5083 6328 5109
rect 672 5066 6328 5083
rect 672 4717 6408 4734
rect 672 4691 2021 4717
rect 2047 4691 2073 4717
rect 2099 4691 2125 4717
rect 2151 4691 3435 4717
rect 3461 4691 3487 4717
rect 3513 4691 3539 4717
rect 3565 4691 4849 4717
rect 4875 4691 4901 4717
rect 4927 4691 4953 4717
rect 4979 4691 6263 4717
rect 6289 4691 6315 4717
rect 6341 4691 6367 4717
rect 6393 4691 6408 4717
rect 672 4674 6408 4691
rect 2703 4521 2729 4527
rect 2703 4489 2729 4495
rect 2983 4521 3009 4527
rect 2983 4489 3009 4495
rect 3039 4521 3065 4527
rect 3039 4489 3065 4495
rect 2647 4409 2673 4415
rect 2647 4377 2673 4383
rect 672 4325 6328 4342
rect 672 4299 1314 4325
rect 1340 4299 1366 4325
rect 1392 4299 1418 4325
rect 1444 4299 2728 4325
rect 2754 4299 2780 4325
rect 2806 4299 2832 4325
rect 2858 4299 4142 4325
rect 4168 4299 4194 4325
rect 4220 4299 4246 4325
rect 4272 4299 5556 4325
rect 5582 4299 5608 4325
rect 5634 4299 5660 4325
rect 5686 4299 6328 4325
rect 672 4282 6328 4299
rect 2423 4073 2449 4079
rect 2423 4041 2449 4047
rect 2871 4073 2897 4079
rect 2871 4041 2897 4047
rect 3375 4073 3401 4079
rect 3375 4041 3401 4047
rect 3655 4073 3681 4079
rect 3655 4041 3681 4047
rect 2479 4017 2505 4023
rect 2479 3985 2505 3991
rect 2927 4017 2953 4023
rect 2927 3985 2953 3991
rect 3319 4017 3345 4023
rect 3319 3985 3345 3991
rect 3711 4017 3737 4023
rect 3711 3985 3737 3991
rect 672 3933 6408 3950
rect 672 3907 2021 3933
rect 2047 3907 2073 3933
rect 2099 3907 2125 3933
rect 2151 3907 3435 3933
rect 3461 3907 3487 3933
rect 3513 3907 3539 3933
rect 3565 3907 4849 3933
rect 4875 3907 4901 3933
rect 4927 3907 4953 3933
rect 4979 3907 6263 3933
rect 6289 3907 6315 3933
rect 6341 3907 6367 3933
rect 6393 3907 6408 3933
rect 672 3890 6408 3907
rect 1807 3737 1833 3743
rect 1807 3705 1833 3711
rect 2143 3737 2169 3743
rect 2143 3705 2169 3711
rect 2479 3737 2505 3743
rect 2479 3705 2505 3711
rect 2815 3737 2841 3743
rect 2815 3705 2841 3711
rect 3151 3737 3177 3743
rect 3151 3705 3177 3711
rect 3487 3737 3513 3743
rect 3487 3705 3513 3711
rect 4103 3737 4129 3743
rect 4103 3705 4129 3711
rect 1863 3625 1889 3631
rect 1863 3593 1889 3599
rect 2199 3625 2225 3631
rect 2199 3593 2225 3599
rect 2535 3625 2561 3631
rect 2535 3593 2561 3599
rect 2871 3625 2897 3631
rect 2871 3593 2897 3599
rect 3207 3625 3233 3631
rect 3207 3593 3233 3599
rect 3543 3625 3569 3631
rect 3543 3593 3569 3599
rect 4047 3625 4073 3631
rect 4047 3593 4073 3599
rect 672 3541 6328 3558
rect 672 3515 1314 3541
rect 1340 3515 1366 3541
rect 1392 3515 1418 3541
rect 1444 3515 2728 3541
rect 2754 3515 2780 3541
rect 2806 3515 2832 3541
rect 2858 3515 4142 3541
rect 4168 3515 4194 3541
rect 4220 3515 4246 3541
rect 4272 3515 5556 3541
rect 5582 3515 5608 3541
rect 5634 3515 5660 3541
rect 5686 3515 6328 3541
rect 672 3498 6328 3515
rect 1079 3289 1105 3295
rect 1079 3257 1105 3263
rect 1415 3289 1441 3295
rect 1415 3257 1441 3263
rect 1471 3289 1497 3295
rect 1471 3257 1497 3263
rect 1751 3289 1777 3295
rect 1751 3257 1777 3263
rect 2087 3289 2113 3295
rect 2087 3257 2113 3263
rect 2423 3289 2449 3295
rect 2423 3257 2449 3263
rect 2927 3289 2953 3295
rect 2927 3257 2953 3263
rect 3263 3289 3289 3295
rect 3263 3257 3289 3263
rect 3599 3289 3625 3295
rect 3599 3257 3625 3263
rect 3935 3289 3961 3295
rect 3935 3257 3961 3263
rect 4271 3289 4297 3295
rect 4271 3257 4297 3263
rect 4607 3289 4633 3295
rect 4607 3257 4633 3263
rect 4663 3289 4689 3295
rect 4663 3257 4689 3263
rect 1135 3233 1161 3239
rect 1135 3201 1161 3207
rect 1807 3233 1833 3239
rect 1807 3201 1833 3207
rect 2143 3233 2169 3239
rect 2143 3201 2169 3207
rect 2479 3233 2505 3239
rect 2479 3201 2505 3207
rect 2983 3233 3009 3239
rect 2983 3201 3009 3207
rect 3319 3233 3345 3239
rect 3319 3201 3345 3207
rect 3655 3233 3681 3239
rect 3655 3201 3681 3207
rect 3991 3233 4017 3239
rect 3991 3201 4017 3207
rect 4327 3233 4353 3239
rect 4327 3201 4353 3207
rect 672 3149 6408 3166
rect 672 3123 2021 3149
rect 2047 3123 2073 3149
rect 2099 3123 2125 3149
rect 2151 3123 3435 3149
rect 3461 3123 3487 3149
rect 3513 3123 3539 3149
rect 3565 3123 4849 3149
rect 4875 3123 4901 3149
rect 4927 3123 4953 3149
rect 4979 3123 6263 3149
rect 6289 3123 6315 3149
rect 6341 3123 6367 3149
rect 6393 3123 6408 3149
rect 672 3106 6408 3123
rect 1303 3009 1329 3015
rect 1303 2977 1329 2983
rect 3263 3009 3289 3015
rect 3263 2977 3289 2983
rect 3599 3009 3625 3015
rect 3599 2977 3625 2983
rect 4271 3009 4297 3015
rect 4271 2977 4297 2983
rect 4943 3009 4969 3015
rect 4943 2977 4969 2983
rect 911 2953 937 2959
rect 911 2921 937 2927
rect 1583 2953 1609 2959
rect 1583 2921 1609 2927
rect 1919 2953 1945 2959
rect 1919 2921 1945 2927
rect 1975 2953 2001 2959
rect 1975 2921 2001 2927
rect 2255 2953 2281 2959
rect 2255 2921 2281 2927
rect 2591 2953 2617 2959
rect 2591 2921 2617 2927
rect 2927 2953 2953 2959
rect 2927 2921 2953 2927
rect 3935 2953 3961 2959
rect 3935 2921 3961 2927
rect 3991 2953 4017 2959
rect 3991 2921 4017 2927
rect 4887 2953 4913 2959
rect 4887 2921 4913 2927
rect 967 2841 993 2847
rect 967 2809 993 2815
rect 1247 2841 1273 2847
rect 1247 2809 1273 2815
rect 1639 2841 1665 2847
rect 1639 2809 1665 2815
rect 2311 2841 2337 2847
rect 2311 2809 2337 2815
rect 2647 2841 2673 2847
rect 2647 2809 2673 2815
rect 2983 2841 3009 2847
rect 2983 2809 3009 2815
rect 3319 2841 3345 2847
rect 3319 2809 3345 2815
rect 3655 2841 3681 2847
rect 3655 2809 3681 2815
rect 4327 2841 4353 2847
rect 4327 2809 4353 2815
rect 672 2757 6328 2774
rect 672 2731 1314 2757
rect 1340 2731 1366 2757
rect 1392 2731 1418 2757
rect 1444 2731 2728 2757
rect 2754 2731 2780 2757
rect 2806 2731 2832 2757
rect 2858 2731 4142 2757
rect 4168 2731 4194 2757
rect 4220 2731 4246 2757
rect 4272 2731 5556 2757
rect 5582 2731 5608 2757
rect 5634 2731 5660 2757
rect 5686 2731 6328 2757
rect 672 2714 6328 2731
rect 3263 2673 3289 2679
rect 3263 2641 3289 2647
rect 3599 2673 3625 2679
rect 3599 2641 3625 2647
rect 4943 2673 4969 2679
rect 4943 2641 4969 2647
rect 5223 2673 5249 2679
rect 5223 2641 5249 2647
rect 1135 2561 1161 2567
rect 1135 2529 1161 2535
rect 1415 2561 1441 2567
rect 1415 2529 1441 2535
rect 1751 2561 1777 2567
rect 1751 2529 1777 2535
rect 2143 2561 2169 2567
rect 2143 2529 2169 2535
rect 2479 2561 2505 2567
rect 2479 2529 2505 2535
rect 3543 2561 3569 2567
rect 3543 2529 3569 2535
rect 3879 2561 3905 2567
rect 3879 2529 3905 2535
rect 4551 2561 4577 2567
rect 4551 2529 4577 2535
rect 5559 2561 5585 2567
rect 5559 2529 5585 2535
rect 2087 2505 2113 2511
rect 2087 2473 2113 2479
rect 2423 2505 2449 2511
rect 2423 2473 2449 2479
rect 2871 2505 2897 2511
rect 2871 2473 2897 2479
rect 3207 2505 3233 2511
rect 3207 2473 3233 2479
rect 3935 2505 3961 2511
rect 3935 2473 3961 2479
rect 4215 2505 4241 2511
rect 4215 2473 4241 2479
rect 4887 2505 4913 2511
rect 4887 2473 4913 2479
rect 5279 2505 5305 2511
rect 5279 2473 5305 2479
rect 1079 2449 1105 2455
rect 1079 2417 1105 2423
rect 1471 2449 1497 2455
rect 1471 2417 1497 2423
rect 1807 2449 1833 2455
rect 1807 2417 1833 2423
rect 2927 2449 2953 2455
rect 2927 2417 2953 2423
rect 4271 2449 4297 2455
rect 4271 2417 4297 2423
rect 4607 2449 4633 2455
rect 4607 2417 4633 2423
rect 5615 2449 5641 2455
rect 5615 2417 5641 2423
rect 672 2365 6408 2382
rect 672 2339 2021 2365
rect 2047 2339 2073 2365
rect 2099 2339 2125 2365
rect 2151 2339 3435 2365
rect 3461 2339 3487 2365
rect 3513 2339 3539 2365
rect 3565 2339 4849 2365
rect 4875 2339 4901 2365
rect 4927 2339 4953 2365
rect 4979 2339 6263 2365
rect 6289 2339 6315 2365
rect 6341 2339 6367 2365
rect 6393 2339 6408 2365
rect 672 2322 6408 2339
rect 3543 2281 3569 2287
rect 3543 2249 3569 2255
rect 3935 2281 3961 2287
rect 3935 2249 3961 2255
rect 1807 2225 1833 2231
rect 1807 2193 1833 2199
rect 2143 2225 2169 2231
rect 2143 2193 2169 2199
rect 2479 2225 2505 2231
rect 2479 2193 2505 2199
rect 2815 2225 2841 2231
rect 2815 2193 2841 2199
rect 3151 2225 3177 2231
rect 3151 2193 3177 2199
rect 3879 2225 3905 2231
rect 3879 2193 3905 2199
rect 4271 2225 4297 2231
rect 4271 2193 4297 2199
rect 1135 2169 1161 2175
rect 1135 2137 1161 2143
rect 1471 2169 1497 2175
rect 1471 2137 1497 2143
rect 3487 2169 3513 2175
rect 3487 2137 3513 2143
rect 4215 2169 4241 2175
rect 4215 2137 4241 2143
rect 4887 2169 4913 2175
rect 4887 2137 4913 2143
rect 5223 2169 5249 2175
rect 5223 2137 5249 2143
rect 5559 2169 5585 2175
rect 5559 2137 5585 2143
rect 5895 2169 5921 2175
rect 5895 2137 5921 2143
rect 1191 2057 1217 2063
rect 1191 2025 1217 2031
rect 1527 2057 1553 2063
rect 1527 2025 1553 2031
rect 1863 2057 1889 2063
rect 1863 2025 1889 2031
rect 2199 2057 2225 2063
rect 2199 2025 2225 2031
rect 2535 2057 2561 2063
rect 2535 2025 2561 2031
rect 2871 2057 2897 2063
rect 2871 2025 2897 2031
rect 3207 2057 3233 2063
rect 3207 2025 3233 2031
rect 4943 2057 4969 2063
rect 4943 2025 4969 2031
rect 5279 2057 5305 2063
rect 5279 2025 5305 2031
rect 5615 2057 5641 2063
rect 5615 2025 5641 2031
rect 5951 2057 5977 2063
rect 5951 2025 5977 2031
rect 672 1973 6328 1990
rect 672 1947 1314 1973
rect 1340 1947 1366 1973
rect 1392 1947 1418 1973
rect 1444 1947 2728 1973
rect 2754 1947 2780 1973
rect 2806 1947 2832 1973
rect 2858 1947 4142 1973
rect 4168 1947 4194 1973
rect 4220 1947 4246 1973
rect 4272 1947 5556 1973
rect 5582 1947 5608 1973
rect 5634 1947 5660 1973
rect 5686 1947 6328 1973
rect 672 1930 6328 1947
rect 1471 1889 1497 1895
rect 1471 1857 1497 1863
rect 1807 1889 1833 1895
rect 1807 1857 1833 1863
rect 2143 1889 2169 1895
rect 2143 1857 2169 1863
rect 3767 1889 3793 1895
rect 3767 1857 3793 1863
rect 4271 1889 4297 1895
rect 4271 1857 4297 1863
rect 4887 1889 4913 1895
rect 4887 1857 4913 1863
rect 5223 1889 5249 1895
rect 5223 1857 5249 1863
rect 2423 1777 2449 1783
rect 2423 1745 2449 1751
rect 3375 1777 3401 1783
rect 3375 1745 3401 1751
rect 3711 1777 3737 1783
rect 3711 1745 3737 1751
rect 4215 1777 4241 1783
rect 4215 1745 4241 1751
rect 5559 1777 5585 1783
rect 5559 1745 5585 1751
rect 1079 1721 1105 1727
rect 1079 1689 1105 1695
rect 1135 1721 1161 1727
rect 1135 1689 1161 1695
rect 1415 1721 1441 1727
rect 1415 1689 1441 1695
rect 1751 1721 1777 1727
rect 1751 1689 1777 1695
rect 2087 1721 2113 1727
rect 2087 1689 2113 1695
rect 2479 1721 2505 1727
rect 2479 1689 2505 1695
rect 2927 1721 2953 1727
rect 2927 1689 2953 1695
rect 2983 1721 3009 1727
rect 2983 1689 3009 1695
rect 3431 1721 3457 1727
rect 3431 1689 3457 1695
rect 4831 1721 4857 1727
rect 4831 1689 4857 1695
rect 5167 1721 5193 1727
rect 5167 1689 5193 1695
rect 5503 1721 5529 1727
rect 5503 1689 5529 1695
rect 672 1581 6408 1598
rect 672 1555 2021 1581
rect 2047 1555 2073 1581
rect 2099 1555 2125 1581
rect 2151 1555 3435 1581
rect 3461 1555 3487 1581
rect 3513 1555 3539 1581
rect 3565 1555 4849 1581
rect 4875 1555 4901 1581
rect 4927 1555 4953 1581
rect 4979 1555 6263 1581
rect 6289 1555 6315 1581
rect 6341 1555 6367 1581
rect 6393 1555 6408 1581
rect 672 1538 6408 1555
<< via1 >>
rect 1314 5083 1340 5109
rect 1366 5083 1392 5109
rect 1418 5083 1444 5109
rect 2728 5083 2754 5109
rect 2780 5083 2806 5109
rect 2832 5083 2858 5109
rect 4142 5083 4168 5109
rect 4194 5083 4220 5109
rect 4246 5083 4272 5109
rect 5556 5083 5582 5109
rect 5608 5083 5634 5109
rect 5660 5083 5686 5109
rect 2021 4691 2047 4717
rect 2073 4691 2099 4717
rect 2125 4691 2151 4717
rect 3435 4691 3461 4717
rect 3487 4691 3513 4717
rect 3539 4691 3565 4717
rect 4849 4691 4875 4717
rect 4901 4691 4927 4717
rect 4953 4691 4979 4717
rect 6263 4691 6289 4717
rect 6315 4691 6341 4717
rect 6367 4691 6393 4717
rect 2703 4495 2729 4521
rect 2983 4495 3009 4521
rect 3039 4495 3065 4521
rect 2647 4383 2673 4409
rect 1314 4299 1340 4325
rect 1366 4299 1392 4325
rect 1418 4299 1444 4325
rect 2728 4299 2754 4325
rect 2780 4299 2806 4325
rect 2832 4299 2858 4325
rect 4142 4299 4168 4325
rect 4194 4299 4220 4325
rect 4246 4299 4272 4325
rect 5556 4299 5582 4325
rect 5608 4299 5634 4325
rect 5660 4299 5686 4325
rect 2423 4047 2449 4073
rect 2871 4047 2897 4073
rect 3375 4047 3401 4073
rect 3655 4047 3681 4073
rect 2479 3991 2505 4017
rect 2927 3991 2953 4017
rect 3319 3991 3345 4017
rect 3711 3991 3737 4017
rect 2021 3907 2047 3933
rect 2073 3907 2099 3933
rect 2125 3907 2151 3933
rect 3435 3907 3461 3933
rect 3487 3907 3513 3933
rect 3539 3907 3565 3933
rect 4849 3907 4875 3933
rect 4901 3907 4927 3933
rect 4953 3907 4979 3933
rect 6263 3907 6289 3933
rect 6315 3907 6341 3933
rect 6367 3907 6393 3933
rect 1807 3711 1833 3737
rect 2143 3711 2169 3737
rect 2479 3711 2505 3737
rect 2815 3711 2841 3737
rect 3151 3711 3177 3737
rect 3487 3711 3513 3737
rect 4103 3711 4129 3737
rect 1863 3599 1889 3625
rect 2199 3599 2225 3625
rect 2535 3599 2561 3625
rect 2871 3599 2897 3625
rect 3207 3599 3233 3625
rect 3543 3599 3569 3625
rect 4047 3599 4073 3625
rect 1314 3515 1340 3541
rect 1366 3515 1392 3541
rect 1418 3515 1444 3541
rect 2728 3515 2754 3541
rect 2780 3515 2806 3541
rect 2832 3515 2858 3541
rect 4142 3515 4168 3541
rect 4194 3515 4220 3541
rect 4246 3515 4272 3541
rect 5556 3515 5582 3541
rect 5608 3515 5634 3541
rect 5660 3515 5686 3541
rect 1079 3263 1105 3289
rect 1415 3263 1441 3289
rect 1471 3263 1497 3289
rect 1751 3263 1777 3289
rect 2087 3263 2113 3289
rect 2423 3263 2449 3289
rect 2927 3263 2953 3289
rect 3263 3263 3289 3289
rect 3599 3263 3625 3289
rect 3935 3263 3961 3289
rect 4271 3263 4297 3289
rect 4607 3263 4633 3289
rect 4663 3263 4689 3289
rect 1135 3207 1161 3233
rect 1807 3207 1833 3233
rect 2143 3207 2169 3233
rect 2479 3207 2505 3233
rect 2983 3207 3009 3233
rect 3319 3207 3345 3233
rect 3655 3207 3681 3233
rect 3991 3207 4017 3233
rect 4327 3207 4353 3233
rect 2021 3123 2047 3149
rect 2073 3123 2099 3149
rect 2125 3123 2151 3149
rect 3435 3123 3461 3149
rect 3487 3123 3513 3149
rect 3539 3123 3565 3149
rect 4849 3123 4875 3149
rect 4901 3123 4927 3149
rect 4953 3123 4979 3149
rect 6263 3123 6289 3149
rect 6315 3123 6341 3149
rect 6367 3123 6393 3149
rect 1303 2983 1329 3009
rect 3263 2983 3289 3009
rect 3599 2983 3625 3009
rect 4271 2983 4297 3009
rect 4943 2983 4969 3009
rect 911 2927 937 2953
rect 1583 2927 1609 2953
rect 1919 2927 1945 2953
rect 1975 2927 2001 2953
rect 2255 2927 2281 2953
rect 2591 2927 2617 2953
rect 2927 2927 2953 2953
rect 3935 2927 3961 2953
rect 3991 2927 4017 2953
rect 4887 2927 4913 2953
rect 967 2815 993 2841
rect 1247 2815 1273 2841
rect 1639 2815 1665 2841
rect 2311 2815 2337 2841
rect 2647 2815 2673 2841
rect 2983 2815 3009 2841
rect 3319 2815 3345 2841
rect 3655 2815 3681 2841
rect 4327 2815 4353 2841
rect 1314 2731 1340 2757
rect 1366 2731 1392 2757
rect 1418 2731 1444 2757
rect 2728 2731 2754 2757
rect 2780 2731 2806 2757
rect 2832 2731 2858 2757
rect 4142 2731 4168 2757
rect 4194 2731 4220 2757
rect 4246 2731 4272 2757
rect 5556 2731 5582 2757
rect 5608 2731 5634 2757
rect 5660 2731 5686 2757
rect 3263 2647 3289 2673
rect 3599 2647 3625 2673
rect 4943 2647 4969 2673
rect 5223 2647 5249 2673
rect 1135 2535 1161 2561
rect 1415 2535 1441 2561
rect 1751 2535 1777 2561
rect 2143 2535 2169 2561
rect 2479 2535 2505 2561
rect 3543 2535 3569 2561
rect 3879 2535 3905 2561
rect 4551 2535 4577 2561
rect 5559 2535 5585 2561
rect 2087 2479 2113 2505
rect 2423 2479 2449 2505
rect 2871 2479 2897 2505
rect 3207 2479 3233 2505
rect 3935 2479 3961 2505
rect 4215 2479 4241 2505
rect 4887 2479 4913 2505
rect 5279 2479 5305 2505
rect 1079 2423 1105 2449
rect 1471 2423 1497 2449
rect 1807 2423 1833 2449
rect 2927 2423 2953 2449
rect 4271 2423 4297 2449
rect 4607 2423 4633 2449
rect 5615 2423 5641 2449
rect 2021 2339 2047 2365
rect 2073 2339 2099 2365
rect 2125 2339 2151 2365
rect 3435 2339 3461 2365
rect 3487 2339 3513 2365
rect 3539 2339 3565 2365
rect 4849 2339 4875 2365
rect 4901 2339 4927 2365
rect 4953 2339 4979 2365
rect 6263 2339 6289 2365
rect 6315 2339 6341 2365
rect 6367 2339 6393 2365
rect 3543 2255 3569 2281
rect 3935 2255 3961 2281
rect 1807 2199 1833 2225
rect 2143 2199 2169 2225
rect 2479 2199 2505 2225
rect 2815 2199 2841 2225
rect 3151 2199 3177 2225
rect 3879 2199 3905 2225
rect 4271 2199 4297 2225
rect 1135 2143 1161 2169
rect 1471 2143 1497 2169
rect 3487 2143 3513 2169
rect 4215 2143 4241 2169
rect 4887 2143 4913 2169
rect 5223 2143 5249 2169
rect 5559 2143 5585 2169
rect 5895 2143 5921 2169
rect 1191 2031 1217 2057
rect 1527 2031 1553 2057
rect 1863 2031 1889 2057
rect 2199 2031 2225 2057
rect 2535 2031 2561 2057
rect 2871 2031 2897 2057
rect 3207 2031 3233 2057
rect 4943 2031 4969 2057
rect 5279 2031 5305 2057
rect 5615 2031 5641 2057
rect 5951 2031 5977 2057
rect 1314 1947 1340 1973
rect 1366 1947 1392 1973
rect 1418 1947 1444 1973
rect 2728 1947 2754 1973
rect 2780 1947 2806 1973
rect 2832 1947 2858 1973
rect 4142 1947 4168 1973
rect 4194 1947 4220 1973
rect 4246 1947 4272 1973
rect 5556 1947 5582 1973
rect 5608 1947 5634 1973
rect 5660 1947 5686 1973
rect 1471 1863 1497 1889
rect 1807 1863 1833 1889
rect 2143 1863 2169 1889
rect 3767 1863 3793 1889
rect 4271 1863 4297 1889
rect 4887 1863 4913 1889
rect 5223 1863 5249 1889
rect 2423 1751 2449 1777
rect 3375 1751 3401 1777
rect 3711 1751 3737 1777
rect 4215 1751 4241 1777
rect 5559 1751 5585 1777
rect 1079 1695 1105 1721
rect 1135 1695 1161 1721
rect 1415 1695 1441 1721
rect 1751 1695 1777 1721
rect 2087 1695 2113 1721
rect 2479 1695 2505 1721
rect 2927 1695 2953 1721
rect 2983 1695 3009 1721
rect 3431 1695 3457 1721
rect 4831 1695 4857 1721
rect 5167 1695 5193 1721
rect 5503 1695 5529 1721
rect 2021 1555 2047 1581
rect 2073 1555 2099 1581
rect 2125 1555 2151 1581
rect 3435 1555 3461 1581
rect 3487 1555 3513 1581
rect 3539 1555 3565 1581
rect 4849 1555 4875 1581
rect 4901 1555 4927 1581
rect 4953 1555 4979 1581
rect 6263 1555 6289 1581
rect 6315 1555 6341 1581
rect 6367 1555 6393 1581
<< metal2 >>
rect 1313 5110 1445 5115
rect 1341 5082 1365 5110
rect 1393 5082 1417 5110
rect 1313 5077 1445 5082
rect 2727 5110 2859 5115
rect 2755 5082 2779 5110
rect 2807 5082 2831 5110
rect 2727 5077 2859 5082
rect 4141 5110 4273 5115
rect 4169 5082 4193 5110
rect 4221 5082 4245 5110
rect 4141 5077 4273 5082
rect 5555 5110 5687 5115
rect 5583 5082 5607 5110
rect 5635 5082 5659 5110
rect 5555 5077 5687 5082
rect 2020 4718 2152 4723
rect 2048 4690 2072 4718
rect 2100 4690 2124 4718
rect 2020 4685 2152 4690
rect 3434 4718 3566 4723
rect 3462 4690 3486 4718
rect 3514 4690 3538 4718
rect 3434 4685 3566 4690
rect 4848 4718 4980 4723
rect 4876 4690 4900 4718
rect 4928 4690 4952 4718
rect 4848 4685 4980 4690
rect 6262 4718 6394 4723
rect 6290 4690 6314 4718
rect 6342 4690 6366 4718
rect 6262 4685 6394 4690
rect 2702 4522 2730 4527
rect 2982 4522 3010 4527
rect 3038 4522 3066 4527
rect 2702 4521 3066 4522
rect 2702 4495 2703 4521
rect 2729 4495 2983 4521
rect 3009 4495 3039 4521
rect 3065 4495 3066 4521
rect 2702 4494 3066 4495
rect 2702 4489 2730 4494
rect 2646 4409 2674 4415
rect 2646 4383 2647 4409
rect 2673 4383 2674 4409
rect 1313 4326 1445 4331
rect 1341 4298 1365 4326
rect 1393 4298 1417 4326
rect 1313 4293 1445 4298
rect 2422 4073 2450 4079
rect 2422 4047 2423 4073
rect 2449 4047 2450 4073
rect 2422 4018 2450 4047
rect 2020 3934 2152 3939
rect 2048 3906 2072 3934
rect 2100 3906 2124 3934
rect 2020 3901 2152 3906
rect 1806 3737 1834 3743
rect 1806 3711 1807 3737
rect 1833 3711 1834 3737
rect 1313 3542 1445 3547
rect 1341 3514 1365 3542
rect 1393 3514 1417 3542
rect 1313 3509 1445 3514
rect 1078 3290 1106 3295
rect 1302 3290 1330 3295
rect 1078 3289 1162 3290
rect 1078 3263 1079 3289
rect 1105 3263 1162 3289
rect 1078 3262 1162 3263
rect 1078 3257 1106 3262
rect 1134 3233 1162 3262
rect 1134 3207 1135 3233
rect 1161 3207 1162 3233
rect 910 2954 938 2959
rect 910 2953 994 2954
rect 910 2927 911 2953
rect 937 2927 994 2953
rect 910 2926 994 2927
rect 910 2921 938 2926
rect 966 2841 994 2926
rect 966 2815 967 2841
rect 993 2815 994 2841
rect 966 2450 994 2815
rect 1134 2842 1162 3207
rect 1302 3009 1330 3262
rect 1414 3289 1442 3295
rect 1414 3263 1415 3289
rect 1441 3263 1442 3289
rect 1414 3234 1442 3263
rect 1470 3290 1498 3295
rect 1470 3243 1498 3262
rect 1750 3290 1778 3295
rect 1750 3243 1778 3262
rect 1414 3201 1442 3206
rect 1806 3234 1834 3711
rect 2142 3737 2170 3743
rect 2142 3711 2143 3737
rect 2169 3711 2170 3737
rect 1862 3625 1890 3631
rect 1862 3599 1863 3625
rect 1889 3599 1890 3625
rect 1862 3290 1890 3599
rect 2142 3626 2170 3711
rect 1862 3257 1890 3262
rect 2086 3290 2114 3295
rect 2086 3243 2114 3262
rect 1302 2983 1303 3009
rect 1329 2983 1330 3009
rect 1302 2977 1330 2983
rect 1582 2953 1610 2959
rect 1582 2927 1583 2953
rect 1609 2927 1610 2953
rect 1246 2842 1274 2847
rect 1134 2841 1274 2842
rect 1134 2815 1247 2841
rect 1273 2815 1274 2841
rect 1134 2814 1274 2815
rect 1134 2562 1162 2567
rect 1134 2515 1162 2534
rect 1078 2450 1106 2455
rect 1246 2450 1274 2814
rect 1313 2758 1445 2763
rect 1341 2730 1365 2758
rect 1393 2730 1417 2758
rect 1313 2725 1445 2730
rect 1414 2562 1442 2567
rect 1414 2515 1442 2534
rect 1582 2562 1610 2927
rect 1582 2529 1610 2534
rect 1638 2841 1666 2847
rect 1638 2815 1639 2841
rect 1665 2815 1666 2841
rect 966 2449 1274 2450
rect 966 2423 1079 2449
rect 1105 2423 1274 2449
rect 966 2422 1274 2423
rect 1470 2450 1498 2455
rect 1078 2417 1106 2422
rect 1134 2170 1162 2422
rect 1078 1722 1106 1727
rect 1134 1722 1162 2142
rect 1470 2170 1498 2422
rect 1638 2450 1666 2815
rect 1638 2417 1666 2422
rect 1750 2562 1778 2567
rect 1750 2226 1778 2534
rect 1806 2450 1834 3206
rect 2142 3234 2170 3598
rect 2198 3625 2226 3631
rect 2198 3599 2199 3625
rect 2225 3599 2226 3625
rect 2198 3290 2226 3599
rect 2422 3626 2450 3990
rect 2422 3593 2450 3598
rect 2478 4017 2506 4023
rect 2478 3991 2479 4017
rect 2505 3991 2506 4017
rect 2478 3738 2506 3991
rect 2646 3738 2674 4383
rect 2727 4326 2859 4331
rect 2755 4298 2779 4326
rect 2807 4298 2831 4326
rect 2727 4293 2859 4298
rect 2870 4073 2898 4079
rect 2870 4047 2871 4073
rect 2897 4047 2898 4073
rect 2814 3738 2842 3743
rect 2870 3738 2898 4047
rect 2926 4018 2954 4494
rect 2982 4489 3010 4494
rect 3038 4489 3066 4494
rect 4141 4326 4273 4331
rect 4169 4298 4193 4326
rect 4221 4298 4245 4326
rect 4141 4293 4273 4298
rect 5555 4326 5687 4331
rect 5583 4298 5607 4326
rect 5635 4298 5659 4326
rect 5555 4293 5687 4298
rect 3374 4073 3402 4079
rect 3374 4047 3375 4073
rect 3401 4047 3402 4073
rect 2926 3971 2954 3990
rect 3318 4017 3346 4023
rect 3318 3991 3319 4017
rect 3345 3991 3346 4017
rect 2478 3737 2898 3738
rect 2478 3711 2479 3737
rect 2505 3711 2815 3737
rect 2841 3711 2898 3737
rect 2478 3710 2898 3711
rect 3150 3737 3178 3743
rect 3150 3711 3151 3737
rect 3177 3711 3178 3737
rect 2198 3257 2226 3262
rect 2422 3290 2450 3295
rect 2422 3234 2450 3262
rect 2478 3234 2506 3710
rect 2814 3705 2842 3710
rect 2534 3626 2562 3631
rect 2534 3579 2562 3598
rect 2870 3626 2898 3631
rect 2870 3625 2954 3626
rect 2870 3599 2871 3625
rect 2897 3599 2954 3625
rect 2870 3598 2954 3599
rect 2870 3593 2898 3598
rect 2727 3542 2859 3547
rect 2755 3514 2779 3542
rect 2807 3514 2831 3542
rect 2727 3509 2859 3514
rect 2926 3458 2954 3598
rect 2926 3430 3010 3458
rect 2422 3233 2506 3234
rect 2422 3207 2479 3233
rect 2505 3207 2506 3233
rect 2422 3206 2506 3207
rect 2142 3201 2170 3206
rect 2020 3150 2152 3155
rect 2048 3122 2072 3150
rect 2100 3122 2124 3150
rect 2020 3117 2152 3122
rect 1918 2954 1946 2959
rect 1974 2954 2002 2959
rect 1918 2953 1974 2954
rect 1918 2927 1919 2953
rect 1945 2927 1974 2953
rect 1918 2926 1974 2927
rect 1918 2921 1946 2926
rect 1974 2907 2002 2926
rect 2254 2954 2282 2959
rect 2310 2954 2338 2959
rect 2254 2953 2310 2954
rect 2254 2927 2255 2953
rect 2281 2927 2310 2953
rect 2254 2926 2310 2927
rect 2254 2921 2282 2926
rect 2310 2841 2338 2926
rect 2478 2954 2506 3206
rect 2926 3290 2954 3295
rect 2478 2921 2506 2926
rect 2590 2954 2618 2959
rect 2590 2907 2618 2926
rect 2926 2953 2954 3262
rect 2926 2927 2927 2953
rect 2953 2927 2954 2953
rect 2646 2842 2674 2847
rect 2310 2815 2311 2841
rect 2337 2815 2338 2841
rect 2142 2562 2170 2567
rect 2142 2515 2170 2534
rect 2310 2562 2338 2815
rect 2534 2814 2646 2842
rect 2310 2529 2338 2534
rect 2478 2562 2506 2567
rect 2478 2515 2506 2534
rect 2086 2506 2114 2511
rect 2086 2459 2114 2478
rect 2254 2506 2282 2511
rect 1806 2403 1834 2422
rect 2020 2366 2152 2371
rect 2048 2338 2072 2366
rect 2100 2338 2124 2366
rect 2020 2333 2152 2338
rect 1806 2226 1834 2231
rect 2142 2226 2170 2231
rect 1750 2225 2142 2226
rect 1750 2199 1807 2225
rect 1833 2199 2142 2225
rect 1750 2198 2142 2199
rect 1806 2193 1834 2198
rect 2142 2160 2170 2198
rect 1470 2123 1498 2142
rect 1190 2057 1218 2063
rect 1190 2031 1191 2057
rect 1217 2031 1218 2057
rect 1190 1890 1218 2031
rect 1526 2057 1554 2063
rect 1526 2031 1527 2057
rect 1553 2031 1554 2057
rect 1313 1974 1445 1979
rect 1341 1946 1365 1974
rect 1393 1946 1417 1974
rect 1313 1941 1445 1946
rect 1190 1857 1218 1862
rect 1470 1890 1498 1895
rect 1526 1890 1554 2031
rect 1862 2057 1890 2063
rect 1862 2031 1863 2057
rect 1889 2031 1890 2057
rect 1470 1889 1526 1890
rect 1470 1863 1471 1889
rect 1497 1863 1526 1889
rect 1470 1862 1526 1863
rect 1470 1857 1498 1862
rect 1526 1857 1554 1862
rect 1806 1890 1834 1895
rect 1806 1843 1834 1862
rect 1078 1721 1134 1722
rect 1078 1695 1079 1721
rect 1105 1695 1134 1721
rect 1078 1694 1134 1695
rect 1078 1666 1106 1694
rect 854 1638 1106 1666
rect 1134 1656 1162 1694
rect 1414 1722 1442 1727
rect 1414 1675 1442 1694
rect 1750 1722 1778 1727
rect 1750 1675 1778 1694
rect 1862 1722 1890 2031
rect 2198 2057 2226 2063
rect 2198 2031 2199 2057
rect 2225 2031 2226 2057
rect 2198 2002 2226 2031
rect 1862 1689 1890 1694
rect 2086 1974 2226 2002
rect 2086 1722 2114 1974
rect 2254 1946 2282 2478
rect 2422 2506 2450 2511
rect 2422 2459 2450 2478
rect 2534 2338 2562 2814
rect 2646 2776 2674 2814
rect 2727 2758 2859 2763
rect 2755 2730 2779 2758
rect 2807 2730 2831 2758
rect 2727 2725 2859 2730
rect 2926 2562 2954 2927
rect 2982 3234 3010 3430
rect 3150 3290 3178 3711
rect 3150 3257 3178 3262
rect 3206 3626 3234 3631
rect 3318 3626 3346 3991
rect 3374 3738 3402 4047
rect 3654 4073 3682 4079
rect 3654 4047 3655 4073
rect 3681 4047 3682 4073
rect 3434 3934 3566 3939
rect 3462 3906 3486 3934
rect 3514 3906 3538 3934
rect 3434 3901 3566 3906
rect 3486 3738 3514 3743
rect 3374 3737 3514 3738
rect 3374 3711 3487 3737
rect 3513 3711 3514 3737
rect 3374 3710 3514 3711
rect 3206 3625 3346 3626
rect 3206 3599 3207 3625
rect 3233 3599 3346 3625
rect 3206 3598 3346 3599
rect 2982 2842 3010 3206
rect 3206 3234 3234 3598
rect 3262 3290 3290 3295
rect 3262 3243 3290 3262
rect 3486 3290 3514 3710
rect 3542 3626 3570 3631
rect 3654 3626 3682 4047
rect 3710 4018 3738 4023
rect 3710 3971 3738 3990
rect 4848 3934 4980 3939
rect 4876 3906 4900 3934
rect 4928 3906 4952 3934
rect 4848 3901 4980 3906
rect 6262 3934 6394 3939
rect 6290 3906 6314 3934
rect 6342 3906 6366 3934
rect 6262 3901 6394 3906
rect 4102 3738 4130 3743
rect 3542 3625 3682 3626
rect 3542 3599 3543 3625
rect 3569 3599 3682 3625
rect 3542 3598 3682 3599
rect 3710 3737 4130 3738
rect 3710 3711 4103 3737
rect 4129 3711 4130 3737
rect 3710 3710 4130 3711
rect 3542 3593 3570 3598
rect 3486 3257 3514 3262
rect 3598 3289 3626 3598
rect 3598 3263 3599 3289
rect 3625 3263 3626 3289
rect 3206 3201 3234 3206
rect 3318 3234 3346 3239
rect 3318 3187 3346 3206
rect 3598 3234 3626 3263
rect 3654 3234 3682 3239
rect 3626 3233 3682 3234
rect 3626 3207 3655 3233
rect 3681 3207 3682 3233
rect 3626 3206 3682 3207
rect 3598 3201 3626 3206
rect 3654 3201 3682 3206
rect 3434 3150 3566 3155
rect 3462 3122 3486 3150
rect 3514 3122 3538 3150
rect 3434 3117 3566 3122
rect 3710 3066 3738 3710
rect 4102 3705 4130 3710
rect 4046 3625 4074 3631
rect 4046 3599 4047 3625
rect 4073 3599 4074 3625
rect 3598 3038 3738 3066
rect 3934 3289 3962 3295
rect 3934 3263 3935 3289
rect 3961 3263 3962 3289
rect 3934 3234 3962 3263
rect 3990 3234 4018 3239
rect 4046 3234 4074 3599
rect 4141 3542 4273 3547
rect 4169 3514 4193 3542
rect 4221 3514 4245 3542
rect 4141 3509 4273 3514
rect 5555 3542 5687 3547
rect 5583 3514 5607 3542
rect 5635 3514 5659 3542
rect 5555 3509 5687 3514
rect 3934 3233 4074 3234
rect 3934 3207 3991 3233
rect 4017 3207 4074 3233
rect 3934 3206 4074 3207
rect 4270 3289 4298 3295
rect 4270 3263 4271 3289
rect 4297 3263 4298 3289
rect 4270 3234 4298 3263
rect 4606 3289 4634 3295
rect 4606 3263 4607 3289
rect 4633 3263 4634 3289
rect 4326 3234 4354 3239
rect 4270 3233 4354 3234
rect 4270 3207 4327 3233
rect 4353 3207 4354 3233
rect 4270 3206 4354 3207
rect 3262 3010 3290 3015
rect 3598 3010 3626 3038
rect 3262 3009 3626 3010
rect 3262 2983 3263 3009
rect 3289 2983 3599 3009
rect 3625 2983 3626 3009
rect 3262 2982 3626 2983
rect 3262 2977 3290 2982
rect 2982 2795 3010 2814
rect 3262 2842 3290 2847
rect 3318 2842 3346 2847
rect 3290 2841 3346 2842
rect 3290 2815 3319 2841
rect 3345 2815 3346 2841
rect 3290 2814 3346 2815
rect 3262 2673 3290 2814
rect 3318 2809 3346 2814
rect 3262 2647 3263 2673
rect 3289 2647 3290 2673
rect 3262 2641 3290 2647
rect 2478 2310 2562 2338
rect 2870 2506 2898 2511
rect 2478 2226 2506 2310
rect 2142 1918 2282 1946
rect 2422 2198 2478 2226
rect 2142 1890 2170 1918
rect 2142 1824 2170 1862
rect 2422 1777 2450 2198
rect 2478 2179 2506 2198
rect 2814 2226 2842 2231
rect 2870 2226 2898 2478
rect 2814 2225 2898 2226
rect 2814 2199 2815 2225
rect 2841 2199 2898 2225
rect 2814 2198 2898 2199
rect 2926 2449 2954 2534
rect 3542 2561 3570 2982
rect 3598 2977 3626 2982
rect 3934 2954 3962 3206
rect 3990 3201 4018 3206
rect 4270 3010 4298 3206
rect 4326 3201 4354 3206
rect 4270 2963 4298 2982
rect 3990 2954 4018 2959
rect 3878 2953 3990 2954
rect 3878 2927 3935 2953
rect 3961 2927 3990 2953
rect 3878 2926 3990 2927
rect 3542 2535 3543 2561
rect 3569 2535 3570 2561
rect 2926 2423 2927 2449
rect 2953 2423 2954 2449
rect 2814 2193 2842 2198
rect 2534 2058 2562 2063
rect 2422 1751 2423 1777
rect 2449 1751 2450 1777
rect 2422 1745 2450 1751
rect 2478 2057 2562 2058
rect 2478 2031 2535 2057
rect 2561 2031 2562 2057
rect 2478 2030 2562 2031
rect 2086 1675 2114 1694
rect 2478 1722 2506 2030
rect 2534 2025 2562 2030
rect 2870 2058 2898 2063
rect 2926 2058 2954 2423
rect 3150 2506 3178 2511
rect 3150 2225 3178 2478
rect 3150 2199 3151 2225
rect 3177 2199 3178 2225
rect 3150 2193 3178 2199
rect 3206 2505 3234 2511
rect 3206 2479 3207 2505
rect 3233 2479 3234 2505
rect 3206 2058 3234 2479
rect 3374 2506 3402 2511
rect 2870 2057 3346 2058
rect 2870 2031 2871 2057
rect 2897 2031 3207 2057
rect 3233 2031 3346 2057
rect 2870 2030 3346 2031
rect 2870 2025 2898 2030
rect 2727 1974 2859 1979
rect 2755 1946 2779 1974
rect 2807 1946 2831 1974
rect 2727 1941 2859 1946
rect 2478 1675 2506 1694
rect 2926 1722 2954 2030
rect 3206 2025 3234 2030
rect 2982 1722 3010 1727
rect 2926 1721 3010 1722
rect 2926 1695 2927 1721
rect 2953 1695 2983 1721
rect 3009 1695 3010 1721
rect 2926 1694 3010 1695
rect 854 400 882 1638
rect 2020 1582 2152 1587
rect 2048 1554 2072 1582
rect 2100 1554 2124 1582
rect 2020 1549 2152 1554
rect 2590 462 2786 490
rect 2590 400 2618 462
rect 840 0 896 400
rect 2576 0 2632 400
rect 2758 378 2786 462
rect 2926 378 2954 1694
rect 2982 1689 3010 1694
rect 3318 1666 3346 2030
rect 3374 1778 3402 2478
rect 3542 2506 3570 2535
rect 3542 2473 3570 2478
rect 3598 2842 3626 2847
rect 3654 2842 3682 2847
rect 3626 2841 3682 2842
rect 3626 2815 3655 2841
rect 3681 2815 3682 2841
rect 3626 2814 3682 2815
rect 3598 2673 3626 2814
rect 3654 2809 3682 2814
rect 3598 2647 3599 2673
rect 3625 2647 3626 2673
rect 3598 2562 3626 2647
rect 3434 2366 3566 2371
rect 3462 2338 3486 2366
rect 3514 2338 3538 2366
rect 3434 2333 3566 2338
rect 3542 2282 3570 2287
rect 3598 2282 3626 2534
rect 3878 2562 3906 2926
rect 3934 2921 3962 2926
rect 3990 2888 4018 2926
rect 4326 2841 4354 2847
rect 4326 2815 4327 2841
rect 4353 2815 4354 2841
rect 4141 2758 4273 2763
rect 4169 2730 4193 2758
rect 4221 2730 4245 2758
rect 4141 2725 4273 2730
rect 3878 2515 3906 2534
rect 4214 2562 4242 2567
rect 3542 2281 3626 2282
rect 3542 2255 3543 2281
rect 3569 2255 3626 2281
rect 3542 2254 3626 2255
rect 3934 2506 3962 2511
rect 3934 2281 3962 2478
rect 3934 2255 3935 2281
rect 3961 2255 3962 2281
rect 3542 2249 3570 2254
rect 3878 2226 3906 2231
rect 3934 2226 3962 2255
rect 3878 2225 3934 2226
rect 3878 2199 3879 2225
rect 3905 2199 3934 2225
rect 3878 2198 3934 2199
rect 3878 2193 3906 2198
rect 3486 2170 3514 2175
rect 3374 1712 3402 1750
rect 3430 2169 3514 2170
rect 3430 2143 3487 2169
rect 3513 2143 3514 2169
rect 3934 2160 3962 2198
rect 4214 2505 4242 2534
rect 4214 2479 4215 2505
rect 4241 2479 4242 2505
rect 4214 2169 4242 2479
rect 4270 2450 4298 2455
rect 4326 2450 4354 2815
rect 4550 2562 4578 2567
rect 4550 2515 4578 2534
rect 4298 2422 4354 2450
rect 4606 2450 4634 3263
rect 4662 3290 4690 3295
rect 4662 2674 4690 3262
rect 4848 3150 4980 3155
rect 4876 3122 4900 3150
rect 4928 3122 4952 3150
rect 4848 3117 4980 3122
rect 6262 3150 6394 3155
rect 6290 3122 6314 3150
rect 6342 3122 6366 3150
rect 6262 3117 6394 3122
rect 4942 3010 4970 3015
rect 4942 2963 4970 2982
rect 4662 2641 4690 2646
rect 4886 2953 4914 2959
rect 4886 2927 4887 2953
rect 4913 2927 4914 2953
rect 4270 2226 4298 2422
rect 4606 2403 4634 2422
rect 4886 2505 4914 2927
rect 5555 2758 5687 2763
rect 5583 2730 5607 2758
rect 5635 2730 5659 2758
rect 5555 2725 5687 2730
rect 4942 2674 4970 2679
rect 4942 2627 4970 2646
rect 5222 2674 5250 2679
rect 5222 2627 5250 2646
rect 5558 2562 5586 2567
rect 5558 2515 5586 2534
rect 4886 2479 4887 2505
rect 4913 2479 4914 2505
rect 4886 2450 4914 2479
rect 4886 2417 4914 2422
rect 5278 2505 5306 2511
rect 5278 2479 5279 2505
rect 5305 2479 5306 2505
rect 4848 2366 4980 2371
rect 4876 2338 4900 2366
rect 4928 2338 4952 2366
rect 4848 2333 4980 2338
rect 4270 2179 4298 2198
rect 3430 2142 3514 2143
rect 3430 1890 3458 2142
rect 3486 2137 3514 2142
rect 4214 2143 4215 2169
rect 4241 2143 4242 2169
rect 4214 2058 4242 2143
rect 4886 2169 4914 2175
rect 4886 2143 4887 2169
rect 4913 2143 4914 2169
rect 4214 2030 4354 2058
rect 4141 1974 4273 1979
rect 4169 1946 4193 1974
rect 4221 1946 4245 1974
rect 4141 1941 4273 1946
rect 3766 1890 3794 1895
rect 3430 1889 3794 1890
rect 3430 1863 3767 1889
rect 3793 1863 3794 1889
rect 3430 1862 3794 1863
rect 3430 1721 3458 1862
rect 3766 1857 3794 1862
rect 4270 1890 4298 1895
rect 3710 1778 3738 1783
rect 3710 1731 3738 1750
rect 4214 1778 4242 1783
rect 4270 1778 4298 1862
rect 4242 1750 4298 1778
rect 3430 1695 3431 1721
rect 3457 1695 3458 1721
rect 4214 1712 4242 1750
rect 3430 1666 3458 1695
rect 3318 1638 3458 1666
rect 3434 1582 3566 1587
rect 3462 1554 3486 1582
rect 3514 1554 3538 1582
rect 3434 1549 3566 1554
rect 4326 400 4354 2030
rect 4886 1890 4914 2143
rect 5222 2169 5250 2175
rect 5222 2143 5223 2169
rect 5249 2143 5250 2169
rect 4942 2058 4970 2063
rect 4942 1890 4970 2030
rect 4914 1862 4970 1890
rect 5222 1890 5250 2143
rect 5278 2058 5306 2479
rect 5614 2449 5642 2455
rect 5614 2423 5615 2449
rect 5641 2423 5642 2449
rect 5558 2170 5586 2175
rect 5614 2170 5642 2423
rect 6262 2366 6394 2371
rect 6290 2338 6314 2366
rect 6342 2338 6366 2366
rect 6262 2333 6394 2338
rect 5558 2169 5614 2170
rect 5558 2143 5559 2169
rect 5585 2143 5614 2169
rect 5558 2142 5614 2143
rect 5558 2058 5586 2142
rect 5614 2137 5642 2142
rect 5894 2170 5922 2175
rect 5894 2123 5922 2142
rect 5278 1890 5306 2030
rect 5222 1889 5306 1890
rect 5222 1863 5223 1889
rect 5249 1863 5306 1889
rect 5222 1862 5306 1863
rect 5446 2030 5586 2058
rect 5614 2058 5642 2096
rect 5642 2030 5754 2058
rect 4886 1824 4914 1862
rect 5222 1857 5250 1862
rect 4830 1722 4858 1727
rect 4830 1675 4858 1694
rect 5166 1722 5194 1727
rect 5446 1722 5474 2030
rect 5614 2025 5642 2030
rect 5555 1974 5687 1979
rect 5583 1946 5607 1974
rect 5635 1946 5659 1974
rect 5555 1941 5687 1946
rect 5558 1778 5586 1783
rect 5558 1731 5586 1750
rect 5726 1778 5754 2030
rect 5726 1745 5754 1750
rect 5950 2057 5978 2063
rect 5950 2031 5951 2057
rect 5977 2031 5978 2057
rect 5950 1778 5978 2031
rect 5950 1745 5978 1750
rect 6062 1778 6090 1783
rect 5502 1722 5530 1727
rect 5446 1694 5502 1722
rect 5166 1675 5194 1694
rect 5502 1675 5530 1694
rect 4848 1582 4980 1587
rect 4876 1554 4900 1582
rect 4928 1554 4952 1582
rect 4848 1549 4980 1554
rect 6062 400 6090 1750
rect 6262 1582 6394 1587
rect 6290 1554 6314 1582
rect 6342 1554 6366 1582
rect 6262 1549 6394 1554
rect 2758 350 2954 378
rect 4312 0 4368 400
rect 6048 0 6104 400
<< via2 >>
rect 1313 5109 1341 5110
rect 1313 5083 1314 5109
rect 1314 5083 1340 5109
rect 1340 5083 1341 5109
rect 1313 5082 1341 5083
rect 1365 5109 1393 5110
rect 1365 5083 1366 5109
rect 1366 5083 1392 5109
rect 1392 5083 1393 5109
rect 1365 5082 1393 5083
rect 1417 5109 1445 5110
rect 1417 5083 1418 5109
rect 1418 5083 1444 5109
rect 1444 5083 1445 5109
rect 1417 5082 1445 5083
rect 2727 5109 2755 5110
rect 2727 5083 2728 5109
rect 2728 5083 2754 5109
rect 2754 5083 2755 5109
rect 2727 5082 2755 5083
rect 2779 5109 2807 5110
rect 2779 5083 2780 5109
rect 2780 5083 2806 5109
rect 2806 5083 2807 5109
rect 2779 5082 2807 5083
rect 2831 5109 2859 5110
rect 2831 5083 2832 5109
rect 2832 5083 2858 5109
rect 2858 5083 2859 5109
rect 2831 5082 2859 5083
rect 4141 5109 4169 5110
rect 4141 5083 4142 5109
rect 4142 5083 4168 5109
rect 4168 5083 4169 5109
rect 4141 5082 4169 5083
rect 4193 5109 4221 5110
rect 4193 5083 4194 5109
rect 4194 5083 4220 5109
rect 4220 5083 4221 5109
rect 4193 5082 4221 5083
rect 4245 5109 4273 5110
rect 4245 5083 4246 5109
rect 4246 5083 4272 5109
rect 4272 5083 4273 5109
rect 4245 5082 4273 5083
rect 5555 5109 5583 5110
rect 5555 5083 5556 5109
rect 5556 5083 5582 5109
rect 5582 5083 5583 5109
rect 5555 5082 5583 5083
rect 5607 5109 5635 5110
rect 5607 5083 5608 5109
rect 5608 5083 5634 5109
rect 5634 5083 5635 5109
rect 5607 5082 5635 5083
rect 5659 5109 5687 5110
rect 5659 5083 5660 5109
rect 5660 5083 5686 5109
rect 5686 5083 5687 5109
rect 5659 5082 5687 5083
rect 2020 4717 2048 4718
rect 2020 4691 2021 4717
rect 2021 4691 2047 4717
rect 2047 4691 2048 4717
rect 2020 4690 2048 4691
rect 2072 4717 2100 4718
rect 2072 4691 2073 4717
rect 2073 4691 2099 4717
rect 2099 4691 2100 4717
rect 2072 4690 2100 4691
rect 2124 4717 2152 4718
rect 2124 4691 2125 4717
rect 2125 4691 2151 4717
rect 2151 4691 2152 4717
rect 2124 4690 2152 4691
rect 3434 4717 3462 4718
rect 3434 4691 3435 4717
rect 3435 4691 3461 4717
rect 3461 4691 3462 4717
rect 3434 4690 3462 4691
rect 3486 4717 3514 4718
rect 3486 4691 3487 4717
rect 3487 4691 3513 4717
rect 3513 4691 3514 4717
rect 3486 4690 3514 4691
rect 3538 4717 3566 4718
rect 3538 4691 3539 4717
rect 3539 4691 3565 4717
rect 3565 4691 3566 4717
rect 3538 4690 3566 4691
rect 4848 4717 4876 4718
rect 4848 4691 4849 4717
rect 4849 4691 4875 4717
rect 4875 4691 4876 4717
rect 4848 4690 4876 4691
rect 4900 4717 4928 4718
rect 4900 4691 4901 4717
rect 4901 4691 4927 4717
rect 4927 4691 4928 4717
rect 4900 4690 4928 4691
rect 4952 4717 4980 4718
rect 4952 4691 4953 4717
rect 4953 4691 4979 4717
rect 4979 4691 4980 4717
rect 4952 4690 4980 4691
rect 6262 4717 6290 4718
rect 6262 4691 6263 4717
rect 6263 4691 6289 4717
rect 6289 4691 6290 4717
rect 6262 4690 6290 4691
rect 6314 4717 6342 4718
rect 6314 4691 6315 4717
rect 6315 4691 6341 4717
rect 6341 4691 6342 4717
rect 6314 4690 6342 4691
rect 6366 4717 6394 4718
rect 6366 4691 6367 4717
rect 6367 4691 6393 4717
rect 6393 4691 6394 4717
rect 6366 4690 6394 4691
rect 1313 4325 1341 4326
rect 1313 4299 1314 4325
rect 1314 4299 1340 4325
rect 1340 4299 1341 4325
rect 1313 4298 1341 4299
rect 1365 4325 1393 4326
rect 1365 4299 1366 4325
rect 1366 4299 1392 4325
rect 1392 4299 1393 4325
rect 1365 4298 1393 4299
rect 1417 4325 1445 4326
rect 1417 4299 1418 4325
rect 1418 4299 1444 4325
rect 1444 4299 1445 4325
rect 1417 4298 1445 4299
rect 2422 3990 2450 4018
rect 2020 3933 2048 3934
rect 2020 3907 2021 3933
rect 2021 3907 2047 3933
rect 2047 3907 2048 3933
rect 2020 3906 2048 3907
rect 2072 3933 2100 3934
rect 2072 3907 2073 3933
rect 2073 3907 2099 3933
rect 2099 3907 2100 3933
rect 2072 3906 2100 3907
rect 2124 3933 2152 3934
rect 2124 3907 2125 3933
rect 2125 3907 2151 3933
rect 2151 3907 2152 3933
rect 2124 3906 2152 3907
rect 1313 3541 1341 3542
rect 1313 3515 1314 3541
rect 1314 3515 1340 3541
rect 1340 3515 1341 3541
rect 1313 3514 1341 3515
rect 1365 3541 1393 3542
rect 1365 3515 1366 3541
rect 1366 3515 1392 3541
rect 1392 3515 1393 3541
rect 1365 3514 1393 3515
rect 1417 3541 1445 3542
rect 1417 3515 1418 3541
rect 1418 3515 1444 3541
rect 1444 3515 1445 3541
rect 1417 3514 1445 3515
rect 1302 3262 1330 3290
rect 1470 3289 1498 3290
rect 1470 3263 1471 3289
rect 1471 3263 1497 3289
rect 1497 3263 1498 3289
rect 1470 3262 1498 3263
rect 1750 3289 1778 3290
rect 1750 3263 1751 3289
rect 1751 3263 1777 3289
rect 1777 3263 1778 3289
rect 1750 3262 1778 3263
rect 1414 3206 1442 3234
rect 2142 3598 2170 3626
rect 1862 3262 1890 3290
rect 2086 3289 2114 3290
rect 2086 3263 2087 3289
rect 2087 3263 2113 3289
rect 2113 3263 2114 3289
rect 2086 3262 2114 3263
rect 1806 3233 1834 3234
rect 1806 3207 1807 3233
rect 1807 3207 1833 3233
rect 1833 3207 1834 3233
rect 1806 3206 1834 3207
rect 1134 2561 1162 2562
rect 1134 2535 1135 2561
rect 1135 2535 1161 2561
rect 1161 2535 1162 2561
rect 1134 2534 1162 2535
rect 1313 2757 1341 2758
rect 1313 2731 1314 2757
rect 1314 2731 1340 2757
rect 1340 2731 1341 2757
rect 1313 2730 1341 2731
rect 1365 2757 1393 2758
rect 1365 2731 1366 2757
rect 1366 2731 1392 2757
rect 1392 2731 1393 2757
rect 1365 2730 1393 2731
rect 1417 2757 1445 2758
rect 1417 2731 1418 2757
rect 1418 2731 1444 2757
rect 1444 2731 1445 2757
rect 1417 2730 1445 2731
rect 1414 2561 1442 2562
rect 1414 2535 1415 2561
rect 1415 2535 1441 2561
rect 1441 2535 1442 2561
rect 1414 2534 1442 2535
rect 1582 2534 1610 2562
rect 1470 2449 1498 2450
rect 1470 2423 1471 2449
rect 1471 2423 1497 2449
rect 1497 2423 1498 2449
rect 1470 2422 1498 2423
rect 1134 2169 1162 2170
rect 1134 2143 1135 2169
rect 1135 2143 1161 2169
rect 1161 2143 1162 2169
rect 1134 2142 1162 2143
rect 1638 2422 1666 2450
rect 1750 2561 1778 2562
rect 1750 2535 1751 2561
rect 1751 2535 1777 2561
rect 1777 2535 1778 2561
rect 1750 2534 1778 2535
rect 2422 3598 2450 3626
rect 2727 4325 2755 4326
rect 2727 4299 2728 4325
rect 2728 4299 2754 4325
rect 2754 4299 2755 4325
rect 2727 4298 2755 4299
rect 2779 4325 2807 4326
rect 2779 4299 2780 4325
rect 2780 4299 2806 4325
rect 2806 4299 2807 4325
rect 2779 4298 2807 4299
rect 2831 4325 2859 4326
rect 2831 4299 2832 4325
rect 2832 4299 2858 4325
rect 2858 4299 2859 4325
rect 2831 4298 2859 4299
rect 4141 4325 4169 4326
rect 4141 4299 4142 4325
rect 4142 4299 4168 4325
rect 4168 4299 4169 4325
rect 4141 4298 4169 4299
rect 4193 4325 4221 4326
rect 4193 4299 4194 4325
rect 4194 4299 4220 4325
rect 4220 4299 4221 4325
rect 4193 4298 4221 4299
rect 4245 4325 4273 4326
rect 4245 4299 4246 4325
rect 4246 4299 4272 4325
rect 4272 4299 4273 4325
rect 4245 4298 4273 4299
rect 5555 4325 5583 4326
rect 5555 4299 5556 4325
rect 5556 4299 5582 4325
rect 5582 4299 5583 4325
rect 5555 4298 5583 4299
rect 5607 4325 5635 4326
rect 5607 4299 5608 4325
rect 5608 4299 5634 4325
rect 5634 4299 5635 4325
rect 5607 4298 5635 4299
rect 5659 4325 5687 4326
rect 5659 4299 5660 4325
rect 5660 4299 5686 4325
rect 5686 4299 5687 4325
rect 5659 4298 5687 4299
rect 2926 4017 2954 4018
rect 2926 3991 2927 4017
rect 2927 3991 2953 4017
rect 2953 3991 2954 4017
rect 2926 3990 2954 3991
rect 2198 3262 2226 3290
rect 2422 3289 2450 3290
rect 2422 3263 2423 3289
rect 2423 3263 2449 3289
rect 2449 3263 2450 3289
rect 2422 3262 2450 3263
rect 2142 3233 2170 3234
rect 2142 3207 2143 3233
rect 2143 3207 2169 3233
rect 2169 3207 2170 3233
rect 2142 3206 2170 3207
rect 2534 3625 2562 3626
rect 2534 3599 2535 3625
rect 2535 3599 2561 3625
rect 2561 3599 2562 3625
rect 2534 3598 2562 3599
rect 2727 3541 2755 3542
rect 2727 3515 2728 3541
rect 2728 3515 2754 3541
rect 2754 3515 2755 3541
rect 2727 3514 2755 3515
rect 2779 3541 2807 3542
rect 2779 3515 2780 3541
rect 2780 3515 2806 3541
rect 2806 3515 2807 3541
rect 2779 3514 2807 3515
rect 2831 3541 2859 3542
rect 2831 3515 2832 3541
rect 2832 3515 2858 3541
rect 2858 3515 2859 3541
rect 2831 3514 2859 3515
rect 2020 3149 2048 3150
rect 2020 3123 2021 3149
rect 2021 3123 2047 3149
rect 2047 3123 2048 3149
rect 2020 3122 2048 3123
rect 2072 3149 2100 3150
rect 2072 3123 2073 3149
rect 2073 3123 2099 3149
rect 2099 3123 2100 3149
rect 2072 3122 2100 3123
rect 2124 3149 2152 3150
rect 2124 3123 2125 3149
rect 2125 3123 2151 3149
rect 2151 3123 2152 3149
rect 2124 3122 2152 3123
rect 1974 2953 2002 2954
rect 1974 2927 1975 2953
rect 1975 2927 2001 2953
rect 2001 2927 2002 2953
rect 1974 2926 2002 2927
rect 2310 2926 2338 2954
rect 2926 3289 2954 3290
rect 2926 3263 2927 3289
rect 2927 3263 2953 3289
rect 2953 3263 2954 3289
rect 2926 3262 2954 3263
rect 2478 2926 2506 2954
rect 2590 2953 2618 2954
rect 2590 2927 2591 2953
rect 2591 2927 2617 2953
rect 2617 2927 2618 2953
rect 2590 2926 2618 2927
rect 2142 2561 2170 2562
rect 2142 2535 2143 2561
rect 2143 2535 2169 2561
rect 2169 2535 2170 2561
rect 2142 2534 2170 2535
rect 2646 2841 2674 2842
rect 2646 2815 2647 2841
rect 2647 2815 2673 2841
rect 2673 2815 2674 2841
rect 2646 2814 2674 2815
rect 2310 2534 2338 2562
rect 2478 2561 2506 2562
rect 2478 2535 2479 2561
rect 2479 2535 2505 2561
rect 2505 2535 2506 2561
rect 2478 2534 2506 2535
rect 2086 2505 2114 2506
rect 2086 2479 2087 2505
rect 2087 2479 2113 2505
rect 2113 2479 2114 2505
rect 2086 2478 2114 2479
rect 2254 2478 2282 2506
rect 1806 2449 1834 2450
rect 1806 2423 1807 2449
rect 1807 2423 1833 2449
rect 1833 2423 1834 2449
rect 1806 2422 1834 2423
rect 2020 2365 2048 2366
rect 2020 2339 2021 2365
rect 2021 2339 2047 2365
rect 2047 2339 2048 2365
rect 2020 2338 2048 2339
rect 2072 2365 2100 2366
rect 2072 2339 2073 2365
rect 2073 2339 2099 2365
rect 2099 2339 2100 2365
rect 2072 2338 2100 2339
rect 2124 2365 2152 2366
rect 2124 2339 2125 2365
rect 2125 2339 2151 2365
rect 2151 2339 2152 2365
rect 2124 2338 2152 2339
rect 2142 2225 2170 2226
rect 2142 2199 2143 2225
rect 2143 2199 2169 2225
rect 2169 2199 2170 2225
rect 2142 2198 2170 2199
rect 1470 2169 1498 2170
rect 1470 2143 1471 2169
rect 1471 2143 1497 2169
rect 1497 2143 1498 2169
rect 1470 2142 1498 2143
rect 1313 1973 1341 1974
rect 1313 1947 1314 1973
rect 1314 1947 1340 1973
rect 1340 1947 1341 1973
rect 1313 1946 1341 1947
rect 1365 1973 1393 1974
rect 1365 1947 1366 1973
rect 1366 1947 1392 1973
rect 1392 1947 1393 1973
rect 1365 1946 1393 1947
rect 1417 1973 1445 1974
rect 1417 1947 1418 1973
rect 1418 1947 1444 1973
rect 1444 1947 1445 1973
rect 1417 1946 1445 1947
rect 1190 1862 1218 1890
rect 1526 1862 1554 1890
rect 1806 1889 1834 1890
rect 1806 1863 1807 1889
rect 1807 1863 1833 1889
rect 1833 1863 1834 1889
rect 1806 1862 1834 1863
rect 1134 1721 1162 1722
rect 1134 1695 1135 1721
rect 1135 1695 1161 1721
rect 1161 1695 1162 1721
rect 1134 1694 1162 1695
rect 1414 1721 1442 1722
rect 1414 1695 1415 1721
rect 1415 1695 1441 1721
rect 1441 1695 1442 1721
rect 1414 1694 1442 1695
rect 1750 1721 1778 1722
rect 1750 1695 1751 1721
rect 1751 1695 1777 1721
rect 1777 1695 1778 1721
rect 1750 1694 1778 1695
rect 1862 1694 1890 1722
rect 2422 2505 2450 2506
rect 2422 2479 2423 2505
rect 2423 2479 2449 2505
rect 2449 2479 2450 2505
rect 2422 2478 2450 2479
rect 2727 2757 2755 2758
rect 2727 2731 2728 2757
rect 2728 2731 2754 2757
rect 2754 2731 2755 2757
rect 2727 2730 2755 2731
rect 2779 2757 2807 2758
rect 2779 2731 2780 2757
rect 2780 2731 2806 2757
rect 2806 2731 2807 2757
rect 2779 2730 2807 2731
rect 2831 2757 2859 2758
rect 2831 2731 2832 2757
rect 2832 2731 2858 2757
rect 2858 2731 2859 2757
rect 2831 2730 2859 2731
rect 3150 3262 3178 3290
rect 3434 3933 3462 3934
rect 3434 3907 3435 3933
rect 3435 3907 3461 3933
rect 3461 3907 3462 3933
rect 3434 3906 3462 3907
rect 3486 3933 3514 3934
rect 3486 3907 3487 3933
rect 3487 3907 3513 3933
rect 3513 3907 3514 3933
rect 3486 3906 3514 3907
rect 3538 3933 3566 3934
rect 3538 3907 3539 3933
rect 3539 3907 3565 3933
rect 3565 3907 3566 3933
rect 3538 3906 3566 3907
rect 2982 3233 3010 3234
rect 2982 3207 2983 3233
rect 2983 3207 3009 3233
rect 3009 3207 3010 3233
rect 2982 3206 3010 3207
rect 3262 3289 3290 3290
rect 3262 3263 3263 3289
rect 3263 3263 3289 3289
rect 3289 3263 3290 3289
rect 3262 3262 3290 3263
rect 3710 4017 3738 4018
rect 3710 3991 3711 4017
rect 3711 3991 3737 4017
rect 3737 3991 3738 4017
rect 3710 3990 3738 3991
rect 4848 3933 4876 3934
rect 4848 3907 4849 3933
rect 4849 3907 4875 3933
rect 4875 3907 4876 3933
rect 4848 3906 4876 3907
rect 4900 3933 4928 3934
rect 4900 3907 4901 3933
rect 4901 3907 4927 3933
rect 4927 3907 4928 3933
rect 4900 3906 4928 3907
rect 4952 3933 4980 3934
rect 4952 3907 4953 3933
rect 4953 3907 4979 3933
rect 4979 3907 4980 3933
rect 4952 3906 4980 3907
rect 6262 3933 6290 3934
rect 6262 3907 6263 3933
rect 6263 3907 6289 3933
rect 6289 3907 6290 3933
rect 6262 3906 6290 3907
rect 6314 3933 6342 3934
rect 6314 3907 6315 3933
rect 6315 3907 6341 3933
rect 6341 3907 6342 3933
rect 6314 3906 6342 3907
rect 6366 3933 6394 3934
rect 6366 3907 6367 3933
rect 6367 3907 6393 3933
rect 6393 3907 6394 3933
rect 6366 3906 6394 3907
rect 3486 3262 3514 3290
rect 3206 3206 3234 3234
rect 3318 3233 3346 3234
rect 3318 3207 3319 3233
rect 3319 3207 3345 3233
rect 3345 3207 3346 3233
rect 3318 3206 3346 3207
rect 3598 3206 3626 3234
rect 3434 3149 3462 3150
rect 3434 3123 3435 3149
rect 3435 3123 3461 3149
rect 3461 3123 3462 3149
rect 3434 3122 3462 3123
rect 3486 3149 3514 3150
rect 3486 3123 3487 3149
rect 3487 3123 3513 3149
rect 3513 3123 3514 3149
rect 3486 3122 3514 3123
rect 3538 3149 3566 3150
rect 3538 3123 3539 3149
rect 3539 3123 3565 3149
rect 3565 3123 3566 3149
rect 3538 3122 3566 3123
rect 4141 3541 4169 3542
rect 4141 3515 4142 3541
rect 4142 3515 4168 3541
rect 4168 3515 4169 3541
rect 4141 3514 4169 3515
rect 4193 3541 4221 3542
rect 4193 3515 4194 3541
rect 4194 3515 4220 3541
rect 4220 3515 4221 3541
rect 4193 3514 4221 3515
rect 4245 3541 4273 3542
rect 4245 3515 4246 3541
rect 4246 3515 4272 3541
rect 4272 3515 4273 3541
rect 4245 3514 4273 3515
rect 5555 3541 5583 3542
rect 5555 3515 5556 3541
rect 5556 3515 5582 3541
rect 5582 3515 5583 3541
rect 5555 3514 5583 3515
rect 5607 3541 5635 3542
rect 5607 3515 5608 3541
rect 5608 3515 5634 3541
rect 5634 3515 5635 3541
rect 5607 3514 5635 3515
rect 5659 3541 5687 3542
rect 5659 3515 5660 3541
rect 5660 3515 5686 3541
rect 5686 3515 5687 3541
rect 5659 3514 5687 3515
rect 2982 2841 3010 2842
rect 2982 2815 2983 2841
rect 2983 2815 3009 2841
rect 3009 2815 3010 2841
rect 2982 2814 3010 2815
rect 3262 2814 3290 2842
rect 2926 2534 2954 2562
rect 2870 2505 2898 2506
rect 2870 2479 2871 2505
rect 2871 2479 2897 2505
rect 2897 2479 2898 2505
rect 2870 2478 2898 2479
rect 2478 2225 2506 2226
rect 2478 2199 2479 2225
rect 2479 2199 2505 2225
rect 2505 2199 2506 2225
rect 2478 2198 2506 2199
rect 2142 1889 2170 1890
rect 2142 1863 2143 1889
rect 2143 1863 2169 1889
rect 2169 1863 2170 1889
rect 2142 1862 2170 1863
rect 4270 3009 4298 3010
rect 4270 2983 4271 3009
rect 4271 2983 4297 3009
rect 4297 2983 4298 3009
rect 4270 2982 4298 2983
rect 3990 2953 4018 2954
rect 3990 2927 3991 2953
rect 3991 2927 4017 2953
rect 4017 2927 4018 2953
rect 3990 2926 4018 2927
rect 2086 1721 2114 1722
rect 2086 1695 2087 1721
rect 2087 1695 2113 1721
rect 2113 1695 2114 1721
rect 2086 1694 2114 1695
rect 3150 2478 3178 2506
rect 3374 2478 3402 2506
rect 2727 1973 2755 1974
rect 2727 1947 2728 1973
rect 2728 1947 2754 1973
rect 2754 1947 2755 1973
rect 2727 1946 2755 1947
rect 2779 1973 2807 1974
rect 2779 1947 2780 1973
rect 2780 1947 2806 1973
rect 2806 1947 2807 1973
rect 2779 1946 2807 1947
rect 2831 1973 2859 1974
rect 2831 1947 2832 1973
rect 2832 1947 2858 1973
rect 2858 1947 2859 1973
rect 2831 1946 2859 1947
rect 2478 1721 2506 1722
rect 2478 1695 2479 1721
rect 2479 1695 2505 1721
rect 2505 1695 2506 1721
rect 2478 1694 2506 1695
rect 2020 1581 2048 1582
rect 2020 1555 2021 1581
rect 2021 1555 2047 1581
rect 2047 1555 2048 1581
rect 2020 1554 2048 1555
rect 2072 1581 2100 1582
rect 2072 1555 2073 1581
rect 2073 1555 2099 1581
rect 2099 1555 2100 1581
rect 2072 1554 2100 1555
rect 2124 1581 2152 1582
rect 2124 1555 2125 1581
rect 2125 1555 2151 1581
rect 2151 1555 2152 1581
rect 2124 1554 2152 1555
rect 3542 2478 3570 2506
rect 3598 2814 3626 2842
rect 3598 2534 3626 2562
rect 3434 2365 3462 2366
rect 3434 2339 3435 2365
rect 3435 2339 3461 2365
rect 3461 2339 3462 2365
rect 3434 2338 3462 2339
rect 3486 2365 3514 2366
rect 3486 2339 3487 2365
rect 3487 2339 3513 2365
rect 3513 2339 3514 2365
rect 3486 2338 3514 2339
rect 3538 2365 3566 2366
rect 3538 2339 3539 2365
rect 3539 2339 3565 2365
rect 3565 2339 3566 2365
rect 3538 2338 3566 2339
rect 4141 2757 4169 2758
rect 4141 2731 4142 2757
rect 4142 2731 4168 2757
rect 4168 2731 4169 2757
rect 4141 2730 4169 2731
rect 4193 2757 4221 2758
rect 4193 2731 4194 2757
rect 4194 2731 4220 2757
rect 4220 2731 4221 2757
rect 4193 2730 4221 2731
rect 4245 2757 4273 2758
rect 4245 2731 4246 2757
rect 4246 2731 4272 2757
rect 4272 2731 4273 2757
rect 4245 2730 4273 2731
rect 3878 2561 3906 2562
rect 3878 2535 3879 2561
rect 3879 2535 3905 2561
rect 3905 2535 3906 2561
rect 3878 2534 3906 2535
rect 4214 2534 4242 2562
rect 3934 2505 3962 2506
rect 3934 2479 3935 2505
rect 3935 2479 3961 2505
rect 3961 2479 3962 2505
rect 3934 2478 3962 2479
rect 3934 2198 3962 2226
rect 3374 1777 3402 1778
rect 3374 1751 3375 1777
rect 3375 1751 3401 1777
rect 3401 1751 3402 1777
rect 3374 1750 3402 1751
rect 4550 2561 4578 2562
rect 4550 2535 4551 2561
rect 4551 2535 4577 2561
rect 4577 2535 4578 2561
rect 4550 2534 4578 2535
rect 4270 2449 4298 2450
rect 4270 2423 4271 2449
rect 4271 2423 4297 2449
rect 4297 2423 4298 2449
rect 4270 2422 4298 2423
rect 4662 3289 4690 3290
rect 4662 3263 4663 3289
rect 4663 3263 4689 3289
rect 4689 3263 4690 3289
rect 4662 3262 4690 3263
rect 4848 3149 4876 3150
rect 4848 3123 4849 3149
rect 4849 3123 4875 3149
rect 4875 3123 4876 3149
rect 4848 3122 4876 3123
rect 4900 3149 4928 3150
rect 4900 3123 4901 3149
rect 4901 3123 4927 3149
rect 4927 3123 4928 3149
rect 4900 3122 4928 3123
rect 4952 3149 4980 3150
rect 4952 3123 4953 3149
rect 4953 3123 4979 3149
rect 4979 3123 4980 3149
rect 4952 3122 4980 3123
rect 6262 3149 6290 3150
rect 6262 3123 6263 3149
rect 6263 3123 6289 3149
rect 6289 3123 6290 3149
rect 6262 3122 6290 3123
rect 6314 3149 6342 3150
rect 6314 3123 6315 3149
rect 6315 3123 6341 3149
rect 6341 3123 6342 3149
rect 6314 3122 6342 3123
rect 6366 3149 6394 3150
rect 6366 3123 6367 3149
rect 6367 3123 6393 3149
rect 6393 3123 6394 3149
rect 6366 3122 6394 3123
rect 4942 3009 4970 3010
rect 4942 2983 4943 3009
rect 4943 2983 4969 3009
rect 4969 2983 4970 3009
rect 4942 2982 4970 2983
rect 4662 2646 4690 2674
rect 4606 2449 4634 2450
rect 4606 2423 4607 2449
rect 4607 2423 4633 2449
rect 4633 2423 4634 2449
rect 4606 2422 4634 2423
rect 5555 2757 5583 2758
rect 5555 2731 5556 2757
rect 5556 2731 5582 2757
rect 5582 2731 5583 2757
rect 5555 2730 5583 2731
rect 5607 2757 5635 2758
rect 5607 2731 5608 2757
rect 5608 2731 5634 2757
rect 5634 2731 5635 2757
rect 5607 2730 5635 2731
rect 5659 2757 5687 2758
rect 5659 2731 5660 2757
rect 5660 2731 5686 2757
rect 5686 2731 5687 2757
rect 5659 2730 5687 2731
rect 4942 2673 4970 2674
rect 4942 2647 4943 2673
rect 4943 2647 4969 2673
rect 4969 2647 4970 2673
rect 4942 2646 4970 2647
rect 5222 2673 5250 2674
rect 5222 2647 5223 2673
rect 5223 2647 5249 2673
rect 5249 2647 5250 2673
rect 5222 2646 5250 2647
rect 5558 2561 5586 2562
rect 5558 2535 5559 2561
rect 5559 2535 5585 2561
rect 5585 2535 5586 2561
rect 5558 2534 5586 2535
rect 4886 2422 4914 2450
rect 4848 2365 4876 2366
rect 4848 2339 4849 2365
rect 4849 2339 4875 2365
rect 4875 2339 4876 2365
rect 4848 2338 4876 2339
rect 4900 2365 4928 2366
rect 4900 2339 4901 2365
rect 4901 2339 4927 2365
rect 4927 2339 4928 2365
rect 4900 2338 4928 2339
rect 4952 2365 4980 2366
rect 4952 2339 4953 2365
rect 4953 2339 4979 2365
rect 4979 2339 4980 2365
rect 4952 2338 4980 2339
rect 4270 2225 4298 2226
rect 4270 2199 4271 2225
rect 4271 2199 4297 2225
rect 4297 2199 4298 2225
rect 4270 2198 4298 2199
rect 4141 1973 4169 1974
rect 4141 1947 4142 1973
rect 4142 1947 4168 1973
rect 4168 1947 4169 1973
rect 4141 1946 4169 1947
rect 4193 1973 4221 1974
rect 4193 1947 4194 1973
rect 4194 1947 4220 1973
rect 4220 1947 4221 1973
rect 4193 1946 4221 1947
rect 4245 1973 4273 1974
rect 4245 1947 4246 1973
rect 4246 1947 4272 1973
rect 4272 1947 4273 1973
rect 4245 1946 4273 1947
rect 4270 1889 4298 1890
rect 4270 1863 4271 1889
rect 4271 1863 4297 1889
rect 4297 1863 4298 1889
rect 4270 1862 4298 1863
rect 3710 1777 3738 1778
rect 3710 1751 3711 1777
rect 3711 1751 3737 1777
rect 3737 1751 3738 1777
rect 3710 1750 3738 1751
rect 4214 1777 4242 1778
rect 4214 1751 4215 1777
rect 4215 1751 4241 1777
rect 4241 1751 4242 1777
rect 4214 1750 4242 1751
rect 3434 1581 3462 1582
rect 3434 1555 3435 1581
rect 3435 1555 3461 1581
rect 3461 1555 3462 1581
rect 3434 1554 3462 1555
rect 3486 1581 3514 1582
rect 3486 1555 3487 1581
rect 3487 1555 3513 1581
rect 3513 1555 3514 1581
rect 3486 1554 3514 1555
rect 3538 1581 3566 1582
rect 3538 1555 3539 1581
rect 3539 1555 3565 1581
rect 3565 1555 3566 1581
rect 3538 1554 3566 1555
rect 4942 2057 4970 2058
rect 4942 2031 4943 2057
rect 4943 2031 4969 2057
rect 4969 2031 4970 2057
rect 4942 2030 4970 2031
rect 4886 1889 4914 1890
rect 4886 1863 4887 1889
rect 4887 1863 4913 1889
rect 4913 1863 4914 1889
rect 4886 1862 4914 1863
rect 6262 2365 6290 2366
rect 6262 2339 6263 2365
rect 6263 2339 6289 2365
rect 6289 2339 6290 2365
rect 6262 2338 6290 2339
rect 6314 2365 6342 2366
rect 6314 2339 6315 2365
rect 6315 2339 6341 2365
rect 6341 2339 6342 2365
rect 6314 2338 6342 2339
rect 6366 2365 6394 2366
rect 6366 2339 6367 2365
rect 6367 2339 6393 2365
rect 6393 2339 6394 2365
rect 6366 2338 6394 2339
rect 5614 2142 5642 2170
rect 5894 2169 5922 2170
rect 5894 2143 5895 2169
rect 5895 2143 5921 2169
rect 5921 2143 5922 2169
rect 5894 2142 5922 2143
rect 5278 2057 5306 2058
rect 5278 2031 5279 2057
rect 5279 2031 5305 2057
rect 5305 2031 5306 2057
rect 5278 2030 5306 2031
rect 5614 2057 5642 2058
rect 5614 2031 5615 2057
rect 5615 2031 5641 2057
rect 5641 2031 5642 2057
rect 5614 2030 5642 2031
rect 4830 1721 4858 1722
rect 4830 1695 4831 1721
rect 4831 1695 4857 1721
rect 4857 1695 4858 1721
rect 4830 1694 4858 1695
rect 5166 1721 5194 1722
rect 5166 1695 5167 1721
rect 5167 1695 5193 1721
rect 5193 1695 5194 1721
rect 5166 1694 5194 1695
rect 5555 1973 5583 1974
rect 5555 1947 5556 1973
rect 5556 1947 5582 1973
rect 5582 1947 5583 1973
rect 5555 1946 5583 1947
rect 5607 1973 5635 1974
rect 5607 1947 5608 1973
rect 5608 1947 5634 1973
rect 5634 1947 5635 1973
rect 5607 1946 5635 1947
rect 5659 1973 5687 1974
rect 5659 1947 5660 1973
rect 5660 1947 5686 1973
rect 5686 1947 5687 1973
rect 5659 1946 5687 1947
rect 5558 1777 5586 1778
rect 5558 1751 5559 1777
rect 5559 1751 5585 1777
rect 5585 1751 5586 1777
rect 5558 1750 5586 1751
rect 5726 1750 5754 1778
rect 5950 1750 5978 1778
rect 6062 1750 6090 1778
rect 5502 1721 5530 1722
rect 5502 1695 5503 1721
rect 5503 1695 5529 1721
rect 5529 1695 5530 1721
rect 5502 1694 5530 1695
rect 4848 1581 4876 1582
rect 4848 1555 4849 1581
rect 4849 1555 4875 1581
rect 4875 1555 4876 1581
rect 4848 1554 4876 1555
rect 4900 1581 4928 1582
rect 4900 1555 4901 1581
rect 4901 1555 4927 1581
rect 4927 1555 4928 1581
rect 4900 1554 4928 1555
rect 4952 1581 4980 1582
rect 4952 1555 4953 1581
rect 4953 1555 4979 1581
rect 4979 1555 4980 1581
rect 4952 1554 4980 1555
rect 6262 1581 6290 1582
rect 6262 1555 6263 1581
rect 6263 1555 6289 1581
rect 6289 1555 6290 1581
rect 6262 1554 6290 1555
rect 6314 1581 6342 1582
rect 6314 1555 6315 1581
rect 6315 1555 6341 1581
rect 6341 1555 6342 1581
rect 6314 1554 6342 1555
rect 6366 1581 6394 1582
rect 6366 1555 6367 1581
rect 6367 1555 6393 1581
rect 6393 1555 6394 1581
rect 6366 1554 6394 1555
<< metal3 >>
rect 1308 5082 1313 5110
rect 1341 5082 1365 5110
rect 1393 5082 1417 5110
rect 1445 5082 1450 5110
rect 2722 5082 2727 5110
rect 2755 5082 2779 5110
rect 2807 5082 2831 5110
rect 2859 5082 2864 5110
rect 4136 5082 4141 5110
rect 4169 5082 4193 5110
rect 4221 5082 4245 5110
rect 4273 5082 4278 5110
rect 5550 5082 5555 5110
rect 5583 5082 5607 5110
rect 5635 5082 5659 5110
rect 5687 5082 5692 5110
rect 2015 4690 2020 4718
rect 2048 4690 2072 4718
rect 2100 4690 2124 4718
rect 2152 4690 2157 4718
rect 3429 4690 3434 4718
rect 3462 4690 3486 4718
rect 3514 4690 3538 4718
rect 3566 4690 3571 4718
rect 4843 4690 4848 4718
rect 4876 4690 4900 4718
rect 4928 4690 4952 4718
rect 4980 4690 4985 4718
rect 6257 4690 6262 4718
rect 6290 4690 6314 4718
rect 6342 4690 6366 4718
rect 6394 4690 6399 4718
rect 1308 4298 1313 4326
rect 1341 4298 1365 4326
rect 1393 4298 1417 4326
rect 1445 4298 1450 4326
rect 2722 4298 2727 4326
rect 2755 4298 2779 4326
rect 2807 4298 2831 4326
rect 2859 4298 2864 4326
rect 4136 4298 4141 4326
rect 4169 4298 4193 4326
rect 4221 4298 4245 4326
rect 4273 4298 4278 4326
rect 5550 4298 5555 4326
rect 5583 4298 5607 4326
rect 5635 4298 5659 4326
rect 5687 4298 5692 4326
rect 2417 3990 2422 4018
rect 2450 3990 2926 4018
rect 2954 3990 3710 4018
rect 3738 3990 3743 4018
rect 2015 3906 2020 3934
rect 2048 3906 2072 3934
rect 2100 3906 2124 3934
rect 2152 3906 2157 3934
rect 3429 3906 3434 3934
rect 3462 3906 3486 3934
rect 3514 3906 3538 3934
rect 3566 3906 3571 3934
rect 4843 3906 4848 3934
rect 4876 3906 4900 3934
rect 4928 3906 4952 3934
rect 4980 3906 4985 3934
rect 6257 3906 6262 3934
rect 6290 3906 6314 3934
rect 6342 3906 6366 3934
rect 6394 3906 6399 3934
rect 2137 3598 2142 3626
rect 2170 3598 2422 3626
rect 2450 3598 2534 3626
rect 2562 3598 2567 3626
rect 1308 3514 1313 3542
rect 1341 3514 1365 3542
rect 1393 3514 1417 3542
rect 1445 3514 1450 3542
rect 2722 3514 2727 3542
rect 2755 3514 2779 3542
rect 2807 3514 2831 3542
rect 2859 3514 2864 3542
rect 4136 3514 4141 3542
rect 4169 3514 4193 3542
rect 4221 3514 4245 3542
rect 4273 3514 4278 3542
rect 5550 3514 5555 3542
rect 5583 3514 5607 3542
rect 5635 3514 5659 3542
rect 5687 3514 5692 3542
rect 1297 3262 1302 3290
rect 1330 3262 1470 3290
rect 1498 3262 1750 3290
rect 1778 3262 1862 3290
rect 1890 3262 2086 3290
rect 2114 3262 2198 3290
rect 2226 3262 2422 3290
rect 2450 3262 2455 3290
rect 2921 3262 2926 3290
rect 2954 3262 3150 3290
rect 3178 3262 3262 3290
rect 3290 3262 3486 3290
rect 3514 3262 4662 3290
rect 4690 3262 4695 3290
rect 1409 3206 1414 3234
rect 1442 3206 1806 3234
rect 1834 3206 2142 3234
rect 2170 3206 2175 3234
rect 2977 3206 2982 3234
rect 3010 3206 3206 3234
rect 3234 3206 3318 3234
rect 3346 3206 3598 3234
rect 3626 3206 3631 3234
rect 2015 3122 2020 3150
rect 2048 3122 2072 3150
rect 2100 3122 2124 3150
rect 2152 3122 2157 3150
rect 3429 3122 3434 3150
rect 3462 3122 3486 3150
rect 3514 3122 3538 3150
rect 3566 3122 3571 3150
rect 4843 3122 4848 3150
rect 4876 3122 4900 3150
rect 4928 3122 4952 3150
rect 4980 3122 4985 3150
rect 6257 3122 6262 3150
rect 6290 3122 6314 3150
rect 6342 3122 6366 3150
rect 6394 3122 6399 3150
rect 4186 2982 4270 3010
rect 4298 2982 4942 3010
rect 4970 2982 4975 3010
rect 4186 2954 4214 2982
rect 1969 2926 1974 2954
rect 2002 2926 2310 2954
rect 2338 2926 2478 2954
rect 2506 2926 2590 2954
rect 2618 2926 2623 2954
rect 3985 2926 3990 2954
rect 4018 2926 4214 2954
rect 2641 2814 2646 2842
rect 2674 2814 2982 2842
rect 3010 2814 3262 2842
rect 3290 2814 3598 2842
rect 3626 2814 3631 2842
rect 1308 2730 1313 2758
rect 1341 2730 1365 2758
rect 1393 2730 1417 2758
rect 1445 2730 1450 2758
rect 2722 2730 2727 2758
rect 2755 2730 2779 2758
rect 2807 2730 2831 2758
rect 2859 2730 2864 2758
rect 4136 2730 4141 2758
rect 4169 2730 4193 2758
rect 4221 2730 4245 2758
rect 4273 2730 4278 2758
rect 5550 2730 5555 2758
rect 5583 2730 5607 2758
rect 5635 2730 5659 2758
rect 5687 2730 5692 2758
rect 4657 2646 4662 2674
rect 4690 2646 4942 2674
rect 4970 2646 5222 2674
rect 5250 2646 5255 2674
rect 1129 2534 1134 2562
rect 1162 2534 1414 2562
rect 1442 2534 1582 2562
rect 1610 2534 1750 2562
rect 1778 2534 1783 2562
rect 2137 2534 2142 2562
rect 2170 2534 2310 2562
rect 2338 2534 2478 2562
rect 2506 2534 2926 2562
rect 2954 2534 2959 2562
rect 3593 2534 3598 2562
rect 3626 2534 3878 2562
rect 3906 2534 4214 2562
rect 4242 2534 4550 2562
rect 4578 2534 5558 2562
rect 5586 2534 5591 2562
rect 2081 2478 2086 2506
rect 2114 2478 2254 2506
rect 2282 2478 2422 2506
rect 2450 2478 2870 2506
rect 2898 2478 3150 2506
rect 3178 2478 3374 2506
rect 3402 2478 3542 2506
rect 3570 2478 3934 2506
rect 3962 2478 3967 2506
rect 1465 2422 1470 2450
rect 1498 2422 1638 2450
rect 1666 2422 1806 2450
rect 1834 2422 1839 2450
rect 4265 2422 4270 2450
rect 4298 2422 4606 2450
rect 4634 2422 4886 2450
rect 4914 2422 4919 2450
rect 2015 2338 2020 2366
rect 2048 2338 2072 2366
rect 2100 2338 2124 2366
rect 2152 2338 2157 2366
rect 3429 2338 3434 2366
rect 3462 2338 3486 2366
rect 3514 2338 3538 2366
rect 3566 2338 3571 2366
rect 4843 2338 4848 2366
rect 4876 2338 4900 2366
rect 4928 2338 4952 2366
rect 4980 2338 4985 2366
rect 6257 2338 6262 2366
rect 6290 2338 6314 2366
rect 6342 2338 6366 2366
rect 6394 2338 6399 2366
rect 2137 2198 2142 2226
rect 2170 2198 2478 2226
rect 2506 2198 2511 2226
rect 3929 2198 3934 2226
rect 3962 2198 4270 2226
rect 4298 2198 4303 2226
rect 1129 2142 1134 2170
rect 1162 2142 1470 2170
rect 1498 2142 1503 2170
rect 5609 2142 5614 2170
rect 5642 2142 5894 2170
rect 5922 2142 5927 2170
rect 4937 2030 4942 2058
rect 4970 2030 5278 2058
rect 5306 2030 5614 2058
rect 5642 2030 5647 2058
rect 1308 1946 1313 1974
rect 1341 1946 1365 1974
rect 1393 1946 1417 1974
rect 1445 1946 1450 1974
rect 2722 1946 2727 1974
rect 2755 1946 2779 1974
rect 2807 1946 2831 1974
rect 2859 1946 2864 1974
rect 4136 1946 4141 1974
rect 4169 1946 4193 1974
rect 4221 1946 4245 1974
rect 4273 1946 4278 1974
rect 5550 1946 5555 1974
rect 5583 1946 5607 1974
rect 5635 1946 5659 1974
rect 5687 1946 5692 1974
rect 1185 1862 1190 1890
rect 1218 1862 1526 1890
rect 1554 1862 1806 1890
rect 1834 1862 2142 1890
rect 2170 1862 2175 1890
rect 4265 1862 4270 1890
rect 4298 1862 4886 1890
rect 4914 1862 4919 1890
rect 3369 1750 3374 1778
rect 3402 1750 3710 1778
rect 3738 1750 4214 1778
rect 4242 1750 4247 1778
rect 5553 1750 5558 1778
rect 5586 1750 5726 1778
rect 5754 1750 5950 1778
rect 5978 1750 6062 1778
rect 6090 1750 6095 1778
rect 1129 1694 1134 1722
rect 1162 1694 1414 1722
rect 1442 1694 1750 1722
rect 1778 1694 1862 1722
rect 1890 1694 2086 1722
rect 2114 1694 2478 1722
rect 2506 1694 4830 1722
rect 4858 1694 5166 1722
rect 5194 1694 5502 1722
rect 5530 1694 5535 1722
rect 2015 1554 2020 1582
rect 2048 1554 2072 1582
rect 2100 1554 2124 1582
rect 2152 1554 2157 1582
rect 3429 1554 3434 1582
rect 3462 1554 3486 1582
rect 3514 1554 3538 1582
rect 3566 1554 3571 1582
rect 4843 1554 4848 1582
rect 4876 1554 4900 1582
rect 4928 1554 4952 1582
rect 4980 1554 4985 1582
rect 6257 1554 6262 1582
rect 6290 1554 6314 1582
rect 6342 1554 6366 1582
rect 6394 1554 6399 1582
<< via3 >>
rect 1313 5082 1341 5110
rect 1365 5082 1393 5110
rect 1417 5082 1445 5110
rect 2727 5082 2755 5110
rect 2779 5082 2807 5110
rect 2831 5082 2859 5110
rect 4141 5082 4169 5110
rect 4193 5082 4221 5110
rect 4245 5082 4273 5110
rect 5555 5082 5583 5110
rect 5607 5082 5635 5110
rect 5659 5082 5687 5110
rect 2020 4690 2048 4718
rect 2072 4690 2100 4718
rect 2124 4690 2152 4718
rect 3434 4690 3462 4718
rect 3486 4690 3514 4718
rect 3538 4690 3566 4718
rect 4848 4690 4876 4718
rect 4900 4690 4928 4718
rect 4952 4690 4980 4718
rect 6262 4690 6290 4718
rect 6314 4690 6342 4718
rect 6366 4690 6394 4718
rect 1313 4298 1341 4326
rect 1365 4298 1393 4326
rect 1417 4298 1445 4326
rect 2727 4298 2755 4326
rect 2779 4298 2807 4326
rect 2831 4298 2859 4326
rect 4141 4298 4169 4326
rect 4193 4298 4221 4326
rect 4245 4298 4273 4326
rect 5555 4298 5583 4326
rect 5607 4298 5635 4326
rect 5659 4298 5687 4326
rect 2020 3906 2048 3934
rect 2072 3906 2100 3934
rect 2124 3906 2152 3934
rect 3434 3906 3462 3934
rect 3486 3906 3514 3934
rect 3538 3906 3566 3934
rect 4848 3906 4876 3934
rect 4900 3906 4928 3934
rect 4952 3906 4980 3934
rect 6262 3906 6290 3934
rect 6314 3906 6342 3934
rect 6366 3906 6394 3934
rect 1313 3514 1341 3542
rect 1365 3514 1393 3542
rect 1417 3514 1445 3542
rect 2727 3514 2755 3542
rect 2779 3514 2807 3542
rect 2831 3514 2859 3542
rect 4141 3514 4169 3542
rect 4193 3514 4221 3542
rect 4245 3514 4273 3542
rect 5555 3514 5583 3542
rect 5607 3514 5635 3542
rect 5659 3514 5687 3542
rect 2020 3122 2048 3150
rect 2072 3122 2100 3150
rect 2124 3122 2152 3150
rect 3434 3122 3462 3150
rect 3486 3122 3514 3150
rect 3538 3122 3566 3150
rect 4848 3122 4876 3150
rect 4900 3122 4928 3150
rect 4952 3122 4980 3150
rect 6262 3122 6290 3150
rect 6314 3122 6342 3150
rect 6366 3122 6394 3150
rect 1313 2730 1341 2758
rect 1365 2730 1393 2758
rect 1417 2730 1445 2758
rect 2727 2730 2755 2758
rect 2779 2730 2807 2758
rect 2831 2730 2859 2758
rect 4141 2730 4169 2758
rect 4193 2730 4221 2758
rect 4245 2730 4273 2758
rect 5555 2730 5583 2758
rect 5607 2730 5635 2758
rect 5659 2730 5687 2758
rect 2020 2338 2048 2366
rect 2072 2338 2100 2366
rect 2124 2338 2152 2366
rect 3434 2338 3462 2366
rect 3486 2338 3514 2366
rect 3538 2338 3566 2366
rect 4848 2338 4876 2366
rect 4900 2338 4928 2366
rect 4952 2338 4980 2366
rect 6262 2338 6290 2366
rect 6314 2338 6342 2366
rect 6366 2338 6394 2366
rect 1313 1946 1341 1974
rect 1365 1946 1393 1974
rect 1417 1946 1445 1974
rect 2727 1946 2755 1974
rect 2779 1946 2807 1974
rect 2831 1946 2859 1974
rect 4141 1946 4169 1974
rect 4193 1946 4221 1974
rect 4245 1946 4273 1974
rect 5555 1946 5583 1974
rect 5607 1946 5635 1974
rect 5659 1946 5687 1974
rect 2020 1554 2048 1582
rect 2072 1554 2100 1582
rect 2124 1554 2152 1582
rect 3434 1554 3462 1582
rect 3486 1554 3514 1582
rect 3538 1554 3566 1582
rect 4848 1554 4876 1582
rect 4900 1554 4928 1582
rect 4952 1554 4980 1582
rect 6262 1554 6290 1582
rect 6314 1554 6342 1582
rect 6366 1554 6394 1582
<< metal4 >>
rect 1299 5110 1459 5126
rect 1299 5082 1313 5110
rect 1341 5082 1365 5110
rect 1393 5082 1417 5110
rect 1445 5082 1459 5110
rect 1299 4326 1459 5082
rect 1299 4298 1313 4326
rect 1341 4298 1365 4326
rect 1393 4298 1417 4326
rect 1445 4298 1459 4326
rect 1299 3542 1459 4298
rect 1299 3514 1313 3542
rect 1341 3514 1365 3542
rect 1393 3514 1417 3542
rect 1445 3514 1459 3542
rect 1299 2758 1459 3514
rect 1299 2730 1313 2758
rect 1341 2730 1365 2758
rect 1393 2730 1417 2758
rect 1445 2730 1459 2758
rect 1299 1974 1459 2730
rect 1299 1946 1313 1974
rect 1341 1946 1365 1974
rect 1393 1946 1417 1974
rect 1445 1946 1459 1974
rect 1299 1538 1459 1946
rect 2006 4718 2166 5126
rect 2006 4690 2020 4718
rect 2048 4690 2072 4718
rect 2100 4690 2124 4718
rect 2152 4690 2166 4718
rect 2006 3934 2166 4690
rect 2006 3906 2020 3934
rect 2048 3906 2072 3934
rect 2100 3906 2124 3934
rect 2152 3906 2166 3934
rect 2006 3150 2166 3906
rect 2006 3122 2020 3150
rect 2048 3122 2072 3150
rect 2100 3122 2124 3150
rect 2152 3122 2166 3150
rect 2006 2366 2166 3122
rect 2006 2338 2020 2366
rect 2048 2338 2072 2366
rect 2100 2338 2124 2366
rect 2152 2338 2166 2366
rect 2006 1582 2166 2338
rect 2006 1554 2020 1582
rect 2048 1554 2072 1582
rect 2100 1554 2124 1582
rect 2152 1554 2166 1582
rect 2006 1538 2166 1554
rect 2713 5110 2873 5126
rect 2713 5082 2727 5110
rect 2755 5082 2779 5110
rect 2807 5082 2831 5110
rect 2859 5082 2873 5110
rect 2713 4326 2873 5082
rect 2713 4298 2727 4326
rect 2755 4298 2779 4326
rect 2807 4298 2831 4326
rect 2859 4298 2873 4326
rect 2713 3542 2873 4298
rect 2713 3514 2727 3542
rect 2755 3514 2779 3542
rect 2807 3514 2831 3542
rect 2859 3514 2873 3542
rect 2713 2758 2873 3514
rect 2713 2730 2727 2758
rect 2755 2730 2779 2758
rect 2807 2730 2831 2758
rect 2859 2730 2873 2758
rect 2713 1974 2873 2730
rect 2713 1946 2727 1974
rect 2755 1946 2779 1974
rect 2807 1946 2831 1974
rect 2859 1946 2873 1974
rect 2713 1538 2873 1946
rect 3420 4718 3580 5126
rect 3420 4690 3434 4718
rect 3462 4690 3486 4718
rect 3514 4690 3538 4718
rect 3566 4690 3580 4718
rect 3420 3934 3580 4690
rect 3420 3906 3434 3934
rect 3462 3906 3486 3934
rect 3514 3906 3538 3934
rect 3566 3906 3580 3934
rect 3420 3150 3580 3906
rect 3420 3122 3434 3150
rect 3462 3122 3486 3150
rect 3514 3122 3538 3150
rect 3566 3122 3580 3150
rect 3420 2366 3580 3122
rect 3420 2338 3434 2366
rect 3462 2338 3486 2366
rect 3514 2338 3538 2366
rect 3566 2338 3580 2366
rect 3420 1582 3580 2338
rect 3420 1554 3434 1582
rect 3462 1554 3486 1582
rect 3514 1554 3538 1582
rect 3566 1554 3580 1582
rect 3420 1538 3580 1554
rect 4127 5110 4287 5126
rect 4127 5082 4141 5110
rect 4169 5082 4193 5110
rect 4221 5082 4245 5110
rect 4273 5082 4287 5110
rect 4127 4326 4287 5082
rect 4127 4298 4141 4326
rect 4169 4298 4193 4326
rect 4221 4298 4245 4326
rect 4273 4298 4287 4326
rect 4127 3542 4287 4298
rect 4127 3514 4141 3542
rect 4169 3514 4193 3542
rect 4221 3514 4245 3542
rect 4273 3514 4287 3542
rect 4127 2758 4287 3514
rect 4127 2730 4141 2758
rect 4169 2730 4193 2758
rect 4221 2730 4245 2758
rect 4273 2730 4287 2758
rect 4127 1974 4287 2730
rect 4127 1946 4141 1974
rect 4169 1946 4193 1974
rect 4221 1946 4245 1974
rect 4273 1946 4287 1974
rect 4127 1538 4287 1946
rect 4834 4718 4994 5126
rect 4834 4690 4848 4718
rect 4876 4690 4900 4718
rect 4928 4690 4952 4718
rect 4980 4690 4994 4718
rect 4834 3934 4994 4690
rect 4834 3906 4848 3934
rect 4876 3906 4900 3934
rect 4928 3906 4952 3934
rect 4980 3906 4994 3934
rect 4834 3150 4994 3906
rect 4834 3122 4848 3150
rect 4876 3122 4900 3150
rect 4928 3122 4952 3150
rect 4980 3122 4994 3150
rect 4834 2366 4994 3122
rect 4834 2338 4848 2366
rect 4876 2338 4900 2366
rect 4928 2338 4952 2366
rect 4980 2338 4994 2366
rect 4834 1582 4994 2338
rect 4834 1554 4848 1582
rect 4876 1554 4900 1582
rect 4928 1554 4952 1582
rect 4980 1554 4994 1582
rect 4834 1538 4994 1554
rect 5541 5110 5701 5126
rect 5541 5082 5555 5110
rect 5583 5082 5607 5110
rect 5635 5082 5659 5110
rect 5687 5082 5701 5110
rect 5541 4326 5701 5082
rect 5541 4298 5555 4326
rect 5583 4298 5607 4326
rect 5635 4298 5659 4326
rect 5687 4298 5701 4326
rect 5541 3542 5701 4298
rect 5541 3514 5555 3542
rect 5583 3514 5607 3542
rect 5635 3514 5659 3542
rect 5687 3514 5701 3542
rect 5541 2758 5701 3514
rect 5541 2730 5555 2758
rect 5583 2730 5607 2758
rect 5635 2730 5659 2758
rect 5687 2730 5701 2758
rect 5541 1974 5701 2730
rect 5541 1946 5555 1974
rect 5583 1946 5607 1974
rect 5635 1946 5659 1974
rect 5687 1946 5701 1974
rect 5541 1538 5701 1946
rect 6248 4718 6408 5126
rect 6248 4690 6262 4718
rect 6290 4690 6314 4718
rect 6342 4690 6366 4718
rect 6394 4690 6408 4718
rect 6248 3934 6408 4690
rect 6248 3906 6262 3934
rect 6290 3906 6314 3934
rect 6342 3906 6366 3934
rect 6394 3906 6408 3934
rect 6248 3150 6408 3906
rect 6248 3122 6262 3150
rect 6290 3122 6314 3150
rect 6342 3122 6366 3150
rect 6394 3122 6408 3150
rect 6248 2366 6408 3122
rect 6248 2338 6262 2366
rect 6290 2338 6314 2366
rect 6342 2338 6366 2366
rect 6394 2338 6408 2366
rect 6248 1582 6408 2338
rect 6248 1554 6262 1582
rect 6290 1554 6314 1582
rect 6342 1554 6366 1582
rect 6394 1554 6408 1582
rect 6248 1538 6408 1554
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1232 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16
timestamp 1667941163
transform 1 0 1568 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22
timestamp 1667941163
transform 1 0 1904 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28
timestamp 1667941163
transform 1 0 2240 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43
timestamp 1667941163
transform 1 0 3080 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51
timestamp 1667941163
transform 1 0 3528 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57
timestamp 1667941163
transform 1 0 3864 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61
timestamp 1667941163
transform 1 0 4088 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66
timestamp 1667941163
transform 1 0 4368 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77
timestamp 1667941163
transform 1 0 4984 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83
timestamp 1667941163
transform 1 0 5320 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5656 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97
timestamp 1667941163
transform 1 0 6104 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1667941163
transform 1 0 784 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_6
timestamp 1667941163
transform 1 0 1008 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_11
timestamp 1667941163
transform 1 0 1288 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_17
timestamp 1667941163
transform 1 0 1624 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_23
timestamp 1667941163
transform 1 0 1960 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_29
timestamp 1667941163
transform 1 0 2296 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_35
timestamp 1667941163
transform 1 0 2632 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_41
timestamp 1667941163
transform 1 0 2968 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_47
timestamp 1667941163
transform 1 0 3304 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_53
timestamp 1667941163
transform 1 0 3640 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 3752 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_60
timestamp 1667941163
transform 1 0 4032 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_78
timestamp 1667941163
transform 1 0 5040 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_84
timestamp 1667941163
transform 1 0 5376 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_90
timestamp 1667941163
transform 1 0 5712 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_96
timestamp 1667941163
transform 1 0 6048 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_98
timestamp 1667941163
transform 1 0 6160 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_10
timestamp 1667941163
transform 1 0 1232 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_16
timestamp 1667941163
transform 1 0 1568 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_22
timestamp 1667941163
transform 1 0 1904 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_28
timestamp 1667941163
transform 1 0 2240 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_42
timestamp 1667941163
transform 1 0 3024 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_48
timestamp 1667941163
transform 1 0 3360 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_54
timestamp 1667941163
transform 1 0 3696 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_60
timestamp 1667941163
transform 1 0 4032 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_66
timestamp 1667941163
transform 1 0 4368 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_72
timestamp 1667941163
transform 1 0 4704 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_78
timestamp 1667941163
transform 1 0 5040 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_84
timestamp 1667941163
transform 1 0 5376 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_90
timestamp 1667941163
transform 1 0 5712 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_98
timestamp 1667941163
transform 1 0 6160 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_7
timestamp 1667941163
transform 1 0 1064 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_13
timestamp 1667941163
transform 1 0 1400 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_19
timestamp 1667941163
transform 1 0 1736 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_25
timestamp 1667941163
transform 1 0 2072 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_31
timestamp 1667941163
transform 1 0 2408 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_37
timestamp 1667941163
transform 1 0 2744 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_43
timestamp 1667941163
transform 1 0 3080 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_49
timestamp 1667941163
transform 1 0 3416 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_55
timestamp 1667941163
transform 1 0 3752 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_61
timestamp 1667941163
transform 1 0 4088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_67
timestamp 1667941163
transform 1 0 4424 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_78 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5040 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_94
timestamp 1667941163
transform 1 0 5936 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_98
timestamp 1667941163
transform 1 0 6160 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_10
timestamp 1667941163
transform 1 0 1232 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_16
timestamp 1667941163
transform 1 0 1568 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_22
timestamp 1667941163
transform 1 0 1904 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_28
timestamp 1667941163
transform 1 0 2240 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_43
timestamp 1667941163
transform 1 0 3080 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_49
timestamp 1667941163
transform 1 0 3416 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_55
timestamp 1667941163
transform 1 0 3752 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_61
timestamp 1667941163
transform 1 0 4088 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_67
timestamp 1667941163
transform 1 0 4424 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_73
timestamp 1667941163
transform 1 0 4760 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_89
timestamp 1667941163
transform 1 0 5656 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_97
timestamp 1667941163
transform 1 0 6104 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_18
timestamp 1667941163
transform 1 0 1680 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_23
timestamp 1667941163
transform 1 0 1960 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_29
timestamp 1667941163
transform 1 0 2296 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_35
timestamp 1667941163
transform 1 0 2632 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_41
timestamp 1667941163
transform 1 0 2968 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_47
timestamp 1667941163
transform 1 0 3304 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_53
timestamp 1667941163
transform 1 0 3640 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 3864 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_63
timestamp 1667941163
transform 1 0 4200 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_89
timestamp 1667941163
transform 1 0 5656 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_97
timestamp 1667941163
transform 1 0 6104 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_18
timestamp 1667941163
transform 1 0 1680 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_26
timestamp 1667941163
transform 1 0 2128 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_42
timestamp 1667941163
transform 1 0 3024 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_50
timestamp 1667941163
transform 1 0 3472 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_56 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 3808 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_88
timestamp 1667941163
transform 1 0 5600 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_96
timestamp 1667941163
transform 1 0 6048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_98
timestamp 1667941163
transform 1 0 6160 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1667941163
transform 1 0 784 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_38
timestamp 1667941163
transform 1 0 2800 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_44
timestamp 1667941163
transform 1 0 3136 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_60
timestamp 1667941163
transform 1 0 4032 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_68
timestamp 1667941163
transform 1 0 4480 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 4592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1667941163
transform 1 0 4760 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_89
timestamp 1667941163
transform 1 0 5656 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_97
timestamp 1667941163
transform 1 0 6104 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1667941163
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1667941163
transform 1 0 2744 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_69
timestamp 1667941163
transform 1 0 4536 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_72
timestamp 1667941163
transform 1 0 4704 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_88
timestamp 1667941163
transform 1 0 5600 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_96
timestamp 1667941163
transform 1 0 6048 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_98
timestamp 1667941163
transform 1 0 6160 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 6328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 6328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 6328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 6328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 6328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 6328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 6328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 6328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 6328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_23
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1667941163
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1667941163
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1667941163
transform 1 0 4592 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[0\].fbn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 4144 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 3864 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 3808 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 3864 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 4816 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 4200 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 5152 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 3528 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 5096 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 3416 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 5824 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 2744 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 1344 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 3136 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 5488 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 2856 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 4760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 3416 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 1680 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 3192 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 1064 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 2520 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 2016 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 2856 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 5432 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 3080 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 1400 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_T\[9\].thrup
timestamp 1667941163
transform -1 0 3472 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 3808 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 3192 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 4480 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 4816 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 4144 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 3472 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 4144 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[3\].crossp
timestamp 1667941163
transform -1 0 4200 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 4200 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_f.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 3528 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 2352 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[0\].fbp
timestamp 1667941163
transform -1 0 3136 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 1848 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 1008 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 2184 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 1008 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 2856 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 840 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 4816 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 1736 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 2800 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 5488 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[2\].thrun
timestamp 1667941163
transform -1 0 5376 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 1680 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 3080 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 2408 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 2352 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 1512 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 4536 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 1344 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 2744 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 3584 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 3640 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 2352 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 2016 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[8\].thrup
timestamp 1667941163
transform -1 0 1232 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 3304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 2072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 2352 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 2800 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[1\].crossn
timestamp 1667941163
transform -1 0 2800 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[1\].crossp
timestamp 1667941163
transform -1 0 1400 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 1736 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 1680 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 2072 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 2016 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_r.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 2408 0 -1 3920
box -43 -43 267 435
<< labels >>
flabel metal2 s 2576 0 2632 400 0 FreeSans 224 90 0 0 nbus
port 0 nsew signal bidirectional
flabel metal2 s 6048 0 6104 400 0 FreeSans 224 90 0 0 nload
port 1 nsew signal bidirectional
flabel metal2 s 840 0 896 400 0 FreeSans 224 90 0 0 pbus
port 2 nsew signal bidirectional
flabel metal2 s 4312 0 4368 400 0 FreeSans 224 90 0 0 pload
port 3 nsew signal bidirectional
flabel metal4 s 1299 1538 1459 5126 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 2713 1538 2873 5126 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 4127 1538 4287 5126 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 5541 1538 5701 5126 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 2006 1538 2166 5126 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 3420 1538 3580 5126 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 4834 1538 4994 5126 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 6248 1538 6408 5126 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
rlabel metal1 3500 5096 3500 5096 0 vdd
rlabel via1 3540 4704 3540 4704 0 vss
rlabel metal2 2940 1036 2940 1036 0 nbus
rlabel metal2 3612 3024 3612 3024 0 nload
rlabel metal2 1092 1680 1092 1680 0 pbus
rlabel metal3 1288 2548 1288 2548 0 pload
<< properties >>
string FIXED_BBOX 0 0 7000 7000
<< end >>
