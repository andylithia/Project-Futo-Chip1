module caparray_s2 (cap_series_gygyn,
    cap_series_gygyp,
    cap_series_gyn,
    cap_series_gyp,
    cap_shunt_gyn,
    cap_shunt_gyp,
    cap_shunt_n,
    cap_shunt_p,
    vdd,
    vss,
    tune_series_gy,
    tune_series_gygy,
    tune_shunt,
    tune_shunt_gy);
 inout cap_series_gygyn;
 inout cap_series_gygyp;
 inout cap_series_gyn;
 inout cap_series_gyp;
 inout cap_shunt_gyn;
 inout cap_shunt_gyp;
 inout cap_shunt_n;
 inout cap_shunt_p;
 input vdd;
 input vss;
 input [7:0] tune_series_gy;
 input [7:0] tune_series_gygy;
 input [10:0] tune_shunt;
 input [4:0] tune_shunt_gy;

 wire \gen_series_gy_g1[0].d1 ;
 wire \gen_series_gy_g1[0].d2 ;
 wire \gen_series_gy_g1[10].d1 ;
 wire \gen_series_gy_g1[10].d2 ;
 wire \gen_series_gy_g1[11].d1 ;
 wire \gen_series_gy_g1[11].d2 ;
 wire \gen_series_gy_g1[12].d1 ;
 wire \gen_series_gy_g1[12].d2 ;
 wire \gen_series_gy_g1[13].d1 ;
 wire \gen_series_gy_g1[13].d2 ;
 wire \gen_series_gy_g1[14].d1 ;
 wire \gen_series_gy_g1[14].d2 ;
 wire \gen_series_gy_g1[15].d1 ;
 wire \gen_series_gy_g1[15].d2 ;
 wire \gen_series_gy_g1[16].d1 ;
 wire \gen_series_gy_g1[16].d2 ;
 wire \gen_series_gy_g1[17].d1 ;
 wire \gen_series_gy_g1[17].d2 ;
 wire \gen_series_gy_g1[18].d1 ;
 wire \gen_series_gy_g1[18].d2 ;
 wire \gen_series_gy_g1[19].d1 ;
 wire \gen_series_gy_g1[19].d2 ;
 wire \gen_series_gy_g1[1].d1 ;
 wire \gen_series_gy_g1[1].d2 ;
 wire \gen_series_gy_g1[20].d1 ;
 wire \gen_series_gy_g1[20].d2 ;
 wire \gen_series_gy_g1[21].d1 ;
 wire \gen_series_gy_g1[21].d2 ;
 wire \gen_series_gy_g1[22].d1 ;
 wire \gen_series_gy_g1[22].d2 ;
 wire \gen_series_gy_g1[23].d1 ;
 wire \gen_series_gy_g1[23].d2 ;
 wire \gen_series_gy_g1[24].d1 ;
 wire \gen_series_gy_g1[24].d2 ;
 wire \gen_series_gy_g1[25].d1 ;
 wire \gen_series_gy_g1[25].d2 ;
 wire \gen_series_gy_g1[26].d1 ;
 wire \gen_series_gy_g1[26].d2 ;
 wire \gen_series_gy_g1[27].d1 ;
 wire \gen_series_gy_g1[27].d2 ;
 wire \gen_series_gy_g1[28].d1 ;
 wire \gen_series_gy_g1[28].d2 ;
 wire \gen_series_gy_g1[29].d1 ;
 wire \gen_series_gy_g1[29].d2 ;
 wire \gen_series_gy_g1[2].d1 ;
 wire \gen_series_gy_g1[2].d2 ;
 wire \gen_series_gy_g1[30].d1 ;
 wire \gen_series_gy_g1[30].d2 ;
 wire \gen_series_gy_g1[31].d1 ;
 wire \gen_series_gy_g1[31].d2 ;
 wire \gen_series_gy_g1[3].d1 ;
 wire \gen_series_gy_g1[3].d2 ;
 wire \gen_series_gy_g1[4].d1 ;
 wire \gen_series_gy_g1[4].d2 ;
 wire \gen_series_gy_g1[5].d1 ;
 wire \gen_series_gy_g1[5].d2 ;
 wire \gen_series_gy_g1[6].d1 ;
 wire \gen_series_gy_g1[6].d2 ;
 wire \gen_series_gy_g1[7].d1 ;
 wire \gen_series_gy_g1[7].d2 ;
 wire \gen_series_gy_g1[8].d1 ;
 wire \gen_series_gy_g1[8].d2 ;
 wire \gen_series_gy_g1[9].d1 ;
 wire \gen_series_gy_g1[9].d2 ;
 wire \gen_series_gy_g2[0].d1 ;
 wire \gen_series_gy_g2[0].d2 ;
 wire \gen_series_gy_g2[10].d1 ;
 wire \gen_series_gy_g2[10].d2 ;
 wire \gen_series_gy_g2[11].d1 ;
 wire \gen_series_gy_g2[11].d2 ;
 wire \gen_series_gy_g2[12].d1 ;
 wire \gen_series_gy_g2[12].d2 ;
 wire \gen_series_gy_g2[13].d1 ;
 wire \gen_series_gy_g2[13].d2 ;
 wire \gen_series_gy_g2[14].d1 ;
 wire \gen_series_gy_g2[14].d2 ;
 wire \gen_series_gy_g2[15].d1 ;
 wire \gen_series_gy_g2[15].d2 ;
 wire \gen_series_gy_g2[1].d1 ;
 wire \gen_series_gy_g2[1].d2 ;
 wire \gen_series_gy_g2[2].d1 ;
 wire \gen_series_gy_g2[2].d2 ;
 wire \gen_series_gy_g2[3].d1 ;
 wire \gen_series_gy_g2[3].d2 ;
 wire \gen_series_gy_g2[4].d1 ;
 wire \gen_series_gy_g2[4].d2 ;
 wire \gen_series_gy_g2[5].d1 ;
 wire \gen_series_gy_g2[5].d2 ;
 wire \gen_series_gy_g2[6].d1 ;
 wire \gen_series_gy_g2[6].d2 ;
 wire \gen_series_gy_g2[7].d1 ;
 wire \gen_series_gy_g2[7].d2 ;
 wire \gen_series_gy_g2[8].d1 ;
 wire \gen_series_gy_g2[8].d2 ;
 wire \gen_series_gy_g2[9].d1 ;
 wire \gen_series_gy_g2[9].d2 ;
 wire \gen_series_gy_g3[0].d1 ;
 wire \gen_series_gy_g3[0].d2 ;
 wire \gen_series_gy_g3[0].d3 ;
 wire \gen_series_gy_g3[0].d4 ;
 wire \gen_series_gy_g3[1].d1 ;
 wire \gen_series_gy_g3[1].d2 ;
 wire \gen_series_gy_g3[1].d3 ;
 wire \gen_series_gy_g3[1].d4 ;
 wire \gen_series_gy_g3[2].d1 ;
 wire \gen_series_gy_g3[2].d2 ;
 wire \gen_series_gy_g3[2].d3 ;
 wire \gen_series_gy_g3[2].d4 ;
 wire \gen_series_gy_g3[3].d1 ;
 wire \gen_series_gy_g3[3].d2 ;
 wire \gen_series_gy_g3[3].d3 ;
 wire \gen_series_gy_g3[3].d4 ;
 wire \gen_series_gy_g3[4].d1 ;
 wire \gen_series_gy_g3[4].d2 ;
 wire \gen_series_gy_g3[4].d3 ;
 wire \gen_series_gy_g3[4].d4 ;
 wire \gen_series_gy_g3[5].d1 ;
 wire \gen_series_gy_g3[5].d2 ;
 wire \gen_series_gy_g3[5].d3 ;
 wire \gen_series_gy_g3[5].d4 ;
 wire \gen_series_gy_g3[6].d1 ;
 wire \gen_series_gy_g3[6].d2 ;
 wire \gen_series_gy_g3[6].d3 ;
 wire \gen_series_gy_g3[6].d4 ;
 wire \gen_series_gy_g3[7].d1 ;
 wire \gen_series_gy_g3[7].d2 ;
 wire \gen_series_gy_g3[7].d3 ;
 wire \gen_series_gy_g3[7].d4 ;
 wire \gen_series_gy_g4[0].d1 ;
 wire \gen_series_gy_g4[0].d2 ;
 wire \gen_series_gy_g4[0].d3 ;
 wire \gen_series_gy_g4[0].d4 ;
 wire \gen_series_gy_g4[1].d1 ;
 wire \gen_series_gy_g4[1].d2 ;
 wire \gen_series_gy_g4[1].d3 ;
 wire \gen_series_gy_g4[1].d4 ;
 wire \gen_series_gy_g4[2].d1 ;
 wire \gen_series_gy_g4[2].d2 ;
 wire \gen_series_gy_g4[2].d3 ;
 wire \gen_series_gy_g4[2].d4 ;
 wire \gen_series_gy_g4[3].d1 ;
 wire \gen_series_gy_g4[3].d2 ;
 wire \gen_series_gy_g4[3].d3 ;
 wire \gen_series_gy_g4[3].d4 ;
 wire \gen_series_gy_g5[0].d1 ;
 wire \gen_series_gy_g5[0].d2 ;
 wire \gen_series_gy_g5[1].d1 ;
 wire \gen_series_gy_g5[1].d2 ;
 wire \gen_series_gy_g6[0].d1 ;
 wire \gen_series_gy_g6[0].d2 ;
 wire \gen_shunt_g1[0].d1 ;
 wire \gen_shunt_g1[0].d2 ;
 wire \gen_shunt_g1[10].d1 ;
 wire \gen_shunt_g1[10].d2 ;
 wire \gen_shunt_g1[11].d1 ;
 wire \gen_shunt_g1[11].d2 ;
 wire \gen_shunt_g1[12].d1 ;
 wire \gen_shunt_g1[12].d2 ;
 wire \gen_shunt_g1[13].d1 ;
 wire \gen_shunt_g1[13].d2 ;
 wire \gen_shunt_g1[14].d1 ;
 wire \gen_shunt_g1[14].d2 ;
 wire \gen_shunt_g1[15].d1 ;
 wire \gen_shunt_g1[15].d2 ;
 wire \gen_shunt_g1[16].d1 ;
 wire \gen_shunt_g1[16].d2 ;
 wire \gen_shunt_g1[17].d1 ;
 wire \gen_shunt_g1[17].d2 ;
 wire \gen_shunt_g1[18].d1 ;
 wire \gen_shunt_g1[18].d2 ;
 wire \gen_shunt_g1[19].d1 ;
 wire \gen_shunt_g1[19].d2 ;
 wire \gen_shunt_g1[1].d1 ;
 wire \gen_shunt_g1[1].d2 ;
 wire \gen_shunt_g1[20].d1 ;
 wire \gen_shunt_g1[20].d2 ;
 wire \gen_shunt_g1[21].d1 ;
 wire \gen_shunt_g1[21].d2 ;
 wire \gen_shunt_g1[22].d1 ;
 wire \gen_shunt_g1[22].d2 ;
 wire \gen_shunt_g1[23].d1 ;
 wire \gen_shunt_g1[23].d2 ;
 wire \gen_shunt_g1[24].d1 ;
 wire \gen_shunt_g1[24].d2 ;
 wire \gen_shunt_g1[25].d1 ;
 wire \gen_shunt_g1[25].d2 ;
 wire \gen_shunt_g1[26].d1 ;
 wire \gen_shunt_g1[26].d2 ;
 wire \gen_shunt_g1[27].d1 ;
 wire \gen_shunt_g1[27].d2 ;
 wire \gen_shunt_g1[28].d1 ;
 wire \gen_shunt_g1[28].d2 ;
 wire \gen_shunt_g1[29].d1 ;
 wire \gen_shunt_g1[29].d2 ;
 wire \gen_shunt_g1[2].d1 ;
 wire \gen_shunt_g1[2].d2 ;
 wire \gen_shunt_g1[30].d1 ;
 wire \gen_shunt_g1[30].d2 ;
 wire \gen_shunt_g1[31].d1 ;
 wire \gen_shunt_g1[31].d2 ;
 wire \gen_shunt_g1[32].d1 ;
 wire \gen_shunt_g1[32].d2 ;
 wire \gen_shunt_g1[33].d1 ;
 wire \gen_shunt_g1[33].d2 ;
 wire \gen_shunt_g1[34].d1 ;
 wire \gen_shunt_g1[34].d2 ;
 wire \gen_shunt_g1[35].d1 ;
 wire \gen_shunt_g1[35].d2 ;
 wire \gen_shunt_g1[36].d1 ;
 wire \gen_shunt_g1[36].d2 ;
 wire \gen_shunt_g1[37].d1 ;
 wire \gen_shunt_g1[37].d2 ;
 wire \gen_shunt_g1[38].d1 ;
 wire \gen_shunt_g1[38].d2 ;
 wire \gen_shunt_g1[39].d1 ;
 wire \gen_shunt_g1[39].d2 ;
 wire \gen_shunt_g1[3].d1 ;
 wire \gen_shunt_g1[3].d2 ;
 wire \gen_shunt_g1[40].d1 ;
 wire \gen_shunt_g1[40].d2 ;
 wire \gen_shunt_g1[41].d1 ;
 wire \gen_shunt_g1[41].d2 ;
 wire \gen_shunt_g1[42].d1 ;
 wire \gen_shunt_g1[42].d2 ;
 wire \gen_shunt_g1[43].d1 ;
 wire \gen_shunt_g1[43].d2 ;
 wire \gen_shunt_g1[44].d1 ;
 wire \gen_shunt_g1[44].d2 ;
 wire \gen_shunt_g1[45].d1 ;
 wire \gen_shunt_g1[45].d2 ;
 wire \gen_shunt_g1[46].d1 ;
 wire \gen_shunt_g1[46].d2 ;
 wire \gen_shunt_g1[47].d1 ;
 wire \gen_shunt_g1[47].d2 ;
 wire \gen_shunt_g1[48].d1 ;
 wire \gen_shunt_g1[48].d2 ;
 wire \gen_shunt_g1[49].d1 ;
 wire \gen_shunt_g1[49].d2 ;
 wire \gen_shunt_g1[4].d1 ;
 wire \gen_shunt_g1[4].d2 ;
 wire \gen_shunt_g1[50].d1 ;
 wire \gen_shunt_g1[50].d2 ;
 wire \gen_shunt_g1[51].d1 ;
 wire \gen_shunt_g1[51].d2 ;
 wire \gen_shunt_g1[52].d1 ;
 wire \gen_shunt_g1[52].d2 ;
 wire \gen_shunt_g1[53].d1 ;
 wire \gen_shunt_g1[53].d2 ;
 wire \gen_shunt_g1[54].d1 ;
 wire \gen_shunt_g1[54].d2 ;
 wire \gen_shunt_g1[55].d1 ;
 wire \gen_shunt_g1[55].d2 ;
 wire \gen_shunt_g1[56].d1 ;
 wire \gen_shunt_g1[56].d2 ;
 wire \gen_shunt_g1[57].d1 ;
 wire \gen_shunt_g1[57].d2 ;
 wire \gen_shunt_g1[58].d1 ;
 wire \gen_shunt_g1[58].d2 ;
 wire \gen_shunt_g1[59].d1 ;
 wire \gen_shunt_g1[59].d2 ;
 wire \gen_shunt_g1[5].d1 ;
 wire \gen_shunt_g1[5].d2 ;
 wire \gen_shunt_g1[60].d1 ;
 wire \gen_shunt_g1[60].d2 ;
 wire \gen_shunt_g1[61].d1 ;
 wire \gen_shunt_g1[61].d2 ;
 wire \gen_shunt_g1[62].d1 ;
 wire \gen_shunt_g1[62].d2 ;
 wire \gen_shunt_g1[63].d1 ;
 wire \gen_shunt_g1[63].d2 ;
 wire \gen_shunt_g1[6].d1 ;
 wire \gen_shunt_g1[6].d2 ;
 wire \gen_shunt_g1[7].d1 ;
 wire \gen_shunt_g1[7].d2 ;
 wire \gen_shunt_g1[8].d1 ;
 wire \gen_shunt_g1[8].d2 ;
 wire \gen_shunt_g1[9].d1 ;
 wire \gen_shunt_g1[9].d2 ;
 wire \gen_shunt_g2[0].d1 ;
 wire \gen_shunt_g2[0].d2 ;
 wire \gen_shunt_g2[0].d3 ;
 wire \gen_shunt_g2[0].d4 ;
 wire \gen_shunt_g2[10].d1 ;
 wire \gen_shunt_g2[10].d2 ;
 wire \gen_shunt_g2[10].d3 ;
 wire \gen_shunt_g2[10].d4 ;
 wire \gen_shunt_g2[11].d1 ;
 wire \gen_shunt_g2[11].d2 ;
 wire \gen_shunt_g2[11].d3 ;
 wire \gen_shunt_g2[11].d4 ;
 wire \gen_shunt_g2[12].d1 ;
 wire \gen_shunt_g2[12].d2 ;
 wire \gen_shunt_g2[12].d3 ;
 wire \gen_shunt_g2[12].d4 ;
 wire \gen_shunt_g2[13].d1 ;
 wire \gen_shunt_g2[13].d2 ;
 wire \gen_shunt_g2[13].d3 ;
 wire \gen_shunt_g2[13].d4 ;
 wire \gen_shunt_g2[14].d1 ;
 wire \gen_shunt_g2[14].d2 ;
 wire \gen_shunt_g2[14].d3 ;
 wire \gen_shunt_g2[14].d4 ;
 wire \gen_shunt_g2[15].d1 ;
 wire \gen_shunt_g2[15].d2 ;
 wire \gen_shunt_g2[15].d3 ;
 wire \gen_shunt_g2[15].d4 ;
 wire \gen_shunt_g2[16].d1 ;
 wire \gen_shunt_g2[16].d2 ;
 wire \gen_shunt_g2[16].d3 ;
 wire \gen_shunt_g2[16].d4 ;
 wire \gen_shunt_g2[17].d1 ;
 wire \gen_shunt_g2[17].d2 ;
 wire \gen_shunt_g2[17].d3 ;
 wire \gen_shunt_g2[17].d4 ;
 wire \gen_shunt_g2[18].d1 ;
 wire \gen_shunt_g2[18].d2 ;
 wire \gen_shunt_g2[18].d3 ;
 wire \gen_shunt_g2[18].d4 ;
 wire \gen_shunt_g2[19].d1 ;
 wire \gen_shunt_g2[19].d2 ;
 wire \gen_shunt_g2[19].d3 ;
 wire \gen_shunt_g2[19].d4 ;
 wire \gen_shunt_g2[1].d1 ;
 wire \gen_shunt_g2[1].d2 ;
 wire \gen_shunt_g2[1].d3 ;
 wire \gen_shunt_g2[1].d4 ;
 wire \gen_shunt_g2[20].d1 ;
 wire \gen_shunt_g2[20].d2 ;
 wire \gen_shunt_g2[20].d3 ;
 wire \gen_shunt_g2[20].d4 ;
 wire \gen_shunt_g2[21].d1 ;
 wire \gen_shunt_g2[21].d2 ;
 wire \gen_shunt_g2[21].d3 ;
 wire \gen_shunt_g2[21].d4 ;
 wire \gen_shunt_g2[22].d1 ;
 wire \gen_shunt_g2[22].d2 ;
 wire \gen_shunt_g2[22].d3 ;
 wire \gen_shunt_g2[22].d4 ;
 wire \gen_shunt_g2[23].d1 ;
 wire \gen_shunt_g2[23].d2 ;
 wire \gen_shunt_g2[23].d3 ;
 wire \gen_shunt_g2[23].d4 ;
 wire \gen_shunt_g2[24].d1 ;
 wire \gen_shunt_g2[24].d2 ;
 wire \gen_shunt_g2[24].d3 ;
 wire \gen_shunt_g2[24].d4 ;
 wire \gen_shunt_g2[25].d1 ;
 wire \gen_shunt_g2[25].d2 ;
 wire \gen_shunt_g2[25].d3 ;
 wire \gen_shunt_g2[25].d4 ;
 wire \gen_shunt_g2[26].d1 ;
 wire \gen_shunt_g2[26].d2 ;
 wire \gen_shunt_g2[26].d3 ;
 wire \gen_shunt_g2[26].d4 ;
 wire \gen_shunt_g2[27].d1 ;
 wire \gen_shunt_g2[27].d2 ;
 wire \gen_shunt_g2[27].d3 ;
 wire \gen_shunt_g2[27].d4 ;
 wire \gen_shunt_g2[28].d1 ;
 wire \gen_shunt_g2[28].d2 ;
 wire \gen_shunt_g2[28].d3 ;
 wire \gen_shunt_g2[28].d4 ;
 wire \gen_shunt_g2[29].d1 ;
 wire \gen_shunt_g2[29].d2 ;
 wire \gen_shunt_g2[29].d3 ;
 wire \gen_shunt_g2[29].d4 ;
 wire \gen_shunt_g2[2].d1 ;
 wire \gen_shunt_g2[2].d2 ;
 wire \gen_shunt_g2[2].d3 ;
 wire \gen_shunt_g2[2].d4 ;
 wire \gen_shunt_g2[30].d1 ;
 wire \gen_shunt_g2[30].d2 ;
 wire \gen_shunt_g2[30].d3 ;
 wire \gen_shunt_g2[30].d4 ;
 wire \gen_shunt_g2[31].d1 ;
 wire \gen_shunt_g2[31].d2 ;
 wire \gen_shunt_g2[31].d3 ;
 wire \gen_shunt_g2[31].d4 ;
 wire \gen_shunt_g2[3].d1 ;
 wire \gen_shunt_g2[3].d2 ;
 wire \gen_shunt_g2[3].d3 ;
 wire \gen_shunt_g2[3].d4 ;
 wire \gen_shunt_g2[4].d1 ;
 wire \gen_shunt_g2[4].d2 ;
 wire \gen_shunt_g2[4].d3 ;
 wire \gen_shunt_g2[4].d4 ;
 wire \gen_shunt_g2[5].d1 ;
 wire \gen_shunt_g2[5].d2 ;
 wire \gen_shunt_g2[5].d3 ;
 wire \gen_shunt_g2[5].d4 ;
 wire \gen_shunt_g2[6].d1 ;
 wire \gen_shunt_g2[6].d2 ;
 wire \gen_shunt_g2[6].d3 ;
 wire \gen_shunt_g2[6].d4 ;
 wire \gen_shunt_g2[7].d1 ;
 wire \gen_shunt_g2[7].d2 ;
 wire \gen_shunt_g2[7].d3 ;
 wire \gen_shunt_g2[7].d4 ;
 wire \gen_shunt_g2[8].d1 ;
 wire \gen_shunt_g2[8].d2 ;
 wire \gen_shunt_g2[8].d3 ;
 wire \gen_shunt_g2[8].d4 ;
 wire \gen_shunt_g2[9].d1 ;
 wire \gen_shunt_g2[9].d2 ;
 wire \gen_shunt_g2[9].d3 ;
 wire \gen_shunt_g2[9].d4 ;
 wire \gen_shunt_g3[0].d1 ;
 wire \gen_shunt_g3[0].d2 ;
 wire \gen_shunt_g3[0].d3 ;
 wire \gen_shunt_g3[0].d4 ;
 wire \gen_shunt_g3[10].d1 ;
 wire \gen_shunt_g3[10].d2 ;
 wire \gen_shunt_g3[10].d3 ;
 wire \gen_shunt_g3[10].d4 ;
 wire \gen_shunt_g3[11].d1 ;
 wire \gen_shunt_g3[11].d2 ;
 wire \gen_shunt_g3[11].d3 ;
 wire \gen_shunt_g3[11].d4 ;
 wire \gen_shunt_g3[12].d1 ;
 wire \gen_shunt_g3[12].d2 ;
 wire \gen_shunt_g3[12].d3 ;
 wire \gen_shunt_g3[12].d4 ;
 wire \gen_shunt_g3[13].d1 ;
 wire \gen_shunt_g3[13].d2 ;
 wire \gen_shunt_g3[13].d3 ;
 wire \gen_shunt_g3[13].d4 ;
 wire \gen_shunt_g3[14].d1 ;
 wire \gen_shunt_g3[14].d2 ;
 wire \gen_shunt_g3[14].d3 ;
 wire \gen_shunt_g3[14].d4 ;
 wire \gen_shunt_g3[15].d1 ;
 wire \gen_shunt_g3[15].d2 ;
 wire \gen_shunt_g3[15].d3 ;
 wire \gen_shunt_g3[15].d4 ;
 wire \gen_shunt_g3[1].d1 ;
 wire \gen_shunt_g3[1].d2 ;
 wire \gen_shunt_g3[1].d3 ;
 wire \gen_shunt_g3[1].d4 ;
 wire \gen_shunt_g3[2].d1 ;
 wire \gen_shunt_g3[2].d2 ;
 wire \gen_shunt_g3[2].d3 ;
 wire \gen_shunt_g3[2].d4 ;
 wire \gen_shunt_g3[3].d1 ;
 wire \gen_shunt_g3[3].d2 ;
 wire \gen_shunt_g3[3].d3 ;
 wire \gen_shunt_g3[3].d4 ;
 wire \gen_shunt_g3[4].d1 ;
 wire \gen_shunt_g3[4].d2 ;
 wire \gen_shunt_g3[4].d3 ;
 wire \gen_shunt_g3[4].d4 ;
 wire \gen_shunt_g3[5].d1 ;
 wire \gen_shunt_g3[5].d2 ;
 wire \gen_shunt_g3[5].d3 ;
 wire \gen_shunt_g3[5].d4 ;
 wire \gen_shunt_g3[6].d1 ;
 wire \gen_shunt_g3[6].d2 ;
 wire \gen_shunt_g3[6].d3 ;
 wire \gen_shunt_g3[6].d4 ;
 wire \gen_shunt_g3[7].d1 ;
 wire \gen_shunt_g3[7].d2 ;
 wire \gen_shunt_g3[7].d3 ;
 wire \gen_shunt_g3[7].d4 ;
 wire \gen_shunt_g3[8].d1 ;
 wire \gen_shunt_g3[8].d2 ;
 wire \gen_shunt_g3[8].d3 ;
 wire \gen_shunt_g3[8].d4 ;
 wire \gen_shunt_g3[9].d1 ;
 wire \gen_shunt_g3[9].d2 ;
 wire \gen_shunt_g3[9].d3 ;
 wire \gen_shunt_g3[9].d4 ;
 wire \gen_shunt_g4[0].d1 ;
 wire \gen_shunt_g4[0].d2 ;
 wire \gen_shunt_g4[0].d3 ;
 wire \gen_shunt_g4[0].d4 ;
 wire \gen_shunt_g4[1].d1 ;
 wire \gen_shunt_g4[1].d2 ;
 wire \gen_shunt_g4[1].d3 ;
 wire \gen_shunt_g4[1].d4 ;
 wire \gen_shunt_g4[2].d1 ;
 wire \gen_shunt_g4[2].d2 ;
 wire \gen_shunt_g4[2].d3 ;
 wire \gen_shunt_g4[2].d4 ;
 wire \gen_shunt_g4[3].d1 ;
 wire \gen_shunt_g4[3].d2 ;
 wire \gen_shunt_g4[3].d3 ;
 wire \gen_shunt_g4[3].d4 ;
 wire \gen_shunt_g4[4].d1 ;
 wire \gen_shunt_g4[4].d2 ;
 wire \gen_shunt_g4[4].d3 ;
 wire \gen_shunt_g4[4].d4 ;
 wire \gen_shunt_g4[5].d1 ;
 wire \gen_shunt_g4[5].d2 ;
 wire \gen_shunt_g4[5].d3 ;
 wire \gen_shunt_g4[5].d4 ;
 wire \gen_shunt_g4[6].d1 ;
 wire \gen_shunt_g4[6].d2 ;
 wire \gen_shunt_g4[6].d3 ;
 wire \gen_shunt_g4[6].d4 ;
 wire \gen_shunt_g4[7].d1 ;
 wire \gen_shunt_g4[7].d2 ;
 wire \gen_shunt_g4[7].d3 ;
 wire \gen_shunt_g4[7].d4 ;
 wire \gen_shunt_g5[0].d1 ;
 wire \gen_shunt_g5[0].d2 ;
 wire \gen_shunt_g5[1].d1 ;
 wire \gen_shunt_g5[1].d2 ;
 wire \gen_shunt_g5[2].d1 ;
 wire \gen_shunt_g5[2].d2 ;
 wire \gen_shunt_g5[3].d1 ;
 wire \gen_shunt_g5[3].d2 ;
 wire \gen_shunt_g6[0].d1 ;
 wire \gen_shunt_g6[0].d2 ;
 wire \gen_shunt_g6[0].d3 ;
 wire \gen_shunt_g6[0].d4 ;
 wire \gen_shunt_g6[1].d1 ;
 wire \gen_shunt_g6[1].d2 ;
 wire \gen_shunt_g6[1].d3 ;
 wire \gen_shunt_g6[1].d4 ;
 wire \gen_shunt_g7[0].d1 ;
 wire \gen_shunt_g7[0].d2 ;
 wire \gen_shunt_gy_g1[0].d1 ;
 wire \gen_shunt_gy_g1[0].d2 ;
 wire \gen_shunt_gy_g1[0].d3 ;
 wire \gen_shunt_gy_g1[0].d4 ;
 wire \gen_shunt_gy_g1[1].d1 ;
 wire \gen_shunt_gy_g1[1].d2 ;
 wire \gen_shunt_gy_g1[1].d3 ;
 wire \gen_shunt_gy_g1[1].d4 ;
 wire \gen_shunt_gy_g1[2].d1 ;
 wire \gen_shunt_gy_g1[2].d2 ;
 wire \gen_shunt_gy_g1[2].d3 ;
 wire \gen_shunt_gy_g1[2].d4 ;
 wire \gen_shunt_gy_g1[3].d1 ;
 wire \gen_shunt_gy_g1[3].d2 ;
 wire \gen_shunt_gy_g1[3].d3 ;
 wire \gen_shunt_gy_g1[3].d4 ;
 wire \gen_shunt_gy_g1[4].d1 ;
 wire \gen_shunt_gy_g1[4].d2 ;
 wire \gen_shunt_gy_g1[4].d3 ;
 wire \gen_shunt_gy_g1[4].d4 ;
 wire \gen_shunt_gy_g1[5].d1 ;
 wire \gen_shunt_gy_g1[5].d2 ;
 wire \gen_shunt_gy_g1[5].d3 ;
 wire \gen_shunt_gy_g1[5].d4 ;
 wire \gen_shunt_gy_g1[6].d1 ;
 wire \gen_shunt_gy_g1[6].d2 ;
 wire \gen_shunt_gy_g1[6].d3 ;
 wire \gen_shunt_gy_g1[6].d4 ;
 wire \gen_shunt_gy_g1[7].d1 ;
 wire \gen_shunt_gy_g1[7].d2 ;
 wire \gen_shunt_gy_g1[7].d3 ;
 wire \gen_shunt_gy_g1[7].d4 ;
 wire \gen_shunt_gy_g2[0].d1 ;
 wire \gen_shunt_gy_g2[0].d2 ;
 wire \gen_shunt_gy_g2[0].d3 ;
 wire \gen_shunt_gy_g2[0].d4 ;
 wire \gen_shunt_gy_g2[1].d1 ;
 wire \gen_shunt_gy_g2[1].d2 ;
 wire \gen_shunt_gy_g2[1].d3 ;
 wire \gen_shunt_gy_g2[1].d4 ;
 wire \gen_shunt_gy_g2[2].d1 ;
 wire \gen_shunt_gy_g2[2].d2 ;
 wire \gen_shunt_gy_g2[2].d3 ;
 wire \gen_shunt_gy_g2[2].d4 ;
 wire \gen_shunt_gy_g2[3].d1 ;
 wire \gen_shunt_gy_g2[3].d2 ;
 wire \gen_shunt_gy_g2[3].d3 ;
 wire \gen_shunt_gy_g2[3].d4 ;
 wire \gen_shunt_gy_g3[0].d1 ;
 wire \gen_shunt_gy_g3[0].d2 ;
 wire \gen_shunt_gy_g3[1].d1 ;
 wire \gen_shunt_gy_g3[1].d2 ;
 wire \gen_shunt_gy_g4[0].d1 ;
 wire \gen_shunt_gy_g4[0].d2 ;
 wire \gen_shunt_gygy_g1[0].d1 ;
 wire \gen_shunt_gygy_g1[0].d2 ;
 wire \gen_shunt_gygy_g1[0].d3 ;
 wire \gen_shunt_gygy_g1[0].d4 ;
 wire \gen_shunt_gygy_g1[10].d1 ;
 wire \gen_shunt_gygy_g1[10].d2 ;
 wire \gen_shunt_gygy_g1[10].d3 ;
 wire \gen_shunt_gygy_g1[10].d4 ;
 wire \gen_shunt_gygy_g1[11].d1 ;
 wire \gen_shunt_gygy_g1[11].d2 ;
 wire \gen_shunt_gygy_g1[11].d3 ;
 wire \gen_shunt_gygy_g1[11].d4 ;
 wire \gen_shunt_gygy_g1[12].d1 ;
 wire \gen_shunt_gygy_g1[12].d2 ;
 wire \gen_shunt_gygy_g1[12].d3 ;
 wire \gen_shunt_gygy_g1[12].d4 ;
 wire \gen_shunt_gygy_g1[13].d1 ;
 wire \gen_shunt_gygy_g1[13].d2 ;
 wire \gen_shunt_gygy_g1[13].d3 ;
 wire \gen_shunt_gygy_g1[13].d4 ;
 wire \gen_shunt_gygy_g1[14].d1 ;
 wire \gen_shunt_gygy_g1[14].d2 ;
 wire \gen_shunt_gygy_g1[14].d3 ;
 wire \gen_shunt_gygy_g1[14].d4 ;
 wire \gen_shunt_gygy_g1[15].d1 ;
 wire \gen_shunt_gygy_g1[15].d2 ;
 wire \gen_shunt_gygy_g1[15].d3 ;
 wire \gen_shunt_gygy_g1[15].d4 ;
 wire \gen_shunt_gygy_g1[1].d1 ;
 wire \gen_shunt_gygy_g1[1].d2 ;
 wire \gen_shunt_gygy_g1[1].d3 ;
 wire \gen_shunt_gygy_g1[1].d4 ;
 wire \gen_shunt_gygy_g1[2].d1 ;
 wire \gen_shunt_gygy_g1[2].d2 ;
 wire \gen_shunt_gygy_g1[2].d3 ;
 wire \gen_shunt_gygy_g1[2].d4 ;
 wire \gen_shunt_gygy_g1[3].d1 ;
 wire \gen_shunt_gygy_g1[3].d2 ;
 wire \gen_shunt_gygy_g1[3].d3 ;
 wire \gen_shunt_gygy_g1[3].d4 ;
 wire \gen_shunt_gygy_g1[4].d1 ;
 wire \gen_shunt_gygy_g1[4].d2 ;
 wire \gen_shunt_gygy_g1[4].d3 ;
 wire \gen_shunt_gygy_g1[4].d4 ;
 wire \gen_shunt_gygy_g1[5].d1 ;
 wire \gen_shunt_gygy_g1[5].d2 ;
 wire \gen_shunt_gygy_g1[5].d3 ;
 wire \gen_shunt_gygy_g1[5].d4 ;
 wire \gen_shunt_gygy_g1[6].d1 ;
 wire \gen_shunt_gygy_g1[6].d2 ;
 wire \gen_shunt_gygy_g1[6].d3 ;
 wire \gen_shunt_gygy_g1[6].d4 ;
 wire \gen_shunt_gygy_g1[7].d1 ;
 wire \gen_shunt_gygy_g1[7].d2 ;
 wire \gen_shunt_gygy_g1[7].d3 ;
 wire \gen_shunt_gygy_g1[7].d4 ;
 wire \gen_shunt_gygy_g1[8].d1 ;
 wire \gen_shunt_gygy_g1[8].d2 ;
 wire \gen_shunt_gygy_g1[8].d3 ;
 wire \gen_shunt_gygy_g1[8].d4 ;
 wire \gen_shunt_gygy_g1[9].d1 ;
 wire \gen_shunt_gygy_g1[9].d2 ;
 wire \gen_shunt_gygy_g1[9].d3 ;
 wire \gen_shunt_gygy_g1[9].d4 ;
 wire \gen_shunt_gygy_g2[0].d1 ;
 wire \gen_shunt_gygy_g2[0].d2 ;
 wire \gen_shunt_gygy_g2[0].d3 ;
 wire \gen_shunt_gygy_g2[0].d4 ;
 wire \gen_shunt_gygy_g2[1].d1 ;
 wire \gen_shunt_gygy_g2[1].d2 ;
 wire \gen_shunt_gygy_g2[1].d3 ;
 wire \gen_shunt_gygy_g2[1].d4 ;
 wire \gen_shunt_gygy_g2[2].d1 ;
 wire \gen_shunt_gygy_g2[2].d2 ;
 wire \gen_shunt_gygy_g2[2].d3 ;
 wire \gen_shunt_gygy_g2[2].d4 ;
 wire \gen_shunt_gygy_g2[3].d1 ;
 wire \gen_shunt_gygy_g2[3].d2 ;
 wire \gen_shunt_gygy_g2[3].d3 ;
 wire \gen_shunt_gygy_g2[3].d4 ;
 wire \gen_shunt_gygy_g2[4].d1 ;
 wire \gen_shunt_gygy_g2[4].d2 ;
 wire \gen_shunt_gygy_g2[4].d3 ;
 wire \gen_shunt_gygy_g2[4].d4 ;
 wire \gen_shunt_gygy_g2[5].d1 ;
 wire \gen_shunt_gygy_g2[5].d2 ;
 wire \gen_shunt_gygy_g2[5].d3 ;
 wire \gen_shunt_gygy_g2[5].d4 ;
 wire \gen_shunt_gygy_g2[6].d1 ;
 wire \gen_shunt_gygy_g2[6].d2 ;
 wire \gen_shunt_gygy_g2[6].d3 ;
 wire \gen_shunt_gygy_g2[6].d4 ;
 wire \gen_shunt_gygy_g2[7].d1 ;
 wire \gen_shunt_gygy_g2[7].d2 ;
 wire \gen_shunt_gygy_g2[7].d3 ;
 wire \gen_shunt_gygy_g2[7].d4 ;
 wire \gen_shunt_gygy_g3[0].d1 ;
 wire \gen_shunt_gygy_g3[0].d2 ;
 wire \gen_shunt_gygy_g3[1].d1 ;
 wire \gen_shunt_gygy_g3[1].d2 ;
 wire \gen_shunt_gygy_g3[2].d1 ;
 wire \gen_shunt_gygy_g3[2].d2 ;
 wire \gen_shunt_gygy_g3[3].d1 ;
 wire \gen_shunt_gygy_g3[3].d2 ;
 wire \gen_shunt_gygy_g4[0].d1 ;
 wire \gen_shunt_gygy_g4[0].d2 ;
 wire \gen_shunt_gygy_g4[0].d3 ;
 wire \gen_shunt_gygy_g4[0].d4 ;
 wire \gen_shunt_gygy_g4[1].d1 ;
 wire \gen_shunt_gygy_g4[1].d2 ;
 wire \gen_shunt_gygy_g4[1].d3 ;
 wire \gen_shunt_gygy_g4[1].d4 ;
 wire \gen_shunt_gygy_g5[0].d1 ;
 wire \gen_shunt_gygy_g5[0].d2 ;

 gf180mcu_fd_sc_mcu7t5v0__tiel _0_ (.ZN(\gen_shunt_gy_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1_ (.ZN(\gen_shunt_gy_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2_ (.ZN(\gen_shunt_gy_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3_ (.ZN(\gen_shunt_gy_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _4_ (.ZN(\gen_shunt_gy_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _5_ (.ZN(\gen_shunt_gy_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _6_ (.ZN(\gen_shunt_gy_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel _7_ (.ZN(\gen_shunt_gy_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[16].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[16].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[16].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[16].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[17].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[17].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[17].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[17].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[18].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[18].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[18].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[18].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[19].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[19].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[19].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[19].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[20].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[20].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[20].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[20].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[21].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[21].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[21].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[21].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[22].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[22].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[22].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[22].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[23].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[23].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[23].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[23].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[24].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[24].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[24].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[24].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[25].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[25].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[25].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[25].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[26].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[26].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[26].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[26].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[27].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[27].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[27].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[27].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[28].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[28].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[28].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[28].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[29].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[29].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[29].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[29].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[30].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[30].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[30].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[30].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[31].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[31].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[31].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[31].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[10].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[10].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[11].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[11].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[12].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[12].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[13].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[13].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[14].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[14].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[15].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[15].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[8].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[8].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[9].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[9].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g6[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[0]),
    .ZN(\gen_series_gy_g6[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g6[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[0]),
    .ZN(\gen_series_gy_g6[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[10].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[10].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[11].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[11].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[12].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[12].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[13].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[13].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[14].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[14].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[15].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[15].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[16].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[16].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[16].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[16].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[17].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[17].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[17].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[17].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[18].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[18].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[18].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[18].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[19].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[19].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[19].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[19].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[20].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[20].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[20].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[20].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[21].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[21].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[21].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[21].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[22].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[22].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[22].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[22].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[23].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[23].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[23].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[23].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[24].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[24].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[24].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[24].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[25].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[25].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[25].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[25].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[26].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[26].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[26].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[26].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[27].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[27].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[27].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[27].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[28].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[28].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[28].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[28].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[29].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[29].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[29].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[29].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[30].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[30].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[30].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[30].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[31].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[31].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[31].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[31].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[32].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[32].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[32].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[32].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[33].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[33].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[33].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[33].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[34].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[34].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[34].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[34].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[35].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[35].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[35].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[35].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[36].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[36].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[36].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[36].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[37].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[37].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[37].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[37].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[38].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[38].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[38].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[38].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[39].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[39].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[39].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[39].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[40].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[40].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[40].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[40].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[41].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[41].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[41].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[41].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[42].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[42].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[42].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[42].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[43].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[43].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[43].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[43].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[44].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[44].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[44].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[44].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[45].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[45].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[45].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[45].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[46].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[46].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[46].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[46].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[47].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[47].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[47].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[47].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[48].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[48].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[48].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[48].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[49].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[49].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[49].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[49].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[50].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[50].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[50].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[50].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[51].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[51].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[51].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[51].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[52].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[52].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[52].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[52].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[53].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[53].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[53].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[53].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[54].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[54].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[54].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[54].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[55].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[55].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[55].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[55].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[56].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[56].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[56].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[56].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[57].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[57].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[57].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[57].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[58].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[58].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[58].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[58].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[59].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[59].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[59].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[59].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[60].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[60].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[60].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[60].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[61].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[61].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[61].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[61].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[62].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[62].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[62].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[62].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[63].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[63].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[63].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[63].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[6].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[6].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[7].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[7].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[8].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[8].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[9].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[9].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[10].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[10].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[11].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[11].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[12].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[12].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[13].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[13].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[14].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[14].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[15].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[15].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[16].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[16].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[16].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[16].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[17].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[17].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[17].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[17].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[18].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[18].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[18].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[18].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[19].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[19].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[19].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[19].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[20].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[20].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[20].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[20].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[21].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[21].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[21].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[21].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[22].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[22].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[22].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[22].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[23].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[23].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[23].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[23].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[24].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[24].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[24].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[24].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[25].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[25].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[25].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[25].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[26].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[26].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[26].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[26].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[27].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[27].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[27].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[27].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[28].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[28].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[28].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[28].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[29].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[29].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[29].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[29].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[30].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[30].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[30].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[30].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[31].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[31].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[31].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[31].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[8].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[8].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[9].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[9].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[10].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[10].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[11].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[11].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[12].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[12].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[13].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[13].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[14].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[14].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[15].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[15].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[8].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[8].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[9].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[9].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[0]),
    .ZN(\gen_shunt_g7[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[0]),
    .ZN(\gen_shunt_g7[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g4[0].u_shunt_n  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[0]),
    .ZN(\gen_shunt_gy_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g4[0].u_shunt_p  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[0]),
    .ZN(\gen_shunt_gy_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[10].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[10].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[10].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[10].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[11].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[11].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[11].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[11].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[12].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[12].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[12].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[12].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[13].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[13].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[13].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[13].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[14].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[14].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[14].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[14].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[15].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[15].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[15].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[15].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[8].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[8].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[8].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[8].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[9].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[9].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[9].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[9].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[2].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[2].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[3].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[3].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[4].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[4].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[4].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[4].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[5].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[5].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[5].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[5].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[6].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[6].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[6].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[6].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[7].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[7].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[7].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[7].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[2].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[2].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[2].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[2].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[3].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[3].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[3].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[3].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[0].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[0].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[1].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[1].d4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[1].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[1].d3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g5[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[0]),
    .ZN(\gen_shunt_gygy_g5[0].d2 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g5[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[0]),
    .ZN(\gen_shunt_gygy_g5[0].d1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_687 (.VDD(vdd),
    .VSS(vss));
endmodule
