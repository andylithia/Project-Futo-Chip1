magic
tech gf180mcuC
magscale 1 10
timestamp 1669736112
<< nwell >>
rect 1258 16032 22710 16550
rect 1258 14464 22710 15328
rect 1258 12896 22710 13760
rect 1258 11328 22710 12192
rect 1258 9760 22710 10624
rect 1258 8192 22710 9056
rect 1258 6624 22710 7488
rect 1258 5056 22710 5920
rect 1258 3488 22710 4352
<< pwell >>
rect 1258 15328 22710 16032
rect 1258 13760 22710 14464
rect 1258 12192 22710 12896
rect 1258 10624 22710 11328
rect 1258 9056 22710 9760
rect 1258 7488 22710 8192
rect 1258 5920 22710 6624
rect 1258 4352 22710 5056
rect 1258 3050 22710 3488
<< mvnmos >>
rect 1692 15748 1892 15912
rect 2140 15748 2340 15912
rect 2588 15748 2788 15912
rect 3036 15748 3236 15912
rect 3484 15748 3684 15912
rect 3932 15748 4132 15912
rect 4380 15748 4580 15912
rect 4828 15748 5028 15912
rect 5612 15748 5812 15912
rect 6060 15748 6260 15912
rect 6508 15748 6708 15912
rect 6956 15748 7156 15912
rect 7404 15748 7604 15912
rect 7852 15748 8052 15912
rect 8300 15748 8500 15912
rect 8748 15748 8948 15912
rect 9532 15748 9732 15912
rect 9980 15748 10180 15912
rect 10428 15748 10628 15912
rect 10876 15748 11076 15912
rect 11324 15748 11524 15912
rect 11772 15748 11972 15912
rect 12220 15748 12420 15912
rect 12668 15748 12868 15912
rect 13452 15748 13652 15912
rect 13900 15748 14100 15912
rect 14348 15748 14548 15912
rect 14796 15748 14996 15912
rect 15244 15748 15444 15912
rect 15692 15748 15892 15912
rect 16140 15748 16340 15912
rect 16588 15748 16788 15912
rect 17372 15748 17572 15912
rect 17820 15748 18020 15912
rect 18268 15748 18468 15912
rect 18716 15748 18916 15912
rect 19164 15748 19364 15912
rect 19612 15748 19812 15912
rect 20060 15748 20260 15912
rect 20508 15748 20708 15912
rect 21292 15748 21492 15912
rect 21740 15748 21940 15912
rect 1692 15448 1892 15612
rect 2140 15448 2340 15612
rect 2588 15448 2788 15612
rect 3036 15448 3236 15612
rect 3484 15448 3684 15612
rect 3932 15448 4132 15612
rect 4380 15448 4580 15612
rect 4828 15448 5028 15612
rect 5276 15448 5476 15612
rect 5724 15448 5924 15612
rect 6172 15448 6372 15612
rect 6620 15448 6820 15612
rect 7068 15448 7268 15612
rect 7516 15448 7716 15612
rect 7964 15448 8164 15612
rect 8412 15448 8612 15612
rect 8860 15448 9060 15612
rect 9644 15448 9844 15612
rect 10092 15448 10292 15612
rect 10540 15448 10740 15612
rect 10988 15448 11188 15612
rect 11436 15448 11636 15612
rect 11884 15448 12084 15612
rect 12332 15448 12532 15612
rect 12780 15448 12980 15612
rect 13228 15448 13428 15612
rect 13676 15448 13876 15612
rect 14124 15448 14324 15612
rect 14572 15448 14772 15612
rect 15020 15448 15220 15612
rect 15468 15448 15668 15612
rect 15916 15448 16116 15612
rect 16364 15448 16564 15612
rect 16812 15448 17012 15612
rect 17596 15448 17796 15612
rect 18044 15448 18244 15612
rect 18492 15448 18692 15612
rect 18940 15448 19140 15612
rect 19388 15448 19588 15612
rect 19836 15448 20036 15612
rect 20284 15448 20484 15612
rect 20732 15448 20932 15612
rect 21180 15448 21380 15612
rect 21628 15448 21828 15612
rect 22076 15448 22276 15612
rect 1692 14180 1892 14344
rect 2140 14180 2340 14344
rect 2588 14180 2788 14344
rect 3036 14180 3236 14344
rect 3484 14180 3684 14344
rect 3932 14180 4132 14344
rect 4380 14180 4580 14344
rect 4828 14180 5028 14344
rect 5612 14180 5812 14344
rect 6060 14180 6260 14344
rect 6508 14180 6708 14344
rect 6956 14180 7156 14344
rect 7404 14180 7604 14344
rect 7852 14180 8052 14344
rect 8300 14180 8500 14344
rect 8748 14180 8948 14344
rect 9196 14180 9396 14344
rect 9644 14180 9844 14344
rect 10092 14180 10292 14344
rect 10540 14180 10740 14344
rect 10988 14180 11188 14344
rect 11436 14180 11636 14344
rect 11884 14180 12084 14344
rect 12332 14180 12532 14344
rect 12780 14180 12980 14344
rect 13564 14180 13764 14344
rect 14012 14180 14212 14344
rect 14460 14180 14660 14344
rect 14908 14180 15108 14344
rect 15356 14180 15556 14344
rect 15804 14180 16004 14344
rect 16252 14180 16452 14344
rect 16892 14180 17012 14344
rect 17564 14180 17684 14344
rect 17932 14180 18132 14344
rect 18380 14180 18580 14344
rect 18828 14180 19028 14344
rect 19276 14180 19476 14344
rect 19724 14180 19924 14344
rect 20172 14180 20372 14344
rect 20620 14180 20820 14344
rect 21516 14180 21716 14344
rect 21964 14180 22164 14344
rect 1692 13880 1892 14044
rect 2140 13880 2340 14044
rect 2588 13880 2788 14044
rect 3036 13880 3236 14044
rect 3484 13880 3684 14044
rect 3932 13880 4132 14044
rect 4380 13880 4580 14044
rect 4828 13880 5028 14044
rect 5276 13880 5476 14044
rect 5724 13880 5924 14044
rect 6172 13880 6372 14044
rect 6620 13880 6820 14044
rect 7068 13880 7268 14044
rect 7516 13880 7716 14044
rect 7964 13880 8164 14044
rect 8412 13880 8612 14044
rect 8860 13880 9060 14044
rect 9644 13880 9844 14044
rect 10092 13880 10292 14044
rect 10540 13880 10740 14044
rect 10988 13880 11188 14044
rect 11436 13880 11636 14044
rect 11884 13880 12084 14044
rect 12332 13880 12532 14044
rect 12780 13880 12980 14044
rect 13228 13880 13428 14044
rect 13676 13880 13876 14044
rect 14124 13880 14324 14044
rect 14572 13880 14772 14044
rect 15020 13880 15220 14044
rect 15468 13880 15668 14044
rect 16140 13880 16260 14044
rect 16812 13880 16932 14044
rect 17708 13880 17828 14044
rect 18380 13880 18500 14044
rect 18828 13880 19028 14044
rect 19276 13880 19476 14044
rect 19724 13880 19924 14044
rect 20172 13880 20372 14044
rect 20620 13880 20820 14044
rect 21068 13880 21268 14044
rect 21516 13880 21716 14044
rect 21964 13880 22164 14044
rect 1692 12612 1892 12776
rect 2140 12612 2340 12776
rect 2588 12612 2788 12776
rect 3036 12612 3236 12776
rect 3484 12612 3684 12776
rect 3932 12612 4132 12776
rect 4380 12612 4580 12776
rect 4828 12612 5028 12776
rect 5612 12612 5812 12776
rect 6060 12612 6260 12776
rect 6508 12612 6708 12776
rect 6956 12612 7156 12776
rect 7404 12612 7604 12776
rect 7852 12612 8052 12776
rect 8300 12612 8500 12776
rect 8748 12612 8948 12776
rect 9196 12612 9396 12776
rect 9644 12612 9844 12776
rect 10092 12612 10292 12776
rect 10540 12612 10740 12776
rect 10988 12612 11188 12776
rect 11436 12612 11636 12776
rect 11884 12612 12084 12776
rect 12332 12612 12532 12776
rect 12780 12612 12980 12776
rect 13564 12612 13764 12776
rect 14012 12612 14212 12776
rect 14796 12612 14916 12776
rect 15468 12612 15588 12776
rect 16140 12612 16260 12776
rect 16812 12612 16932 12776
rect 17484 12612 17604 12776
rect 18156 12612 18276 12776
rect 18828 12612 18948 12776
rect 19500 12612 19620 12776
rect 19948 12612 20148 12776
rect 20396 12612 20596 12776
rect 20844 12612 21044 12776
rect 21516 12612 21716 12776
rect 21964 12612 22164 12776
rect 1692 12312 1892 12476
rect 2140 12312 2340 12476
rect 2588 12312 2788 12476
rect 3036 12312 3236 12476
rect 3484 12312 3684 12476
rect 3932 12312 4132 12476
rect 4380 12312 4580 12476
rect 4828 12312 5028 12476
rect 5276 12312 5476 12476
rect 5724 12312 5924 12476
rect 6172 12312 6372 12476
rect 6620 12312 6820 12476
rect 7068 12312 7268 12476
rect 7516 12312 7716 12476
rect 7964 12312 8164 12476
rect 8412 12312 8612 12476
rect 8860 12312 9060 12476
rect 9644 12312 9844 12476
rect 10092 12312 10292 12476
rect 10540 12312 10740 12476
rect 10988 12312 11188 12476
rect 11436 12312 11636 12476
rect 11884 12312 12084 12476
rect 12332 12312 12532 12476
rect 12780 12312 12980 12476
rect 13228 12312 13428 12476
rect 13676 12312 13876 12476
rect 14124 12312 14244 12476
rect 14796 12312 14916 12476
rect 15468 12312 15588 12476
rect 16140 12312 16260 12476
rect 16812 12312 16932 12476
rect 17708 12312 17828 12476
rect 18380 12312 18500 12476
rect 19052 12312 19172 12476
rect 19724 12312 19844 12476
rect 20396 12312 20516 12476
rect 20844 12312 21044 12476
rect 21292 12312 21492 12476
rect 21740 12312 21940 12476
rect 1692 11044 1892 11208
rect 2140 11044 2340 11208
rect 2588 11044 2788 11208
rect 3036 11044 3236 11208
rect 3484 11044 3684 11208
rect 3932 11044 4132 11208
rect 4380 11044 4580 11208
rect 4828 11044 5028 11208
rect 5612 11044 5812 11208
rect 6140 11044 6260 11208
rect 6924 11044 7044 11208
rect 7596 11044 7716 11208
rect 8268 11044 8388 11208
rect 8636 11044 8836 11208
rect 9196 11044 9316 11208
rect 9868 11044 9988 11208
rect 10540 11044 10660 11208
rect 10988 11044 11188 11208
rect 11436 11044 11636 11208
rect 12108 11044 12228 11208
rect 12780 11044 12900 11208
rect 13676 11044 13796 11208
rect 14124 11044 14324 11208
rect 14796 11044 14916 11208
rect 15468 11044 15588 11208
rect 16140 11044 16260 11208
rect 16812 11044 16932 11208
rect 17484 11044 17604 11208
rect 18156 11044 18276 11208
rect 18828 11044 18948 11208
rect 19500 11044 19620 11208
rect 20172 11044 20292 11208
rect 20620 11044 20820 11208
rect 21516 11044 21716 11208
rect 21964 11044 22164 11208
rect 1692 10744 1892 10908
rect 2140 10744 2340 10908
rect 2588 10744 2788 10908
rect 3036 10744 3236 10908
rect 3484 10744 3684 10908
rect 3932 10744 4132 10908
rect 4380 10744 4580 10908
rect 4828 10744 5028 10908
rect 5388 10744 5508 10908
rect 6060 10744 6180 10908
rect 6732 10744 6852 10908
rect 7404 10744 7524 10908
rect 8076 10744 8196 10908
rect 8860 10744 8980 10908
rect 9868 10744 9988 10908
rect 10540 10744 10660 10908
rect 11212 10744 11332 10908
rect 11996 10744 12116 10908
rect 12668 10744 12788 10908
rect 13340 10744 13460 10908
rect 14012 10744 14132 10908
rect 14684 10744 14804 10908
rect 15356 10744 15476 10908
rect 16028 10744 16148 10908
rect 16700 10744 16820 10908
rect 17708 10744 17828 10908
rect 18380 10744 18500 10908
rect 19052 10744 19172 10908
rect 19724 10744 19844 10908
rect 20396 10744 20516 10908
rect 21068 10744 21188 10908
rect 21740 10744 21860 10908
rect 1692 9476 1892 9640
rect 2140 9476 2340 9640
rect 2588 9476 2788 9640
rect 3036 9476 3236 9640
rect 3484 9476 3684 9640
rect 4156 9476 4276 9640
rect 4828 9476 4948 9640
rect 5836 9476 5956 9640
rect 6508 9476 6628 9640
rect 7180 9476 7300 9640
rect 7852 9476 7972 9640
rect 8524 9476 8644 9640
rect 9196 9476 9316 9640
rect 9868 9476 9988 9640
rect 10540 9476 10660 9640
rect 10988 9476 11188 9640
rect 11436 9476 11556 9640
rect 12108 9476 12228 9640
rect 12780 9476 12900 9640
rect 13676 9476 13796 9640
rect 14348 9476 14468 9640
rect 15020 9476 15140 9640
rect 15692 9476 15812 9640
rect 16364 9476 16484 9640
rect 17036 9476 17156 9640
rect 17788 9476 17908 9640
rect 18380 9476 18500 9640
rect 19052 9476 19172 9640
rect 19724 9476 19844 9640
rect 20396 9476 20516 9640
rect 20844 9476 21044 9640
rect 21628 9476 21748 9640
rect 22076 9476 22276 9640
rect 1692 9176 1892 9340
rect 2140 9176 2340 9340
rect 2588 9176 2788 9340
rect 3372 9176 3492 9340
rect 4044 9176 4164 9340
rect 4716 9176 4836 9340
rect 5388 9176 5508 9340
rect 6060 9176 6180 9340
rect 6732 9176 6852 9340
rect 7404 9176 7524 9340
rect 8188 9176 8308 9340
rect 8860 9176 8980 9340
rect 9644 9176 9844 9340
rect 10316 9176 10436 9340
rect 10988 9176 11108 9340
rect 11660 9176 11780 9340
rect 12332 9176 12452 9340
rect 13004 9176 13124 9340
rect 13676 9176 13796 9340
rect 14348 9176 14468 9340
rect 15020 9176 15140 9340
rect 15692 9176 15812 9340
rect 16364 9176 16484 9340
rect 16812 9176 17012 9340
rect 17708 9176 17828 9340
rect 18380 9176 18500 9340
rect 19052 9176 19172 9340
rect 19724 9176 19844 9340
rect 20396 9176 20516 9340
rect 20844 9176 21044 9340
rect 21292 9176 21492 9340
rect 21740 9176 21940 9340
rect 1692 7908 1892 8072
rect 2140 7908 2340 8072
rect 2892 7908 3012 8072
rect 3484 7908 3604 8072
rect 4156 7908 4276 8072
rect 4828 7908 4948 8072
rect 5836 7908 5956 8072
rect 6508 7908 6628 8072
rect 7180 7908 7300 8072
rect 7852 7908 7972 8072
rect 8524 7908 8644 8072
rect 9196 7908 9316 8072
rect 9868 7908 9988 8072
rect 10540 7908 10660 8072
rect 11292 7908 11412 8072
rect 11660 7908 11860 8072
rect 12108 7908 12228 8072
rect 12780 7908 12900 8072
rect 13676 7908 13796 8072
rect 14348 7908 14468 8072
rect 15020 7908 15140 8072
rect 15692 7908 15812 8072
rect 16364 7908 16484 8072
rect 17036 7908 17156 8072
rect 17708 7908 17828 8072
rect 18380 7908 18500 8072
rect 19052 7908 19172 8072
rect 19724 7908 19844 8072
rect 20476 7908 20596 8072
rect 20844 7908 21044 8072
rect 21516 7908 21716 8072
rect 21964 7908 22164 8072
rect 2108 7608 2228 7772
rect 2700 7608 2820 7772
rect 3372 7608 3492 7772
rect 4044 7608 4164 7772
rect 4716 7608 4836 7772
rect 5388 7608 5508 7772
rect 6060 7608 6180 7772
rect 6732 7608 6852 7772
rect 7404 7608 7524 7772
rect 8188 7608 8308 7772
rect 8860 7608 8980 7772
rect 9868 7608 9988 7772
rect 10540 7608 10660 7772
rect 11292 7608 11412 7772
rect 11884 7608 12004 7772
rect 12556 7608 12676 7772
rect 13228 7608 13348 7772
rect 13900 7608 14020 7772
rect 14572 7608 14692 7772
rect 15244 7608 15364 7772
rect 15916 7608 16036 7772
rect 16588 7608 16708 7772
rect 17708 7608 17828 7772
rect 18380 7608 18500 7772
rect 19052 7608 19172 7772
rect 19724 7608 19844 7772
rect 20396 7608 20516 7772
rect 21068 7608 21188 7772
rect 21516 7608 21716 7772
rect 21964 7608 22164 7772
rect 1692 6340 1892 6504
rect 2140 6340 2260 6504
rect 2812 6340 2932 6504
rect 3484 6340 3604 6504
rect 4156 6340 4276 6504
rect 4828 6340 4948 6504
rect 5724 6340 5844 6504
rect 6396 6340 6516 6504
rect 7068 6340 7188 6504
rect 7740 6340 7860 6504
rect 8412 6340 8532 6504
rect 9084 6340 9204 6504
rect 9756 6340 9876 6504
rect 10428 6340 10548 6504
rect 11100 6340 11220 6504
rect 11772 6340 11892 6504
rect 12444 6340 12564 6504
rect 12892 6340 13092 6504
rect 13564 6340 13764 6504
rect 14124 6340 14244 6504
rect 14796 6340 14916 6504
rect 15468 6340 15588 6504
rect 16140 6340 16260 6504
rect 16812 6340 16932 6504
rect 17484 6340 17604 6504
rect 18156 6340 18276 6504
rect 18828 6340 18948 6504
rect 19500 6340 19620 6504
rect 20252 6340 20372 6504
rect 20620 6340 20820 6504
rect 21628 6340 21748 6504
rect 22076 6340 22276 6504
rect 2028 6040 2148 6204
rect 2700 6040 2820 6204
rect 3372 6040 3492 6204
rect 4044 6040 4164 6204
rect 4716 6040 4836 6204
rect 5388 6040 5508 6204
rect 6060 6040 6180 6204
rect 6732 6040 6852 6204
rect 7404 6040 7524 6204
rect 8076 6040 8196 6204
rect 8748 6040 8868 6204
rect 9756 6040 9876 6204
rect 10428 6040 10548 6204
rect 11100 6040 11220 6204
rect 11772 6040 11892 6204
rect 12556 6040 12676 6204
rect 13228 6040 13348 6204
rect 13900 6040 14020 6204
rect 14572 6040 14692 6204
rect 15244 6040 15364 6204
rect 15916 6040 16036 6204
rect 16588 6040 16708 6204
rect 17708 6040 17828 6204
rect 18380 6040 18500 6204
rect 19052 6040 19172 6204
rect 19724 6040 19844 6204
rect 20396 6040 20516 6204
rect 21068 6040 21188 6204
rect 21820 6040 21940 6204
rect 1692 4772 1892 4936
rect 2140 4772 2260 4936
rect 2812 4772 2932 4936
rect 3484 4772 3604 4936
rect 4156 4772 4276 4936
rect 4828 4772 4948 4936
rect 5724 4772 5844 4936
rect 6396 4772 6516 4936
rect 7068 4772 7188 4936
rect 7740 4772 7860 4936
rect 8412 4772 8532 4936
rect 9084 4772 9204 4936
rect 9756 4772 9876 4936
rect 10428 4772 10548 4936
rect 10876 4772 11076 4936
rect 11436 4772 11556 4936
rect 12108 4772 12228 4936
rect 12780 4772 12900 4936
rect 13564 4772 13764 4936
rect 14012 4772 14132 4936
rect 14684 4772 14804 4936
rect 15356 4772 15476 4936
rect 16028 4772 16148 4936
rect 16700 4772 16820 4936
rect 17372 4772 17492 4936
rect 18044 4772 18164 4936
rect 18716 4772 18836 4936
rect 19388 4772 19508 4936
rect 20060 4772 20180 4936
rect 20732 4772 20852 4936
rect 21628 4772 21748 4936
rect 22076 4772 22276 4936
rect 1692 4472 1892 4636
rect 2364 4472 2484 4636
rect 3036 4472 3156 4636
rect 3708 4472 3828 4636
rect 4380 4472 4500 4636
rect 5052 4472 5172 4636
rect 5724 4472 5844 4636
rect 6396 4472 6516 4636
rect 7068 4472 7188 4636
rect 7740 4472 7860 4636
rect 8412 4472 8532 4636
rect 8860 4472 9060 4636
rect 9756 4472 9876 4636
rect 10428 4472 10548 4636
rect 11100 4472 11220 4636
rect 11548 4472 11748 4636
rect 12332 4472 12452 4636
rect 13004 4472 13124 4636
rect 13676 4472 13796 4636
rect 14348 4472 14468 4636
rect 15020 4472 15140 4636
rect 15692 4472 15812 4636
rect 16364 4472 16484 4636
rect 16812 4472 17012 4636
rect 17708 4472 17828 4636
rect 18380 4472 18500 4636
rect 19052 4472 19172 4636
rect 19724 4472 19844 4636
rect 20396 4472 20516 4636
rect 21068 4472 21188 4636
rect 21820 4472 21940 4636
rect 1692 3204 1892 3368
rect 2140 3204 2340 3368
rect 2812 3204 2932 3368
rect 3484 3204 3604 3368
rect 4156 3204 4276 3368
rect 4828 3204 4948 3368
rect 5804 3204 5924 3368
rect 6476 3204 6596 3368
rect 7148 3204 7268 3368
rect 7740 3204 7860 3368
rect 8492 3204 8612 3368
rect 8860 3204 9060 3368
rect 9724 3204 9844 3368
rect 10316 3204 10436 3368
rect 10988 3204 11108 3368
rect 11740 3204 11860 3368
rect 12108 3204 12308 3368
rect 12556 3204 12756 3368
rect 13452 3204 13652 3368
rect 13900 3204 14020 3368
rect 14572 3204 14692 3368
rect 15244 3204 15364 3368
rect 15916 3204 16036 3368
rect 16588 3204 16708 3368
rect 17484 3204 17604 3368
rect 18156 3204 18276 3368
rect 18828 3204 18948 3368
rect 19500 3204 19620 3368
rect 20172 3204 20292 3368
rect 20620 3204 20820 3368
rect 21292 3204 21492 3368
rect 21740 3204 21940 3368
<< mvpmos >>
rect 1692 16152 1892 16396
rect 2140 16152 2340 16396
rect 2588 16152 2788 16396
rect 3036 16152 3236 16396
rect 3484 16152 3684 16396
rect 3932 16152 4132 16396
rect 4380 16152 4580 16396
rect 4828 16152 5028 16396
rect 5612 16152 5812 16396
rect 6060 16152 6260 16396
rect 6508 16152 6708 16396
rect 6956 16152 7156 16396
rect 7404 16152 7604 16396
rect 7852 16152 8052 16396
rect 8300 16152 8500 16396
rect 8748 16152 8948 16396
rect 9532 16152 9732 16396
rect 9980 16152 10180 16396
rect 10428 16152 10628 16396
rect 10876 16152 11076 16396
rect 11324 16152 11524 16396
rect 11772 16152 11972 16396
rect 12220 16152 12420 16396
rect 12668 16152 12868 16396
rect 13452 16152 13652 16396
rect 13900 16152 14100 16396
rect 14348 16152 14548 16396
rect 14796 16152 14996 16396
rect 15244 16152 15444 16396
rect 15692 16152 15892 16396
rect 16140 16152 16340 16396
rect 16588 16152 16788 16396
rect 17372 16152 17572 16396
rect 17820 16152 18020 16396
rect 18268 16152 18468 16396
rect 18716 16152 18916 16396
rect 19164 16152 19364 16396
rect 19612 16152 19812 16396
rect 20060 16152 20260 16396
rect 20508 16152 20708 16396
rect 21292 16152 21492 16396
rect 21740 16152 21940 16396
rect 1692 14964 1892 15208
rect 2140 14964 2340 15208
rect 2588 14964 2788 15208
rect 3036 14964 3236 15208
rect 3484 14964 3684 15208
rect 3932 14964 4132 15208
rect 4380 14964 4580 15208
rect 4828 14964 5028 15208
rect 5276 14964 5476 15208
rect 5724 14964 5924 15208
rect 6172 14964 6372 15208
rect 6620 14964 6820 15208
rect 7068 14964 7268 15208
rect 7516 14964 7716 15208
rect 7964 14964 8164 15208
rect 8412 14964 8612 15208
rect 8860 14964 9060 15208
rect 9644 14964 9844 15208
rect 10092 14964 10292 15208
rect 10540 14964 10740 15208
rect 10988 14964 11188 15208
rect 11436 14964 11636 15208
rect 11884 14964 12084 15208
rect 12332 14964 12532 15208
rect 12780 14964 12980 15208
rect 13228 14964 13428 15208
rect 13676 14964 13876 15208
rect 14124 14964 14324 15208
rect 14572 14964 14772 15208
rect 15020 14964 15220 15208
rect 15468 14964 15668 15208
rect 15916 14964 16116 15208
rect 16364 14964 16564 15208
rect 16812 14964 17012 15208
rect 17596 14964 17796 15208
rect 18044 14964 18244 15208
rect 18492 14964 18692 15208
rect 18940 14964 19140 15208
rect 19388 14964 19588 15208
rect 19836 14964 20036 15208
rect 20284 14964 20484 15208
rect 20732 14964 20932 15208
rect 21180 14964 21380 15208
rect 21628 14964 21828 15208
rect 22076 14964 22276 15208
rect 1692 14584 1892 14828
rect 2140 14584 2340 14828
rect 2588 14584 2788 14828
rect 3036 14584 3236 14828
rect 3484 14584 3684 14828
rect 3932 14584 4132 14828
rect 4380 14584 4580 14828
rect 4828 14584 5028 14828
rect 5612 14584 5812 14828
rect 6060 14584 6260 14828
rect 6508 14584 6708 14828
rect 6956 14584 7156 14828
rect 7404 14584 7604 14828
rect 7852 14584 8052 14828
rect 8300 14584 8500 14828
rect 8748 14584 8948 14828
rect 9196 14584 9396 14828
rect 9644 14584 9844 14828
rect 10092 14584 10292 14828
rect 10540 14584 10740 14828
rect 10988 14584 11188 14828
rect 11436 14584 11636 14828
rect 11884 14584 12084 14828
rect 12332 14584 12532 14828
rect 12780 14584 12980 14828
rect 13564 14584 13764 14828
rect 14012 14584 14212 14828
rect 14460 14584 14660 14828
rect 14908 14584 15108 14828
rect 15356 14584 15556 14828
rect 15804 14584 16004 14828
rect 16252 14584 16452 14828
rect 16892 14584 16992 14828
rect 17564 14584 17664 14828
rect 17932 14584 18132 14828
rect 18380 14584 18580 14828
rect 18828 14584 19028 14828
rect 19276 14584 19476 14828
rect 19724 14584 19924 14828
rect 20172 14584 20372 14828
rect 20620 14584 20820 14828
rect 21516 14584 21716 14828
rect 21964 14584 22164 14828
rect 1692 13396 1892 13640
rect 2140 13396 2340 13640
rect 2588 13396 2788 13640
rect 3036 13396 3236 13640
rect 3484 13396 3684 13640
rect 3932 13396 4132 13640
rect 4380 13396 4580 13640
rect 4828 13396 5028 13640
rect 5276 13396 5476 13640
rect 5724 13396 5924 13640
rect 6172 13396 6372 13640
rect 6620 13396 6820 13640
rect 7068 13396 7268 13640
rect 7516 13396 7716 13640
rect 7964 13396 8164 13640
rect 8412 13396 8612 13640
rect 8860 13396 9060 13640
rect 9644 13396 9844 13640
rect 10092 13396 10292 13640
rect 10540 13396 10740 13640
rect 10988 13396 11188 13640
rect 11436 13396 11636 13640
rect 11884 13396 12084 13640
rect 12332 13396 12532 13640
rect 12780 13396 12980 13640
rect 13228 13396 13428 13640
rect 13676 13396 13876 13640
rect 14124 13396 14324 13640
rect 14572 13396 14772 13640
rect 15020 13396 15220 13640
rect 15468 13396 15668 13640
rect 16160 13396 16260 13640
rect 16832 13396 16932 13640
rect 17728 13396 17828 13640
rect 18400 13396 18500 13640
rect 18828 13396 19028 13640
rect 19276 13396 19476 13640
rect 19724 13396 19924 13640
rect 20172 13396 20372 13640
rect 20620 13396 20820 13640
rect 21068 13396 21268 13640
rect 21516 13396 21716 13640
rect 21964 13396 22164 13640
rect 1692 13016 1892 13260
rect 2140 13016 2340 13260
rect 2588 13016 2788 13260
rect 3036 13016 3236 13260
rect 3484 13016 3684 13260
rect 3932 13016 4132 13260
rect 4380 13016 4580 13260
rect 4828 13016 5028 13260
rect 5612 13016 5812 13260
rect 6060 13016 6260 13260
rect 6508 13016 6708 13260
rect 6956 13016 7156 13260
rect 7404 13016 7604 13260
rect 7852 13016 8052 13260
rect 8300 13016 8500 13260
rect 8748 13016 8948 13260
rect 9196 13016 9396 13260
rect 9644 13016 9844 13260
rect 10092 13016 10292 13260
rect 10540 13016 10740 13260
rect 10988 13016 11188 13260
rect 11436 13016 11636 13260
rect 11884 13016 12084 13260
rect 12332 13016 12532 13260
rect 12780 13016 12980 13260
rect 13564 13016 13764 13260
rect 14012 13016 14212 13260
rect 14816 13016 14916 13260
rect 15488 13016 15588 13260
rect 16160 13016 16260 13260
rect 16832 13016 16932 13260
rect 17504 13016 17604 13260
rect 18176 13016 18276 13260
rect 18848 13016 18948 13260
rect 19520 13016 19620 13260
rect 19948 13016 20148 13260
rect 20396 13016 20596 13260
rect 20844 13016 21044 13260
rect 21516 13016 21716 13260
rect 21964 13016 22164 13260
rect 1692 11828 1892 12072
rect 2140 11828 2340 12072
rect 2588 11828 2788 12072
rect 3036 11828 3236 12072
rect 3484 11828 3684 12072
rect 3932 11828 4132 12072
rect 4380 11828 4580 12072
rect 4828 11828 5028 12072
rect 5276 11828 5476 12072
rect 5724 11828 5924 12072
rect 6172 11828 6372 12072
rect 6620 11828 6820 12072
rect 7068 11828 7268 12072
rect 7516 11828 7716 12072
rect 7964 11828 8164 12072
rect 8412 11828 8612 12072
rect 8860 11828 9060 12072
rect 9644 11828 9844 12072
rect 10092 11828 10292 12072
rect 10540 11828 10740 12072
rect 10988 11828 11188 12072
rect 11436 11828 11636 12072
rect 11884 11828 12084 12072
rect 12332 11828 12532 12072
rect 12780 11828 12980 12072
rect 13228 11828 13428 12072
rect 13676 11828 13876 12072
rect 14144 11828 14244 12072
rect 14816 11828 14916 12072
rect 15488 11828 15588 12072
rect 16160 11828 16260 12072
rect 16832 11828 16932 12072
rect 17728 11828 17828 12072
rect 18400 11828 18500 12072
rect 19072 11828 19172 12072
rect 19744 11828 19844 12072
rect 20416 11828 20516 12072
rect 20844 11828 21044 12072
rect 21292 11828 21492 12072
rect 21740 11828 21940 12072
rect 1692 11448 1892 11692
rect 2140 11448 2340 11692
rect 2588 11448 2788 11692
rect 3036 11448 3236 11692
rect 3484 11448 3684 11692
rect 3932 11448 4132 11692
rect 4380 11448 4580 11692
rect 4828 11448 5028 11692
rect 5612 11448 5812 11692
rect 6140 11448 6240 11692
rect 6924 11448 7024 11692
rect 7596 11448 7696 11692
rect 8268 11448 8368 11692
rect 8636 11448 8836 11692
rect 9216 11448 9316 11692
rect 9888 11448 9988 11692
rect 10560 11448 10660 11692
rect 10988 11448 11188 11692
rect 11436 11448 11636 11692
rect 12128 11448 12228 11692
rect 12800 11448 12900 11692
rect 13696 11448 13796 11692
rect 14124 11448 14324 11692
rect 14816 11448 14916 11692
rect 15488 11448 15588 11692
rect 16160 11448 16260 11692
rect 16832 11448 16932 11692
rect 17504 11448 17604 11692
rect 18176 11448 18276 11692
rect 18848 11448 18948 11692
rect 19520 11448 19620 11692
rect 20192 11448 20292 11692
rect 20620 11448 20820 11692
rect 21516 11448 21716 11692
rect 21964 11448 22164 11692
rect 1692 10260 1892 10504
rect 2140 10260 2340 10504
rect 2588 10260 2788 10504
rect 3036 10260 3236 10504
rect 3484 10260 3684 10504
rect 3932 10260 4132 10504
rect 4380 10260 4580 10504
rect 4828 10260 5028 10504
rect 5408 10260 5508 10504
rect 6080 10260 6180 10504
rect 6752 10260 6852 10504
rect 7424 10260 7524 10504
rect 8096 10260 8196 10504
rect 8880 10260 8980 10504
rect 9888 10260 9988 10504
rect 10560 10260 10660 10504
rect 11232 10260 11332 10504
rect 12016 10260 12116 10504
rect 12688 10260 12788 10504
rect 13360 10260 13460 10504
rect 14032 10260 14132 10504
rect 14704 10260 14804 10504
rect 15376 10260 15476 10504
rect 16048 10260 16148 10504
rect 16720 10260 16820 10504
rect 17728 10260 17828 10504
rect 18400 10260 18500 10504
rect 19072 10260 19172 10504
rect 19744 10260 19844 10504
rect 20416 10260 20516 10504
rect 21088 10260 21188 10504
rect 21760 10260 21860 10504
rect 1692 9880 1892 10124
rect 2140 9880 2340 10124
rect 2588 9880 2788 10124
rect 3036 9880 3236 10124
rect 3484 9880 3684 10124
rect 4176 9880 4276 10124
rect 4848 9880 4948 10124
rect 5856 9880 5956 10124
rect 6528 9880 6628 10124
rect 7200 9880 7300 10124
rect 7872 9880 7972 10124
rect 8544 9880 8644 10124
rect 9216 9880 9316 10124
rect 9888 9880 9988 10124
rect 10560 9880 10660 10124
rect 10988 9880 11188 10124
rect 11456 9880 11556 10124
rect 12128 9880 12228 10124
rect 12800 9880 12900 10124
rect 13696 9880 13796 10124
rect 14368 9880 14468 10124
rect 15040 9880 15140 10124
rect 15712 9880 15812 10124
rect 16384 9880 16484 10124
rect 17056 9880 17156 10124
rect 17788 9880 17888 10124
rect 18400 9880 18500 10124
rect 19072 9880 19172 10124
rect 19744 9880 19844 10124
rect 20416 9880 20516 10124
rect 20844 9880 21044 10124
rect 21648 9880 21748 10124
rect 22076 9880 22276 10124
rect 1692 8692 1892 8936
rect 2140 8692 2340 8936
rect 2588 8692 2788 8936
rect 3392 8692 3492 8936
rect 4064 8692 4164 8936
rect 4736 8692 4836 8936
rect 5408 8692 5508 8936
rect 6080 8692 6180 8936
rect 6752 8692 6852 8936
rect 7424 8692 7524 8936
rect 8208 8692 8308 8936
rect 8880 8692 8980 8936
rect 9644 8692 9844 8936
rect 10336 8692 10436 8936
rect 11008 8692 11108 8936
rect 11680 8692 11780 8936
rect 12352 8692 12452 8936
rect 13024 8692 13124 8936
rect 13696 8692 13796 8936
rect 14368 8692 14468 8936
rect 15040 8692 15140 8936
rect 15712 8692 15812 8936
rect 16384 8692 16484 8936
rect 16812 8692 17012 8936
rect 17728 8692 17828 8936
rect 18400 8692 18500 8936
rect 19072 8692 19172 8936
rect 19744 8692 19844 8936
rect 20416 8692 20516 8936
rect 20844 8692 21044 8936
rect 21292 8692 21492 8936
rect 21740 8692 21940 8936
rect 1692 8312 1892 8556
rect 2140 8312 2340 8556
rect 2892 8312 2992 8556
rect 3504 8312 3604 8556
rect 4176 8312 4276 8556
rect 4848 8312 4948 8556
rect 5856 8312 5956 8556
rect 6528 8312 6628 8556
rect 7200 8312 7300 8556
rect 7872 8312 7972 8556
rect 8544 8312 8644 8556
rect 9216 8312 9316 8556
rect 9888 8312 9988 8556
rect 10560 8312 10660 8556
rect 11292 8312 11392 8556
rect 11660 8312 11860 8556
rect 12128 8312 12228 8556
rect 12800 8312 12900 8556
rect 13696 8312 13796 8556
rect 14368 8312 14468 8556
rect 15040 8312 15140 8556
rect 15712 8312 15812 8556
rect 16384 8312 16484 8556
rect 17056 8312 17156 8556
rect 17728 8312 17828 8556
rect 18400 8312 18500 8556
rect 19072 8312 19172 8556
rect 19744 8312 19844 8556
rect 20476 8312 20576 8556
rect 20844 8312 21044 8556
rect 21516 8312 21716 8556
rect 21964 8312 22164 8556
rect 2108 7124 2208 7368
rect 2720 7124 2820 7368
rect 3392 7124 3492 7368
rect 4064 7124 4164 7368
rect 4736 7124 4836 7368
rect 5408 7124 5508 7368
rect 6080 7124 6180 7368
rect 6752 7124 6852 7368
rect 7424 7124 7524 7368
rect 8208 7124 8308 7368
rect 8880 7124 8980 7368
rect 9888 7124 9988 7368
rect 10560 7124 10660 7368
rect 11292 7124 11392 7368
rect 11904 7124 12004 7368
rect 12576 7124 12676 7368
rect 13248 7124 13348 7368
rect 13920 7124 14020 7368
rect 14592 7124 14692 7368
rect 15264 7124 15364 7368
rect 15936 7124 16036 7368
rect 16608 7124 16708 7368
rect 17728 7124 17828 7368
rect 18400 7124 18500 7368
rect 19072 7124 19172 7368
rect 19744 7124 19844 7368
rect 20416 7124 20516 7368
rect 21088 7124 21188 7368
rect 21516 7124 21716 7368
rect 21964 7124 22164 7368
rect 1692 6744 1892 6988
rect 2160 6744 2260 6988
rect 2832 6744 2932 6988
rect 3504 6744 3604 6988
rect 4176 6744 4276 6988
rect 4848 6744 4948 6988
rect 5744 6744 5844 6988
rect 6416 6744 6516 6988
rect 7088 6744 7188 6988
rect 7760 6744 7860 6988
rect 8432 6744 8532 6988
rect 9104 6744 9204 6988
rect 9776 6744 9876 6988
rect 10448 6744 10548 6988
rect 11120 6744 11220 6988
rect 11792 6744 11892 6988
rect 12464 6744 12564 6988
rect 12892 6744 13092 6988
rect 13564 6744 13764 6988
rect 14144 6744 14244 6988
rect 14816 6744 14916 6988
rect 15488 6744 15588 6988
rect 16160 6744 16260 6988
rect 16832 6744 16932 6988
rect 17504 6744 17604 6988
rect 18176 6744 18276 6988
rect 18848 6744 18948 6988
rect 19520 6744 19620 6988
rect 20252 6744 20352 6988
rect 20620 6744 20820 6988
rect 21648 6744 21748 6988
rect 22076 6744 22276 6988
rect 2048 5556 2148 5800
rect 2720 5556 2820 5800
rect 3392 5556 3492 5800
rect 4064 5556 4164 5800
rect 4736 5556 4836 5800
rect 5408 5556 5508 5800
rect 6080 5556 6180 5800
rect 6752 5556 6852 5800
rect 7424 5556 7524 5800
rect 8096 5556 8196 5800
rect 8768 5556 8868 5800
rect 9776 5556 9876 5800
rect 10448 5556 10548 5800
rect 11120 5556 11220 5800
rect 11792 5556 11892 5800
rect 12576 5556 12676 5800
rect 13248 5556 13348 5800
rect 13920 5556 14020 5800
rect 14592 5556 14692 5800
rect 15264 5556 15364 5800
rect 15936 5556 16036 5800
rect 16608 5556 16708 5800
rect 17728 5556 17828 5800
rect 18400 5556 18500 5800
rect 19072 5556 19172 5800
rect 19744 5556 19844 5800
rect 20416 5556 20516 5800
rect 21088 5556 21188 5800
rect 21820 5556 21920 5800
rect 1692 5176 1892 5420
rect 2160 5176 2260 5420
rect 2832 5176 2932 5420
rect 3504 5176 3604 5420
rect 4176 5176 4276 5420
rect 4848 5176 4948 5420
rect 5744 5176 5844 5420
rect 6416 5176 6516 5420
rect 7088 5176 7188 5420
rect 7760 5176 7860 5420
rect 8432 5176 8532 5420
rect 9104 5176 9204 5420
rect 9776 5176 9876 5420
rect 10448 5176 10548 5420
rect 10876 5176 11076 5420
rect 11456 5176 11556 5420
rect 12128 5176 12228 5420
rect 12800 5176 12900 5420
rect 13564 5176 13764 5420
rect 14032 5176 14132 5420
rect 14704 5176 14804 5420
rect 15376 5176 15476 5420
rect 16048 5176 16148 5420
rect 16720 5176 16820 5420
rect 17392 5176 17492 5420
rect 18064 5176 18164 5420
rect 18736 5176 18836 5420
rect 19408 5176 19508 5420
rect 20080 5176 20180 5420
rect 20752 5176 20852 5420
rect 21648 5176 21748 5420
rect 22076 5176 22276 5420
rect 1692 3988 1892 4232
rect 2384 3988 2484 4232
rect 3056 3988 3156 4232
rect 3728 3988 3828 4232
rect 4400 3988 4500 4232
rect 5072 3988 5172 4232
rect 5744 3988 5844 4232
rect 6416 3988 6516 4232
rect 7088 3988 7188 4232
rect 7760 3988 7860 4232
rect 8432 3988 8532 4232
rect 8860 3988 9060 4232
rect 9776 3988 9876 4232
rect 10448 3988 10548 4232
rect 11120 3988 11220 4232
rect 11548 3988 11748 4232
rect 12352 3988 12452 4232
rect 13024 3988 13124 4232
rect 13696 3988 13796 4232
rect 14368 3988 14468 4232
rect 15040 3988 15140 4232
rect 15712 3988 15812 4232
rect 16384 3988 16484 4232
rect 16812 3988 17012 4232
rect 17728 3988 17828 4232
rect 18400 3988 18500 4232
rect 19072 3988 19172 4232
rect 19744 3988 19844 4232
rect 20416 3988 20516 4232
rect 21088 3988 21188 4232
rect 21820 3988 21920 4232
rect 1692 3608 1892 3852
rect 2140 3608 2340 3852
rect 2832 3608 2932 3852
rect 3504 3608 3604 3852
rect 4176 3608 4276 3852
rect 4848 3608 4948 3852
rect 5804 3608 5904 3852
rect 6476 3608 6576 3852
rect 7148 3608 7248 3852
rect 7760 3608 7860 3852
rect 8492 3608 8592 3852
rect 8860 3608 9060 3852
rect 9724 3608 9824 3852
rect 10336 3608 10436 3852
rect 11008 3608 11108 3852
rect 11740 3608 11840 3852
rect 12108 3608 12308 3852
rect 12556 3608 12756 3852
rect 13452 3608 13652 3852
rect 13920 3608 14020 3852
rect 14592 3608 14692 3852
rect 15264 3608 15364 3852
rect 15936 3608 16036 3852
rect 16608 3608 16708 3852
rect 17504 3608 17604 3852
rect 18176 3608 18276 3852
rect 18848 3608 18948 3852
rect 19520 3608 19620 3852
rect 20192 3608 20292 3852
rect 20620 3608 20820 3852
rect 21292 3608 21492 3852
rect 21740 3608 21940 3852
<< mvndiff >>
rect 1604 15872 1692 15912
rect 1604 15826 1617 15872
rect 1663 15826 1692 15872
rect 1604 15748 1692 15826
rect 1892 15872 1980 15912
rect 1892 15826 1921 15872
rect 1967 15826 1980 15872
rect 1892 15748 1980 15826
rect 2052 15872 2140 15912
rect 2052 15826 2065 15872
rect 2111 15826 2140 15872
rect 2052 15748 2140 15826
rect 2340 15872 2428 15912
rect 2340 15826 2369 15872
rect 2415 15826 2428 15872
rect 2340 15748 2428 15826
rect 2500 15872 2588 15912
rect 2500 15826 2513 15872
rect 2559 15826 2588 15872
rect 2500 15748 2588 15826
rect 2788 15872 2876 15912
rect 2788 15826 2817 15872
rect 2863 15826 2876 15872
rect 2788 15748 2876 15826
rect 2948 15872 3036 15912
rect 2948 15826 2961 15872
rect 3007 15826 3036 15872
rect 2948 15748 3036 15826
rect 3236 15872 3324 15912
rect 3236 15826 3265 15872
rect 3311 15826 3324 15872
rect 3236 15748 3324 15826
rect 3396 15872 3484 15912
rect 3396 15826 3409 15872
rect 3455 15826 3484 15872
rect 3396 15748 3484 15826
rect 3684 15872 3772 15912
rect 3684 15826 3713 15872
rect 3759 15826 3772 15872
rect 3684 15748 3772 15826
rect 3844 15872 3932 15912
rect 3844 15826 3857 15872
rect 3903 15826 3932 15872
rect 3844 15748 3932 15826
rect 4132 15872 4220 15912
rect 4132 15826 4161 15872
rect 4207 15826 4220 15872
rect 4132 15748 4220 15826
rect 4292 15872 4380 15912
rect 4292 15826 4305 15872
rect 4351 15826 4380 15872
rect 4292 15748 4380 15826
rect 4580 15872 4668 15912
rect 4580 15826 4609 15872
rect 4655 15826 4668 15872
rect 4580 15748 4668 15826
rect 4740 15872 4828 15912
rect 4740 15826 4753 15872
rect 4799 15826 4828 15872
rect 4740 15748 4828 15826
rect 5028 15872 5116 15912
rect 5028 15826 5057 15872
rect 5103 15826 5116 15872
rect 5028 15748 5116 15826
rect 5524 15872 5612 15912
rect 5524 15826 5537 15872
rect 5583 15826 5612 15872
rect 5524 15748 5612 15826
rect 5812 15872 5900 15912
rect 5812 15826 5841 15872
rect 5887 15826 5900 15872
rect 5812 15748 5900 15826
rect 5972 15872 6060 15912
rect 5972 15826 5985 15872
rect 6031 15826 6060 15872
rect 5972 15748 6060 15826
rect 6260 15872 6348 15912
rect 6260 15826 6289 15872
rect 6335 15826 6348 15872
rect 6260 15748 6348 15826
rect 6420 15872 6508 15912
rect 6420 15826 6433 15872
rect 6479 15826 6508 15872
rect 6420 15748 6508 15826
rect 6708 15872 6796 15912
rect 6708 15826 6737 15872
rect 6783 15826 6796 15872
rect 6708 15748 6796 15826
rect 6868 15872 6956 15912
rect 6868 15826 6881 15872
rect 6927 15826 6956 15872
rect 6868 15748 6956 15826
rect 7156 15872 7244 15912
rect 7156 15826 7185 15872
rect 7231 15826 7244 15872
rect 7156 15748 7244 15826
rect 7316 15872 7404 15912
rect 7316 15826 7329 15872
rect 7375 15826 7404 15872
rect 7316 15748 7404 15826
rect 7604 15872 7692 15912
rect 7604 15826 7633 15872
rect 7679 15826 7692 15872
rect 7604 15748 7692 15826
rect 7764 15872 7852 15912
rect 7764 15826 7777 15872
rect 7823 15826 7852 15872
rect 7764 15748 7852 15826
rect 8052 15872 8140 15912
rect 8052 15826 8081 15872
rect 8127 15826 8140 15872
rect 8052 15748 8140 15826
rect 8212 15872 8300 15912
rect 8212 15826 8225 15872
rect 8271 15826 8300 15872
rect 8212 15748 8300 15826
rect 8500 15872 8588 15912
rect 8500 15826 8529 15872
rect 8575 15826 8588 15872
rect 8500 15748 8588 15826
rect 8660 15872 8748 15912
rect 8660 15826 8673 15872
rect 8719 15826 8748 15872
rect 8660 15748 8748 15826
rect 8948 15872 9036 15912
rect 8948 15826 8977 15872
rect 9023 15826 9036 15872
rect 8948 15748 9036 15826
rect 9444 15872 9532 15912
rect 9444 15826 9457 15872
rect 9503 15826 9532 15872
rect 9444 15748 9532 15826
rect 9732 15872 9820 15912
rect 9732 15826 9761 15872
rect 9807 15826 9820 15872
rect 9732 15748 9820 15826
rect 9892 15872 9980 15912
rect 9892 15826 9905 15872
rect 9951 15826 9980 15872
rect 9892 15748 9980 15826
rect 10180 15872 10268 15912
rect 10180 15826 10209 15872
rect 10255 15826 10268 15872
rect 10180 15748 10268 15826
rect 10340 15872 10428 15912
rect 10340 15826 10353 15872
rect 10399 15826 10428 15872
rect 10340 15748 10428 15826
rect 10628 15872 10716 15912
rect 10628 15826 10657 15872
rect 10703 15826 10716 15872
rect 10628 15748 10716 15826
rect 10788 15872 10876 15912
rect 10788 15826 10801 15872
rect 10847 15826 10876 15872
rect 10788 15748 10876 15826
rect 11076 15872 11164 15912
rect 11076 15826 11105 15872
rect 11151 15826 11164 15872
rect 11076 15748 11164 15826
rect 11236 15872 11324 15912
rect 11236 15826 11249 15872
rect 11295 15826 11324 15872
rect 11236 15748 11324 15826
rect 11524 15872 11612 15912
rect 11524 15826 11553 15872
rect 11599 15826 11612 15872
rect 11524 15748 11612 15826
rect 11684 15872 11772 15912
rect 11684 15826 11697 15872
rect 11743 15826 11772 15872
rect 11684 15748 11772 15826
rect 11972 15872 12060 15912
rect 11972 15826 12001 15872
rect 12047 15826 12060 15872
rect 11972 15748 12060 15826
rect 12132 15872 12220 15912
rect 12132 15826 12145 15872
rect 12191 15826 12220 15872
rect 12132 15748 12220 15826
rect 12420 15872 12508 15912
rect 12420 15826 12449 15872
rect 12495 15826 12508 15872
rect 12420 15748 12508 15826
rect 12580 15872 12668 15912
rect 12580 15826 12593 15872
rect 12639 15826 12668 15872
rect 12580 15748 12668 15826
rect 12868 15872 12956 15912
rect 12868 15826 12897 15872
rect 12943 15826 12956 15872
rect 12868 15748 12956 15826
rect 13364 15872 13452 15912
rect 13364 15826 13377 15872
rect 13423 15826 13452 15872
rect 13364 15748 13452 15826
rect 13652 15872 13740 15912
rect 13652 15826 13681 15872
rect 13727 15826 13740 15872
rect 13652 15748 13740 15826
rect 13812 15872 13900 15912
rect 13812 15826 13825 15872
rect 13871 15826 13900 15872
rect 13812 15748 13900 15826
rect 14100 15872 14188 15912
rect 14100 15826 14129 15872
rect 14175 15826 14188 15872
rect 14100 15748 14188 15826
rect 14260 15872 14348 15912
rect 14260 15826 14273 15872
rect 14319 15826 14348 15872
rect 14260 15748 14348 15826
rect 14548 15872 14636 15912
rect 14548 15826 14577 15872
rect 14623 15826 14636 15872
rect 14548 15748 14636 15826
rect 14708 15872 14796 15912
rect 14708 15826 14721 15872
rect 14767 15826 14796 15872
rect 14708 15748 14796 15826
rect 14996 15872 15084 15912
rect 14996 15826 15025 15872
rect 15071 15826 15084 15872
rect 14996 15748 15084 15826
rect 15156 15872 15244 15912
rect 15156 15826 15169 15872
rect 15215 15826 15244 15872
rect 15156 15748 15244 15826
rect 15444 15872 15532 15912
rect 15444 15826 15473 15872
rect 15519 15826 15532 15872
rect 15444 15748 15532 15826
rect 15604 15872 15692 15912
rect 15604 15826 15617 15872
rect 15663 15826 15692 15872
rect 15604 15748 15692 15826
rect 15892 15872 15980 15912
rect 15892 15826 15921 15872
rect 15967 15826 15980 15872
rect 15892 15748 15980 15826
rect 16052 15872 16140 15912
rect 16052 15826 16065 15872
rect 16111 15826 16140 15872
rect 16052 15748 16140 15826
rect 16340 15872 16428 15912
rect 16340 15826 16369 15872
rect 16415 15826 16428 15872
rect 16340 15748 16428 15826
rect 16500 15872 16588 15912
rect 16500 15826 16513 15872
rect 16559 15826 16588 15872
rect 16500 15748 16588 15826
rect 16788 15872 16876 15912
rect 16788 15826 16817 15872
rect 16863 15826 16876 15872
rect 16788 15748 16876 15826
rect 17284 15872 17372 15912
rect 17284 15826 17297 15872
rect 17343 15826 17372 15872
rect 17284 15748 17372 15826
rect 17572 15872 17660 15912
rect 17572 15826 17601 15872
rect 17647 15826 17660 15872
rect 17572 15748 17660 15826
rect 17732 15872 17820 15912
rect 17732 15826 17745 15872
rect 17791 15826 17820 15872
rect 17732 15748 17820 15826
rect 18020 15872 18108 15912
rect 18020 15826 18049 15872
rect 18095 15826 18108 15872
rect 18020 15748 18108 15826
rect 18180 15872 18268 15912
rect 18180 15826 18193 15872
rect 18239 15826 18268 15872
rect 18180 15748 18268 15826
rect 18468 15872 18556 15912
rect 18468 15826 18497 15872
rect 18543 15826 18556 15872
rect 18468 15748 18556 15826
rect 18628 15872 18716 15912
rect 18628 15826 18641 15872
rect 18687 15826 18716 15872
rect 18628 15748 18716 15826
rect 18916 15872 19004 15912
rect 18916 15826 18945 15872
rect 18991 15826 19004 15872
rect 18916 15748 19004 15826
rect 19076 15872 19164 15912
rect 19076 15826 19089 15872
rect 19135 15826 19164 15872
rect 19076 15748 19164 15826
rect 19364 15872 19452 15912
rect 19364 15826 19393 15872
rect 19439 15826 19452 15872
rect 19364 15748 19452 15826
rect 19524 15872 19612 15912
rect 19524 15826 19537 15872
rect 19583 15826 19612 15872
rect 19524 15748 19612 15826
rect 19812 15872 19900 15912
rect 19812 15826 19841 15872
rect 19887 15826 19900 15872
rect 19812 15748 19900 15826
rect 19972 15872 20060 15912
rect 19972 15826 19985 15872
rect 20031 15826 20060 15872
rect 19972 15748 20060 15826
rect 20260 15872 20348 15912
rect 20260 15826 20289 15872
rect 20335 15826 20348 15872
rect 20260 15748 20348 15826
rect 20420 15872 20508 15912
rect 20420 15826 20433 15872
rect 20479 15826 20508 15872
rect 20420 15748 20508 15826
rect 20708 15872 20796 15912
rect 20708 15826 20737 15872
rect 20783 15826 20796 15872
rect 20708 15748 20796 15826
rect 21204 15872 21292 15912
rect 21204 15826 21217 15872
rect 21263 15826 21292 15872
rect 21204 15748 21292 15826
rect 21492 15872 21580 15912
rect 21492 15826 21521 15872
rect 21567 15826 21580 15872
rect 21492 15748 21580 15826
rect 21652 15872 21740 15912
rect 21652 15826 21665 15872
rect 21711 15826 21740 15872
rect 21652 15748 21740 15826
rect 21940 15872 22028 15912
rect 21940 15826 21969 15872
rect 22015 15826 22028 15872
rect 21940 15748 22028 15826
rect 1604 15534 1692 15612
rect 1604 15488 1617 15534
rect 1663 15488 1692 15534
rect 1604 15448 1692 15488
rect 1892 15534 1980 15612
rect 1892 15488 1921 15534
rect 1967 15488 1980 15534
rect 1892 15448 1980 15488
rect 2052 15534 2140 15612
rect 2052 15488 2065 15534
rect 2111 15488 2140 15534
rect 2052 15448 2140 15488
rect 2340 15534 2428 15612
rect 2340 15488 2369 15534
rect 2415 15488 2428 15534
rect 2340 15448 2428 15488
rect 2500 15534 2588 15612
rect 2500 15488 2513 15534
rect 2559 15488 2588 15534
rect 2500 15448 2588 15488
rect 2788 15534 2876 15612
rect 2788 15488 2817 15534
rect 2863 15488 2876 15534
rect 2788 15448 2876 15488
rect 2948 15534 3036 15612
rect 2948 15488 2961 15534
rect 3007 15488 3036 15534
rect 2948 15448 3036 15488
rect 3236 15534 3324 15612
rect 3236 15488 3265 15534
rect 3311 15488 3324 15534
rect 3236 15448 3324 15488
rect 3396 15534 3484 15612
rect 3396 15488 3409 15534
rect 3455 15488 3484 15534
rect 3396 15448 3484 15488
rect 3684 15534 3772 15612
rect 3684 15488 3713 15534
rect 3759 15488 3772 15534
rect 3684 15448 3772 15488
rect 3844 15534 3932 15612
rect 3844 15488 3857 15534
rect 3903 15488 3932 15534
rect 3844 15448 3932 15488
rect 4132 15534 4220 15612
rect 4132 15488 4161 15534
rect 4207 15488 4220 15534
rect 4132 15448 4220 15488
rect 4292 15534 4380 15612
rect 4292 15488 4305 15534
rect 4351 15488 4380 15534
rect 4292 15448 4380 15488
rect 4580 15534 4668 15612
rect 4580 15488 4609 15534
rect 4655 15488 4668 15534
rect 4580 15448 4668 15488
rect 4740 15534 4828 15612
rect 4740 15488 4753 15534
rect 4799 15488 4828 15534
rect 4740 15448 4828 15488
rect 5028 15534 5116 15612
rect 5028 15488 5057 15534
rect 5103 15488 5116 15534
rect 5028 15448 5116 15488
rect 5188 15534 5276 15612
rect 5188 15488 5201 15534
rect 5247 15488 5276 15534
rect 5188 15448 5276 15488
rect 5476 15534 5564 15612
rect 5476 15488 5505 15534
rect 5551 15488 5564 15534
rect 5476 15448 5564 15488
rect 5636 15534 5724 15612
rect 5636 15488 5649 15534
rect 5695 15488 5724 15534
rect 5636 15448 5724 15488
rect 5924 15534 6012 15612
rect 5924 15488 5953 15534
rect 5999 15488 6012 15534
rect 5924 15448 6012 15488
rect 6084 15534 6172 15612
rect 6084 15488 6097 15534
rect 6143 15488 6172 15534
rect 6084 15448 6172 15488
rect 6372 15534 6460 15612
rect 6372 15488 6401 15534
rect 6447 15488 6460 15534
rect 6372 15448 6460 15488
rect 6532 15534 6620 15612
rect 6532 15488 6545 15534
rect 6591 15488 6620 15534
rect 6532 15448 6620 15488
rect 6820 15534 6908 15612
rect 6820 15488 6849 15534
rect 6895 15488 6908 15534
rect 6820 15448 6908 15488
rect 6980 15534 7068 15612
rect 6980 15488 6993 15534
rect 7039 15488 7068 15534
rect 6980 15448 7068 15488
rect 7268 15534 7356 15612
rect 7268 15488 7297 15534
rect 7343 15488 7356 15534
rect 7268 15448 7356 15488
rect 7428 15534 7516 15612
rect 7428 15488 7441 15534
rect 7487 15488 7516 15534
rect 7428 15448 7516 15488
rect 7716 15534 7804 15612
rect 7716 15488 7745 15534
rect 7791 15488 7804 15534
rect 7716 15448 7804 15488
rect 7876 15534 7964 15612
rect 7876 15488 7889 15534
rect 7935 15488 7964 15534
rect 7876 15448 7964 15488
rect 8164 15534 8252 15612
rect 8164 15488 8193 15534
rect 8239 15488 8252 15534
rect 8164 15448 8252 15488
rect 8324 15534 8412 15612
rect 8324 15488 8337 15534
rect 8383 15488 8412 15534
rect 8324 15448 8412 15488
rect 8612 15534 8700 15612
rect 8612 15488 8641 15534
rect 8687 15488 8700 15534
rect 8612 15448 8700 15488
rect 8772 15534 8860 15612
rect 8772 15488 8785 15534
rect 8831 15488 8860 15534
rect 8772 15448 8860 15488
rect 9060 15534 9148 15612
rect 9060 15488 9089 15534
rect 9135 15488 9148 15534
rect 9060 15448 9148 15488
rect 9556 15534 9644 15612
rect 9556 15488 9569 15534
rect 9615 15488 9644 15534
rect 9556 15448 9644 15488
rect 9844 15534 9932 15612
rect 9844 15488 9873 15534
rect 9919 15488 9932 15534
rect 9844 15448 9932 15488
rect 10004 15534 10092 15612
rect 10004 15488 10017 15534
rect 10063 15488 10092 15534
rect 10004 15448 10092 15488
rect 10292 15534 10380 15612
rect 10292 15488 10321 15534
rect 10367 15488 10380 15534
rect 10292 15448 10380 15488
rect 10452 15534 10540 15612
rect 10452 15488 10465 15534
rect 10511 15488 10540 15534
rect 10452 15448 10540 15488
rect 10740 15534 10828 15612
rect 10740 15488 10769 15534
rect 10815 15488 10828 15534
rect 10740 15448 10828 15488
rect 10900 15534 10988 15612
rect 10900 15488 10913 15534
rect 10959 15488 10988 15534
rect 10900 15448 10988 15488
rect 11188 15534 11276 15612
rect 11188 15488 11217 15534
rect 11263 15488 11276 15534
rect 11188 15448 11276 15488
rect 11348 15534 11436 15612
rect 11348 15488 11361 15534
rect 11407 15488 11436 15534
rect 11348 15448 11436 15488
rect 11636 15534 11724 15612
rect 11636 15488 11665 15534
rect 11711 15488 11724 15534
rect 11636 15448 11724 15488
rect 11796 15534 11884 15612
rect 11796 15488 11809 15534
rect 11855 15488 11884 15534
rect 11796 15448 11884 15488
rect 12084 15534 12172 15612
rect 12084 15488 12113 15534
rect 12159 15488 12172 15534
rect 12084 15448 12172 15488
rect 12244 15534 12332 15612
rect 12244 15488 12257 15534
rect 12303 15488 12332 15534
rect 12244 15448 12332 15488
rect 12532 15534 12620 15612
rect 12532 15488 12561 15534
rect 12607 15488 12620 15534
rect 12532 15448 12620 15488
rect 12692 15534 12780 15612
rect 12692 15488 12705 15534
rect 12751 15488 12780 15534
rect 12692 15448 12780 15488
rect 12980 15534 13068 15612
rect 12980 15488 13009 15534
rect 13055 15488 13068 15534
rect 12980 15448 13068 15488
rect 13140 15534 13228 15612
rect 13140 15488 13153 15534
rect 13199 15488 13228 15534
rect 13140 15448 13228 15488
rect 13428 15534 13516 15612
rect 13428 15488 13457 15534
rect 13503 15488 13516 15534
rect 13428 15448 13516 15488
rect 13588 15534 13676 15612
rect 13588 15488 13601 15534
rect 13647 15488 13676 15534
rect 13588 15448 13676 15488
rect 13876 15534 13964 15612
rect 13876 15488 13905 15534
rect 13951 15488 13964 15534
rect 13876 15448 13964 15488
rect 14036 15534 14124 15612
rect 14036 15488 14049 15534
rect 14095 15488 14124 15534
rect 14036 15448 14124 15488
rect 14324 15534 14412 15612
rect 14324 15488 14353 15534
rect 14399 15488 14412 15534
rect 14324 15448 14412 15488
rect 14484 15534 14572 15612
rect 14484 15488 14497 15534
rect 14543 15488 14572 15534
rect 14484 15448 14572 15488
rect 14772 15534 14860 15612
rect 14772 15488 14801 15534
rect 14847 15488 14860 15534
rect 14772 15448 14860 15488
rect 14932 15534 15020 15612
rect 14932 15488 14945 15534
rect 14991 15488 15020 15534
rect 14932 15448 15020 15488
rect 15220 15534 15308 15612
rect 15220 15488 15249 15534
rect 15295 15488 15308 15534
rect 15220 15448 15308 15488
rect 15380 15534 15468 15612
rect 15380 15488 15393 15534
rect 15439 15488 15468 15534
rect 15380 15448 15468 15488
rect 15668 15534 15756 15612
rect 15668 15488 15697 15534
rect 15743 15488 15756 15534
rect 15668 15448 15756 15488
rect 15828 15534 15916 15612
rect 15828 15488 15841 15534
rect 15887 15488 15916 15534
rect 15828 15448 15916 15488
rect 16116 15534 16204 15612
rect 16116 15488 16145 15534
rect 16191 15488 16204 15534
rect 16116 15448 16204 15488
rect 16276 15534 16364 15612
rect 16276 15488 16289 15534
rect 16335 15488 16364 15534
rect 16276 15448 16364 15488
rect 16564 15534 16652 15612
rect 16564 15488 16593 15534
rect 16639 15488 16652 15534
rect 16564 15448 16652 15488
rect 16724 15534 16812 15612
rect 16724 15488 16737 15534
rect 16783 15488 16812 15534
rect 16724 15448 16812 15488
rect 17012 15534 17100 15612
rect 17012 15488 17041 15534
rect 17087 15488 17100 15534
rect 17012 15448 17100 15488
rect 17508 15534 17596 15612
rect 17508 15488 17521 15534
rect 17567 15488 17596 15534
rect 17508 15448 17596 15488
rect 17796 15534 17884 15612
rect 17796 15488 17825 15534
rect 17871 15488 17884 15534
rect 17796 15448 17884 15488
rect 17956 15534 18044 15612
rect 17956 15488 17969 15534
rect 18015 15488 18044 15534
rect 17956 15448 18044 15488
rect 18244 15534 18332 15612
rect 18244 15488 18273 15534
rect 18319 15488 18332 15534
rect 18244 15448 18332 15488
rect 18404 15534 18492 15612
rect 18404 15488 18417 15534
rect 18463 15488 18492 15534
rect 18404 15448 18492 15488
rect 18692 15534 18780 15612
rect 18692 15488 18721 15534
rect 18767 15488 18780 15534
rect 18692 15448 18780 15488
rect 18852 15534 18940 15612
rect 18852 15488 18865 15534
rect 18911 15488 18940 15534
rect 18852 15448 18940 15488
rect 19140 15534 19228 15612
rect 19140 15488 19169 15534
rect 19215 15488 19228 15534
rect 19140 15448 19228 15488
rect 19300 15534 19388 15612
rect 19300 15488 19313 15534
rect 19359 15488 19388 15534
rect 19300 15448 19388 15488
rect 19588 15534 19676 15612
rect 19588 15488 19617 15534
rect 19663 15488 19676 15534
rect 19588 15448 19676 15488
rect 19748 15534 19836 15612
rect 19748 15488 19761 15534
rect 19807 15488 19836 15534
rect 19748 15448 19836 15488
rect 20036 15534 20124 15612
rect 20036 15488 20065 15534
rect 20111 15488 20124 15534
rect 20036 15448 20124 15488
rect 20196 15534 20284 15612
rect 20196 15488 20209 15534
rect 20255 15488 20284 15534
rect 20196 15448 20284 15488
rect 20484 15534 20572 15612
rect 20484 15488 20513 15534
rect 20559 15488 20572 15534
rect 20484 15448 20572 15488
rect 20644 15534 20732 15612
rect 20644 15488 20657 15534
rect 20703 15488 20732 15534
rect 20644 15448 20732 15488
rect 20932 15534 21020 15612
rect 20932 15488 20961 15534
rect 21007 15488 21020 15534
rect 20932 15448 21020 15488
rect 21092 15534 21180 15612
rect 21092 15488 21105 15534
rect 21151 15488 21180 15534
rect 21092 15448 21180 15488
rect 21380 15534 21468 15612
rect 21380 15488 21409 15534
rect 21455 15488 21468 15534
rect 21380 15448 21468 15488
rect 21540 15534 21628 15612
rect 21540 15488 21553 15534
rect 21599 15488 21628 15534
rect 21540 15448 21628 15488
rect 21828 15534 21916 15612
rect 21828 15488 21857 15534
rect 21903 15488 21916 15534
rect 21828 15448 21916 15488
rect 21988 15534 22076 15612
rect 21988 15488 22001 15534
rect 22047 15488 22076 15534
rect 21988 15448 22076 15488
rect 22276 15534 22364 15612
rect 22276 15488 22305 15534
rect 22351 15488 22364 15534
rect 22276 15448 22364 15488
rect 1604 14304 1692 14344
rect 1604 14258 1617 14304
rect 1663 14258 1692 14304
rect 1604 14180 1692 14258
rect 1892 14304 1980 14344
rect 1892 14258 1921 14304
rect 1967 14258 1980 14304
rect 1892 14180 1980 14258
rect 2052 14304 2140 14344
rect 2052 14258 2065 14304
rect 2111 14258 2140 14304
rect 2052 14180 2140 14258
rect 2340 14304 2428 14344
rect 2340 14258 2369 14304
rect 2415 14258 2428 14304
rect 2340 14180 2428 14258
rect 2500 14304 2588 14344
rect 2500 14258 2513 14304
rect 2559 14258 2588 14304
rect 2500 14180 2588 14258
rect 2788 14304 2876 14344
rect 2788 14258 2817 14304
rect 2863 14258 2876 14304
rect 2788 14180 2876 14258
rect 2948 14304 3036 14344
rect 2948 14258 2961 14304
rect 3007 14258 3036 14304
rect 2948 14180 3036 14258
rect 3236 14304 3324 14344
rect 3236 14258 3265 14304
rect 3311 14258 3324 14304
rect 3236 14180 3324 14258
rect 3396 14304 3484 14344
rect 3396 14258 3409 14304
rect 3455 14258 3484 14304
rect 3396 14180 3484 14258
rect 3684 14304 3772 14344
rect 3684 14258 3713 14304
rect 3759 14258 3772 14304
rect 3684 14180 3772 14258
rect 3844 14304 3932 14344
rect 3844 14258 3857 14304
rect 3903 14258 3932 14304
rect 3844 14180 3932 14258
rect 4132 14304 4220 14344
rect 4132 14258 4161 14304
rect 4207 14258 4220 14304
rect 4132 14180 4220 14258
rect 4292 14304 4380 14344
rect 4292 14258 4305 14304
rect 4351 14258 4380 14304
rect 4292 14180 4380 14258
rect 4580 14304 4668 14344
rect 4580 14258 4609 14304
rect 4655 14258 4668 14304
rect 4580 14180 4668 14258
rect 4740 14304 4828 14344
rect 4740 14258 4753 14304
rect 4799 14258 4828 14304
rect 4740 14180 4828 14258
rect 5028 14304 5116 14344
rect 5028 14258 5057 14304
rect 5103 14258 5116 14304
rect 5028 14180 5116 14258
rect 5524 14304 5612 14344
rect 5524 14258 5537 14304
rect 5583 14258 5612 14304
rect 5524 14180 5612 14258
rect 5812 14304 5900 14344
rect 5812 14258 5841 14304
rect 5887 14258 5900 14304
rect 5812 14180 5900 14258
rect 5972 14304 6060 14344
rect 5972 14258 5985 14304
rect 6031 14258 6060 14304
rect 5972 14180 6060 14258
rect 6260 14304 6348 14344
rect 6260 14258 6289 14304
rect 6335 14258 6348 14304
rect 6260 14180 6348 14258
rect 6420 14304 6508 14344
rect 6420 14258 6433 14304
rect 6479 14258 6508 14304
rect 6420 14180 6508 14258
rect 6708 14304 6796 14344
rect 6708 14258 6737 14304
rect 6783 14258 6796 14304
rect 6708 14180 6796 14258
rect 6868 14304 6956 14344
rect 6868 14258 6881 14304
rect 6927 14258 6956 14304
rect 6868 14180 6956 14258
rect 7156 14304 7244 14344
rect 7156 14258 7185 14304
rect 7231 14258 7244 14304
rect 7156 14180 7244 14258
rect 7316 14304 7404 14344
rect 7316 14258 7329 14304
rect 7375 14258 7404 14304
rect 7316 14180 7404 14258
rect 7604 14304 7692 14344
rect 7604 14258 7633 14304
rect 7679 14258 7692 14304
rect 7604 14180 7692 14258
rect 7764 14304 7852 14344
rect 7764 14258 7777 14304
rect 7823 14258 7852 14304
rect 7764 14180 7852 14258
rect 8052 14304 8140 14344
rect 8052 14258 8081 14304
rect 8127 14258 8140 14304
rect 8052 14180 8140 14258
rect 8212 14304 8300 14344
rect 8212 14258 8225 14304
rect 8271 14258 8300 14304
rect 8212 14180 8300 14258
rect 8500 14304 8588 14344
rect 8500 14258 8529 14304
rect 8575 14258 8588 14304
rect 8500 14180 8588 14258
rect 8660 14304 8748 14344
rect 8660 14258 8673 14304
rect 8719 14258 8748 14304
rect 8660 14180 8748 14258
rect 8948 14304 9036 14344
rect 8948 14258 8977 14304
rect 9023 14258 9036 14304
rect 8948 14180 9036 14258
rect 9108 14304 9196 14344
rect 9108 14258 9121 14304
rect 9167 14258 9196 14304
rect 9108 14180 9196 14258
rect 9396 14304 9484 14344
rect 9396 14258 9425 14304
rect 9471 14258 9484 14304
rect 9396 14180 9484 14258
rect 9556 14304 9644 14344
rect 9556 14258 9569 14304
rect 9615 14258 9644 14304
rect 9556 14180 9644 14258
rect 9844 14304 9932 14344
rect 9844 14258 9873 14304
rect 9919 14258 9932 14304
rect 9844 14180 9932 14258
rect 10004 14304 10092 14344
rect 10004 14258 10017 14304
rect 10063 14258 10092 14304
rect 10004 14180 10092 14258
rect 10292 14304 10380 14344
rect 10292 14258 10321 14304
rect 10367 14258 10380 14304
rect 10292 14180 10380 14258
rect 10452 14304 10540 14344
rect 10452 14258 10465 14304
rect 10511 14258 10540 14304
rect 10452 14180 10540 14258
rect 10740 14304 10828 14344
rect 10740 14258 10769 14304
rect 10815 14258 10828 14304
rect 10740 14180 10828 14258
rect 10900 14304 10988 14344
rect 10900 14258 10913 14304
rect 10959 14258 10988 14304
rect 10900 14180 10988 14258
rect 11188 14304 11276 14344
rect 11188 14258 11217 14304
rect 11263 14258 11276 14304
rect 11188 14180 11276 14258
rect 11348 14304 11436 14344
rect 11348 14258 11361 14304
rect 11407 14258 11436 14304
rect 11348 14180 11436 14258
rect 11636 14304 11724 14344
rect 11636 14258 11665 14304
rect 11711 14258 11724 14304
rect 11636 14180 11724 14258
rect 11796 14304 11884 14344
rect 11796 14258 11809 14304
rect 11855 14258 11884 14304
rect 11796 14180 11884 14258
rect 12084 14304 12172 14344
rect 12084 14258 12113 14304
rect 12159 14258 12172 14304
rect 12084 14180 12172 14258
rect 12244 14304 12332 14344
rect 12244 14258 12257 14304
rect 12303 14258 12332 14304
rect 12244 14180 12332 14258
rect 12532 14304 12620 14344
rect 12532 14258 12561 14304
rect 12607 14258 12620 14304
rect 12532 14180 12620 14258
rect 12692 14304 12780 14344
rect 12692 14258 12705 14304
rect 12751 14258 12780 14304
rect 12692 14180 12780 14258
rect 12980 14304 13068 14344
rect 12980 14258 13009 14304
rect 13055 14258 13068 14304
rect 12980 14180 13068 14258
rect 13476 14304 13564 14344
rect 13476 14258 13489 14304
rect 13535 14258 13564 14304
rect 13476 14180 13564 14258
rect 13764 14304 13852 14344
rect 13764 14258 13793 14304
rect 13839 14258 13852 14304
rect 13764 14180 13852 14258
rect 13924 14304 14012 14344
rect 13924 14258 13937 14304
rect 13983 14258 14012 14304
rect 13924 14180 14012 14258
rect 14212 14304 14300 14344
rect 14212 14258 14241 14304
rect 14287 14258 14300 14304
rect 14212 14180 14300 14258
rect 14372 14304 14460 14344
rect 14372 14258 14385 14304
rect 14431 14258 14460 14304
rect 14372 14180 14460 14258
rect 14660 14304 14748 14344
rect 14660 14258 14689 14304
rect 14735 14258 14748 14304
rect 14660 14180 14748 14258
rect 14820 14304 14908 14344
rect 14820 14258 14833 14304
rect 14879 14258 14908 14304
rect 14820 14180 14908 14258
rect 15108 14304 15196 14344
rect 15108 14258 15137 14304
rect 15183 14258 15196 14304
rect 15108 14180 15196 14258
rect 15268 14304 15356 14344
rect 15268 14258 15281 14304
rect 15327 14258 15356 14304
rect 15268 14180 15356 14258
rect 15556 14304 15644 14344
rect 15556 14258 15585 14304
rect 15631 14258 15644 14304
rect 15556 14180 15644 14258
rect 15716 14304 15804 14344
rect 15716 14258 15729 14304
rect 15775 14258 15804 14304
rect 15716 14180 15804 14258
rect 16004 14304 16092 14344
rect 16004 14258 16033 14304
rect 16079 14258 16092 14304
rect 16004 14180 16092 14258
rect 16164 14304 16252 14344
rect 16164 14258 16177 14304
rect 16223 14258 16252 14304
rect 16164 14180 16252 14258
rect 16452 14304 16540 14344
rect 16452 14258 16481 14304
rect 16527 14258 16540 14304
rect 16452 14180 16540 14258
rect 16804 14304 16892 14344
rect 16804 14258 16817 14304
rect 16863 14258 16892 14304
rect 16804 14180 16892 14258
rect 17012 14304 17100 14344
rect 17012 14258 17041 14304
rect 17087 14258 17100 14304
rect 17012 14180 17100 14258
rect 17476 14304 17564 14344
rect 17476 14258 17489 14304
rect 17535 14258 17564 14304
rect 17476 14180 17564 14258
rect 17684 14304 17772 14344
rect 17684 14258 17713 14304
rect 17759 14258 17772 14304
rect 17684 14180 17772 14258
rect 17844 14304 17932 14344
rect 17844 14258 17857 14304
rect 17903 14258 17932 14304
rect 17844 14180 17932 14258
rect 18132 14304 18220 14344
rect 18132 14258 18161 14304
rect 18207 14258 18220 14304
rect 18132 14180 18220 14258
rect 18292 14304 18380 14344
rect 18292 14258 18305 14304
rect 18351 14258 18380 14304
rect 18292 14180 18380 14258
rect 18580 14304 18668 14344
rect 18580 14258 18609 14304
rect 18655 14258 18668 14304
rect 18580 14180 18668 14258
rect 18740 14304 18828 14344
rect 18740 14258 18753 14304
rect 18799 14258 18828 14304
rect 18740 14180 18828 14258
rect 19028 14304 19116 14344
rect 19028 14258 19057 14304
rect 19103 14258 19116 14304
rect 19028 14180 19116 14258
rect 19188 14304 19276 14344
rect 19188 14258 19201 14304
rect 19247 14258 19276 14304
rect 19188 14180 19276 14258
rect 19476 14304 19564 14344
rect 19476 14258 19505 14304
rect 19551 14258 19564 14304
rect 19476 14180 19564 14258
rect 19636 14304 19724 14344
rect 19636 14258 19649 14304
rect 19695 14258 19724 14304
rect 19636 14180 19724 14258
rect 19924 14304 20012 14344
rect 19924 14258 19953 14304
rect 19999 14258 20012 14304
rect 19924 14180 20012 14258
rect 20084 14304 20172 14344
rect 20084 14258 20097 14304
rect 20143 14258 20172 14304
rect 20084 14180 20172 14258
rect 20372 14304 20460 14344
rect 20372 14258 20401 14304
rect 20447 14258 20460 14304
rect 20372 14180 20460 14258
rect 20532 14304 20620 14344
rect 20532 14258 20545 14304
rect 20591 14258 20620 14304
rect 20532 14180 20620 14258
rect 20820 14304 20908 14344
rect 20820 14258 20849 14304
rect 20895 14258 20908 14304
rect 20820 14180 20908 14258
rect 21428 14304 21516 14344
rect 21428 14258 21441 14304
rect 21487 14258 21516 14304
rect 21428 14180 21516 14258
rect 21716 14304 21804 14344
rect 21716 14258 21745 14304
rect 21791 14258 21804 14304
rect 21716 14180 21804 14258
rect 21876 14304 21964 14344
rect 21876 14258 21889 14304
rect 21935 14258 21964 14304
rect 21876 14180 21964 14258
rect 22164 14304 22252 14344
rect 22164 14258 22193 14304
rect 22239 14258 22252 14304
rect 22164 14180 22252 14258
rect 1604 13966 1692 14044
rect 1604 13920 1617 13966
rect 1663 13920 1692 13966
rect 1604 13880 1692 13920
rect 1892 13966 1980 14044
rect 1892 13920 1921 13966
rect 1967 13920 1980 13966
rect 1892 13880 1980 13920
rect 2052 13966 2140 14044
rect 2052 13920 2065 13966
rect 2111 13920 2140 13966
rect 2052 13880 2140 13920
rect 2340 13966 2428 14044
rect 2340 13920 2369 13966
rect 2415 13920 2428 13966
rect 2340 13880 2428 13920
rect 2500 13966 2588 14044
rect 2500 13920 2513 13966
rect 2559 13920 2588 13966
rect 2500 13880 2588 13920
rect 2788 13966 2876 14044
rect 2788 13920 2817 13966
rect 2863 13920 2876 13966
rect 2788 13880 2876 13920
rect 2948 13966 3036 14044
rect 2948 13920 2961 13966
rect 3007 13920 3036 13966
rect 2948 13880 3036 13920
rect 3236 13966 3324 14044
rect 3236 13920 3265 13966
rect 3311 13920 3324 13966
rect 3236 13880 3324 13920
rect 3396 13966 3484 14044
rect 3396 13920 3409 13966
rect 3455 13920 3484 13966
rect 3396 13880 3484 13920
rect 3684 13966 3772 14044
rect 3684 13920 3713 13966
rect 3759 13920 3772 13966
rect 3684 13880 3772 13920
rect 3844 13966 3932 14044
rect 3844 13920 3857 13966
rect 3903 13920 3932 13966
rect 3844 13880 3932 13920
rect 4132 13966 4220 14044
rect 4132 13920 4161 13966
rect 4207 13920 4220 13966
rect 4132 13880 4220 13920
rect 4292 13966 4380 14044
rect 4292 13920 4305 13966
rect 4351 13920 4380 13966
rect 4292 13880 4380 13920
rect 4580 13966 4668 14044
rect 4580 13920 4609 13966
rect 4655 13920 4668 13966
rect 4580 13880 4668 13920
rect 4740 13966 4828 14044
rect 4740 13920 4753 13966
rect 4799 13920 4828 13966
rect 4740 13880 4828 13920
rect 5028 13966 5116 14044
rect 5028 13920 5057 13966
rect 5103 13920 5116 13966
rect 5028 13880 5116 13920
rect 5188 13966 5276 14044
rect 5188 13920 5201 13966
rect 5247 13920 5276 13966
rect 5188 13880 5276 13920
rect 5476 13966 5564 14044
rect 5476 13920 5505 13966
rect 5551 13920 5564 13966
rect 5476 13880 5564 13920
rect 5636 13966 5724 14044
rect 5636 13920 5649 13966
rect 5695 13920 5724 13966
rect 5636 13880 5724 13920
rect 5924 13966 6012 14044
rect 5924 13920 5953 13966
rect 5999 13920 6012 13966
rect 5924 13880 6012 13920
rect 6084 13966 6172 14044
rect 6084 13920 6097 13966
rect 6143 13920 6172 13966
rect 6084 13880 6172 13920
rect 6372 13966 6460 14044
rect 6372 13920 6401 13966
rect 6447 13920 6460 13966
rect 6372 13880 6460 13920
rect 6532 13966 6620 14044
rect 6532 13920 6545 13966
rect 6591 13920 6620 13966
rect 6532 13880 6620 13920
rect 6820 13966 6908 14044
rect 6820 13920 6849 13966
rect 6895 13920 6908 13966
rect 6820 13880 6908 13920
rect 6980 13966 7068 14044
rect 6980 13920 6993 13966
rect 7039 13920 7068 13966
rect 6980 13880 7068 13920
rect 7268 13966 7356 14044
rect 7268 13920 7297 13966
rect 7343 13920 7356 13966
rect 7268 13880 7356 13920
rect 7428 13966 7516 14044
rect 7428 13920 7441 13966
rect 7487 13920 7516 13966
rect 7428 13880 7516 13920
rect 7716 13966 7804 14044
rect 7716 13920 7745 13966
rect 7791 13920 7804 13966
rect 7716 13880 7804 13920
rect 7876 13966 7964 14044
rect 7876 13920 7889 13966
rect 7935 13920 7964 13966
rect 7876 13880 7964 13920
rect 8164 13966 8252 14044
rect 8164 13920 8193 13966
rect 8239 13920 8252 13966
rect 8164 13880 8252 13920
rect 8324 13966 8412 14044
rect 8324 13920 8337 13966
rect 8383 13920 8412 13966
rect 8324 13880 8412 13920
rect 8612 13966 8700 14044
rect 8612 13920 8641 13966
rect 8687 13920 8700 13966
rect 8612 13880 8700 13920
rect 8772 13966 8860 14044
rect 8772 13920 8785 13966
rect 8831 13920 8860 13966
rect 8772 13880 8860 13920
rect 9060 13966 9148 14044
rect 9060 13920 9089 13966
rect 9135 13920 9148 13966
rect 9060 13880 9148 13920
rect 9556 13966 9644 14044
rect 9556 13920 9569 13966
rect 9615 13920 9644 13966
rect 9556 13880 9644 13920
rect 9844 13966 9932 14044
rect 9844 13920 9873 13966
rect 9919 13920 9932 13966
rect 9844 13880 9932 13920
rect 10004 13966 10092 14044
rect 10004 13920 10017 13966
rect 10063 13920 10092 13966
rect 10004 13880 10092 13920
rect 10292 13966 10380 14044
rect 10292 13920 10321 13966
rect 10367 13920 10380 13966
rect 10292 13880 10380 13920
rect 10452 13966 10540 14044
rect 10452 13920 10465 13966
rect 10511 13920 10540 13966
rect 10452 13880 10540 13920
rect 10740 13966 10828 14044
rect 10740 13920 10769 13966
rect 10815 13920 10828 13966
rect 10740 13880 10828 13920
rect 10900 13966 10988 14044
rect 10900 13920 10913 13966
rect 10959 13920 10988 13966
rect 10900 13880 10988 13920
rect 11188 13966 11276 14044
rect 11188 13920 11217 13966
rect 11263 13920 11276 13966
rect 11188 13880 11276 13920
rect 11348 13966 11436 14044
rect 11348 13920 11361 13966
rect 11407 13920 11436 13966
rect 11348 13880 11436 13920
rect 11636 13966 11724 14044
rect 11636 13920 11665 13966
rect 11711 13920 11724 13966
rect 11636 13880 11724 13920
rect 11796 13966 11884 14044
rect 11796 13920 11809 13966
rect 11855 13920 11884 13966
rect 11796 13880 11884 13920
rect 12084 13966 12172 14044
rect 12084 13920 12113 13966
rect 12159 13920 12172 13966
rect 12084 13880 12172 13920
rect 12244 13966 12332 14044
rect 12244 13920 12257 13966
rect 12303 13920 12332 13966
rect 12244 13880 12332 13920
rect 12532 13966 12620 14044
rect 12532 13920 12561 13966
rect 12607 13920 12620 13966
rect 12532 13880 12620 13920
rect 12692 13966 12780 14044
rect 12692 13920 12705 13966
rect 12751 13920 12780 13966
rect 12692 13880 12780 13920
rect 12980 13966 13068 14044
rect 12980 13920 13009 13966
rect 13055 13920 13068 13966
rect 12980 13880 13068 13920
rect 13140 13966 13228 14044
rect 13140 13920 13153 13966
rect 13199 13920 13228 13966
rect 13140 13880 13228 13920
rect 13428 13966 13516 14044
rect 13428 13920 13457 13966
rect 13503 13920 13516 13966
rect 13428 13880 13516 13920
rect 13588 13966 13676 14044
rect 13588 13920 13601 13966
rect 13647 13920 13676 13966
rect 13588 13880 13676 13920
rect 13876 13966 13964 14044
rect 13876 13920 13905 13966
rect 13951 13920 13964 13966
rect 13876 13880 13964 13920
rect 14036 13966 14124 14044
rect 14036 13920 14049 13966
rect 14095 13920 14124 13966
rect 14036 13880 14124 13920
rect 14324 13966 14412 14044
rect 14324 13920 14353 13966
rect 14399 13920 14412 13966
rect 14324 13880 14412 13920
rect 14484 13966 14572 14044
rect 14484 13920 14497 13966
rect 14543 13920 14572 13966
rect 14484 13880 14572 13920
rect 14772 13966 14860 14044
rect 14772 13920 14801 13966
rect 14847 13920 14860 13966
rect 14772 13880 14860 13920
rect 14932 13966 15020 14044
rect 14932 13920 14945 13966
rect 14991 13920 15020 13966
rect 14932 13880 15020 13920
rect 15220 13966 15308 14044
rect 15220 13920 15249 13966
rect 15295 13920 15308 13966
rect 15220 13880 15308 13920
rect 15380 13966 15468 14044
rect 15380 13920 15393 13966
rect 15439 13920 15468 13966
rect 15380 13880 15468 13920
rect 15668 13966 15756 14044
rect 15668 13920 15697 13966
rect 15743 13920 15756 13966
rect 15668 13880 15756 13920
rect 16052 13966 16140 14044
rect 16052 13920 16065 13966
rect 16111 13920 16140 13966
rect 16052 13880 16140 13920
rect 16260 13966 16348 14044
rect 16260 13920 16289 13966
rect 16335 13920 16348 13966
rect 16260 13880 16348 13920
rect 16724 13966 16812 14044
rect 16724 13920 16737 13966
rect 16783 13920 16812 13966
rect 16724 13880 16812 13920
rect 16932 13966 17020 14044
rect 16932 13920 16961 13966
rect 17007 13920 17020 13966
rect 16932 13880 17020 13920
rect 17620 13966 17708 14044
rect 17620 13920 17633 13966
rect 17679 13920 17708 13966
rect 17620 13880 17708 13920
rect 17828 13966 17916 14044
rect 17828 13920 17857 13966
rect 17903 13920 17916 13966
rect 17828 13880 17916 13920
rect 18292 13966 18380 14044
rect 18292 13920 18305 13966
rect 18351 13920 18380 13966
rect 18292 13880 18380 13920
rect 18500 13966 18588 14044
rect 18500 13920 18529 13966
rect 18575 13920 18588 13966
rect 18500 13880 18588 13920
rect 18740 13966 18828 14044
rect 18740 13920 18753 13966
rect 18799 13920 18828 13966
rect 18740 13880 18828 13920
rect 19028 13966 19116 14044
rect 19028 13920 19057 13966
rect 19103 13920 19116 13966
rect 19028 13880 19116 13920
rect 19188 13966 19276 14044
rect 19188 13920 19201 13966
rect 19247 13920 19276 13966
rect 19188 13880 19276 13920
rect 19476 13966 19564 14044
rect 19476 13920 19505 13966
rect 19551 13920 19564 13966
rect 19476 13880 19564 13920
rect 19636 13966 19724 14044
rect 19636 13920 19649 13966
rect 19695 13920 19724 13966
rect 19636 13880 19724 13920
rect 19924 13966 20012 14044
rect 19924 13920 19953 13966
rect 19999 13920 20012 13966
rect 19924 13880 20012 13920
rect 20084 13966 20172 14044
rect 20084 13920 20097 13966
rect 20143 13920 20172 13966
rect 20084 13880 20172 13920
rect 20372 13966 20460 14044
rect 20372 13920 20401 13966
rect 20447 13920 20460 13966
rect 20372 13880 20460 13920
rect 20532 13966 20620 14044
rect 20532 13920 20545 13966
rect 20591 13920 20620 13966
rect 20532 13880 20620 13920
rect 20820 13966 20908 14044
rect 20820 13920 20849 13966
rect 20895 13920 20908 13966
rect 20820 13880 20908 13920
rect 20980 13966 21068 14044
rect 20980 13920 20993 13966
rect 21039 13920 21068 13966
rect 20980 13880 21068 13920
rect 21268 13966 21356 14044
rect 21268 13920 21297 13966
rect 21343 13920 21356 13966
rect 21268 13880 21356 13920
rect 21428 13966 21516 14044
rect 21428 13920 21441 13966
rect 21487 13920 21516 13966
rect 21428 13880 21516 13920
rect 21716 13966 21804 14044
rect 21716 13920 21745 13966
rect 21791 13920 21804 13966
rect 21716 13880 21804 13920
rect 21876 13966 21964 14044
rect 21876 13920 21889 13966
rect 21935 13920 21964 13966
rect 21876 13880 21964 13920
rect 22164 13966 22252 14044
rect 22164 13920 22193 13966
rect 22239 13920 22252 13966
rect 22164 13880 22252 13920
rect 1604 12736 1692 12776
rect 1604 12690 1617 12736
rect 1663 12690 1692 12736
rect 1604 12612 1692 12690
rect 1892 12736 1980 12776
rect 1892 12690 1921 12736
rect 1967 12690 1980 12736
rect 1892 12612 1980 12690
rect 2052 12736 2140 12776
rect 2052 12690 2065 12736
rect 2111 12690 2140 12736
rect 2052 12612 2140 12690
rect 2340 12736 2428 12776
rect 2340 12690 2369 12736
rect 2415 12690 2428 12736
rect 2340 12612 2428 12690
rect 2500 12736 2588 12776
rect 2500 12690 2513 12736
rect 2559 12690 2588 12736
rect 2500 12612 2588 12690
rect 2788 12736 2876 12776
rect 2788 12690 2817 12736
rect 2863 12690 2876 12736
rect 2788 12612 2876 12690
rect 2948 12736 3036 12776
rect 2948 12690 2961 12736
rect 3007 12690 3036 12736
rect 2948 12612 3036 12690
rect 3236 12736 3324 12776
rect 3236 12690 3265 12736
rect 3311 12690 3324 12736
rect 3236 12612 3324 12690
rect 3396 12736 3484 12776
rect 3396 12690 3409 12736
rect 3455 12690 3484 12736
rect 3396 12612 3484 12690
rect 3684 12736 3772 12776
rect 3684 12690 3713 12736
rect 3759 12690 3772 12736
rect 3684 12612 3772 12690
rect 3844 12736 3932 12776
rect 3844 12690 3857 12736
rect 3903 12690 3932 12736
rect 3844 12612 3932 12690
rect 4132 12736 4220 12776
rect 4132 12690 4161 12736
rect 4207 12690 4220 12736
rect 4132 12612 4220 12690
rect 4292 12736 4380 12776
rect 4292 12690 4305 12736
rect 4351 12690 4380 12736
rect 4292 12612 4380 12690
rect 4580 12736 4668 12776
rect 4580 12690 4609 12736
rect 4655 12690 4668 12736
rect 4580 12612 4668 12690
rect 4740 12736 4828 12776
rect 4740 12690 4753 12736
rect 4799 12690 4828 12736
rect 4740 12612 4828 12690
rect 5028 12736 5116 12776
rect 5028 12690 5057 12736
rect 5103 12690 5116 12736
rect 5028 12612 5116 12690
rect 5524 12736 5612 12776
rect 5524 12690 5537 12736
rect 5583 12690 5612 12736
rect 5524 12612 5612 12690
rect 5812 12736 5900 12776
rect 5812 12690 5841 12736
rect 5887 12690 5900 12736
rect 5812 12612 5900 12690
rect 5972 12736 6060 12776
rect 5972 12690 5985 12736
rect 6031 12690 6060 12736
rect 5972 12612 6060 12690
rect 6260 12736 6348 12776
rect 6260 12690 6289 12736
rect 6335 12690 6348 12736
rect 6260 12612 6348 12690
rect 6420 12736 6508 12776
rect 6420 12690 6433 12736
rect 6479 12690 6508 12736
rect 6420 12612 6508 12690
rect 6708 12736 6796 12776
rect 6708 12690 6737 12736
rect 6783 12690 6796 12736
rect 6708 12612 6796 12690
rect 6868 12736 6956 12776
rect 6868 12690 6881 12736
rect 6927 12690 6956 12736
rect 6868 12612 6956 12690
rect 7156 12736 7244 12776
rect 7156 12690 7185 12736
rect 7231 12690 7244 12736
rect 7156 12612 7244 12690
rect 7316 12736 7404 12776
rect 7316 12690 7329 12736
rect 7375 12690 7404 12736
rect 7316 12612 7404 12690
rect 7604 12736 7692 12776
rect 7604 12690 7633 12736
rect 7679 12690 7692 12736
rect 7604 12612 7692 12690
rect 7764 12736 7852 12776
rect 7764 12690 7777 12736
rect 7823 12690 7852 12736
rect 7764 12612 7852 12690
rect 8052 12736 8140 12776
rect 8052 12690 8081 12736
rect 8127 12690 8140 12736
rect 8052 12612 8140 12690
rect 8212 12736 8300 12776
rect 8212 12690 8225 12736
rect 8271 12690 8300 12736
rect 8212 12612 8300 12690
rect 8500 12736 8588 12776
rect 8500 12690 8529 12736
rect 8575 12690 8588 12736
rect 8500 12612 8588 12690
rect 8660 12736 8748 12776
rect 8660 12690 8673 12736
rect 8719 12690 8748 12736
rect 8660 12612 8748 12690
rect 8948 12736 9036 12776
rect 8948 12690 8977 12736
rect 9023 12690 9036 12736
rect 8948 12612 9036 12690
rect 9108 12736 9196 12776
rect 9108 12690 9121 12736
rect 9167 12690 9196 12736
rect 9108 12612 9196 12690
rect 9396 12736 9484 12776
rect 9396 12690 9425 12736
rect 9471 12690 9484 12736
rect 9396 12612 9484 12690
rect 9556 12736 9644 12776
rect 9556 12690 9569 12736
rect 9615 12690 9644 12736
rect 9556 12612 9644 12690
rect 9844 12736 9932 12776
rect 9844 12690 9873 12736
rect 9919 12690 9932 12736
rect 9844 12612 9932 12690
rect 10004 12736 10092 12776
rect 10004 12690 10017 12736
rect 10063 12690 10092 12736
rect 10004 12612 10092 12690
rect 10292 12736 10380 12776
rect 10292 12690 10321 12736
rect 10367 12690 10380 12736
rect 10292 12612 10380 12690
rect 10452 12736 10540 12776
rect 10452 12690 10465 12736
rect 10511 12690 10540 12736
rect 10452 12612 10540 12690
rect 10740 12736 10828 12776
rect 10740 12690 10769 12736
rect 10815 12690 10828 12736
rect 10740 12612 10828 12690
rect 10900 12736 10988 12776
rect 10900 12690 10913 12736
rect 10959 12690 10988 12736
rect 10900 12612 10988 12690
rect 11188 12736 11276 12776
rect 11188 12690 11217 12736
rect 11263 12690 11276 12736
rect 11188 12612 11276 12690
rect 11348 12736 11436 12776
rect 11348 12690 11361 12736
rect 11407 12690 11436 12736
rect 11348 12612 11436 12690
rect 11636 12736 11724 12776
rect 11636 12690 11665 12736
rect 11711 12690 11724 12736
rect 11636 12612 11724 12690
rect 11796 12736 11884 12776
rect 11796 12690 11809 12736
rect 11855 12690 11884 12736
rect 11796 12612 11884 12690
rect 12084 12736 12172 12776
rect 12084 12690 12113 12736
rect 12159 12690 12172 12736
rect 12084 12612 12172 12690
rect 12244 12736 12332 12776
rect 12244 12690 12257 12736
rect 12303 12690 12332 12736
rect 12244 12612 12332 12690
rect 12532 12736 12620 12776
rect 12532 12690 12561 12736
rect 12607 12690 12620 12736
rect 12532 12612 12620 12690
rect 12692 12736 12780 12776
rect 12692 12690 12705 12736
rect 12751 12690 12780 12736
rect 12692 12612 12780 12690
rect 12980 12736 13068 12776
rect 12980 12690 13009 12736
rect 13055 12690 13068 12736
rect 12980 12612 13068 12690
rect 13476 12736 13564 12776
rect 13476 12690 13489 12736
rect 13535 12690 13564 12736
rect 13476 12612 13564 12690
rect 13764 12736 13852 12776
rect 13764 12690 13793 12736
rect 13839 12690 13852 12736
rect 13764 12612 13852 12690
rect 13924 12736 14012 12776
rect 13924 12690 13937 12736
rect 13983 12690 14012 12736
rect 13924 12612 14012 12690
rect 14212 12736 14300 12776
rect 14212 12690 14241 12736
rect 14287 12690 14300 12736
rect 14212 12612 14300 12690
rect 14708 12736 14796 12776
rect 14708 12690 14721 12736
rect 14767 12690 14796 12736
rect 14708 12612 14796 12690
rect 14916 12736 15004 12776
rect 14916 12690 14945 12736
rect 14991 12690 15004 12736
rect 14916 12612 15004 12690
rect 15380 12736 15468 12776
rect 15380 12690 15393 12736
rect 15439 12690 15468 12736
rect 15380 12612 15468 12690
rect 15588 12736 15676 12776
rect 15588 12690 15617 12736
rect 15663 12690 15676 12736
rect 15588 12612 15676 12690
rect 16052 12736 16140 12776
rect 16052 12690 16065 12736
rect 16111 12690 16140 12736
rect 16052 12612 16140 12690
rect 16260 12736 16348 12776
rect 16260 12690 16289 12736
rect 16335 12690 16348 12736
rect 16260 12612 16348 12690
rect 16724 12736 16812 12776
rect 16724 12690 16737 12736
rect 16783 12690 16812 12736
rect 16724 12612 16812 12690
rect 16932 12736 17020 12776
rect 16932 12690 16961 12736
rect 17007 12690 17020 12736
rect 16932 12612 17020 12690
rect 17396 12736 17484 12776
rect 17396 12690 17409 12736
rect 17455 12690 17484 12736
rect 17396 12612 17484 12690
rect 17604 12736 17692 12776
rect 17604 12690 17633 12736
rect 17679 12690 17692 12736
rect 17604 12612 17692 12690
rect 18068 12736 18156 12776
rect 18068 12690 18081 12736
rect 18127 12690 18156 12736
rect 18068 12612 18156 12690
rect 18276 12736 18364 12776
rect 18276 12690 18305 12736
rect 18351 12690 18364 12736
rect 18276 12612 18364 12690
rect 18740 12736 18828 12776
rect 18740 12690 18753 12736
rect 18799 12690 18828 12736
rect 18740 12612 18828 12690
rect 18948 12736 19036 12776
rect 18948 12690 18977 12736
rect 19023 12690 19036 12736
rect 18948 12612 19036 12690
rect 19412 12736 19500 12776
rect 19412 12690 19425 12736
rect 19471 12690 19500 12736
rect 19412 12612 19500 12690
rect 19620 12736 19708 12776
rect 19620 12690 19649 12736
rect 19695 12690 19708 12736
rect 19620 12612 19708 12690
rect 19860 12736 19948 12776
rect 19860 12690 19873 12736
rect 19919 12690 19948 12736
rect 19860 12612 19948 12690
rect 20148 12736 20236 12776
rect 20148 12690 20177 12736
rect 20223 12690 20236 12736
rect 20148 12612 20236 12690
rect 20308 12736 20396 12776
rect 20308 12690 20321 12736
rect 20367 12690 20396 12736
rect 20308 12612 20396 12690
rect 20596 12736 20684 12776
rect 20596 12690 20625 12736
rect 20671 12690 20684 12736
rect 20596 12612 20684 12690
rect 20756 12736 20844 12776
rect 20756 12690 20769 12736
rect 20815 12690 20844 12736
rect 20756 12612 20844 12690
rect 21044 12736 21132 12776
rect 21044 12690 21073 12736
rect 21119 12690 21132 12736
rect 21044 12612 21132 12690
rect 21428 12736 21516 12776
rect 21428 12690 21441 12736
rect 21487 12690 21516 12736
rect 21428 12612 21516 12690
rect 21716 12736 21804 12776
rect 21716 12690 21745 12736
rect 21791 12690 21804 12736
rect 21716 12612 21804 12690
rect 21876 12736 21964 12776
rect 21876 12690 21889 12736
rect 21935 12690 21964 12736
rect 21876 12612 21964 12690
rect 22164 12736 22252 12776
rect 22164 12690 22193 12736
rect 22239 12690 22252 12736
rect 22164 12612 22252 12690
rect 1604 12398 1692 12476
rect 1604 12352 1617 12398
rect 1663 12352 1692 12398
rect 1604 12312 1692 12352
rect 1892 12398 1980 12476
rect 1892 12352 1921 12398
rect 1967 12352 1980 12398
rect 1892 12312 1980 12352
rect 2052 12398 2140 12476
rect 2052 12352 2065 12398
rect 2111 12352 2140 12398
rect 2052 12312 2140 12352
rect 2340 12398 2428 12476
rect 2340 12352 2369 12398
rect 2415 12352 2428 12398
rect 2340 12312 2428 12352
rect 2500 12398 2588 12476
rect 2500 12352 2513 12398
rect 2559 12352 2588 12398
rect 2500 12312 2588 12352
rect 2788 12398 2876 12476
rect 2788 12352 2817 12398
rect 2863 12352 2876 12398
rect 2788 12312 2876 12352
rect 2948 12398 3036 12476
rect 2948 12352 2961 12398
rect 3007 12352 3036 12398
rect 2948 12312 3036 12352
rect 3236 12398 3324 12476
rect 3236 12352 3265 12398
rect 3311 12352 3324 12398
rect 3236 12312 3324 12352
rect 3396 12398 3484 12476
rect 3396 12352 3409 12398
rect 3455 12352 3484 12398
rect 3396 12312 3484 12352
rect 3684 12398 3772 12476
rect 3684 12352 3713 12398
rect 3759 12352 3772 12398
rect 3684 12312 3772 12352
rect 3844 12398 3932 12476
rect 3844 12352 3857 12398
rect 3903 12352 3932 12398
rect 3844 12312 3932 12352
rect 4132 12398 4220 12476
rect 4132 12352 4161 12398
rect 4207 12352 4220 12398
rect 4132 12312 4220 12352
rect 4292 12398 4380 12476
rect 4292 12352 4305 12398
rect 4351 12352 4380 12398
rect 4292 12312 4380 12352
rect 4580 12398 4668 12476
rect 4580 12352 4609 12398
rect 4655 12352 4668 12398
rect 4580 12312 4668 12352
rect 4740 12398 4828 12476
rect 4740 12352 4753 12398
rect 4799 12352 4828 12398
rect 4740 12312 4828 12352
rect 5028 12398 5116 12476
rect 5028 12352 5057 12398
rect 5103 12352 5116 12398
rect 5028 12312 5116 12352
rect 5188 12398 5276 12476
rect 5188 12352 5201 12398
rect 5247 12352 5276 12398
rect 5188 12312 5276 12352
rect 5476 12398 5564 12476
rect 5476 12352 5505 12398
rect 5551 12352 5564 12398
rect 5476 12312 5564 12352
rect 5636 12398 5724 12476
rect 5636 12352 5649 12398
rect 5695 12352 5724 12398
rect 5636 12312 5724 12352
rect 5924 12398 6012 12476
rect 5924 12352 5953 12398
rect 5999 12352 6012 12398
rect 5924 12312 6012 12352
rect 6084 12398 6172 12476
rect 6084 12352 6097 12398
rect 6143 12352 6172 12398
rect 6084 12312 6172 12352
rect 6372 12398 6460 12476
rect 6372 12352 6401 12398
rect 6447 12352 6460 12398
rect 6372 12312 6460 12352
rect 6532 12398 6620 12476
rect 6532 12352 6545 12398
rect 6591 12352 6620 12398
rect 6532 12312 6620 12352
rect 6820 12398 6908 12476
rect 6820 12352 6849 12398
rect 6895 12352 6908 12398
rect 6820 12312 6908 12352
rect 6980 12398 7068 12476
rect 6980 12352 6993 12398
rect 7039 12352 7068 12398
rect 6980 12312 7068 12352
rect 7268 12398 7356 12476
rect 7268 12352 7297 12398
rect 7343 12352 7356 12398
rect 7268 12312 7356 12352
rect 7428 12398 7516 12476
rect 7428 12352 7441 12398
rect 7487 12352 7516 12398
rect 7428 12312 7516 12352
rect 7716 12398 7804 12476
rect 7716 12352 7745 12398
rect 7791 12352 7804 12398
rect 7716 12312 7804 12352
rect 7876 12398 7964 12476
rect 7876 12352 7889 12398
rect 7935 12352 7964 12398
rect 7876 12312 7964 12352
rect 8164 12398 8252 12476
rect 8164 12352 8193 12398
rect 8239 12352 8252 12398
rect 8164 12312 8252 12352
rect 8324 12398 8412 12476
rect 8324 12352 8337 12398
rect 8383 12352 8412 12398
rect 8324 12312 8412 12352
rect 8612 12398 8700 12476
rect 8612 12352 8641 12398
rect 8687 12352 8700 12398
rect 8612 12312 8700 12352
rect 8772 12398 8860 12476
rect 8772 12352 8785 12398
rect 8831 12352 8860 12398
rect 8772 12312 8860 12352
rect 9060 12398 9148 12476
rect 9060 12352 9089 12398
rect 9135 12352 9148 12398
rect 9060 12312 9148 12352
rect 9556 12398 9644 12476
rect 9556 12352 9569 12398
rect 9615 12352 9644 12398
rect 9556 12312 9644 12352
rect 9844 12398 9932 12476
rect 9844 12352 9873 12398
rect 9919 12352 9932 12398
rect 9844 12312 9932 12352
rect 10004 12398 10092 12476
rect 10004 12352 10017 12398
rect 10063 12352 10092 12398
rect 10004 12312 10092 12352
rect 10292 12398 10380 12476
rect 10292 12352 10321 12398
rect 10367 12352 10380 12398
rect 10292 12312 10380 12352
rect 10452 12398 10540 12476
rect 10452 12352 10465 12398
rect 10511 12352 10540 12398
rect 10452 12312 10540 12352
rect 10740 12398 10828 12476
rect 10740 12352 10769 12398
rect 10815 12352 10828 12398
rect 10740 12312 10828 12352
rect 10900 12398 10988 12476
rect 10900 12352 10913 12398
rect 10959 12352 10988 12398
rect 10900 12312 10988 12352
rect 11188 12398 11276 12476
rect 11188 12352 11217 12398
rect 11263 12352 11276 12398
rect 11188 12312 11276 12352
rect 11348 12398 11436 12476
rect 11348 12352 11361 12398
rect 11407 12352 11436 12398
rect 11348 12312 11436 12352
rect 11636 12398 11724 12476
rect 11636 12352 11665 12398
rect 11711 12352 11724 12398
rect 11636 12312 11724 12352
rect 11796 12398 11884 12476
rect 11796 12352 11809 12398
rect 11855 12352 11884 12398
rect 11796 12312 11884 12352
rect 12084 12398 12172 12476
rect 12084 12352 12113 12398
rect 12159 12352 12172 12398
rect 12084 12312 12172 12352
rect 12244 12398 12332 12476
rect 12244 12352 12257 12398
rect 12303 12352 12332 12398
rect 12244 12312 12332 12352
rect 12532 12398 12620 12476
rect 12532 12352 12561 12398
rect 12607 12352 12620 12398
rect 12532 12312 12620 12352
rect 12692 12398 12780 12476
rect 12692 12352 12705 12398
rect 12751 12352 12780 12398
rect 12692 12312 12780 12352
rect 12980 12398 13068 12476
rect 12980 12352 13009 12398
rect 13055 12352 13068 12398
rect 12980 12312 13068 12352
rect 13140 12398 13228 12476
rect 13140 12352 13153 12398
rect 13199 12352 13228 12398
rect 13140 12312 13228 12352
rect 13428 12398 13516 12476
rect 13428 12352 13457 12398
rect 13503 12352 13516 12398
rect 13428 12312 13516 12352
rect 13588 12398 13676 12476
rect 13588 12352 13601 12398
rect 13647 12352 13676 12398
rect 13588 12312 13676 12352
rect 13876 12398 13964 12476
rect 13876 12352 13905 12398
rect 13951 12352 13964 12398
rect 13876 12312 13964 12352
rect 14036 12398 14124 12476
rect 14036 12352 14049 12398
rect 14095 12352 14124 12398
rect 14036 12312 14124 12352
rect 14244 12398 14332 12476
rect 14244 12352 14273 12398
rect 14319 12352 14332 12398
rect 14244 12312 14332 12352
rect 14708 12398 14796 12476
rect 14708 12352 14721 12398
rect 14767 12352 14796 12398
rect 14708 12312 14796 12352
rect 14916 12398 15004 12476
rect 14916 12352 14945 12398
rect 14991 12352 15004 12398
rect 14916 12312 15004 12352
rect 15380 12398 15468 12476
rect 15380 12352 15393 12398
rect 15439 12352 15468 12398
rect 15380 12312 15468 12352
rect 15588 12398 15676 12476
rect 15588 12352 15617 12398
rect 15663 12352 15676 12398
rect 15588 12312 15676 12352
rect 16052 12398 16140 12476
rect 16052 12352 16065 12398
rect 16111 12352 16140 12398
rect 16052 12312 16140 12352
rect 16260 12398 16348 12476
rect 16260 12352 16289 12398
rect 16335 12352 16348 12398
rect 16260 12312 16348 12352
rect 16724 12398 16812 12476
rect 16724 12352 16737 12398
rect 16783 12352 16812 12398
rect 16724 12312 16812 12352
rect 16932 12398 17020 12476
rect 16932 12352 16961 12398
rect 17007 12352 17020 12398
rect 16932 12312 17020 12352
rect 17620 12398 17708 12476
rect 17620 12352 17633 12398
rect 17679 12352 17708 12398
rect 17620 12312 17708 12352
rect 17828 12398 17916 12476
rect 17828 12352 17857 12398
rect 17903 12352 17916 12398
rect 17828 12312 17916 12352
rect 18292 12398 18380 12476
rect 18292 12352 18305 12398
rect 18351 12352 18380 12398
rect 18292 12312 18380 12352
rect 18500 12398 18588 12476
rect 18500 12352 18529 12398
rect 18575 12352 18588 12398
rect 18500 12312 18588 12352
rect 18964 12398 19052 12476
rect 18964 12352 18977 12398
rect 19023 12352 19052 12398
rect 18964 12312 19052 12352
rect 19172 12398 19260 12476
rect 19172 12352 19201 12398
rect 19247 12352 19260 12398
rect 19172 12312 19260 12352
rect 19636 12398 19724 12476
rect 19636 12352 19649 12398
rect 19695 12352 19724 12398
rect 19636 12312 19724 12352
rect 19844 12398 19932 12476
rect 19844 12352 19873 12398
rect 19919 12352 19932 12398
rect 19844 12312 19932 12352
rect 20308 12398 20396 12476
rect 20308 12352 20321 12398
rect 20367 12352 20396 12398
rect 20308 12312 20396 12352
rect 20516 12398 20604 12476
rect 20516 12352 20545 12398
rect 20591 12352 20604 12398
rect 20516 12312 20604 12352
rect 20756 12398 20844 12476
rect 20756 12352 20769 12398
rect 20815 12352 20844 12398
rect 20756 12312 20844 12352
rect 21044 12398 21132 12476
rect 21044 12352 21073 12398
rect 21119 12352 21132 12398
rect 21044 12312 21132 12352
rect 21204 12398 21292 12476
rect 21204 12352 21217 12398
rect 21263 12352 21292 12398
rect 21204 12312 21292 12352
rect 21492 12398 21580 12476
rect 21492 12352 21521 12398
rect 21567 12352 21580 12398
rect 21492 12312 21580 12352
rect 21652 12398 21740 12476
rect 21652 12352 21665 12398
rect 21711 12352 21740 12398
rect 21652 12312 21740 12352
rect 21940 12398 22028 12476
rect 21940 12352 21969 12398
rect 22015 12352 22028 12398
rect 21940 12312 22028 12352
rect 1604 11168 1692 11208
rect 1604 11122 1617 11168
rect 1663 11122 1692 11168
rect 1604 11044 1692 11122
rect 1892 11168 1980 11208
rect 1892 11122 1921 11168
rect 1967 11122 1980 11168
rect 1892 11044 1980 11122
rect 2052 11168 2140 11208
rect 2052 11122 2065 11168
rect 2111 11122 2140 11168
rect 2052 11044 2140 11122
rect 2340 11168 2428 11208
rect 2340 11122 2369 11168
rect 2415 11122 2428 11168
rect 2340 11044 2428 11122
rect 2500 11168 2588 11208
rect 2500 11122 2513 11168
rect 2559 11122 2588 11168
rect 2500 11044 2588 11122
rect 2788 11168 2876 11208
rect 2788 11122 2817 11168
rect 2863 11122 2876 11168
rect 2788 11044 2876 11122
rect 2948 11168 3036 11208
rect 2948 11122 2961 11168
rect 3007 11122 3036 11168
rect 2948 11044 3036 11122
rect 3236 11168 3324 11208
rect 3236 11122 3265 11168
rect 3311 11122 3324 11168
rect 3236 11044 3324 11122
rect 3396 11168 3484 11208
rect 3396 11122 3409 11168
rect 3455 11122 3484 11168
rect 3396 11044 3484 11122
rect 3684 11168 3772 11208
rect 3684 11122 3713 11168
rect 3759 11122 3772 11168
rect 3684 11044 3772 11122
rect 3844 11168 3932 11208
rect 3844 11122 3857 11168
rect 3903 11122 3932 11168
rect 3844 11044 3932 11122
rect 4132 11168 4220 11208
rect 4132 11122 4161 11168
rect 4207 11122 4220 11168
rect 4132 11044 4220 11122
rect 4292 11168 4380 11208
rect 4292 11122 4305 11168
rect 4351 11122 4380 11168
rect 4292 11044 4380 11122
rect 4580 11168 4668 11208
rect 4580 11122 4609 11168
rect 4655 11122 4668 11168
rect 4580 11044 4668 11122
rect 4740 11168 4828 11208
rect 4740 11122 4753 11168
rect 4799 11122 4828 11168
rect 4740 11044 4828 11122
rect 5028 11168 5116 11208
rect 5028 11122 5057 11168
rect 5103 11122 5116 11168
rect 5028 11044 5116 11122
rect 5524 11168 5612 11208
rect 5524 11122 5537 11168
rect 5583 11122 5612 11168
rect 5524 11044 5612 11122
rect 5812 11168 5900 11208
rect 5812 11122 5841 11168
rect 5887 11122 5900 11168
rect 5812 11044 5900 11122
rect 6052 11168 6140 11208
rect 6052 11122 6065 11168
rect 6111 11122 6140 11168
rect 6052 11044 6140 11122
rect 6260 11168 6348 11208
rect 6260 11122 6289 11168
rect 6335 11122 6348 11168
rect 6260 11044 6348 11122
rect 6836 11168 6924 11208
rect 6836 11122 6849 11168
rect 6895 11122 6924 11168
rect 6836 11044 6924 11122
rect 7044 11168 7132 11208
rect 7044 11122 7073 11168
rect 7119 11122 7132 11168
rect 7044 11044 7132 11122
rect 7508 11168 7596 11208
rect 7508 11122 7521 11168
rect 7567 11122 7596 11168
rect 7508 11044 7596 11122
rect 7716 11168 7804 11208
rect 7716 11122 7745 11168
rect 7791 11122 7804 11168
rect 7716 11044 7804 11122
rect 8180 11168 8268 11208
rect 8180 11122 8193 11168
rect 8239 11122 8268 11168
rect 8180 11044 8268 11122
rect 8388 11168 8476 11208
rect 8388 11122 8417 11168
rect 8463 11122 8476 11168
rect 8388 11044 8476 11122
rect 8548 11168 8636 11208
rect 8548 11122 8561 11168
rect 8607 11122 8636 11168
rect 8548 11044 8636 11122
rect 8836 11168 8924 11208
rect 8836 11122 8865 11168
rect 8911 11122 8924 11168
rect 8836 11044 8924 11122
rect 9108 11168 9196 11208
rect 9108 11122 9121 11168
rect 9167 11122 9196 11168
rect 9108 11044 9196 11122
rect 9316 11168 9404 11208
rect 9316 11122 9345 11168
rect 9391 11122 9404 11168
rect 9316 11044 9404 11122
rect 9780 11168 9868 11208
rect 9780 11122 9793 11168
rect 9839 11122 9868 11168
rect 9780 11044 9868 11122
rect 9988 11168 10076 11208
rect 9988 11122 10017 11168
rect 10063 11122 10076 11168
rect 9988 11044 10076 11122
rect 10452 11168 10540 11208
rect 10452 11122 10465 11168
rect 10511 11122 10540 11168
rect 10452 11044 10540 11122
rect 10660 11168 10748 11208
rect 10660 11122 10689 11168
rect 10735 11122 10748 11168
rect 10660 11044 10748 11122
rect 10900 11168 10988 11208
rect 10900 11122 10913 11168
rect 10959 11122 10988 11168
rect 10900 11044 10988 11122
rect 11188 11168 11276 11208
rect 11188 11122 11217 11168
rect 11263 11122 11276 11168
rect 11188 11044 11276 11122
rect 11348 11168 11436 11208
rect 11348 11122 11361 11168
rect 11407 11122 11436 11168
rect 11348 11044 11436 11122
rect 11636 11168 11724 11208
rect 11636 11122 11665 11168
rect 11711 11122 11724 11168
rect 11636 11044 11724 11122
rect 12020 11168 12108 11208
rect 12020 11122 12033 11168
rect 12079 11122 12108 11168
rect 12020 11044 12108 11122
rect 12228 11168 12316 11208
rect 12228 11122 12257 11168
rect 12303 11122 12316 11168
rect 12228 11044 12316 11122
rect 12692 11168 12780 11208
rect 12692 11122 12705 11168
rect 12751 11122 12780 11168
rect 12692 11044 12780 11122
rect 12900 11168 12988 11208
rect 12900 11122 12929 11168
rect 12975 11122 12988 11168
rect 12900 11044 12988 11122
rect 13588 11168 13676 11208
rect 13588 11122 13601 11168
rect 13647 11122 13676 11168
rect 13588 11044 13676 11122
rect 13796 11168 13884 11208
rect 13796 11122 13825 11168
rect 13871 11122 13884 11168
rect 13796 11044 13884 11122
rect 14036 11168 14124 11208
rect 14036 11122 14049 11168
rect 14095 11122 14124 11168
rect 14036 11044 14124 11122
rect 14324 11168 14412 11208
rect 14324 11122 14353 11168
rect 14399 11122 14412 11168
rect 14324 11044 14412 11122
rect 14708 11168 14796 11208
rect 14708 11122 14721 11168
rect 14767 11122 14796 11168
rect 14708 11044 14796 11122
rect 14916 11168 15004 11208
rect 14916 11122 14945 11168
rect 14991 11122 15004 11168
rect 14916 11044 15004 11122
rect 15380 11168 15468 11208
rect 15380 11122 15393 11168
rect 15439 11122 15468 11168
rect 15380 11044 15468 11122
rect 15588 11168 15676 11208
rect 15588 11122 15617 11168
rect 15663 11122 15676 11168
rect 15588 11044 15676 11122
rect 16052 11168 16140 11208
rect 16052 11122 16065 11168
rect 16111 11122 16140 11168
rect 16052 11044 16140 11122
rect 16260 11168 16348 11208
rect 16260 11122 16289 11168
rect 16335 11122 16348 11168
rect 16260 11044 16348 11122
rect 16724 11168 16812 11208
rect 16724 11122 16737 11168
rect 16783 11122 16812 11168
rect 16724 11044 16812 11122
rect 16932 11168 17020 11208
rect 16932 11122 16961 11168
rect 17007 11122 17020 11168
rect 16932 11044 17020 11122
rect 17396 11168 17484 11208
rect 17396 11122 17409 11168
rect 17455 11122 17484 11168
rect 17396 11044 17484 11122
rect 17604 11168 17692 11208
rect 17604 11122 17633 11168
rect 17679 11122 17692 11168
rect 17604 11044 17692 11122
rect 18068 11168 18156 11208
rect 18068 11122 18081 11168
rect 18127 11122 18156 11168
rect 18068 11044 18156 11122
rect 18276 11168 18364 11208
rect 18276 11122 18305 11168
rect 18351 11122 18364 11168
rect 18276 11044 18364 11122
rect 18740 11168 18828 11208
rect 18740 11122 18753 11168
rect 18799 11122 18828 11168
rect 18740 11044 18828 11122
rect 18948 11168 19036 11208
rect 18948 11122 18977 11168
rect 19023 11122 19036 11168
rect 18948 11044 19036 11122
rect 19412 11168 19500 11208
rect 19412 11122 19425 11168
rect 19471 11122 19500 11168
rect 19412 11044 19500 11122
rect 19620 11168 19708 11208
rect 19620 11122 19649 11168
rect 19695 11122 19708 11168
rect 19620 11044 19708 11122
rect 20084 11168 20172 11208
rect 20084 11122 20097 11168
rect 20143 11122 20172 11168
rect 20084 11044 20172 11122
rect 20292 11168 20380 11208
rect 20292 11122 20321 11168
rect 20367 11122 20380 11168
rect 20292 11044 20380 11122
rect 20532 11168 20620 11208
rect 20532 11122 20545 11168
rect 20591 11122 20620 11168
rect 20532 11044 20620 11122
rect 20820 11168 20908 11208
rect 20820 11122 20849 11168
rect 20895 11122 20908 11168
rect 20820 11044 20908 11122
rect 21428 11168 21516 11208
rect 21428 11122 21441 11168
rect 21487 11122 21516 11168
rect 21428 11044 21516 11122
rect 21716 11168 21804 11208
rect 21716 11122 21745 11168
rect 21791 11122 21804 11168
rect 21716 11044 21804 11122
rect 21876 11168 21964 11208
rect 21876 11122 21889 11168
rect 21935 11122 21964 11168
rect 21876 11044 21964 11122
rect 22164 11168 22252 11208
rect 22164 11122 22193 11168
rect 22239 11122 22252 11168
rect 22164 11044 22252 11122
rect 1604 10830 1692 10908
rect 1604 10784 1617 10830
rect 1663 10784 1692 10830
rect 1604 10744 1692 10784
rect 1892 10830 1980 10908
rect 1892 10784 1921 10830
rect 1967 10784 1980 10830
rect 1892 10744 1980 10784
rect 2052 10830 2140 10908
rect 2052 10784 2065 10830
rect 2111 10784 2140 10830
rect 2052 10744 2140 10784
rect 2340 10830 2428 10908
rect 2340 10784 2369 10830
rect 2415 10784 2428 10830
rect 2340 10744 2428 10784
rect 2500 10830 2588 10908
rect 2500 10784 2513 10830
rect 2559 10784 2588 10830
rect 2500 10744 2588 10784
rect 2788 10830 2876 10908
rect 2788 10784 2817 10830
rect 2863 10784 2876 10830
rect 2788 10744 2876 10784
rect 2948 10830 3036 10908
rect 2948 10784 2961 10830
rect 3007 10784 3036 10830
rect 2948 10744 3036 10784
rect 3236 10830 3324 10908
rect 3236 10784 3265 10830
rect 3311 10784 3324 10830
rect 3236 10744 3324 10784
rect 3396 10830 3484 10908
rect 3396 10784 3409 10830
rect 3455 10784 3484 10830
rect 3396 10744 3484 10784
rect 3684 10830 3772 10908
rect 3684 10784 3713 10830
rect 3759 10784 3772 10830
rect 3684 10744 3772 10784
rect 3844 10830 3932 10908
rect 3844 10784 3857 10830
rect 3903 10784 3932 10830
rect 3844 10744 3932 10784
rect 4132 10830 4220 10908
rect 4132 10784 4161 10830
rect 4207 10784 4220 10830
rect 4132 10744 4220 10784
rect 4292 10830 4380 10908
rect 4292 10784 4305 10830
rect 4351 10784 4380 10830
rect 4292 10744 4380 10784
rect 4580 10830 4668 10908
rect 4580 10784 4609 10830
rect 4655 10784 4668 10830
rect 4580 10744 4668 10784
rect 4740 10830 4828 10908
rect 4740 10784 4753 10830
rect 4799 10784 4828 10830
rect 4740 10744 4828 10784
rect 5028 10830 5116 10908
rect 5028 10784 5057 10830
rect 5103 10784 5116 10830
rect 5028 10744 5116 10784
rect 5300 10830 5388 10908
rect 5300 10784 5313 10830
rect 5359 10784 5388 10830
rect 5300 10744 5388 10784
rect 5508 10830 5596 10908
rect 5508 10784 5537 10830
rect 5583 10784 5596 10830
rect 5508 10744 5596 10784
rect 5972 10830 6060 10908
rect 5972 10784 5985 10830
rect 6031 10784 6060 10830
rect 5972 10744 6060 10784
rect 6180 10830 6268 10908
rect 6180 10784 6209 10830
rect 6255 10784 6268 10830
rect 6180 10744 6268 10784
rect 6644 10830 6732 10908
rect 6644 10784 6657 10830
rect 6703 10784 6732 10830
rect 6644 10744 6732 10784
rect 6852 10830 6940 10908
rect 6852 10784 6881 10830
rect 6927 10784 6940 10830
rect 6852 10744 6940 10784
rect 7316 10830 7404 10908
rect 7316 10784 7329 10830
rect 7375 10784 7404 10830
rect 7316 10744 7404 10784
rect 7524 10830 7612 10908
rect 7524 10784 7553 10830
rect 7599 10784 7612 10830
rect 7524 10744 7612 10784
rect 7988 10830 8076 10908
rect 7988 10784 8001 10830
rect 8047 10784 8076 10830
rect 7988 10744 8076 10784
rect 8196 10830 8284 10908
rect 8196 10784 8225 10830
rect 8271 10784 8284 10830
rect 8196 10744 8284 10784
rect 8772 10830 8860 10908
rect 8772 10784 8785 10830
rect 8831 10784 8860 10830
rect 8772 10744 8860 10784
rect 8980 10830 9068 10908
rect 8980 10784 9009 10830
rect 9055 10784 9068 10830
rect 8980 10744 9068 10784
rect 9780 10830 9868 10908
rect 9780 10784 9793 10830
rect 9839 10784 9868 10830
rect 9780 10744 9868 10784
rect 9988 10830 10076 10908
rect 9988 10784 10017 10830
rect 10063 10784 10076 10830
rect 9988 10744 10076 10784
rect 10452 10830 10540 10908
rect 10452 10784 10465 10830
rect 10511 10784 10540 10830
rect 10452 10744 10540 10784
rect 10660 10830 10748 10908
rect 10660 10784 10689 10830
rect 10735 10784 10748 10830
rect 10660 10744 10748 10784
rect 11124 10830 11212 10908
rect 11124 10784 11137 10830
rect 11183 10784 11212 10830
rect 11124 10744 11212 10784
rect 11332 10830 11420 10908
rect 11332 10784 11361 10830
rect 11407 10784 11420 10830
rect 11332 10744 11420 10784
rect 11908 10830 11996 10908
rect 11908 10784 11921 10830
rect 11967 10784 11996 10830
rect 11908 10744 11996 10784
rect 12116 10830 12204 10908
rect 12116 10784 12145 10830
rect 12191 10784 12204 10830
rect 12116 10744 12204 10784
rect 12580 10830 12668 10908
rect 12580 10784 12593 10830
rect 12639 10784 12668 10830
rect 12580 10744 12668 10784
rect 12788 10830 12876 10908
rect 12788 10784 12817 10830
rect 12863 10784 12876 10830
rect 12788 10744 12876 10784
rect 13252 10830 13340 10908
rect 13252 10784 13265 10830
rect 13311 10784 13340 10830
rect 13252 10744 13340 10784
rect 13460 10830 13548 10908
rect 13460 10784 13489 10830
rect 13535 10784 13548 10830
rect 13460 10744 13548 10784
rect 13924 10830 14012 10908
rect 13924 10784 13937 10830
rect 13983 10784 14012 10830
rect 13924 10744 14012 10784
rect 14132 10830 14220 10908
rect 14132 10784 14161 10830
rect 14207 10784 14220 10830
rect 14132 10744 14220 10784
rect 14596 10830 14684 10908
rect 14596 10784 14609 10830
rect 14655 10784 14684 10830
rect 14596 10744 14684 10784
rect 14804 10830 14892 10908
rect 14804 10784 14833 10830
rect 14879 10784 14892 10830
rect 14804 10744 14892 10784
rect 15268 10830 15356 10908
rect 15268 10784 15281 10830
rect 15327 10784 15356 10830
rect 15268 10744 15356 10784
rect 15476 10830 15564 10908
rect 15476 10784 15505 10830
rect 15551 10784 15564 10830
rect 15476 10744 15564 10784
rect 15940 10830 16028 10908
rect 15940 10784 15953 10830
rect 15999 10784 16028 10830
rect 15940 10744 16028 10784
rect 16148 10830 16236 10908
rect 16148 10784 16177 10830
rect 16223 10784 16236 10830
rect 16148 10744 16236 10784
rect 16612 10830 16700 10908
rect 16612 10784 16625 10830
rect 16671 10784 16700 10830
rect 16612 10744 16700 10784
rect 16820 10830 16908 10908
rect 16820 10784 16849 10830
rect 16895 10784 16908 10830
rect 16820 10744 16908 10784
rect 17620 10830 17708 10908
rect 17620 10784 17633 10830
rect 17679 10784 17708 10830
rect 17620 10744 17708 10784
rect 17828 10830 17916 10908
rect 17828 10784 17857 10830
rect 17903 10784 17916 10830
rect 17828 10744 17916 10784
rect 18292 10830 18380 10908
rect 18292 10784 18305 10830
rect 18351 10784 18380 10830
rect 18292 10744 18380 10784
rect 18500 10830 18588 10908
rect 18500 10784 18529 10830
rect 18575 10784 18588 10830
rect 18500 10744 18588 10784
rect 18964 10830 19052 10908
rect 18964 10784 18977 10830
rect 19023 10784 19052 10830
rect 18964 10744 19052 10784
rect 19172 10830 19260 10908
rect 19172 10784 19201 10830
rect 19247 10784 19260 10830
rect 19172 10744 19260 10784
rect 19636 10830 19724 10908
rect 19636 10784 19649 10830
rect 19695 10784 19724 10830
rect 19636 10744 19724 10784
rect 19844 10830 19932 10908
rect 19844 10784 19873 10830
rect 19919 10784 19932 10830
rect 19844 10744 19932 10784
rect 20308 10830 20396 10908
rect 20308 10784 20321 10830
rect 20367 10784 20396 10830
rect 20308 10744 20396 10784
rect 20516 10830 20604 10908
rect 20516 10784 20545 10830
rect 20591 10784 20604 10830
rect 20516 10744 20604 10784
rect 20980 10830 21068 10908
rect 20980 10784 20993 10830
rect 21039 10784 21068 10830
rect 20980 10744 21068 10784
rect 21188 10830 21276 10908
rect 21188 10784 21217 10830
rect 21263 10784 21276 10830
rect 21188 10744 21276 10784
rect 21652 10830 21740 10908
rect 21652 10784 21665 10830
rect 21711 10784 21740 10830
rect 21652 10744 21740 10784
rect 21860 10830 21948 10908
rect 21860 10784 21889 10830
rect 21935 10784 21948 10830
rect 21860 10744 21948 10784
rect 1604 9600 1692 9640
rect 1604 9554 1617 9600
rect 1663 9554 1692 9600
rect 1604 9476 1692 9554
rect 1892 9600 1980 9640
rect 1892 9554 1921 9600
rect 1967 9554 1980 9600
rect 1892 9476 1980 9554
rect 2052 9600 2140 9640
rect 2052 9554 2065 9600
rect 2111 9554 2140 9600
rect 2052 9476 2140 9554
rect 2340 9600 2428 9640
rect 2340 9554 2369 9600
rect 2415 9554 2428 9600
rect 2340 9476 2428 9554
rect 2500 9600 2588 9640
rect 2500 9554 2513 9600
rect 2559 9554 2588 9600
rect 2500 9476 2588 9554
rect 2788 9600 2876 9640
rect 2788 9554 2817 9600
rect 2863 9554 2876 9600
rect 2788 9476 2876 9554
rect 2948 9600 3036 9640
rect 2948 9554 2961 9600
rect 3007 9554 3036 9600
rect 2948 9476 3036 9554
rect 3236 9600 3324 9640
rect 3236 9554 3265 9600
rect 3311 9554 3324 9600
rect 3236 9476 3324 9554
rect 3396 9600 3484 9640
rect 3396 9554 3409 9600
rect 3455 9554 3484 9600
rect 3396 9476 3484 9554
rect 3684 9600 3772 9640
rect 3684 9554 3713 9600
rect 3759 9554 3772 9600
rect 3684 9476 3772 9554
rect 4068 9600 4156 9640
rect 4068 9554 4081 9600
rect 4127 9554 4156 9600
rect 4068 9476 4156 9554
rect 4276 9600 4364 9640
rect 4276 9554 4305 9600
rect 4351 9554 4364 9600
rect 4276 9476 4364 9554
rect 4740 9600 4828 9640
rect 4740 9554 4753 9600
rect 4799 9554 4828 9600
rect 4740 9476 4828 9554
rect 4948 9600 5036 9640
rect 4948 9554 4977 9600
rect 5023 9554 5036 9600
rect 4948 9476 5036 9554
rect 5748 9600 5836 9640
rect 5748 9554 5761 9600
rect 5807 9554 5836 9600
rect 5748 9476 5836 9554
rect 5956 9600 6044 9640
rect 5956 9554 5985 9600
rect 6031 9554 6044 9600
rect 5956 9476 6044 9554
rect 6420 9600 6508 9640
rect 6420 9554 6433 9600
rect 6479 9554 6508 9600
rect 6420 9476 6508 9554
rect 6628 9600 6716 9640
rect 6628 9554 6657 9600
rect 6703 9554 6716 9600
rect 6628 9476 6716 9554
rect 7092 9600 7180 9640
rect 7092 9554 7105 9600
rect 7151 9554 7180 9600
rect 7092 9476 7180 9554
rect 7300 9600 7388 9640
rect 7300 9554 7329 9600
rect 7375 9554 7388 9600
rect 7300 9476 7388 9554
rect 7764 9600 7852 9640
rect 7764 9554 7777 9600
rect 7823 9554 7852 9600
rect 7764 9476 7852 9554
rect 7972 9600 8060 9640
rect 7972 9554 8001 9600
rect 8047 9554 8060 9600
rect 7972 9476 8060 9554
rect 8436 9600 8524 9640
rect 8436 9554 8449 9600
rect 8495 9554 8524 9600
rect 8436 9476 8524 9554
rect 8644 9600 8732 9640
rect 8644 9554 8673 9600
rect 8719 9554 8732 9600
rect 8644 9476 8732 9554
rect 9108 9600 9196 9640
rect 9108 9554 9121 9600
rect 9167 9554 9196 9600
rect 9108 9476 9196 9554
rect 9316 9600 9404 9640
rect 9316 9554 9345 9600
rect 9391 9554 9404 9600
rect 9316 9476 9404 9554
rect 9780 9600 9868 9640
rect 9780 9554 9793 9600
rect 9839 9554 9868 9600
rect 9780 9476 9868 9554
rect 9988 9600 10076 9640
rect 9988 9554 10017 9600
rect 10063 9554 10076 9600
rect 9988 9476 10076 9554
rect 10452 9600 10540 9640
rect 10452 9554 10465 9600
rect 10511 9554 10540 9600
rect 10452 9476 10540 9554
rect 10660 9600 10748 9640
rect 10660 9554 10689 9600
rect 10735 9554 10748 9600
rect 10660 9476 10748 9554
rect 10900 9600 10988 9640
rect 10900 9554 10913 9600
rect 10959 9554 10988 9600
rect 10900 9476 10988 9554
rect 11188 9600 11276 9640
rect 11188 9554 11217 9600
rect 11263 9554 11276 9600
rect 11188 9476 11276 9554
rect 11348 9600 11436 9640
rect 11348 9554 11361 9600
rect 11407 9554 11436 9600
rect 11348 9476 11436 9554
rect 11556 9600 11644 9640
rect 11556 9554 11585 9600
rect 11631 9554 11644 9600
rect 11556 9476 11644 9554
rect 12020 9600 12108 9640
rect 12020 9554 12033 9600
rect 12079 9554 12108 9600
rect 12020 9476 12108 9554
rect 12228 9600 12316 9640
rect 12228 9554 12257 9600
rect 12303 9554 12316 9600
rect 12228 9476 12316 9554
rect 12692 9600 12780 9640
rect 12692 9554 12705 9600
rect 12751 9554 12780 9600
rect 12692 9476 12780 9554
rect 12900 9600 12988 9640
rect 12900 9554 12929 9600
rect 12975 9554 12988 9600
rect 12900 9476 12988 9554
rect 13588 9600 13676 9640
rect 13588 9554 13601 9600
rect 13647 9554 13676 9600
rect 13588 9476 13676 9554
rect 13796 9600 13884 9640
rect 13796 9554 13825 9600
rect 13871 9554 13884 9600
rect 13796 9476 13884 9554
rect 14260 9600 14348 9640
rect 14260 9554 14273 9600
rect 14319 9554 14348 9600
rect 14260 9476 14348 9554
rect 14468 9600 14556 9640
rect 14468 9554 14497 9600
rect 14543 9554 14556 9600
rect 14468 9476 14556 9554
rect 14932 9600 15020 9640
rect 14932 9554 14945 9600
rect 14991 9554 15020 9600
rect 14932 9476 15020 9554
rect 15140 9600 15228 9640
rect 15140 9554 15169 9600
rect 15215 9554 15228 9600
rect 15140 9476 15228 9554
rect 15604 9600 15692 9640
rect 15604 9554 15617 9600
rect 15663 9554 15692 9600
rect 15604 9476 15692 9554
rect 15812 9600 15900 9640
rect 15812 9554 15841 9600
rect 15887 9554 15900 9600
rect 15812 9476 15900 9554
rect 16276 9600 16364 9640
rect 16276 9554 16289 9600
rect 16335 9554 16364 9600
rect 16276 9476 16364 9554
rect 16484 9600 16572 9640
rect 16484 9554 16513 9600
rect 16559 9554 16572 9600
rect 16484 9476 16572 9554
rect 16948 9600 17036 9640
rect 16948 9554 16961 9600
rect 17007 9554 17036 9600
rect 16948 9476 17036 9554
rect 17156 9600 17244 9640
rect 17156 9554 17185 9600
rect 17231 9554 17244 9600
rect 17156 9476 17244 9554
rect 17700 9600 17788 9640
rect 17700 9554 17713 9600
rect 17759 9554 17788 9600
rect 17700 9476 17788 9554
rect 17908 9600 17996 9640
rect 17908 9554 17937 9600
rect 17983 9554 17996 9600
rect 17908 9476 17996 9554
rect 18292 9600 18380 9640
rect 18292 9554 18305 9600
rect 18351 9554 18380 9600
rect 18292 9476 18380 9554
rect 18500 9600 18588 9640
rect 18500 9554 18529 9600
rect 18575 9554 18588 9600
rect 18500 9476 18588 9554
rect 18964 9600 19052 9640
rect 18964 9554 18977 9600
rect 19023 9554 19052 9600
rect 18964 9476 19052 9554
rect 19172 9600 19260 9640
rect 19172 9554 19201 9600
rect 19247 9554 19260 9600
rect 19172 9476 19260 9554
rect 19636 9600 19724 9640
rect 19636 9554 19649 9600
rect 19695 9554 19724 9600
rect 19636 9476 19724 9554
rect 19844 9600 19932 9640
rect 19844 9554 19873 9600
rect 19919 9554 19932 9600
rect 19844 9476 19932 9554
rect 20308 9600 20396 9640
rect 20308 9554 20321 9600
rect 20367 9554 20396 9600
rect 20308 9476 20396 9554
rect 20516 9600 20604 9640
rect 20516 9554 20545 9600
rect 20591 9554 20604 9600
rect 20516 9476 20604 9554
rect 20756 9600 20844 9640
rect 20756 9554 20769 9600
rect 20815 9554 20844 9600
rect 20756 9476 20844 9554
rect 21044 9600 21132 9640
rect 21044 9554 21073 9600
rect 21119 9554 21132 9600
rect 21044 9476 21132 9554
rect 21540 9600 21628 9640
rect 21540 9554 21553 9600
rect 21599 9554 21628 9600
rect 21540 9476 21628 9554
rect 21748 9600 21836 9640
rect 21748 9554 21777 9600
rect 21823 9554 21836 9600
rect 21748 9476 21836 9554
rect 21988 9600 22076 9640
rect 21988 9554 22001 9600
rect 22047 9554 22076 9600
rect 21988 9476 22076 9554
rect 22276 9600 22364 9640
rect 22276 9554 22305 9600
rect 22351 9554 22364 9600
rect 22276 9476 22364 9554
rect 1604 9262 1692 9340
rect 1604 9216 1617 9262
rect 1663 9216 1692 9262
rect 1604 9176 1692 9216
rect 1892 9262 1980 9340
rect 1892 9216 1921 9262
rect 1967 9216 1980 9262
rect 1892 9176 1980 9216
rect 2052 9262 2140 9340
rect 2052 9216 2065 9262
rect 2111 9216 2140 9262
rect 2052 9176 2140 9216
rect 2340 9262 2428 9340
rect 2340 9216 2369 9262
rect 2415 9216 2428 9262
rect 2340 9176 2428 9216
rect 2500 9262 2588 9340
rect 2500 9216 2513 9262
rect 2559 9216 2588 9262
rect 2500 9176 2588 9216
rect 2788 9262 2876 9340
rect 2788 9216 2817 9262
rect 2863 9216 2876 9262
rect 2788 9176 2876 9216
rect 3284 9262 3372 9340
rect 3284 9216 3297 9262
rect 3343 9216 3372 9262
rect 3284 9176 3372 9216
rect 3492 9262 3580 9340
rect 3492 9216 3521 9262
rect 3567 9216 3580 9262
rect 3492 9176 3580 9216
rect 3956 9262 4044 9340
rect 3956 9216 3969 9262
rect 4015 9216 4044 9262
rect 3956 9176 4044 9216
rect 4164 9262 4252 9340
rect 4164 9216 4193 9262
rect 4239 9216 4252 9262
rect 4164 9176 4252 9216
rect 4628 9262 4716 9340
rect 4628 9216 4641 9262
rect 4687 9216 4716 9262
rect 4628 9176 4716 9216
rect 4836 9262 4924 9340
rect 4836 9216 4865 9262
rect 4911 9216 4924 9262
rect 4836 9176 4924 9216
rect 5300 9262 5388 9340
rect 5300 9216 5313 9262
rect 5359 9216 5388 9262
rect 5300 9176 5388 9216
rect 5508 9262 5596 9340
rect 5508 9216 5537 9262
rect 5583 9216 5596 9262
rect 5508 9176 5596 9216
rect 5972 9262 6060 9340
rect 5972 9216 5985 9262
rect 6031 9216 6060 9262
rect 5972 9176 6060 9216
rect 6180 9262 6268 9340
rect 6180 9216 6209 9262
rect 6255 9216 6268 9262
rect 6180 9176 6268 9216
rect 6644 9262 6732 9340
rect 6644 9216 6657 9262
rect 6703 9216 6732 9262
rect 6644 9176 6732 9216
rect 6852 9262 6940 9340
rect 6852 9216 6881 9262
rect 6927 9216 6940 9262
rect 6852 9176 6940 9216
rect 7316 9262 7404 9340
rect 7316 9216 7329 9262
rect 7375 9216 7404 9262
rect 7316 9176 7404 9216
rect 7524 9262 7612 9340
rect 7524 9216 7553 9262
rect 7599 9216 7612 9262
rect 7524 9176 7612 9216
rect 8100 9262 8188 9340
rect 8100 9216 8113 9262
rect 8159 9216 8188 9262
rect 8100 9176 8188 9216
rect 8308 9262 8396 9340
rect 8308 9216 8337 9262
rect 8383 9216 8396 9262
rect 8308 9176 8396 9216
rect 8772 9262 8860 9340
rect 8772 9216 8785 9262
rect 8831 9216 8860 9262
rect 8772 9176 8860 9216
rect 8980 9262 9068 9340
rect 8980 9216 9009 9262
rect 9055 9216 9068 9262
rect 8980 9176 9068 9216
rect 9556 9262 9644 9340
rect 9556 9216 9569 9262
rect 9615 9216 9644 9262
rect 9556 9176 9644 9216
rect 9844 9262 9932 9340
rect 9844 9216 9873 9262
rect 9919 9216 9932 9262
rect 9844 9176 9932 9216
rect 10228 9262 10316 9340
rect 10228 9216 10241 9262
rect 10287 9216 10316 9262
rect 10228 9176 10316 9216
rect 10436 9262 10524 9340
rect 10436 9216 10465 9262
rect 10511 9216 10524 9262
rect 10436 9176 10524 9216
rect 10900 9262 10988 9340
rect 10900 9216 10913 9262
rect 10959 9216 10988 9262
rect 10900 9176 10988 9216
rect 11108 9262 11196 9340
rect 11108 9216 11137 9262
rect 11183 9216 11196 9262
rect 11108 9176 11196 9216
rect 11572 9262 11660 9340
rect 11572 9216 11585 9262
rect 11631 9216 11660 9262
rect 11572 9176 11660 9216
rect 11780 9262 11868 9340
rect 11780 9216 11809 9262
rect 11855 9216 11868 9262
rect 11780 9176 11868 9216
rect 12244 9262 12332 9340
rect 12244 9216 12257 9262
rect 12303 9216 12332 9262
rect 12244 9176 12332 9216
rect 12452 9262 12540 9340
rect 12452 9216 12481 9262
rect 12527 9216 12540 9262
rect 12452 9176 12540 9216
rect 12916 9262 13004 9340
rect 12916 9216 12929 9262
rect 12975 9216 13004 9262
rect 12916 9176 13004 9216
rect 13124 9262 13212 9340
rect 13124 9216 13153 9262
rect 13199 9216 13212 9262
rect 13124 9176 13212 9216
rect 13588 9262 13676 9340
rect 13588 9216 13601 9262
rect 13647 9216 13676 9262
rect 13588 9176 13676 9216
rect 13796 9262 13884 9340
rect 13796 9216 13825 9262
rect 13871 9216 13884 9262
rect 13796 9176 13884 9216
rect 14260 9262 14348 9340
rect 14260 9216 14273 9262
rect 14319 9216 14348 9262
rect 14260 9176 14348 9216
rect 14468 9262 14556 9340
rect 14468 9216 14497 9262
rect 14543 9216 14556 9262
rect 14468 9176 14556 9216
rect 14932 9262 15020 9340
rect 14932 9216 14945 9262
rect 14991 9216 15020 9262
rect 14932 9176 15020 9216
rect 15140 9262 15228 9340
rect 15140 9216 15169 9262
rect 15215 9216 15228 9262
rect 15140 9176 15228 9216
rect 15604 9262 15692 9340
rect 15604 9216 15617 9262
rect 15663 9216 15692 9262
rect 15604 9176 15692 9216
rect 15812 9262 15900 9340
rect 15812 9216 15841 9262
rect 15887 9216 15900 9262
rect 15812 9176 15900 9216
rect 16276 9262 16364 9340
rect 16276 9216 16289 9262
rect 16335 9216 16364 9262
rect 16276 9176 16364 9216
rect 16484 9262 16572 9340
rect 16484 9216 16513 9262
rect 16559 9216 16572 9262
rect 16484 9176 16572 9216
rect 16724 9262 16812 9340
rect 16724 9216 16737 9262
rect 16783 9216 16812 9262
rect 16724 9176 16812 9216
rect 17012 9262 17100 9340
rect 17012 9216 17041 9262
rect 17087 9216 17100 9262
rect 17012 9176 17100 9216
rect 17620 9262 17708 9340
rect 17620 9216 17633 9262
rect 17679 9216 17708 9262
rect 17620 9176 17708 9216
rect 17828 9262 17916 9340
rect 17828 9216 17857 9262
rect 17903 9216 17916 9262
rect 17828 9176 17916 9216
rect 18292 9262 18380 9340
rect 18292 9216 18305 9262
rect 18351 9216 18380 9262
rect 18292 9176 18380 9216
rect 18500 9262 18588 9340
rect 18500 9216 18529 9262
rect 18575 9216 18588 9262
rect 18500 9176 18588 9216
rect 18964 9262 19052 9340
rect 18964 9216 18977 9262
rect 19023 9216 19052 9262
rect 18964 9176 19052 9216
rect 19172 9262 19260 9340
rect 19172 9216 19201 9262
rect 19247 9216 19260 9262
rect 19172 9176 19260 9216
rect 19636 9262 19724 9340
rect 19636 9216 19649 9262
rect 19695 9216 19724 9262
rect 19636 9176 19724 9216
rect 19844 9262 19932 9340
rect 19844 9216 19873 9262
rect 19919 9216 19932 9262
rect 19844 9176 19932 9216
rect 20308 9262 20396 9340
rect 20308 9216 20321 9262
rect 20367 9216 20396 9262
rect 20308 9176 20396 9216
rect 20516 9262 20604 9340
rect 20516 9216 20545 9262
rect 20591 9216 20604 9262
rect 20516 9176 20604 9216
rect 20756 9262 20844 9340
rect 20756 9216 20769 9262
rect 20815 9216 20844 9262
rect 20756 9176 20844 9216
rect 21044 9262 21132 9340
rect 21044 9216 21073 9262
rect 21119 9216 21132 9262
rect 21044 9176 21132 9216
rect 21204 9262 21292 9340
rect 21204 9216 21217 9262
rect 21263 9216 21292 9262
rect 21204 9176 21292 9216
rect 21492 9262 21580 9340
rect 21492 9216 21521 9262
rect 21567 9216 21580 9262
rect 21492 9176 21580 9216
rect 21652 9262 21740 9340
rect 21652 9216 21665 9262
rect 21711 9216 21740 9262
rect 21652 9176 21740 9216
rect 21940 9262 22028 9340
rect 21940 9216 21969 9262
rect 22015 9216 22028 9262
rect 21940 9176 22028 9216
rect 1604 8032 1692 8072
rect 1604 7986 1617 8032
rect 1663 7986 1692 8032
rect 1604 7908 1692 7986
rect 1892 8032 1980 8072
rect 1892 7986 1921 8032
rect 1967 7986 1980 8032
rect 1892 7908 1980 7986
rect 2052 8032 2140 8072
rect 2052 7986 2065 8032
rect 2111 7986 2140 8032
rect 2052 7908 2140 7986
rect 2340 8032 2428 8072
rect 2340 7986 2369 8032
rect 2415 7986 2428 8032
rect 2340 7908 2428 7986
rect 2804 8032 2892 8072
rect 2804 7986 2817 8032
rect 2863 7986 2892 8032
rect 2804 7908 2892 7986
rect 3012 8032 3100 8072
rect 3012 7986 3041 8032
rect 3087 7986 3100 8032
rect 3012 7908 3100 7986
rect 3396 8032 3484 8072
rect 3396 7986 3409 8032
rect 3455 7986 3484 8032
rect 3396 7908 3484 7986
rect 3604 8032 3692 8072
rect 3604 7986 3633 8032
rect 3679 7986 3692 8032
rect 3604 7908 3692 7986
rect 4068 8032 4156 8072
rect 4068 7986 4081 8032
rect 4127 7986 4156 8032
rect 4068 7908 4156 7986
rect 4276 8032 4364 8072
rect 4276 7986 4305 8032
rect 4351 7986 4364 8032
rect 4276 7908 4364 7986
rect 4740 8032 4828 8072
rect 4740 7986 4753 8032
rect 4799 7986 4828 8032
rect 4740 7908 4828 7986
rect 4948 8032 5036 8072
rect 4948 7986 4977 8032
rect 5023 7986 5036 8032
rect 4948 7908 5036 7986
rect 5748 8032 5836 8072
rect 5748 7986 5761 8032
rect 5807 7986 5836 8032
rect 5748 7908 5836 7986
rect 5956 8032 6044 8072
rect 5956 7986 5985 8032
rect 6031 7986 6044 8032
rect 5956 7908 6044 7986
rect 6420 8032 6508 8072
rect 6420 7986 6433 8032
rect 6479 7986 6508 8032
rect 6420 7908 6508 7986
rect 6628 8032 6716 8072
rect 6628 7986 6657 8032
rect 6703 7986 6716 8032
rect 6628 7908 6716 7986
rect 7092 8032 7180 8072
rect 7092 7986 7105 8032
rect 7151 7986 7180 8032
rect 7092 7908 7180 7986
rect 7300 8032 7388 8072
rect 7300 7986 7329 8032
rect 7375 7986 7388 8032
rect 7300 7908 7388 7986
rect 7764 8032 7852 8072
rect 7764 7986 7777 8032
rect 7823 7986 7852 8032
rect 7764 7908 7852 7986
rect 7972 8032 8060 8072
rect 7972 7986 8001 8032
rect 8047 7986 8060 8032
rect 7972 7908 8060 7986
rect 8436 8032 8524 8072
rect 8436 7986 8449 8032
rect 8495 7986 8524 8032
rect 8436 7908 8524 7986
rect 8644 8032 8732 8072
rect 8644 7986 8673 8032
rect 8719 7986 8732 8032
rect 8644 7908 8732 7986
rect 9108 8032 9196 8072
rect 9108 7986 9121 8032
rect 9167 7986 9196 8032
rect 9108 7908 9196 7986
rect 9316 8032 9404 8072
rect 9316 7986 9345 8032
rect 9391 7986 9404 8032
rect 9316 7908 9404 7986
rect 9780 8032 9868 8072
rect 9780 7986 9793 8032
rect 9839 7986 9868 8032
rect 9780 7908 9868 7986
rect 9988 8032 10076 8072
rect 9988 7986 10017 8032
rect 10063 7986 10076 8032
rect 9988 7908 10076 7986
rect 10452 8032 10540 8072
rect 10452 7986 10465 8032
rect 10511 7986 10540 8032
rect 10452 7908 10540 7986
rect 10660 8032 10748 8072
rect 10660 7986 10689 8032
rect 10735 7986 10748 8032
rect 10660 7908 10748 7986
rect 11204 8032 11292 8072
rect 11204 7986 11217 8032
rect 11263 7986 11292 8032
rect 11204 7908 11292 7986
rect 11412 8032 11500 8072
rect 11412 7986 11441 8032
rect 11487 7986 11500 8032
rect 11412 7908 11500 7986
rect 11572 8032 11660 8072
rect 11572 7986 11585 8032
rect 11631 7986 11660 8032
rect 11572 7908 11660 7986
rect 11860 8032 11948 8072
rect 11860 7986 11889 8032
rect 11935 7986 11948 8032
rect 11860 7908 11948 7986
rect 12020 8032 12108 8072
rect 12020 7986 12033 8032
rect 12079 7986 12108 8032
rect 12020 7908 12108 7986
rect 12228 8032 12316 8072
rect 12228 7986 12257 8032
rect 12303 7986 12316 8032
rect 12228 7908 12316 7986
rect 12692 8032 12780 8072
rect 12692 7986 12705 8032
rect 12751 7986 12780 8032
rect 12692 7908 12780 7986
rect 12900 8032 12988 8072
rect 12900 7986 12929 8032
rect 12975 7986 12988 8032
rect 12900 7908 12988 7986
rect 13588 8032 13676 8072
rect 13588 7986 13601 8032
rect 13647 7986 13676 8032
rect 13588 7908 13676 7986
rect 13796 8032 13884 8072
rect 13796 7986 13825 8032
rect 13871 7986 13884 8032
rect 13796 7908 13884 7986
rect 14260 8032 14348 8072
rect 14260 7986 14273 8032
rect 14319 7986 14348 8032
rect 14260 7908 14348 7986
rect 14468 8032 14556 8072
rect 14468 7986 14497 8032
rect 14543 7986 14556 8032
rect 14468 7908 14556 7986
rect 14932 8032 15020 8072
rect 14932 7986 14945 8032
rect 14991 7986 15020 8032
rect 14932 7908 15020 7986
rect 15140 8032 15228 8072
rect 15140 7986 15169 8032
rect 15215 7986 15228 8032
rect 15140 7908 15228 7986
rect 15604 8032 15692 8072
rect 15604 7986 15617 8032
rect 15663 7986 15692 8032
rect 15604 7908 15692 7986
rect 15812 8032 15900 8072
rect 15812 7986 15841 8032
rect 15887 7986 15900 8032
rect 15812 7908 15900 7986
rect 16276 8032 16364 8072
rect 16276 7986 16289 8032
rect 16335 7986 16364 8032
rect 16276 7908 16364 7986
rect 16484 8032 16572 8072
rect 16484 7986 16513 8032
rect 16559 7986 16572 8032
rect 16484 7908 16572 7986
rect 16948 8032 17036 8072
rect 16948 7986 16961 8032
rect 17007 7986 17036 8032
rect 16948 7908 17036 7986
rect 17156 8032 17244 8072
rect 17156 7986 17185 8032
rect 17231 7986 17244 8032
rect 17156 7908 17244 7986
rect 17620 8032 17708 8072
rect 17620 7986 17633 8032
rect 17679 7986 17708 8032
rect 17620 7908 17708 7986
rect 17828 8032 17916 8072
rect 17828 7986 17857 8032
rect 17903 7986 17916 8032
rect 17828 7908 17916 7986
rect 18292 8032 18380 8072
rect 18292 7986 18305 8032
rect 18351 7986 18380 8032
rect 18292 7908 18380 7986
rect 18500 8032 18588 8072
rect 18500 7986 18529 8032
rect 18575 7986 18588 8032
rect 18500 7908 18588 7986
rect 18964 8032 19052 8072
rect 18964 7986 18977 8032
rect 19023 7986 19052 8032
rect 18964 7908 19052 7986
rect 19172 8032 19260 8072
rect 19172 7986 19201 8032
rect 19247 7986 19260 8032
rect 19172 7908 19260 7986
rect 19636 8032 19724 8072
rect 19636 7986 19649 8032
rect 19695 7986 19724 8032
rect 19636 7908 19724 7986
rect 19844 8032 19932 8072
rect 19844 7986 19873 8032
rect 19919 7986 19932 8032
rect 19844 7908 19932 7986
rect 20388 8032 20476 8072
rect 20388 7986 20401 8032
rect 20447 7986 20476 8032
rect 20388 7908 20476 7986
rect 20596 8032 20684 8072
rect 20596 7986 20625 8032
rect 20671 7986 20684 8032
rect 20596 7908 20684 7986
rect 20756 8032 20844 8072
rect 20756 7986 20769 8032
rect 20815 7986 20844 8032
rect 20756 7908 20844 7986
rect 21044 8032 21132 8072
rect 21044 7986 21073 8032
rect 21119 7986 21132 8032
rect 21044 7908 21132 7986
rect 21428 8032 21516 8072
rect 21428 7986 21441 8032
rect 21487 7986 21516 8032
rect 21428 7908 21516 7986
rect 21716 8032 21804 8072
rect 21716 7986 21745 8032
rect 21791 7986 21804 8032
rect 21716 7908 21804 7986
rect 21876 8032 21964 8072
rect 21876 7986 21889 8032
rect 21935 7986 21964 8032
rect 21876 7908 21964 7986
rect 22164 8032 22252 8072
rect 22164 7986 22193 8032
rect 22239 7986 22252 8032
rect 22164 7908 22252 7986
rect 2020 7694 2108 7772
rect 2020 7648 2033 7694
rect 2079 7648 2108 7694
rect 2020 7608 2108 7648
rect 2228 7694 2316 7772
rect 2228 7648 2257 7694
rect 2303 7648 2316 7694
rect 2228 7608 2316 7648
rect 2612 7694 2700 7772
rect 2612 7648 2625 7694
rect 2671 7648 2700 7694
rect 2612 7608 2700 7648
rect 2820 7694 2908 7772
rect 2820 7648 2849 7694
rect 2895 7648 2908 7694
rect 2820 7608 2908 7648
rect 3284 7694 3372 7772
rect 3284 7648 3297 7694
rect 3343 7648 3372 7694
rect 3284 7608 3372 7648
rect 3492 7694 3580 7772
rect 3492 7648 3521 7694
rect 3567 7648 3580 7694
rect 3492 7608 3580 7648
rect 3956 7694 4044 7772
rect 3956 7648 3969 7694
rect 4015 7648 4044 7694
rect 3956 7608 4044 7648
rect 4164 7694 4252 7772
rect 4164 7648 4193 7694
rect 4239 7648 4252 7694
rect 4164 7608 4252 7648
rect 4628 7694 4716 7772
rect 4628 7648 4641 7694
rect 4687 7648 4716 7694
rect 4628 7608 4716 7648
rect 4836 7694 4924 7772
rect 4836 7648 4865 7694
rect 4911 7648 4924 7694
rect 4836 7608 4924 7648
rect 5300 7694 5388 7772
rect 5300 7648 5313 7694
rect 5359 7648 5388 7694
rect 5300 7608 5388 7648
rect 5508 7694 5596 7772
rect 5508 7648 5537 7694
rect 5583 7648 5596 7694
rect 5508 7608 5596 7648
rect 5972 7694 6060 7772
rect 5972 7648 5985 7694
rect 6031 7648 6060 7694
rect 5972 7608 6060 7648
rect 6180 7694 6268 7772
rect 6180 7648 6209 7694
rect 6255 7648 6268 7694
rect 6180 7608 6268 7648
rect 6644 7694 6732 7772
rect 6644 7648 6657 7694
rect 6703 7648 6732 7694
rect 6644 7608 6732 7648
rect 6852 7694 6940 7772
rect 6852 7648 6881 7694
rect 6927 7648 6940 7694
rect 6852 7608 6940 7648
rect 7316 7694 7404 7772
rect 7316 7648 7329 7694
rect 7375 7648 7404 7694
rect 7316 7608 7404 7648
rect 7524 7694 7612 7772
rect 7524 7648 7553 7694
rect 7599 7648 7612 7694
rect 7524 7608 7612 7648
rect 8100 7694 8188 7772
rect 8100 7648 8113 7694
rect 8159 7648 8188 7694
rect 8100 7608 8188 7648
rect 8308 7694 8396 7772
rect 8308 7648 8337 7694
rect 8383 7648 8396 7694
rect 8308 7608 8396 7648
rect 8772 7694 8860 7772
rect 8772 7648 8785 7694
rect 8831 7648 8860 7694
rect 8772 7608 8860 7648
rect 8980 7694 9068 7772
rect 8980 7648 9009 7694
rect 9055 7648 9068 7694
rect 8980 7608 9068 7648
rect 9780 7694 9868 7772
rect 9780 7648 9793 7694
rect 9839 7648 9868 7694
rect 9780 7608 9868 7648
rect 9988 7694 10076 7772
rect 9988 7648 10017 7694
rect 10063 7648 10076 7694
rect 9988 7608 10076 7648
rect 10452 7694 10540 7772
rect 10452 7648 10465 7694
rect 10511 7648 10540 7694
rect 10452 7608 10540 7648
rect 10660 7694 10748 7772
rect 10660 7648 10689 7694
rect 10735 7648 10748 7694
rect 10660 7608 10748 7648
rect 11204 7694 11292 7772
rect 11204 7648 11217 7694
rect 11263 7648 11292 7694
rect 11204 7608 11292 7648
rect 11412 7694 11500 7772
rect 11412 7648 11441 7694
rect 11487 7648 11500 7694
rect 11412 7608 11500 7648
rect 11796 7694 11884 7772
rect 11796 7648 11809 7694
rect 11855 7648 11884 7694
rect 11796 7608 11884 7648
rect 12004 7694 12092 7772
rect 12004 7648 12033 7694
rect 12079 7648 12092 7694
rect 12004 7608 12092 7648
rect 12468 7694 12556 7772
rect 12468 7648 12481 7694
rect 12527 7648 12556 7694
rect 12468 7608 12556 7648
rect 12676 7694 12764 7772
rect 12676 7648 12705 7694
rect 12751 7648 12764 7694
rect 12676 7608 12764 7648
rect 13140 7694 13228 7772
rect 13140 7648 13153 7694
rect 13199 7648 13228 7694
rect 13140 7608 13228 7648
rect 13348 7694 13436 7772
rect 13348 7648 13377 7694
rect 13423 7648 13436 7694
rect 13348 7608 13436 7648
rect 13812 7694 13900 7772
rect 13812 7648 13825 7694
rect 13871 7648 13900 7694
rect 13812 7608 13900 7648
rect 14020 7694 14108 7772
rect 14020 7648 14049 7694
rect 14095 7648 14108 7694
rect 14020 7608 14108 7648
rect 14484 7694 14572 7772
rect 14484 7648 14497 7694
rect 14543 7648 14572 7694
rect 14484 7608 14572 7648
rect 14692 7694 14780 7772
rect 14692 7648 14721 7694
rect 14767 7648 14780 7694
rect 14692 7608 14780 7648
rect 15156 7694 15244 7772
rect 15156 7648 15169 7694
rect 15215 7648 15244 7694
rect 15156 7608 15244 7648
rect 15364 7694 15452 7772
rect 15364 7648 15393 7694
rect 15439 7648 15452 7694
rect 15364 7608 15452 7648
rect 15828 7694 15916 7772
rect 15828 7648 15841 7694
rect 15887 7648 15916 7694
rect 15828 7608 15916 7648
rect 16036 7694 16124 7772
rect 16036 7648 16065 7694
rect 16111 7648 16124 7694
rect 16036 7608 16124 7648
rect 16500 7694 16588 7772
rect 16500 7648 16513 7694
rect 16559 7648 16588 7694
rect 16500 7608 16588 7648
rect 16708 7694 16796 7772
rect 16708 7648 16737 7694
rect 16783 7648 16796 7694
rect 16708 7608 16796 7648
rect 17620 7694 17708 7772
rect 17620 7648 17633 7694
rect 17679 7648 17708 7694
rect 17620 7608 17708 7648
rect 17828 7694 17916 7772
rect 17828 7648 17857 7694
rect 17903 7648 17916 7694
rect 17828 7608 17916 7648
rect 18292 7694 18380 7772
rect 18292 7648 18305 7694
rect 18351 7648 18380 7694
rect 18292 7608 18380 7648
rect 18500 7694 18588 7772
rect 18500 7648 18529 7694
rect 18575 7648 18588 7694
rect 18500 7608 18588 7648
rect 18964 7694 19052 7772
rect 18964 7648 18977 7694
rect 19023 7648 19052 7694
rect 18964 7608 19052 7648
rect 19172 7694 19260 7772
rect 19172 7648 19201 7694
rect 19247 7648 19260 7694
rect 19172 7608 19260 7648
rect 19636 7694 19724 7772
rect 19636 7648 19649 7694
rect 19695 7648 19724 7694
rect 19636 7608 19724 7648
rect 19844 7694 19932 7772
rect 19844 7648 19873 7694
rect 19919 7648 19932 7694
rect 19844 7608 19932 7648
rect 20308 7694 20396 7772
rect 20308 7648 20321 7694
rect 20367 7648 20396 7694
rect 20308 7608 20396 7648
rect 20516 7694 20604 7772
rect 20516 7648 20545 7694
rect 20591 7648 20604 7694
rect 20516 7608 20604 7648
rect 20980 7694 21068 7772
rect 20980 7648 20993 7694
rect 21039 7648 21068 7694
rect 20980 7608 21068 7648
rect 21188 7694 21276 7772
rect 21188 7648 21217 7694
rect 21263 7648 21276 7694
rect 21188 7608 21276 7648
rect 21428 7694 21516 7772
rect 21428 7648 21441 7694
rect 21487 7648 21516 7694
rect 21428 7608 21516 7648
rect 21716 7694 21804 7772
rect 21716 7648 21745 7694
rect 21791 7648 21804 7694
rect 21716 7608 21804 7648
rect 21876 7694 21964 7772
rect 21876 7648 21889 7694
rect 21935 7648 21964 7694
rect 21876 7608 21964 7648
rect 22164 7694 22252 7772
rect 22164 7648 22193 7694
rect 22239 7648 22252 7694
rect 22164 7608 22252 7648
rect 1604 6464 1692 6504
rect 1604 6418 1617 6464
rect 1663 6418 1692 6464
rect 1604 6340 1692 6418
rect 1892 6464 1980 6504
rect 1892 6418 1921 6464
rect 1967 6418 1980 6464
rect 1892 6340 1980 6418
rect 2052 6464 2140 6504
rect 2052 6418 2065 6464
rect 2111 6418 2140 6464
rect 2052 6340 2140 6418
rect 2260 6464 2348 6504
rect 2260 6418 2289 6464
rect 2335 6418 2348 6464
rect 2260 6340 2348 6418
rect 2724 6464 2812 6504
rect 2724 6418 2737 6464
rect 2783 6418 2812 6464
rect 2724 6340 2812 6418
rect 2932 6464 3020 6504
rect 2932 6418 2961 6464
rect 3007 6418 3020 6464
rect 2932 6340 3020 6418
rect 3396 6464 3484 6504
rect 3396 6418 3409 6464
rect 3455 6418 3484 6464
rect 3396 6340 3484 6418
rect 3604 6464 3692 6504
rect 3604 6418 3633 6464
rect 3679 6418 3692 6464
rect 3604 6340 3692 6418
rect 4068 6464 4156 6504
rect 4068 6418 4081 6464
rect 4127 6418 4156 6464
rect 4068 6340 4156 6418
rect 4276 6464 4364 6504
rect 4276 6418 4305 6464
rect 4351 6418 4364 6464
rect 4276 6340 4364 6418
rect 4740 6464 4828 6504
rect 4740 6418 4753 6464
rect 4799 6418 4828 6464
rect 4740 6340 4828 6418
rect 4948 6464 5036 6504
rect 4948 6418 4977 6464
rect 5023 6418 5036 6464
rect 4948 6340 5036 6418
rect 5636 6464 5724 6504
rect 5636 6418 5649 6464
rect 5695 6418 5724 6464
rect 5636 6340 5724 6418
rect 5844 6464 5932 6504
rect 5844 6418 5873 6464
rect 5919 6418 5932 6464
rect 5844 6340 5932 6418
rect 6308 6464 6396 6504
rect 6308 6418 6321 6464
rect 6367 6418 6396 6464
rect 6308 6340 6396 6418
rect 6516 6464 6604 6504
rect 6516 6418 6545 6464
rect 6591 6418 6604 6464
rect 6516 6340 6604 6418
rect 6980 6464 7068 6504
rect 6980 6418 6993 6464
rect 7039 6418 7068 6464
rect 6980 6340 7068 6418
rect 7188 6464 7276 6504
rect 7188 6418 7217 6464
rect 7263 6418 7276 6464
rect 7188 6340 7276 6418
rect 7652 6464 7740 6504
rect 7652 6418 7665 6464
rect 7711 6418 7740 6464
rect 7652 6340 7740 6418
rect 7860 6464 7948 6504
rect 7860 6418 7889 6464
rect 7935 6418 7948 6464
rect 7860 6340 7948 6418
rect 8324 6464 8412 6504
rect 8324 6418 8337 6464
rect 8383 6418 8412 6464
rect 8324 6340 8412 6418
rect 8532 6464 8620 6504
rect 8532 6418 8561 6464
rect 8607 6418 8620 6464
rect 8532 6340 8620 6418
rect 8996 6464 9084 6504
rect 8996 6418 9009 6464
rect 9055 6418 9084 6464
rect 8996 6340 9084 6418
rect 9204 6464 9292 6504
rect 9204 6418 9233 6464
rect 9279 6418 9292 6464
rect 9204 6340 9292 6418
rect 9668 6464 9756 6504
rect 9668 6418 9681 6464
rect 9727 6418 9756 6464
rect 9668 6340 9756 6418
rect 9876 6464 9964 6504
rect 9876 6418 9905 6464
rect 9951 6418 9964 6464
rect 9876 6340 9964 6418
rect 10340 6464 10428 6504
rect 10340 6418 10353 6464
rect 10399 6418 10428 6464
rect 10340 6340 10428 6418
rect 10548 6464 10636 6504
rect 10548 6418 10577 6464
rect 10623 6418 10636 6464
rect 10548 6340 10636 6418
rect 11012 6464 11100 6504
rect 11012 6418 11025 6464
rect 11071 6418 11100 6464
rect 11012 6340 11100 6418
rect 11220 6464 11308 6504
rect 11220 6418 11249 6464
rect 11295 6418 11308 6464
rect 11220 6340 11308 6418
rect 11684 6464 11772 6504
rect 11684 6418 11697 6464
rect 11743 6418 11772 6464
rect 11684 6340 11772 6418
rect 11892 6464 11980 6504
rect 11892 6418 11921 6464
rect 11967 6418 11980 6464
rect 11892 6340 11980 6418
rect 12356 6464 12444 6504
rect 12356 6418 12369 6464
rect 12415 6418 12444 6464
rect 12356 6340 12444 6418
rect 12564 6464 12652 6504
rect 12564 6418 12593 6464
rect 12639 6418 12652 6464
rect 12564 6340 12652 6418
rect 12804 6464 12892 6504
rect 12804 6418 12817 6464
rect 12863 6418 12892 6464
rect 12804 6340 12892 6418
rect 13092 6464 13180 6504
rect 13092 6418 13121 6464
rect 13167 6418 13180 6464
rect 13092 6340 13180 6418
rect 13476 6464 13564 6504
rect 13476 6418 13489 6464
rect 13535 6418 13564 6464
rect 13476 6340 13564 6418
rect 13764 6464 13852 6504
rect 13764 6418 13793 6464
rect 13839 6418 13852 6464
rect 13764 6340 13852 6418
rect 14036 6464 14124 6504
rect 14036 6418 14049 6464
rect 14095 6418 14124 6464
rect 14036 6340 14124 6418
rect 14244 6464 14332 6504
rect 14244 6418 14273 6464
rect 14319 6418 14332 6464
rect 14244 6340 14332 6418
rect 14708 6464 14796 6504
rect 14708 6418 14721 6464
rect 14767 6418 14796 6464
rect 14708 6340 14796 6418
rect 14916 6464 15004 6504
rect 14916 6418 14945 6464
rect 14991 6418 15004 6464
rect 14916 6340 15004 6418
rect 15380 6464 15468 6504
rect 15380 6418 15393 6464
rect 15439 6418 15468 6464
rect 15380 6340 15468 6418
rect 15588 6464 15676 6504
rect 15588 6418 15617 6464
rect 15663 6418 15676 6464
rect 15588 6340 15676 6418
rect 16052 6464 16140 6504
rect 16052 6418 16065 6464
rect 16111 6418 16140 6464
rect 16052 6340 16140 6418
rect 16260 6464 16348 6504
rect 16260 6418 16289 6464
rect 16335 6418 16348 6464
rect 16260 6340 16348 6418
rect 16724 6464 16812 6504
rect 16724 6418 16737 6464
rect 16783 6418 16812 6464
rect 16724 6340 16812 6418
rect 16932 6464 17020 6504
rect 16932 6418 16961 6464
rect 17007 6418 17020 6464
rect 16932 6340 17020 6418
rect 17396 6464 17484 6504
rect 17396 6418 17409 6464
rect 17455 6418 17484 6464
rect 17396 6340 17484 6418
rect 17604 6464 17692 6504
rect 17604 6418 17633 6464
rect 17679 6418 17692 6464
rect 17604 6340 17692 6418
rect 18068 6464 18156 6504
rect 18068 6418 18081 6464
rect 18127 6418 18156 6464
rect 18068 6340 18156 6418
rect 18276 6464 18364 6504
rect 18276 6418 18305 6464
rect 18351 6418 18364 6464
rect 18276 6340 18364 6418
rect 18740 6464 18828 6504
rect 18740 6418 18753 6464
rect 18799 6418 18828 6464
rect 18740 6340 18828 6418
rect 18948 6464 19036 6504
rect 18948 6418 18977 6464
rect 19023 6418 19036 6464
rect 18948 6340 19036 6418
rect 19412 6464 19500 6504
rect 19412 6418 19425 6464
rect 19471 6418 19500 6464
rect 19412 6340 19500 6418
rect 19620 6464 19708 6504
rect 19620 6418 19649 6464
rect 19695 6418 19708 6464
rect 19620 6340 19708 6418
rect 20164 6464 20252 6504
rect 20164 6418 20177 6464
rect 20223 6418 20252 6464
rect 20164 6340 20252 6418
rect 20372 6464 20460 6504
rect 20372 6418 20401 6464
rect 20447 6418 20460 6464
rect 20372 6340 20460 6418
rect 20532 6464 20620 6504
rect 20532 6418 20545 6464
rect 20591 6418 20620 6464
rect 20532 6340 20620 6418
rect 20820 6464 20908 6504
rect 20820 6418 20849 6464
rect 20895 6418 20908 6464
rect 20820 6340 20908 6418
rect 21540 6464 21628 6504
rect 21540 6418 21553 6464
rect 21599 6418 21628 6464
rect 21540 6340 21628 6418
rect 21748 6464 21836 6504
rect 21748 6418 21777 6464
rect 21823 6418 21836 6464
rect 21748 6340 21836 6418
rect 21988 6464 22076 6504
rect 21988 6418 22001 6464
rect 22047 6418 22076 6464
rect 21988 6340 22076 6418
rect 22276 6464 22364 6504
rect 22276 6418 22305 6464
rect 22351 6418 22364 6464
rect 22276 6340 22364 6418
rect 1940 6126 2028 6204
rect 1940 6080 1953 6126
rect 1999 6080 2028 6126
rect 1940 6040 2028 6080
rect 2148 6126 2236 6204
rect 2148 6080 2177 6126
rect 2223 6080 2236 6126
rect 2148 6040 2236 6080
rect 2612 6126 2700 6204
rect 2612 6080 2625 6126
rect 2671 6080 2700 6126
rect 2612 6040 2700 6080
rect 2820 6126 2908 6204
rect 2820 6080 2849 6126
rect 2895 6080 2908 6126
rect 2820 6040 2908 6080
rect 3284 6126 3372 6204
rect 3284 6080 3297 6126
rect 3343 6080 3372 6126
rect 3284 6040 3372 6080
rect 3492 6126 3580 6204
rect 3492 6080 3521 6126
rect 3567 6080 3580 6126
rect 3492 6040 3580 6080
rect 3956 6126 4044 6204
rect 3956 6080 3969 6126
rect 4015 6080 4044 6126
rect 3956 6040 4044 6080
rect 4164 6126 4252 6204
rect 4164 6080 4193 6126
rect 4239 6080 4252 6126
rect 4164 6040 4252 6080
rect 4628 6126 4716 6204
rect 4628 6080 4641 6126
rect 4687 6080 4716 6126
rect 4628 6040 4716 6080
rect 4836 6126 4924 6204
rect 4836 6080 4865 6126
rect 4911 6080 4924 6126
rect 4836 6040 4924 6080
rect 5300 6126 5388 6204
rect 5300 6080 5313 6126
rect 5359 6080 5388 6126
rect 5300 6040 5388 6080
rect 5508 6126 5596 6204
rect 5508 6080 5537 6126
rect 5583 6080 5596 6126
rect 5508 6040 5596 6080
rect 5972 6126 6060 6204
rect 5972 6080 5985 6126
rect 6031 6080 6060 6126
rect 5972 6040 6060 6080
rect 6180 6126 6268 6204
rect 6180 6080 6209 6126
rect 6255 6080 6268 6126
rect 6180 6040 6268 6080
rect 6644 6126 6732 6204
rect 6644 6080 6657 6126
rect 6703 6080 6732 6126
rect 6644 6040 6732 6080
rect 6852 6126 6940 6204
rect 6852 6080 6881 6126
rect 6927 6080 6940 6126
rect 6852 6040 6940 6080
rect 7316 6126 7404 6204
rect 7316 6080 7329 6126
rect 7375 6080 7404 6126
rect 7316 6040 7404 6080
rect 7524 6126 7612 6204
rect 7524 6080 7553 6126
rect 7599 6080 7612 6126
rect 7524 6040 7612 6080
rect 7988 6126 8076 6204
rect 7988 6080 8001 6126
rect 8047 6080 8076 6126
rect 7988 6040 8076 6080
rect 8196 6126 8284 6204
rect 8196 6080 8225 6126
rect 8271 6080 8284 6126
rect 8196 6040 8284 6080
rect 8660 6126 8748 6204
rect 8660 6080 8673 6126
rect 8719 6080 8748 6126
rect 8660 6040 8748 6080
rect 8868 6126 8956 6204
rect 8868 6080 8897 6126
rect 8943 6080 8956 6126
rect 8868 6040 8956 6080
rect 9668 6126 9756 6204
rect 9668 6080 9681 6126
rect 9727 6080 9756 6126
rect 9668 6040 9756 6080
rect 9876 6126 9964 6204
rect 9876 6080 9905 6126
rect 9951 6080 9964 6126
rect 9876 6040 9964 6080
rect 10340 6126 10428 6204
rect 10340 6080 10353 6126
rect 10399 6080 10428 6126
rect 10340 6040 10428 6080
rect 10548 6126 10636 6204
rect 10548 6080 10577 6126
rect 10623 6080 10636 6126
rect 10548 6040 10636 6080
rect 11012 6126 11100 6204
rect 11012 6080 11025 6126
rect 11071 6080 11100 6126
rect 11012 6040 11100 6080
rect 11220 6126 11308 6204
rect 11220 6080 11249 6126
rect 11295 6080 11308 6126
rect 11220 6040 11308 6080
rect 11684 6126 11772 6204
rect 11684 6080 11697 6126
rect 11743 6080 11772 6126
rect 11684 6040 11772 6080
rect 11892 6126 11980 6204
rect 11892 6080 11921 6126
rect 11967 6080 11980 6126
rect 11892 6040 11980 6080
rect 12468 6126 12556 6204
rect 12468 6080 12481 6126
rect 12527 6080 12556 6126
rect 12468 6040 12556 6080
rect 12676 6126 12764 6204
rect 12676 6080 12705 6126
rect 12751 6080 12764 6126
rect 12676 6040 12764 6080
rect 13140 6126 13228 6204
rect 13140 6080 13153 6126
rect 13199 6080 13228 6126
rect 13140 6040 13228 6080
rect 13348 6126 13436 6204
rect 13348 6080 13377 6126
rect 13423 6080 13436 6126
rect 13348 6040 13436 6080
rect 13812 6126 13900 6204
rect 13812 6080 13825 6126
rect 13871 6080 13900 6126
rect 13812 6040 13900 6080
rect 14020 6126 14108 6204
rect 14020 6080 14049 6126
rect 14095 6080 14108 6126
rect 14020 6040 14108 6080
rect 14484 6126 14572 6204
rect 14484 6080 14497 6126
rect 14543 6080 14572 6126
rect 14484 6040 14572 6080
rect 14692 6126 14780 6204
rect 14692 6080 14721 6126
rect 14767 6080 14780 6126
rect 14692 6040 14780 6080
rect 15156 6126 15244 6204
rect 15156 6080 15169 6126
rect 15215 6080 15244 6126
rect 15156 6040 15244 6080
rect 15364 6126 15452 6204
rect 15364 6080 15393 6126
rect 15439 6080 15452 6126
rect 15364 6040 15452 6080
rect 15828 6126 15916 6204
rect 15828 6080 15841 6126
rect 15887 6080 15916 6126
rect 15828 6040 15916 6080
rect 16036 6126 16124 6204
rect 16036 6080 16065 6126
rect 16111 6080 16124 6126
rect 16036 6040 16124 6080
rect 16500 6126 16588 6204
rect 16500 6080 16513 6126
rect 16559 6080 16588 6126
rect 16500 6040 16588 6080
rect 16708 6126 16796 6204
rect 16708 6080 16737 6126
rect 16783 6080 16796 6126
rect 16708 6040 16796 6080
rect 17620 6126 17708 6204
rect 17620 6080 17633 6126
rect 17679 6080 17708 6126
rect 17620 6040 17708 6080
rect 17828 6126 17916 6204
rect 17828 6080 17857 6126
rect 17903 6080 17916 6126
rect 17828 6040 17916 6080
rect 18292 6126 18380 6204
rect 18292 6080 18305 6126
rect 18351 6080 18380 6126
rect 18292 6040 18380 6080
rect 18500 6126 18588 6204
rect 18500 6080 18529 6126
rect 18575 6080 18588 6126
rect 18500 6040 18588 6080
rect 18964 6126 19052 6204
rect 18964 6080 18977 6126
rect 19023 6080 19052 6126
rect 18964 6040 19052 6080
rect 19172 6126 19260 6204
rect 19172 6080 19201 6126
rect 19247 6080 19260 6126
rect 19172 6040 19260 6080
rect 19636 6126 19724 6204
rect 19636 6080 19649 6126
rect 19695 6080 19724 6126
rect 19636 6040 19724 6080
rect 19844 6126 19932 6204
rect 19844 6080 19873 6126
rect 19919 6080 19932 6126
rect 19844 6040 19932 6080
rect 20308 6126 20396 6204
rect 20308 6080 20321 6126
rect 20367 6080 20396 6126
rect 20308 6040 20396 6080
rect 20516 6126 20604 6204
rect 20516 6080 20545 6126
rect 20591 6080 20604 6126
rect 20516 6040 20604 6080
rect 20980 6126 21068 6204
rect 20980 6080 20993 6126
rect 21039 6080 21068 6126
rect 20980 6040 21068 6080
rect 21188 6126 21276 6204
rect 21188 6080 21217 6126
rect 21263 6080 21276 6126
rect 21188 6040 21276 6080
rect 21732 6126 21820 6204
rect 21732 6080 21745 6126
rect 21791 6080 21820 6126
rect 21732 6040 21820 6080
rect 21940 6126 22028 6204
rect 21940 6080 21969 6126
rect 22015 6080 22028 6126
rect 21940 6040 22028 6080
rect 1604 4896 1692 4936
rect 1604 4850 1617 4896
rect 1663 4850 1692 4896
rect 1604 4772 1692 4850
rect 1892 4896 1980 4936
rect 1892 4850 1921 4896
rect 1967 4850 1980 4896
rect 1892 4772 1980 4850
rect 2052 4896 2140 4936
rect 2052 4850 2065 4896
rect 2111 4850 2140 4896
rect 2052 4772 2140 4850
rect 2260 4896 2348 4936
rect 2260 4850 2289 4896
rect 2335 4850 2348 4896
rect 2260 4772 2348 4850
rect 2724 4896 2812 4936
rect 2724 4850 2737 4896
rect 2783 4850 2812 4896
rect 2724 4772 2812 4850
rect 2932 4896 3020 4936
rect 2932 4850 2961 4896
rect 3007 4850 3020 4896
rect 2932 4772 3020 4850
rect 3396 4896 3484 4936
rect 3396 4850 3409 4896
rect 3455 4850 3484 4896
rect 3396 4772 3484 4850
rect 3604 4896 3692 4936
rect 3604 4850 3633 4896
rect 3679 4850 3692 4896
rect 3604 4772 3692 4850
rect 4068 4896 4156 4936
rect 4068 4850 4081 4896
rect 4127 4850 4156 4896
rect 4068 4772 4156 4850
rect 4276 4896 4364 4936
rect 4276 4850 4305 4896
rect 4351 4850 4364 4896
rect 4276 4772 4364 4850
rect 4740 4896 4828 4936
rect 4740 4850 4753 4896
rect 4799 4850 4828 4896
rect 4740 4772 4828 4850
rect 4948 4896 5036 4936
rect 4948 4850 4977 4896
rect 5023 4850 5036 4896
rect 4948 4772 5036 4850
rect 5636 4896 5724 4936
rect 5636 4850 5649 4896
rect 5695 4850 5724 4896
rect 5636 4772 5724 4850
rect 5844 4896 5932 4936
rect 5844 4850 5873 4896
rect 5919 4850 5932 4896
rect 5844 4772 5932 4850
rect 6308 4896 6396 4936
rect 6308 4850 6321 4896
rect 6367 4850 6396 4896
rect 6308 4772 6396 4850
rect 6516 4896 6604 4936
rect 6516 4850 6545 4896
rect 6591 4850 6604 4896
rect 6516 4772 6604 4850
rect 6980 4896 7068 4936
rect 6980 4850 6993 4896
rect 7039 4850 7068 4896
rect 6980 4772 7068 4850
rect 7188 4896 7276 4936
rect 7188 4850 7217 4896
rect 7263 4850 7276 4896
rect 7188 4772 7276 4850
rect 7652 4896 7740 4936
rect 7652 4850 7665 4896
rect 7711 4850 7740 4896
rect 7652 4772 7740 4850
rect 7860 4896 7948 4936
rect 7860 4850 7889 4896
rect 7935 4850 7948 4896
rect 7860 4772 7948 4850
rect 8324 4896 8412 4936
rect 8324 4850 8337 4896
rect 8383 4850 8412 4896
rect 8324 4772 8412 4850
rect 8532 4896 8620 4936
rect 8532 4850 8561 4896
rect 8607 4850 8620 4896
rect 8532 4772 8620 4850
rect 8996 4896 9084 4936
rect 8996 4850 9009 4896
rect 9055 4850 9084 4896
rect 8996 4772 9084 4850
rect 9204 4896 9292 4936
rect 9204 4850 9233 4896
rect 9279 4850 9292 4896
rect 9204 4772 9292 4850
rect 9668 4896 9756 4936
rect 9668 4850 9681 4896
rect 9727 4850 9756 4896
rect 9668 4772 9756 4850
rect 9876 4896 9964 4936
rect 9876 4850 9905 4896
rect 9951 4850 9964 4896
rect 9876 4772 9964 4850
rect 10340 4896 10428 4936
rect 10340 4850 10353 4896
rect 10399 4850 10428 4896
rect 10340 4772 10428 4850
rect 10548 4896 10636 4936
rect 10548 4850 10577 4896
rect 10623 4850 10636 4896
rect 10548 4772 10636 4850
rect 10788 4896 10876 4936
rect 10788 4850 10801 4896
rect 10847 4850 10876 4896
rect 10788 4772 10876 4850
rect 11076 4896 11164 4936
rect 11076 4850 11105 4896
rect 11151 4850 11164 4896
rect 11076 4772 11164 4850
rect 11348 4896 11436 4936
rect 11348 4850 11361 4896
rect 11407 4850 11436 4896
rect 11348 4772 11436 4850
rect 11556 4896 11644 4936
rect 11556 4850 11585 4896
rect 11631 4850 11644 4896
rect 11556 4772 11644 4850
rect 12020 4896 12108 4936
rect 12020 4850 12033 4896
rect 12079 4850 12108 4896
rect 12020 4772 12108 4850
rect 12228 4896 12316 4936
rect 12228 4850 12257 4896
rect 12303 4850 12316 4896
rect 12228 4772 12316 4850
rect 12692 4896 12780 4936
rect 12692 4850 12705 4896
rect 12751 4850 12780 4896
rect 12692 4772 12780 4850
rect 12900 4896 12988 4936
rect 12900 4850 12929 4896
rect 12975 4850 12988 4896
rect 12900 4772 12988 4850
rect 13476 4896 13564 4936
rect 13476 4850 13489 4896
rect 13535 4850 13564 4896
rect 13476 4772 13564 4850
rect 13764 4896 13852 4936
rect 13764 4850 13793 4896
rect 13839 4850 13852 4896
rect 13764 4772 13852 4850
rect 13924 4896 14012 4936
rect 13924 4850 13937 4896
rect 13983 4850 14012 4896
rect 13924 4772 14012 4850
rect 14132 4896 14220 4936
rect 14132 4850 14161 4896
rect 14207 4850 14220 4896
rect 14132 4772 14220 4850
rect 14596 4896 14684 4936
rect 14596 4850 14609 4896
rect 14655 4850 14684 4896
rect 14596 4772 14684 4850
rect 14804 4896 14892 4936
rect 14804 4850 14833 4896
rect 14879 4850 14892 4896
rect 14804 4772 14892 4850
rect 15268 4896 15356 4936
rect 15268 4850 15281 4896
rect 15327 4850 15356 4896
rect 15268 4772 15356 4850
rect 15476 4896 15564 4936
rect 15476 4850 15505 4896
rect 15551 4850 15564 4896
rect 15476 4772 15564 4850
rect 15940 4896 16028 4936
rect 15940 4850 15953 4896
rect 15999 4850 16028 4896
rect 15940 4772 16028 4850
rect 16148 4896 16236 4936
rect 16148 4850 16177 4896
rect 16223 4850 16236 4896
rect 16148 4772 16236 4850
rect 16612 4896 16700 4936
rect 16612 4850 16625 4896
rect 16671 4850 16700 4896
rect 16612 4772 16700 4850
rect 16820 4896 16908 4936
rect 16820 4850 16849 4896
rect 16895 4850 16908 4896
rect 16820 4772 16908 4850
rect 17284 4896 17372 4936
rect 17284 4850 17297 4896
rect 17343 4850 17372 4896
rect 17284 4772 17372 4850
rect 17492 4896 17580 4936
rect 17492 4850 17521 4896
rect 17567 4850 17580 4896
rect 17492 4772 17580 4850
rect 17956 4896 18044 4936
rect 17956 4850 17969 4896
rect 18015 4850 18044 4896
rect 17956 4772 18044 4850
rect 18164 4896 18252 4936
rect 18164 4850 18193 4896
rect 18239 4850 18252 4896
rect 18164 4772 18252 4850
rect 18628 4896 18716 4936
rect 18628 4850 18641 4896
rect 18687 4850 18716 4896
rect 18628 4772 18716 4850
rect 18836 4896 18924 4936
rect 18836 4850 18865 4896
rect 18911 4850 18924 4896
rect 18836 4772 18924 4850
rect 19300 4896 19388 4936
rect 19300 4850 19313 4896
rect 19359 4850 19388 4896
rect 19300 4772 19388 4850
rect 19508 4896 19596 4936
rect 19508 4850 19537 4896
rect 19583 4850 19596 4896
rect 19508 4772 19596 4850
rect 19972 4896 20060 4936
rect 19972 4850 19985 4896
rect 20031 4850 20060 4896
rect 19972 4772 20060 4850
rect 20180 4896 20268 4936
rect 20180 4850 20209 4896
rect 20255 4850 20268 4896
rect 20180 4772 20268 4850
rect 20644 4896 20732 4936
rect 20644 4850 20657 4896
rect 20703 4850 20732 4896
rect 20644 4772 20732 4850
rect 20852 4896 20940 4936
rect 20852 4850 20881 4896
rect 20927 4850 20940 4896
rect 20852 4772 20940 4850
rect 21540 4896 21628 4936
rect 21540 4850 21553 4896
rect 21599 4850 21628 4896
rect 21540 4772 21628 4850
rect 21748 4896 21836 4936
rect 21748 4850 21777 4896
rect 21823 4850 21836 4896
rect 21748 4772 21836 4850
rect 21988 4896 22076 4936
rect 21988 4850 22001 4896
rect 22047 4850 22076 4896
rect 21988 4772 22076 4850
rect 22276 4896 22364 4936
rect 22276 4850 22305 4896
rect 22351 4850 22364 4896
rect 22276 4772 22364 4850
rect 1604 4558 1692 4636
rect 1604 4512 1617 4558
rect 1663 4512 1692 4558
rect 1604 4472 1692 4512
rect 1892 4558 1980 4636
rect 1892 4512 1921 4558
rect 1967 4512 1980 4558
rect 1892 4472 1980 4512
rect 2276 4558 2364 4636
rect 2276 4512 2289 4558
rect 2335 4512 2364 4558
rect 2276 4472 2364 4512
rect 2484 4558 2572 4636
rect 2484 4512 2513 4558
rect 2559 4512 2572 4558
rect 2484 4472 2572 4512
rect 2948 4558 3036 4636
rect 2948 4512 2961 4558
rect 3007 4512 3036 4558
rect 2948 4472 3036 4512
rect 3156 4558 3244 4636
rect 3156 4512 3185 4558
rect 3231 4512 3244 4558
rect 3156 4472 3244 4512
rect 3620 4558 3708 4636
rect 3620 4512 3633 4558
rect 3679 4512 3708 4558
rect 3620 4472 3708 4512
rect 3828 4558 3916 4636
rect 3828 4512 3857 4558
rect 3903 4512 3916 4558
rect 3828 4472 3916 4512
rect 4292 4558 4380 4636
rect 4292 4512 4305 4558
rect 4351 4512 4380 4558
rect 4292 4472 4380 4512
rect 4500 4558 4588 4636
rect 4500 4512 4529 4558
rect 4575 4512 4588 4558
rect 4500 4472 4588 4512
rect 4964 4558 5052 4636
rect 4964 4512 4977 4558
rect 5023 4512 5052 4558
rect 4964 4472 5052 4512
rect 5172 4558 5260 4636
rect 5172 4512 5201 4558
rect 5247 4512 5260 4558
rect 5172 4472 5260 4512
rect 5636 4558 5724 4636
rect 5636 4512 5649 4558
rect 5695 4512 5724 4558
rect 5636 4472 5724 4512
rect 5844 4558 5932 4636
rect 5844 4512 5873 4558
rect 5919 4512 5932 4558
rect 5844 4472 5932 4512
rect 6308 4558 6396 4636
rect 6308 4512 6321 4558
rect 6367 4512 6396 4558
rect 6308 4472 6396 4512
rect 6516 4558 6604 4636
rect 6516 4512 6545 4558
rect 6591 4512 6604 4558
rect 6516 4472 6604 4512
rect 6980 4558 7068 4636
rect 6980 4512 6993 4558
rect 7039 4512 7068 4558
rect 6980 4472 7068 4512
rect 7188 4558 7276 4636
rect 7188 4512 7217 4558
rect 7263 4512 7276 4558
rect 7188 4472 7276 4512
rect 7652 4558 7740 4636
rect 7652 4512 7665 4558
rect 7711 4512 7740 4558
rect 7652 4472 7740 4512
rect 7860 4558 7948 4636
rect 7860 4512 7889 4558
rect 7935 4512 7948 4558
rect 7860 4472 7948 4512
rect 8324 4558 8412 4636
rect 8324 4512 8337 4558
rect 8383 4512 8412 4558
rect 8324 4472 8412 4512
rect 8532 4558 8620 4636
rect 8532 4512 8561 4558
rect 8607 4512 8620 4558
rect 8532 4472 8620 4512
rect 8772 4558 8860 4636
rect 8772 4512 8785 4558
rect 8831 4512 8860 4558
rect 8772 4472 8860 4512
rect 9060 4558 9148 4636
rect 9060 4512 9089 4558
rect 9135 4512 9148 4558
rect 9060 4472 9148 4512
rect 9668 4558 9756 4636
rect 9668 4512 9681 4558
rect 9727 4512 9756 4558
rect 9668 4472 9756 4512
rect 9876 4558 9964 4636
rect 9876 4512 9905 4558
rect 9951 4512 9964 4558
rect 9876 4472 9964 4512
rect 10340 4558 10428 4636
rect 10340 4512 10353 4558
rect 10399 4512 10428 4558
rect 10340 4472 10428 4512
rect 10548 4558 10636 4636
rect 10548 4512 10577 4558
rect 10623 4512 10636 4558
rect 10548 4472 10636 4512
rect 11012 4558 11100 4636
rect 11012 4512 11025 4558
rect 11071 4512 11100 4558
rect 11012 4472 11100 4512
rect 11220 4558 11308 4636
rect 11220 4512 11249 4558
rect 11295 4512 11308 4558
rect 11220 4472 11308 4512
rect 11460 4558 11548 4636
rect 11460 4512 11473 4558
rect 11519 4512 11548 4558
rect 11460 4472 11548 4512
rect 11748 4558 11836 4636
rect 11748 4512 11777 4558
rect 11823 4512 11836 4558
rect 11748 4472 11836 4512
rect 12244 4558 12332 4636
rect 12244 4512 12257 4558
rect 12303 4512 12332 4558
rect 12244 4472 12332 4512
rect 12452 4558 12540 4636
rect 12452 4512 12481 4558
rect 12527 4512 12540 4558
rect 12452 4472 12540 4512
rect 12916 4558 13004 4636
rect 12916 4512 12929 4558
rect 12975 4512 13004 4558
rect 12916 4472 13004 4512
rect 13124 4558 13212 4636
rect 13124 4512 13153 4558
rect 13199 4512 13212 4558
rect 13124 4472 13212 4512
rect 13588 4558 13676 4636
rect 13588 4512 13601 4558
rect 13647 4512 13676 4558
rect 13588 4472 13676 4512
rect 13796 4558 13884 4636
rect 13796 4512 13825 4558
rect 13871 4512 13884 4558
rect 13796 4472 13884 4512
rect 14260 4558 14348 4636
rect 14260 4512 14273 4558
rect 14319 4512 14348 4558
rect 14260 4472 14348 4512
rect 14468 4558 14556 4636
rect 14468 4512 14497 4558
rect 14543 4512 14556 4558
rect 14468 4472 14556 4512
rect 14932 4558 15020 4636
rect 14932 4512 14945 4558
rect 14991 4512 15020 4558
rect 14932 4472 15020 4512
rect 15140 4558 15228 4636
rect 15140 4512 15169 4558
rect 15215 4512 15228 4558
rect 15140 4472 15228 4512
rect 15604 4558 15692 4636
rect 15604 4512 15617 4558
rect 15663 4512 15692 4558
rect 15604 4472 15692 4512
rect 15812 4558 15900 4636
rect 15812 4512 15841 4558
rect 15887 4512 15900 4558
rect 15812 4472 15900 4512
rect 16276 4558 16364 4636
rect 16276 4512 16289 4558
rect 16335 4512 16364 4558
rect 16276 4472 16364 4512
rect 16484 4558 16572 4636
rect 16484 4512 16513 4558
rect 16559 4512 16572 4558
rect 16484 4472 16572 4512
rect 16724 4558 16812 4636
rect 16724 4512 16737 4558
rect 16783 4512 16812 4558
rect 16724 4472 16812 4512
rect 17012 4558 17100 4636
rect 17012 4512 17041 4558
rect 17087 4512 17100 4558
rect 17012 4472 17100 4512
rect 17620 4558 17708 4636
rect 17620 4512 17633 4558
rect 17679 4512 17708 4558
rect 17620 4472 17708 4512
rect 17828 4558 17916 4636
rect 17828 4512 17857 4558
rect 17903 4512 17916 4558
rect 17828 4472 17916 4512
rect 18292 4558 18380 4636
rect 18292 4512 18305 4558
rect 18351 4512 18380 4558
rect 18292 4472 18380 4512
rect 18500 4558 18588 4636
rect 18500 4512 18529 4558
rect 18575 4512 18588 4558
rect 18500 4472 18588 4512
rect 18964 4558 19052 4636
rect 18964 4512 18977 4558
rect 19023 4512 19052 4558
rect 18964 4472 19052 4512
rect 19172 4558 19260 4636
rect 19172 4512 19201 4558
rect 19247 4512 19260 4558
rect 19172 4472 19260 4512
rect 19636 4558 19724 4636
rect 19636 4512 19649 4558
rect 19695 4512 19724 4558
rect 19636 4472 19724 4512
rect 19844 4558 19932 4636
rect 19844 4512 19873 4558
rect 19919 4512 19932 4558
rect 19844 4472 19932 4512
rect 20308 4558 20396 4636
rect 20308 4512 20321 4558
rect 20367 4512 20396 4558
rect 20308 4472 20396 4512
rect 20516 4558 20604 4636
rect 20516 4512 20545 4558
rect 20591 4512 20604 4558
rect 20516 4472 20604 4512
rect 20980 4558 21068 4636
rect 20980 4512 20993 4558
rect 21039 4512 21068 4558
rect 20980 4472 21068 4512
rect 21188 4558 21276 4636
rect 21188 4512 21217 4558
rect 21263 4512 21276 4558
rect 21188 4472 21276 4512
rect 21732 4558 21820 4636
rect 21732 4512 21745 4558
rect 21791 4512 21820 4558
rect 21732 4472 21820 4512
rect 21940 4558 22028 4636
rect 21940 4512 21969 4558
rect 22015 4512 22028 4558
rect 21940 4472 22028 4512
rect 1604 3328 1692 3368
rect 1604 3282 1617 3328
rect 1663 3282 1692 3328
rect 1604 3204 1692 3282
rect 1892 3328 1980 3368
rect 1892 3282 1921 3328
rect 1967 3282 1980 3328
rect 1892 3204 1980 3282
rect 2052 3328 2140 3368
rect 2052 3282 2065 3328
rect 2111 3282 2140 3328
rect 2052 3204 2140 3282
rect 2340 3328 2428 3368
rect 2340 3282 2369 3328
rect 2415 3282 2428 3328
rect 2340 3204 2428 3282
rect 2724 3328 2812 3368
rect 2724 3282 2737 3328
rect 2783 3282 2812 3328
rect 2724 3204 2812 3282
rect 2932 3328 3020 3368
rect 2932 3282 2961 3328
rect 3007 3282 3020 3328
rect 2932 3204 3020 3282
rect 3396 3328 3484 3368
rect 3396 3282 3409 3328
rect 3455 3282 3484 3328
rect 3396 3204 3484 3282
rect 3604 3328 3692 3368
rect 3604 3282 3633 3328
rect 3679 3282 3692 3328
rect 3604 3204 3692 3282
rect 4068 3328 4156 3368
rect 4068 3282 4081 3328
rect 4127 3282 4156 3328
rect 4068 3204 4156 3282
rect 4276 3328 4364 3368
rect 4276 3282 4305 3328
rect 4351 3282 4364 3328
rect 4276 3204 4364 3282
rect 4740 3328 4828 3368
rect 4740 3282 4753 3328
rect 4799 3282 4828 3328
rect 4740 3204 4828 3282
rect 4948 3328 5036 3368
rect 4948 3282 4977 3328
rect 5023 3282 5036 3328
rect 4948 3204 5036 3282
rect 5716 3328 5804 3368
rect 5716 3282 5729 3328
rect 5775 3282 5804 3328
rect 5716 3204 5804 3282
rect 5924 3328 6012 3368
rect 5924 3282 5953 3328
rect 5999 3282 6012 3328
rect 5924 3204 6012 3282
rect 6388 3328 6476 3368
rect 6388 3282 6401 3328
rect 6447 3282 6476 3328
rect 6388 3204 6476 3282
rect 6596 3328 6684 3368
rect 6596 3282 6625 3328
rect 6671 3282 6684 3328
rect 6596 3204 6684 3282
rect 7060 3328 7148 3368
rect 7060 3282 7073 3328
rect 7119 3282 7148 3328
rect 7060 3204 7148 3282
rect 7268 3328 7356 3368
rect 7268 3282 7297 3328
rect 7343 3282 7356 3328
rect 7268 3204 7356 3282
rect 7652 3328 7740 3368
rect 7652 3282 7665 3328
rect 7711 3282 7740 3328
rect 7652 3204 7740 3282
rect 7860 3328 7948 3368
rect 7860 3282 7889 3328
rect 7935 3282 7948 3328
rect 7860 3204 7948 3282
rect 8404 3328 8492 3368
rect 8404 3282 8417 3328
rect 8463 3282 8492 3328
rect 8404 3204 8492 3282
rect 8612 3328 8700 3368
rect 8612 3282 8641 3328
rect 8687 3282 8700 3328
rect 8612 3204 8700 3282
rect 8772 3328 8860 3368
rect 8772 3282 8785 3328
rect 8831 3282 8860 3328
rect 8772 3204 8860 3282
rect 9060 3328 9148 3368
rect 9060 3282 9089 3328
rect 9135 3282 9148 3328
rect 9060 3204 9148 3282
rect 9636 3328 9724 3368
rect 9636 3282 9649 3328
rect 9695 3282 9724 3328
rect 9636 3204 9724 3282
rect 9844 3328 9932 3368
rect 9844 3282 9873 3328
rect 9919 3282 9932 3328
rect 9844 3204 9932 3282
rect 10228 3328 10316 3368
rect 10228 3282 10241 3328
rect 10287 3282 10316 3328
rect 10228 3204 10316 3282
rect 10436 3328 10524 3368
rect 10436 3282 10465 3328
rect 10511 3282 10524 3328
rect 10436 3204 10524 3282
rect 10900 3328 10988 3368
rect 10900 3282 10913 3328
rect 10959 3282 10988 3328
rect 10900 3204 10988 3282
rect 11108 3328 11196 3368
rect 11108 3282 11137 3328
rect 11183 3282 11196 3328
rect 11108 3204 11196 3282
rect 11652 3328 11740 3368
rect 11652 3282 11665 3328
rect 11711 3282 11740 3328
rect 11652 3204 11740 3282
rect 11860 3328 11948 3368
rect 11860 3282 11889 3328
rect 11935 3282 11948 3328
rect 11860 3204 11948 3282
rect 12020 3328 12108 3368
rect 12020 3282 12033 3328
rect 12079 3282 12108 3328
rect 12020 3204 12108 3282
rect 12308 3328 12396 3368
rect 12308 3282 12337 3328
rect 12383 3282 12396 3328
rect 12308 3204 12396 3282
rect 12468 3328 12556 3368
rect 12468 3282 12481 3328
rect 12527 3282 12556 3328
rect 12468 3204 12556 3282
rect 12756 3328 12844 3368
rect 12756 3282 12785 3328
rect 12831 3282 12844 3328
rect 12756 3204 12844 3282
rect 13364 3328 13452 3368
rect 13364 3282 13377 3328
rect 13423 3282 13452 3328
rect 13364 3204 13452 3282
rect 13652 3328 13740 3368
rect 13652 3282 13681 3328
rect 13727 3282 13740 3328
rect 13652 3204 13740 3282
rect 13812 3328 13900 3368
rect 13812 3282 13825 3328
rect 13871 3282 13900 3328
rect 13812 3204 13900 3282
rect 14020 3328 14108 3368
rect 14020 3282 14049 3328
rect 14095 3282 14108 3328
rect 14020 3204 14108 3282
rect 14484 3328 14572 3368
rect 14484 3282 14497 3328
rect 14543 3282 14572 3328
rect 14484 3204 14572 3282
rect 14692 3328 14780 3368
rect 14692 3282 14721 3328
rect 14767 3282 14780 3328
rect 14692 3204 14780 3282
rect 15156 3328 15244 3368
rect 15156 3282 15169 3328
rect 15215 3282 15244 3328
rect 15156 3204 15244 3282
rect 15364 3328 15452 3368
rect 15364 3282 15393 3328
rect 15439 3282 15452 3328
rect 15364 3204 15452 3282
rect 15828 3328 15916 3368
rect 15828 3282 15841 3328
rect 15887 3282 15916 3328
rect 15828 3204 15916 3282
rect 16036 3328 16124 3368
rect 16036 3282 16065 3328
rect 16111 3282 16124 3328
rect 16036 3204 16124 3282
rect 16500 3328 16588 3368
rect 16500 3282 16513 3328
rect 16559 3282 16588 3328
rect 16500 3204 16588 3282
rect 16708 3328 16796 3368
rect 16708 3282 16737 3328
rect 16783 3282 16796 3328
rect 16708 3204 16796 3282
rect 17396 3328 17484 3368
rect 17396 3282 17409 3328
rect 17455 3282 17484 3328
rect 17396 3204 17484 3282
rect 17604 3328 17692 3368
rect 17604 3282 17633 3328
rect 17679 3282 17692 3328
rect 17604 3204 17692 3282
rect 18068 3328 18156 3368
rect 18068 3282 18081 3328
rect 18127 3282 18156 3328
rect 18068 3204 18156 3282
rect 18276 3328 18364 3368
rect 18276 3282 18305 3328
rect 18351 3282 18364 3328
rect 18276 3204 18364 3282
rect 18740 3328 18828 3368
rect 18740 3282 18753 3328
rect 18799 3282 18828 3328
rect 18740 3204 18828 3282
rect 18948 3328 19036 3368
rect 18948 3282 18977 3328
rect 19023 3282 19036 3328
rect 18948 3204 19036 3282
rect 19412 3328 19500 3368
rect 19412 3282 19425 3328
rect 19471 3282 19500 3328
rect 19412 3204 19500 3282
rect 19620 3328 19708 3368
rect 19620 3282 19649 3328
rect 19695 3282 19708 3328
rect 19620 3204 19708 3282
rect 20084 3328 20172 3368
rect 20084 3282 20097 3328
rect 20143 3282 20172 3328
rect 20084 3204 20172 3282
rect 20292 3328 20380 3368
rect 20292 3282 20321 3328
rect 20367 3282 20380 3328
rect 20292 3204 20380 3282
rect 20532 3328 20620 3368
rect 20532 3282 20545 3328
rect 20591 3282 20620 3328
rect 20532 3204 20620 3282
rect 20820 3328 20908 3368
rect 20820 3282 20849 3328
rect 20895 3282 20908 3328
rect 20820 3204 20908 3282
rect 21204 3328 21292 3368
rect 21204 3282 21217 3328
rect 21263 3282 21292 3328
rect 21204 3204 21292 3282
rect 21492 3328 21580 3368
rect 21492 3282 21521 3328
rect 21567 3282 21580 3328
rect 21492 3204 21580 3282
rect 21652 3328 21740 3368
rect 21652 3282 21665 3328
rect 21711 3282 21740 3328
rect 21652 3204 21740 3282
rect 21940 3328 22028 3368
rect 21940 3282 21969 3328
rect 22015 3282 22028 3328
rect 21940 3204 22028 3282
<< mvpdiff >>
rect 1604 16337 1692 16396
rect 1604 16197 1617 16337
rect 1663 16197 1692 16337
rect 1604 16152 1692 16197
rect 1892 16337 1980 16396
rect 1892 16197 1921 16337
rect 1967 16197 1980 16337
rect 1892 16152 1980 16197
rect 2052 16337 2140 16396
rect 2052 16197 2065 16337
rect 2111 16197 2140 16337
rect 2052 16152 2140 16197
rect 2340 16337 2428 16396
rect 2340 16197 2369 16337
rect 2415 16197 2428 16337
rect 2340 16152 2428 16197
rect 2500 16337 2588 16396
rect 2500 16197 2513 16337
rect 2559 16197 2588 16337
rect 2500 16152 2588 16197
rect 2788 16337 2876 16396
rect 2788 16197 2817 16337
rect 2863 16197 2876 16337
rect 2788 16152 2876 16197
rect 2948 16337 3036 16396
rect 2948 16197 2961 16337
rect 3007 16197 3036 16337
rect 2948 16152 3036 16197
rect 3236 16337 3324 16396
rect 3236 16197 3265 16337
rect 3311 16197 3324 16337
rect 3236 16152 3324 16197
rect 3396 16337 3484 16396
rect 3396 16197 3409 16337
rect 3455 16197 3484 16337
rect 3396 16152 3484 16197
rect 3684 16337 3772 16396
rect 3684 16197 3713 16337
rect 3759 16197 3772 16337
rect 3684 16152 3772 16197
rect 3844 16337 3932 16396
rect 3844 16197 3857 16337
rect 3903 16197 3932 16337
rect 3844 16152 3932 16197
rect 4132 16337 4220 16396
rect 4132 16197 4161 16337
rect 4207 16197 4220 16337
rect 4132 16152 4220 16197
rect 4292 16337 4380 16396
rect 4292 16197 4305 16337
rect 4351 16197 4380 16337
rect 4292 16152 4380 16197
rect 4580 16337 4668 16396
rect 4580 16197 4609 16337
rect 4655 16197 4668 16337
rect 4580 16152 4668 16197
rect 4740 16337 4828 16396
rect 4740 16197 4753 16337
rect 4799 16197 4828 16337
rect 4740 16152 4828 16197
rect 5028 16337 5116 16396
rect 5028 16197 5057 16337
rect 5103 16197 5116 16337
rect 5028 16152 5116 16197
rect 5524 16337 5612 16396
rect 5524 16197 5537 16337
rect 5583 16197 5612 16337
rect 5524 16152 5612 16197
rect 5812 16337 5900 16396
rect 5812 16197 5841 16337
rect 5887 16197 5900 16337
rect 5812 16152 5900 16197
rect 5972 16337 6060 16396
rect 5972 16197 5985 16337
rect 6031 16197 6060 16337
rect 5972 16152 6060 16197
rect 6260 16337 6348 16396
rect 6260 16197 6289 16337
rect 6335 16197 6348 16337
rect 6260 16152 6348 16197
rect 6420 16337 6508 16396
rect 6420 16197 6433 16337
rect 6479 16197 6508 16337
rect 6420 16152 6508 16197
rect 6708 16337 6796 16396
rect 6708 16197 6737 16337
rect 6783 16197 6796 16337
rect 6708 16152 6796 16197
rect 6868 16337 6956 16396
rect 6868 16197 6881 16337
rect 6927 16197 6956 16337
rect 6868 16152 6956 16197
rect 7156 16337 7244 16396
rect 7156 16197 7185 16337
rect 7231 16197 7244 16337
rect 7156 16152 7244 16197
rect 7316 16337 7404 16396
rect 7316 16197 7329 16337
rect 7375 16197 7404 16337
rect 7316 16152 7404 16197
rect 7604 16337 7692 16396
rect 7604 16197 7633 16337
rect 7679 16197 7692 16337
rect 7604 16152 7692 16197
rect 7764 16337 7852 16396
rect 7764 16197 7777 16337
rect 7823 16197 7852 16337
rect 7764 16152 7852 16197
rect 8052 16337 8140 16396
rect 8052 16197 8081 16337
rect 8127 16197 8140 16337
rect 8052 16152 8140 16197
rect 8212 16337 8300 16396
rect 8212 16197 8225 16337
rect 8271 16197 8300 16337
rect 8212 16152 8300 16197
rect 8500 16337 8588 16396
rect 8500 16197 8529 16337
rect 8575 16197 8588 16337
rect 8500 16152 8588 16197
rect 8660 16337 8748 16396
rect 8660 16197 8673 16337
rect 8719 16197 8748 16337
rect 8660 16152 8748 16197
rect 8948 16337 9036 16396
rect 8948 16197 8977 16337
rect 9023 16197 9036 16337
rect 8948 16152 9036 16197
rect 9444 16337 9532 16396
rect 9444 16197 9457 16337
rect 9503 16197 9532 16337
rect 9444 16152 9532 16197
rect 9732 16337 9820 16396
rect 9732 16197 9761 16337
rect 9807 16197 9820 16337
rect 9732 16152 9820 16197
rect 9892 16337 9980 16396
rect 9892 16197 9905 16337
rect 9951 16197 9980 16337
rect 9892 16152 9980 16197
rect 10180 16337 10268 16396
rect 10180 16197 10209 16337
rect 10255 16197 10268 16337
rect 10180 16152 10268 16197
rect 10340 16337 10428 16396
rect 10340 16197 10353 16337
rect 10399 16197 10428 16337
rect 10340 16152 10428 16197
rect 10628 16337 10716 16396
rect 10628 16197 10657 16337
rect 10703 16197 10716 16337
rect 10628 16152 10716 16197
rect 10788 16337 10876 16396
rect 10788 16197 10801 16337
rect 10847 16197 10876 16337
rect 10788 16152 10876 16197
rect 11076 16337 11164 16396
rect 11076 16197 11105 16337
rect 11151 16197 11164 16337
rect 11076 16152 11164 16197
rect 11236 16337 11324 16396
rect 11236 16197 11249 16337
rect 11295 16197 11324 16337
rect 11236 16152 11324 16197
rect 11524 16337 11612 16396
rect 11524 16197 11553 16337
rect 11599 16197 11612 16337
rect 11524 16152 11612 16197
rect 11684 16337 11772 16396
rect 11684 16197 11697 16337
rect 11743 16197 11772 16337
rect 11684 16152 11772 16197
rect 11972 16337 12060 16396
rect 11972 16197 12001 16337
rect 12047 16197 12060 16337
rect 11972 16152 12060 16197
rect 12132 16337 12220 16396
rect 12132 16197 12145 16337
rect 12191 16197 12220 16337
rect 12132 16152 12220 16197
rect 12420 16337 12508 16396
rect 12420 16197 12449 16337
rect 12495 16197 12508 16337
rect 12420 16152 12508 16197
rect 12580 16337 12668 16396
rect 12580 16197 12593 16337
rect 12639 16197 12668 16337
rect 12580 16152 12668 16197
rect 12868 16337 12956 16396
rect 12868 16197 12897 16337
rect 12943 16197 12956 16337
rect 12868 16152 12956 16197
rect 13364 16337 13452 16396
rect 13364 16197 13377 16337
rect 13423 16197 13452 16337
rect 13364 16152 13452 16197
rect 13652 16337 13740 16396
rect 13652 16197 13681 16337
rect 13727 16197 13740 16337
rect 13652 16152 13740 16197
rect 13812 16337 13900 16396
rect 13812 16197 13825 16337
rect 13871 16197 13900 16337
rect 13812 16152 13900 16197
rect 14100 16337 14188 16396
rect 14100 16197 14129 16337
rect 14175 16197 14188 16337
rect 14100 16152 14188 16197
rect 14260 16337 14348 16396
rect 14260 16197 14273 16337
rect 14319 16197 14348 16337
rect 14260 16152 14348 16197
rect 14548 16337 14636 16396
rect 14548 16197 14577 16337
rect 14623 16197 14636 16337
rect 14548 16152 14636 16197
rect 14708 16337 14796 16396
rect 14708 16197 14721 16337
rect 14767 16197 14796 16337
rect 14708 16152 14796 16197
rect 14996 16337 15084 16396
rect 14996 16197 15025 16337
rect 15071 16197 15084 16337
rect 14996 16152 15084 16197
rect 15156 16337 15244 16396
rect 15156 16197 15169 16337
rect 15215 16197 15244 16337
rect 15156 16152 15244 16197
rect 15444 16337 15532 16396
rect 15444 16197 15473 16337
rect 15519 16197 15532 16337
rect 15444 16152 15532 16197
rect 15604 16337 15692 16396
rect 15604 16197 15617 16337
rect 15663 16197 15692 16337
rect 15604 16152 15692 16197
rect 15892 16337 15980 16396
rect 15892 16197 15921 16337
rect 15967 16197 15980 16337
rect 15892 16152 15980 16197
rect 16052 16337 16140 16396
rect 16052 16197 16065 16337
rect 16111 16197 16140 16337
rect 16052 16152 16140 16197
rect 16340 16337 16428 16396
rect 16340 16197 16369 16337
rect 16415 16197 16428 16337
rect 16340 16152 16428 16197
rect 16500 16337 16588 16396
rect 16500 16197 16513 16337
rect 16559 16197 16588 16337
rect 16500 16152 16588 16197
rect 16788 16337 16876 16396
rect 16788 16197 16817 16337
rect 16863 16197 16876 16337
rect 16788 16152 16876 16197
rect 17284 16337 17372 16396
rect 17284 16197 17297 16337
rect 17343 16197 17372 16337
rect 17284 16152 17372 16197
rect 17572 16337 17660 16396
rect 17572 16197 17601 16337
rect 17647 16197 17660 16337
rect 17572 16152 17660 16197
rect 17732 16337 17820 16396
rect 17732 16197 17745 16337
rect 17791 16197 17820 16337
rect 17732 16152 17820 16197
rect 18020 16337 18108 16396
rect 18020 16197 18049 16337
rect 18095 16197 18108 16337
rect 18020 16152 18108 16197
rect 18180 16337 18268 16396
rect 18180 16197 18193 16337
rect 18239 16197 18268 16337
rect 18180 16152 18268 16197
rect 18468 16337 18556 16396
rect 18468 16197 18497 16337
rect 18543 16197 18556 16337
rect 18468 16152 18556 16197
rect 18628 16337 18716 16396
rect 18628 16197 18641 16337
rect 18687 16197 18716 16337
rect 18628 16152 18716 16197
rect 18916 16337 19004 16396
rect 18916 16197 18945 16337
rect 18991 16197 19004 16337
rect 18916 16152 19004 16197
rect 19076 16337 19164 16396
rect 19076 16197 19089 16337
rect 19135 16197 19164 16337
rect 19076 16152 19164 16197
rect 19364 16337 19452 16396
rect 19364 16197 19393 16337
rect 19439 16197 19452 16337
rect 19364 16152 19452 16197
rect 19524 16337 19612 16396
rect 19524 16197 19537 16337
rect 19583 16197 19612 16337
rect 19524 16152 19612 16197
rect 19812 16337 19900 16396
rect 19812 16197 19841 16337
rect 19887 16197 19900 16337
rect 19812 16152 19900 16197
rect 19972 16337 20060 16396
rect 19972 16197 19985 16337
rect 20031 16197 20060 16337
rect 19972 16152 20060 16197
rect 20260 16337 20348 16396
rect 20260 16197 20289 16337
rect 20335 16197 20348 16337
rect 20260 16152 20348 16197
rect 20420 16337 20508 16396
rect 20420 16197 20433 16337
rect 20479 16197 20508 16337
rect 20420 16152 20508 16197
rect 20708 16337 20796 16396
rect 20708 16197 20737 16337
rect 20783 16197 20796 16337
rect 20708 16152 20796 16197
rect 21204 16337 21292 16396
rect 21204 16197 21217 16337
rect 21263 16197 21292 16337
rect 21204 16152 21292 16197
rect 21492 16337 21580 16396
rect 21492 16197 21521 16337
rect 21567 16197 21580 16337
rect 21492 16152 21580 16197
rect 21652 16337 21740 16396
rect 21652 16197 21665 16337
rect 21711 16197 21740 16337
rect 21652 16152 21740 16197
rect 21940 16337 22028 16396
rect 21940 16197 21969 16337
rect 22015 16197 22028 16337
rect 21940 16152 22028 16197
rect 1604 15163 1692 15208
rect 1604 15023 1617 15163
rect 1663 15023 1692 15163
rect 1604 14964 1692 15023
rect 1892 15163 1980 15208
rect 1892 15023 1921 15163
rect 1967 15023 1980 15163
rect 1892 14964 1980 15023
rect 2052 15163 2140 15208
rect 2052 15023 2065 15163
rect 2111 15023 2140 15163
rect 2052 14964 2140 15023
rect 2340 15163 2428 15208
rect 2340 15023 2369 15163
rect 2415 15023 2428 15163
rect 2340 14964 2428 15023
rect 2500 15163 2588 15208
rect 2500 15023 2513 15163
rect 2559 15023 2588 15163
rect 2500 14964 2588 15023
rect 2788 15163 2876 15208
rect 2788 15023 2817 15163
rect 2863 15023 2876 15163
rect 2788 14964 2876 15023
rect 2948 15163 3036 15208
rect 2948 15023 2961 15163
rect 3007 15023 3036 15163
rect 2948 14964 3036 15023
rect 3236 15163 3324 15208
rect 3236 15023 3265 15163
rect 3311 15023 3324 15163
rect 3236 14964 3324 15023
rect 3396 15163 3484 15208
rect 3396 15023 3409 15163
rect 3455 15023 3484 15163
rect 3396 14964 3484 15023
rect 3684 15163 3772 15208
rect 3684 15023 3713 15163
rect 3759 15023 3772 15163
rect 3684 14964 3772 15023
rect 3844 15163 3932 15208
rect 3844 15023 3857 15163
rect 3903 15023 3932 15163
rect 3844 14964 3932 15023
rect 4132 15163 4220 15208
rect 4132 15023 4161 15163
rect 4207 15023 4220 15163
rect 4132 14964 4220 15023
rect 4292 15163 4380 15208
rect 4292 15023 4305 15163
rect 4351 15023 4380 15163
rect 4292 14964 4380 15023
rect 4580 15163 4668 15208
rect 4580 15023 4609 15163
rect 4655 15023 4668 15163
rect 4580 14964 4668 15023
rect 4740 15163 4828 15208
rect 4740 15023 4753 15163
rect 4799 15023 4828 15163
rect 4740 14964 4828 15023
rect 5028 15163 5116 15208
rect 5028 15023 5057 15163
rect 5103 15023 5116 15163
rect 5028 14964 5116 15023
rect 5188 15163 5276 15208
rect 5188 15023 5201 15163
rect 5247 15023 5276 15163
rect 5188 14964 5276 15023
rect 5476 15163 5564 15208
rect 5476 15023 5505 15163
rect 5551 15023 5564 15163
rect 5476 14964 5564 15023
rect 5636 15163 5724 15208
rect 5636 15023 5649 15163
rect 5695 15023 5724 15163
rect 5636 14964 5724 15023
rect 5924 15163 6012 15208
rect 5924 15023 5953 15163
rect 5999 15023 6012 15163
rect 5924 14964 6012 15023
rect 6084 15163 6172 15208
rect 6084 15023 6097 15163
rect 6143 15023 6172 15163
rect 6084 14964 6172 15023
rect 6372 15163 6460 15208
rect 6372 15023 6401 15163
rect 6447 15023 6460 15163
rect 6372 14964 6460 15023
rect 6532 15163 6620 15208
rect 6532 15023 6545 15163
rect 6591 15023 6620 15163
rect 6532 14964 6620 15023
rect 6820 15163 6908 15208
rect 6820 15023 6849 15163
rect 6895 15023 6908 15163
rect 6820 14964 6908 15023
rect 6980 15163 7068 15208
rect 6980 15023 6993 15163
rect 7039 15023 7068 15163
rect 6980 14964 7068 15023
rect 7268 15163 7356 15208
rect 7268 15023 7297 15163
rect 7343 15023 7356 15163
rect 7268 14964 7356 15023
rect 7428 15163 7516 15208
rect 7428 15023 7441 15163
rect 7487 15023 7516 15163
rect 7428 14964 7516 15023
rect 7716 15163 7804 15208
rect 7716 15023 7745 15163
rect 7791 15023 7804 15163
rect 7716 14964 7804 15023
rect 7876 15163 7964 15208
rect 7876 15023 7889 15163
rect 7935 15023 7964 15163
rect 7876 14964 7964 15023
rect 8164 15163 8252 15208
rect 8164 15023 8193 15163
rect 8239 15023 8252 15163
rect 8164 14964 8252 15023
rect 8324 15163 8412 15208
rect 8324 15023 8337 15163
rect 8383 15023 8412 15163
rect 8324 14964 8412 15023
rect 8612 15163 8700 15208
rect 8612 15023 8641 15163
rect 8687 15023 8700 15163
rect 8612 14964 8700 15023
rect 8772 15163 8860 15208
rect 8772 15023 8785 15163
rect 8831 15023 8860 15163
rect 8772 14964 8860 15023
rect 9060 15163 9148 15208
rect 9060 15023 9089 15163
rect 9135 15023 9148 15163
rect 9060 14964 9148 15023
rect 9556 15163 9644 15208
rect 9556 15023 9569 15163
rect 9615 15023 9644 15163
rect 9556 14964 9644 15023
rect 9844 15163 9932 15208
rect 9844 15023 9873 15163
rect 9919 15023 9932 15163
rect 9844 14964 9932 15023
rect 10004 15163 10092 15208
rect 10004 15023 10017 15163
rect 10063 15023 10092 15163
rect 10004 14964 10092 15023
rect 10292 15163 10380 15208
rect 10292 15023 10321 15163
rect 10367 15023 10380 15163
rect 10292 14964 10380 15023
rect 10452 15163 10540 15208
rect 10452 15023 10465 15163
rect 10511 15023 10540 15163
rect 10452 14964 10540 15023
rect 10740 15163 10828 15208
rect 10740 15023 10769 15163
rect 10815 15023 10828 15163
rect 10740 14964 10828 15023
rect 10900 15163 10988 15208
rect 10900 15023 10913 15163
rect 10959 15023 10988 15163
rect 10900 14964 10988 15023
rect 11188 15163 11276 15208
rect 11188 15023 11217 15163
rect 11263 15023 11276 15163
rect 11188 14964 11276 15023
rect 11348 15163 11436 15208
rect 11348 15023 11361 15163
rect 11407 15023 11436 15163
rect 11348 14964 11436 15023
rect 11636 15163 11724 15208
rect 11636 15023 11665 15163
rect 11711 15023 11724 15163
rect 11636 14964 11724 15023
rect 11796 15163 11884 15208
rect 11796 15023 11809 15163
rect 11855 15023 11884 15163
rect 11796 14964 11884 15023
rect 12084 15163 12172 15208
rect 12084 15023 12113 15163
rect 12159 15023 12172 15163
rect 12084 14964 12172 15023
rect 12244 15163 12332 15208
rect 12244 15023 12257 15163
rect 12303 15023 12332 15163
rect 12244 14964 12332 15023
rect 12532 15163 12620 15208
rect 12532 15023 12561 15163
rect 12607 15023 12620 15163
rect 12532 14964 12620 15023
rect 12692 15163 12780 15208
rect 12692 15023 12705 15163
rect 12751 15023 12780 15163
rect 12692 14964 12780 15023
rect 12980 15163 13068 15208
rect 12980 15023 13009 15163
rect 13055 15023 13068 15163
rect 12980 14964 13068 15023
rect 13140 15163 13228 15208
rect 13140 15023 13153 15163
rect 13199 15023 13228 15163
rect 13140 14964 13228 15023
rect 13428 15163 13516 15208
rect 13428 15023 13457 15163
rect 13503 15023 13516 15163
rect 13428 14964 13516 15023
rect 13588 15163 13676 15208
rect 13588 15023 13601 15163
rect 13647 15023 13676 15163
rect 13588 14964 13676 15023
rect 13876 15163 13964 15208
rect 13876 15023 13905 15163
rect 13951 15023 13964 15163
rect 13876 14964 13964 15023
rect 14036 15163 14124 15208
rect 14036 15023 14049 15163
rect 14095 15023 14124 15163
rect 14036 14964 14124 15023
rect 14324 15163 14412 15208
rect 14324 15023 14353 15163
rect 14399 15023 14412 15163
rect 14324 14964 14412 15023
rect 14484 15163 14572 15208
rect 14484 15023 14497 15163
rect 14543 15023 14572 15163
rect 14484 14964 14572 15023
rect 14772 15163 14860 15208
rect 14772 15023 14801 15163
rect 14847 15023 14860 15163
rect 14772 14964 14860 15023
rect 14932 15163 15020 15208
rect 14932 15023 14945 15163
rect 14991 15023 15020 15163
rect 14932 14964 15020 15023
rect 15220 15163 15308 15208
rect 15220 15023 15249 15163
rect 15295 15023 15308 15163
rect 15220 14964 15308 15023
rect 15380 15163 15468 15208
rect 15380 15023 15393 15163
rect 15439 15023 15468 15163
rect 15380 14964 15468 15023
rect 15668 15163 15756 15208
rect 15668 15023 15697 15163
rect 15743 15023 15756 15163
rect 15668 14964 15756 15023
rect 15828 15163 15916 15208
rect 15828 15023 15841 15163
rect 15887 15023 15916 15163
rect 15828 14964 15916 15023
rect 16116 15163 16204 15208
rect 16116 15023 16145 15163
rect 16191 15023 16204 15163
rect 16116 14964 16204 15023
rect 16276 15163 16364 15208
rect 16276 15023 16289 15163
rect 16335 15023 16364 15163
rect 16276 14964 16364 15023
rect 16564 15163 16652 15208
rect 16564 15023 16593 15163
rect 16639 15023 16652 15163
rect 16564 14964 16652 15023
rect 16724 15163 16812 15208
rect 16724 15023 16737 15163
rect 16783 15023 16812 15163
rect 16724 14964 16812 15023
rect 17012 15163 17100 15208
rect 17012 15023 17041 15163
rect 17087 15023 17100 15163
rect 17012 14964 17100 15023
rect 17508 15163 17596 15208
rect 17508 15023 17521 15163
rect 17567 15023 17596 15163
rect 17508 14964 17596 15023
rect 17796 15163 17884 15208
rect 17796 15023 17825 15163
rect 17871 15023 17884 15163
rect 17796 14964 17884 15023
rect 17956 15163 18044 15208
rect 17956 15023 17969 15163
rect 18015 15023 18044 15163
rect 17956 14964 18044 15023
rect 18244 15163 18332 15208
rect 18244 15023 18273 15163
rect 18319 15023 18332 15163
rect 18244 14964 18332 15023
rect 18404 15163 18492 15208
rect 18404 15023 18417 15163
rect 18463 15023 18492 15163
rect 18404 14964 18492 15023
rect 18692 15163 18780 15208
rect 18692 15023 18721 15163
rect 18767 15023 18780 15163
rect 18692 14964 18780 15023
rect 18852 15163 18940 15208
rect 18852 15023 18865 15163
rect 18911 15023 18940 15163
rect 18852 14964 18940 15023
rect 19140 15163 19228 15208
rect 19140 15023 19169 15163
rect 19215 15023 19228 15163
rect 19140 14964 19228 15023
rect 19300 15163 19388 15208
rect 19300 15023 19313 15163
rect 19359 15023 19388 15163
rect 19300 14964 19388 15023
rect 19588 15163 19676 15208
rect 19588 15023 19617 15163
rect 19663 15023 19676 15163
rect 19588 14964 19676 15023
rect 19748 15163 19836 15208
rect 19748 15023 19761 15163
rect 19807 15023 19836 15163
rect 19748 14964 19836 15023
rect 20036 15163 20124 15208
rect 20036 15023 20065 15163
rect 20111 15023 20124 15163
rect 20036 14964 20124 15023
rect 20196 15163 20284 15208
rect 20196 15023 20209 15163
rect 20255 15023 20284 15163
rect 20196 14964 20284 15023
rect 20484 15163 20572 15208
rect 20484 15023 20513 15163
rect 20559 15023 20572 15163
rect 20484 14964 20572 15023
rect 20644 15163 20732 15208
rect 20644 15023 20657 15163
rect 20703 15023 20732 15163
rect 20644 14964 20732 15023
rect 20932 15163 21020 15208
rect 20932 15023 20961 15163
rect 21007 15023 21020 15163
rect 20932 14964 21020 15023
rect 21092 15163 21180 15208
rect 21092 15023 21105 15163
rect 21151 15023 21180 15163
rect 21092 14964 21180 15023
rect 21380 15163 21468 15208
rect 21380 15023 21409 15163
rect 21455 15023 21468 15163
rect 21380 14964 21468 15023
rect 21540 15163 21628 15208
rect 21540 15023 21553 15163
rect 21599 15023 21628 15163
rect 21540 14964 21628 15023
rect 21828 15163 21916 15208
rect 21828 15023 21857 15163
rect 21903 15023 21916 15163
rect 21828 14964 21916 15023
rect 21988 15163 22076 15208
rect 21988 15023 22001 15163
rect 22047 15023 22076 15163
rect 21988 14964 22076 15023
rect 22276 15163 22364 15208
rect 22276 15023 22305 15163
rect 22351 15023 22364 15163
rect 22276 14964 22364 15023
rect 1604 14769 1692 14828
rect 1604 14629 1617 14769
rect 1663 14629 1692 14769
rect 1604 14584 1692 14629
rect 1892 14769 1980 14828
rect 1892 14629 1921 14769
rect 1967 14629 1980 14769
rect 1892 14584 1980 14629
rect 2052 14769 2140 14828
rect 2052 14629 2065 14769
rect 2111 14629 2140 14769
rect 2052 14584 2140 14629
rect 2340 14769 2428 14828
rect 2340 14629 2369 14769
rect 2415 14629 2428 14769
rect 2340 14584 2428 14629
rect 2500 14769 2588 14828
rect 2500 14629 2513 14769
rect 2559 14629 2588 14769
rect 2500 14584 2588 14629
rect 2788 14769 2876 14828
rect 2788 14629 2817 14769
rect 2863 14629 2876 14769
rect 2788 14584 2876 14629
rect 2948 14769 3036 14828
rect 2948 14629 2961 14769
rect 3007 14629 3036 14769
rect 2948 14584 3036 14629
rect 3236 14769 3324 14828
rect 3236 14629 3265 14769
rect 3311 14629 3324 14769
rect 3236 14584 3324 14629
rect 3396 14769 3484 14828
rect 3396 14629 3409 14769
rect 3455 14629 3484 14769
rect 3396 14584 3484 14629
rect 3684 14769 3772 14828
rect 3684 14629 3713 14769
rect 3759 14629 3772 14769
rect 3684 14584 3772 14629
rect 3844 14769 3932 14828
rect 3844 14629 3857 14769
rect 3903 14629 3932 14769
rect 3844 14584 3932 14629
rect 4132 14769 4220 14828
rect 4132 14629 4161 14769
rect 4207 14629 4220 14769
rect 4132 14584 4220 14629
rect 4292 14769 4380 14828
rect 4292 14629 4305 14769
rect 4351 14629 4380 14769
rect 4292 14584 4380 14629
rect 4580 14769 4668 14828
rect 4580 14629 4609 14769
rect 4655 14629 4668 14769
rect 4580 14584 4668 14629
rect 4740 14769 4828 14828
rect 4740 14629 4753 14769
rect 4799 14629 4828 14769
rect 4740 14584 4828 14629
rect 5028 14769 5116 14828
rect 5028 14629 5057 14769
rect 5103 14629 5116 14769
rect 5028 14584 5116 14629
rect 5524 14769 5612 14828
rect 5524 14629 5537 14769
rect 5583 14629 5612 14769
rect 5524 14584 5612 14629
rect 5812 14769 5900 14828
rect 5812 14629 5841 14769
rect 5887 14629 5900 14769
rect 5812 14584 5900 14629
rect 5972 14769 6060 14828
rect 5972 14629 5985 14769
rect 6031 14629 6060 14769
rect 5972 14584 6060 14629
rect 6260 14769 6348 14828
rect 6260 14629 6289 14769
rect 6335 14629 6348 14769
rect 6260 14584 6348 14629
rect 6420 14769 6508 14828
rect 6420 14629 6433 14769
rect 6479 14629 6508 14769
rect 6420 14584 6508 14629
rect 6708 14769 6796 14828
rect 6708 14629 6737 14769
rect 6783 14629 6796 14769
rect 6708 14584 6796 14629
rect 6868 14769 6956 14828
rect 6868 14629 6881 14769
rect 6927 14629 6956 14769
rect 6868 14584 6956 14629
rect 7156 14769 7244 14828
rect 7156 14629 7185 14769
rect 7231 14629 7244 14769
rect 7156 14584 7244 14629
rect 7316 14769 7404 14828
rect 7316 14629 7329 14769
rect 7375 14629 7404 14769
rect 7316 14584 7404 14629
rect 7604 14769 7692 14828
rect 7604 14629 7633 14769
rect 7679 14629 7692 14769
rect 7604 14584 7692 14629
rect 7764 14769 7852 14828
rect 7764 14629 7777 14769
rect 7823 14629 7852 14769
rect 7764 14584 7852 14629
rect 8052 14769 8140 14828
rect 8052 14629 8081 14769
rect 8127 14629 8140 14769
rect 8052 14584 8140 14629
rect 8212 14769 8300 14828
rect 8212 14629 8225 14769
rect 8271 14629 8300 14769
rect 8212 14584 8300 14629
rect 8500 14769 8588 14828
rect 8500 14629 8529 14769
rect 8575 14629 8588 14769
rect 8500 14584 8588 14629
rect 8660 14769 8748 14828
rect 8660 14629 8673 14769
rect 8719 14629 8748 14769
rect 8660 14584 8748 14629
rect 8948 14769 9036 14828
rect 8948 14629 8977 14769
rect 9023 14629 9036 14769
rect 8948 14584 9036 14629
rect 9108 14769 9196 14828
rect 9108 14629 9121 14769
rect 9167 14629 9196 14769
rect 9108 14584 9196 14629
rect 9396 14769 9484 14828
rect 9396 14629 9425 14769
rect 9471 14629 9484 14769
rect 9396 14584 9484 14629
rect 9556 14769 9644 14828
rect 9556 14629 9569 14769
rect 9615 14629 9644 14769
rect 9556 14584 9644 14629
rect 9844 14769 9932 14828
rect 9844 14629 9873 14769
rect 9919 14629 9932 14769
rect 9844 14584 9932 14629
rect 10004 14769 10092 14828
rect 10004 14629 10017 14769
rect 10063 14629 10092 14769
rect 10004 14584 10092 14629
rect 10292 14769 10380 14828
rect 10292 14629 10321 14769
rect 10367 14629 10380 14769
rect 10292 14584 10380 14629
rect 10452 14769 10540 14828
rect 10452 14629 10465 14769
rect 10511 14629 10540 14769
rect 10452 14584 10540 14629
rect 10740 14769 10828 14828
rect 10740 14629 10769 14769
rect 10815 14629 10828 14769
rect 10740 14584 10828 14629
rect 10900 14769 10988 14828
rect 10900 14629 10913 14769
rect 10959 14629 10988 14769
rect 10900 14584 10988 14629
rect 11188 14769 11276 14828
rect 11188 14629 11217 14769
rect 11263 14629 11276 14769
rect 11188 14584 11276 14629
rect 11348 14769 11436 14828
rect 11348 14629 11361 14769
rect 11407 14629 11436 14769
rect 11348 14584 11436 14629
rect 11636 14769 11724 14828
rect 11636 14629 11665 14769
rect 11711 14629 11724 14769
rect 11636 14584 11724 14629
rect 11796 14769 11884 14828
rect 11796 14629 11809 14769
rect 11855 14629 11884 14769
rect 11796 14584 11884 14629
rect 12084 14769 12172 14828
rect 12084 14629 12113 14769
rect 12159 14629 12172 14769
rect 12084 14584 12172 14629
rect 12244 14769 12332 14828
rect 12244 14629 12257 14769
rect 12303 14629 12332 14769
rect 12244 14584 12332 14629
rect 12532 14769 12620 14828
rect 12532 14629 12561 14769
rect 12607 14629 12620 14769
rect 12532 14584 12620 14629
rect 12692 14769 12780 14828
rect 12692 14629 12705 14769
rect 12751 14629 12780 14769
rect 12692 14584 12780 14629
rect 12980 14769 13068 14828
rect 12980 14629 13009 14769
rect 13055 14629 13068 14769
rect 12980 14584 13068 14629
rect 13476 14769 13564 14828
rect 13476 14629 13489 14769
rect 13535 14629 13564 14769
rect 13476 14584 13564 14629
rect 13764 14769 13852 14828
rect 13764 14629 13793 14769
rect 13839 14629 13852 14769
rect 13764 14584 13852 14629
rect 13924 14769 14012 14828
rect 13924 14629 13937 14769
rect 13983 14629 14012 14769
rect 13924 14584 14012 14629
rect 14212 14769 14300 14828
rect 14212 14629 14241 14769
rect 14287 14629 14300 14769
rect 14212 14584 14300 14629
rect 14372 14769 14460 14828
rect 14372 14629 14385 14769
rect 14431 14629 14460 14769
rect 14372 14584 14460 14629
rect 14660 14769 14748 14828
rect 14660 14629 14689 14769
rect 14735 14629 14748 14769
rect 14660 14584 14748 14629
rect 14820 14769 14908 14828
rect 14820 14629 14833 14769
rect 14879 14629 14908 14769
rect 14820 14584 14908 14629
rect 15108 14769 15196 14828
rect 15108 14629 15137 14769
rect 15183 14629 15196 14769
rect 15108 14584 15196 14629
rect 15268 14769 15356 14828
rect 15268 14629 15281 14769
rect 15327 14629 15356 14769
rect 15268 14584 15356 14629
rect 15556 14769 15644 14828
rect 15556 14629 15585 14769
rect 15631 14629 15644 14769
rect 15556 14584 15644 14629
rect 15716 14769 15804 14828
rect 15716 14629 15729 14769
rect 15775 14629 15804 14769
rect 15716 14584 15804 14629
rect 16004 14769 16092 14828
rect 16004 14629 16033 14769
rect 16079 14629 16092 14769
rect 16004 14584 16092 14629
rect 16164 14769 16252 14828
rect 16164 14629 16177 14769
rect 16223 14629 16252 14769
rect 16164 14584 16252 14629
rect 16452 14769 16540 14828
rect 16452 14629 16481 14769
rect 16527 14629 16540 14769
rect 16452 14584 16540 14629
rect 16804 14777 16892 14828
rect 16804 14637 16817 14777
rect 16863 14637 16892 14777
rect 16804 14584 16892 14637
rect 16992 14777 17080 14828
rect 16992 14637 17021 14777
rect 17067 14637 17080 14777
rect 16992 14584 17080 14637
rect 17476 14777 17564 14828
rect 17476 14637 17489 14777
rect 17535 14637 17564 14777
rect 17476 14584 17564 14637
rect 17664 14777 17752 14828
rect 17664 14637 17693 14777
rect 17739 14637 17752 14777
rect 17664 14584 17752 14637
rect 17844 14769 17932 14828
rect 17844 14629 17857 14769
rect 17903 14629 17932 14769
rect 17844 14584 17932 14629
rect 18132 14769 18220 14828
rect 18132 14629 18161 14769
rect 18207 14629 18220 14769
rect 18132 14584 18220 14629
rect 18292 14769 18380 14828
rect 18292 14629 18305 14769
rect 18351 14629 18380 14769
rect 18292 14584 18380 14629
rect 18580 14769 18668 14828
rect 18580 14629 18609 14769
rect 18655 14629 18668 14769
rect 18580 14584 18668 14629
rect 18740 14769 18828 14828
rect 18740 14629 18753 14769
rect 18799 14629 18828 14769
rect 18740 14584 18828 14629
rect 19028 14769 19116 14828
rect 19028 14629 19057 14769
rect 19103 14629 19116 14769
rect 19028 14584 19116 14629
rect 19188 14769 19276 14828
rect 19188 14629 19201 14769
rect 19247 14629 19276 14769
rect 19188 14584 19276 14629
rect 19476 14769 19564 14828
rect 19476 14629 19505 14769
rect 19551 14629 19564 14769
rect 19476 14584 19564 14629
rect 19636 14769 19724 14828
rect 19636 14629 19649 14769
rect 19695 14629 19724 14769
rect 19636 14584 19724 14629
rect 19924 14769 20012 14828
rect 19924 14629 19953 14769
rect 19999 14629 20012 14769
rect 19924 14584 20012 14629
rect 20084 14769 20172 14828
rect 20084 14629 20097 14769
rect 20143 14629 20172 14769
rect 20084 14584 20172 14629
rect 20372 14769 20460 14828
rect 20372 14629 20401 14769
rect 20447 14629 20460 14769
rect 20372 14584 20460 14629
rect 20532 14769 20620 14828
rect 20532 14629 20545 14769
rect 20591 14629 20620 14769
rect 20532 14584 20620 14629
rect 20820 14769 20908 14828
rect 20820 14629 20849 14769
rect 20895 14629 20908 14769
rect 20820 14584 20908 14629
rect 21428 14769 21516 14828
rect 21428 14629 21441 14769
rect 21487 14629 21516 14769
rect 21428 14584 21516 14629
rect 21716 14769 21804 14828
rect 21716 14629 21745 14769
rect 21791 14629 21804 14769
rect 21716 14584 21804 14629
rect 21876 14769 21964 14828
rect 21876 14629 21889 14769
rect 21935 14629 21964 14769
rect 21876 14584 21964 14629
rect 22164 14769 22252 14828
rect 22164 14629 22193 14769
rect 22239 14629 22252 14769
rect 22164 14584 22252 14629
rect 1604 13595 1692 13640
rect 1604 13455 1617 13595
rect 1663 13455 1692 13595
rect 1604 13396 1692 13455
rect 1892 13595 1980 13640
rect 1892 13455 1921 13595
rect 1967 13455 1980 13595
rect 1892 13396 1980 13455
rect 2052 13595 2140 13640
rect 2052 13455 2065 13595
rect 2111 13455 2140 13595
rect 2052 13396 2140 13455
rect 2340 13595 2428 13640
rect 2340 13455 2369 13595
rect 2415 13455 2428 13595
rect 2340 13396 2428 13455
rect 2500 13595 2588 13640
rect 2500 13455 2513 13595
rect 2559 13455 2588 13595
rect 2500 13396 2588 13455
rect 2788 13595 2876 13640
rect 2788 13455 2817 13595
rect 2863 13455 2876 13595
rect 2788 13396 2876 13455
rect 2948 13595 3036 13640
rect 2948 13455 2961 13595
rect 3007 13455 3036 13595
rect 2948 13396 3036 13455
rect 3236 13595 3324 13640
rect 3236 13455 3265 13595
rect 3311 13455 3324 13595
rect 3236 13396 3324 13455
rect 3396 13595 3484 13640
rect 3396 13455 3409 13595
rect 3455 13455 3484 13595
rect 3396 13396 3484 13455
rect 3684 13595 3772 13640
rect 3684 13455 3713 13595
rect 3759 13455 3772 13595
rect 3684 13396 3772 13455
rect 3844 13595 3932 13640
rect 3844 13455 3857 13595
rect 3903 13455 3932 13595
rect 3844 13396 3932 13455
rect 4132 13595 4220 13640
rect 4132 13455 4161 13595
rect 4207 13455 4220 13595
rect 4132 13396 4220 13455
rect 4292 13595 4380 13640
rect 4292 13455 4305 13595
rect 4351 13455 4380 13595
rect 4292 13396 4380 13455
rect 4580 13595 4668 13640
rect 4580 13455 4609 13595
rect 4655 13455 4668 13595
rect 4580 13396 4668 13455
rect 4740 13595 4828 13640
rect 4740 13455 4753 13595
rect 4799 13455 4828 13595
rect 4740 13396 4828 13455
rect 5028 13595 5116 13640
rect 5028 13455 5057 13595
rect 5103 13455 5116 13595
rect 5028 13396 5116 13455
rect 5188 13595 5276 13640
rect 5188 13455 5201 13595
rect 5247 13455 5276 13595
rect 5188 13396 5276 13455
rect 5476 13595 5564 13640
rect 5476 13455 5505 13595
rect 5551 13455 5564 13595
rect 5476 13396 5564 13455
rect 5636 13595 5724 13640
rect 5636 13455 5649 13595
rect 5695 13455 5724 13595
rect 5636 13396 5724 13455
rect 5924 13595 6012 13640
rect 5924 13455 5953 13595
rect 5999 13455 6012 13595
rect 5924 13396 6012 13455
rect 6084 13595 6172 13640
rect 6084 13455 6097 13595
rect 6143 13455 6172 13595
rect 6084 13396 6172 13455
rect 6372 13595 6460 13640
rect 6372 13455 6401 13595
rect 6447 13455 6460 13595
rect 6372 13396 6460 13455
rect 6532 13595 6620 13640
rect 6532 13455 6545 13595
rect 6591 13455 6620 13595
rect 6532 13396 6620 13455
rect 6820 13595 6908 13640
rect 6820 13455 6849 13595
rect 6895 13455 6908 13595
rect 6820 13396 6908 13455
rect 6980 13595 7068 13640
rect 6980 13455 6993 13595
rect 7039 13455 7068 13595
rect 6980 13396 7068 13455
rect 7268 13595 7356 13640
rect 7268 13455 7297 13595
rect 7343 13455 7356 13595
rect 7268 13396 7356 13455
rect 7428 13595 7516 13640
rect 7428 13455 7441 13595
rect 7487 13455 7516 13595
rect 7428 13396 7516 13455
rect 7716 13595 7804 13640
rect 7716 13455 7745 13595
rect 7791 13455 7804 13595
rect 7716 13396 7804 13455
rect 7876 13595 7964 13640
rect 7876 13455 7889 13595
rect 7935 13455 7964 13595
rect 7876 13396 7964 13455
rect 8164 13595 8252 13640
rect 8164 13455 8193 13595
rect 8239 13455 8252 13595
rect 8164 13396 8252 13455
rect 8324 13595 8412 13640
rect 8324 13455 8337 13595
rect 8383 13455 8412 13595
rect 8324 13396 8412 13455
rect 8612 13595 8700 13640
rect 8612 13455 8641 13595
rect 8687 13455 8700 13595
rect 8612 13396 8700 13455
rect 8772 13595 8860 13640
rect 8772 13455 8785 13595
rect 8831 13455 8860 13595
rect 8772 13396 8860 13455
rect 9060 13595 9148 13640
rect 9060 13455 9089 13595
rect 9135 13455 9148 13595
rect 9060 13396 9148 13455
rect 9556 13595 9644 13640
rect 9556 13455 9569 13595
rect 9615 13455 9644 13595
rect 9556 13396 9644 13455
rect 9844 13595 9932 13640
rect 9844 13455 9873 13595
rect 9919 13455 9932 13595
rect 9844 13396 9932 13455
rect 10004 13595 10092 13640
rect 10004 13455 10017 13595
rect 10063 13455 10092 13595
rect 10004 13396 10092 13455
rect 10292 13595 10380 13640
rect 10292 13455 10321 13595
rect 10367 13455 10380 13595
rect 10292 13396 10380 13455
rect 10452 13595 10540 13640
rect 10452 13455 10465 13595
rect 10511 13455 10540 13595
rect 10452 13396 10540 13455
rect 10740 13595 10828 13640
rect 10740 13455 10769 13595
rect 10815 13455 10828 13595
rect 10740 13396 10828 13455
rect 10900 13595 10988 13640
rect 10900 13455 10913 13595
rect 10959 13455 10988 13595
rect 10900 13396 10988 13455
rect 11188 13595 11276 13640
rect 11188 13455 11217 13595
rect 11263 13455 11276 13595
rect 11188 13396 11276 13455
rect 11348 13595 11436 13640
rect 11348 13455 11361 13595
rect 11407 13455 11436 13595
rect 11348 13396 11436 13455
rect 11636 13595 11724 13640
rect 11636 13455 11665 13595
rect 11711 13455 11724 13595
rect 11636 13396 11724 13455
rect 11796 13595 11884 13640
rect 11796 13455 11809 13595
rect 11855 13455 11884 13595
rect 11796 13396 11884 13455
rect 12084 13595 12172 13640
rect 12084 13455 12113 13595
rect 12159 13455 12172 13595
rect 12084 13396 12172 13455
rect 12244 13595 12332 13640
rect 12244 13455 12257 13595
rect 12303 13455 12332 13595
rect 12244 13396 12332 13455
rect 12532 13595 12620 13640
rect 12532 13455 12561 13595
rect 12607 13455 12620 13595
rect 12532 13396 12620 13455
rect 12692 13595 12780 13640
rect 12692 13455 12705 13595
rect 12751 13455 12780 13595
rect 12692 13396 12780 13455
rect 12980 13595 13068 13640
rect 12980 13455 13009 13595
rect 13055 13455 13068 13595
rect 12980 13396 13068 13455
rect 13140 13595 13228 13640
rect 13140 13455 13153 13595
rect 13199 13455 13228 13595
rect 13140 13396 13228 13455
rect 13428 13595 13516 13640
rect 13428 13455 13457 13595
rect 13503 13455 13516 13595
rect 13428 13396 13516 13455
rect 13588 13595 13676 13640
rect 13588 13455 13601 13595
rect 13647 13455 13676 13595
rect 13588 13396 13676 13455
rect 13876 13595 13964 13640
rect 13876 13455 13905 13595
rect 13951 13455 13964 13595
rect 13876 13396 13964 13455
rect 14036 13595 14124 13640
rect 14036 13455 14049 13595
rect 14095 13455 14124 13595
rect 14036 13396 14124 13455
rect 14324 13595 14412 13640
rect 14324 13455 14353 13595
rect 14399 13455 14412 13595
rect 14324 13396 14412 13455
rect 14484 13595 14572 13640
rect 14484 13455 14497 13595
rect 14543 13455 14572 13595
rect 14484 13396 14572 13455
rect 14772 13595 14860 13640
rect 14772 13455 14801 13595
rect 14847 13455 14860 13595
rect 14772 13396 14860 13455
rect 14932 13595 15020 13640
rect 14932 13455 14945 13595
rect 14991 13455 15020 13595
rect 14932 13396 15020 13455
rect 15220 13595 15308 13640
rect 15220 13455 15249 13595
rect 15295 13455 15308 13595
rect 15220 13396 15308 13455
rect 15380 13595 15468 13640
rect 15380 13455 15393 13595
rect 15439 13455 15468 13595
rect 15380 13396 15468 13455
rect 15668 13595 15756 13640
rect 15668 13455 15697 13595
rect 15743 13455 15756 13595
rect 15668 13396 15756 13455
rect 16072 13587 16160 13640
rect 16072 13447 16085 13587
rect 16131 13447 16160 13587
rect 16072 13396 16160 13447
rect 16260 13587 16348 13640
rect 16260 13447 16289 13587
rect 16335 13447 16348 13587
rect 16260 13396 16348 13447
rect 16744 13587 16832 13640
rect 16744 13447 16757 13587
rect 16803 13447 16832 13587
rect 16744 13396 16832 13447
rect 16932 13587 17020 13640
rect 16932 13447 16961 13587
rect 17007 13447 17020 13587
rect 16932 13396 17020 13447
rect 17640 13587 17728 13640
rect 17640 13447 17653 13587
rect 17699 13447 17728 13587
rect 17640 13396 17728 13447
rect 17828 13587 17916 13640
rect 17828 13447 17857 13587
rect 17903 13447 17916 13587
rect 17828 13396 17916 13447
rect 18312 13587 18400 13640
rect 18312 13447 18325 13587
rect 18371 13447 18400 13587
rect 18312 13396 18400 13447
rect 18500 13587 18588 13640
rect 18500 13447 18529 13587
rect 18575 13447 18588 13587
rect 18500 13396 18588 13447
rect 18740 13595 18828 13640
rect 18740 13455 18753 13595
rect 18799 13455 18828 13595
rect 18740 13396 18828 13455
rect 19028 13595 19116 13640
rect 19028 13455 19057 13595
rect 19103 13455 19116 13595
rect 19028 13396 19116 13455
rect 19188 13595 19276 13640
rect 19188 13455 19201 13595
rect 19247 13455 19276 13595
rect 19188 13396 19276 13455
rect 19476 13595 19564 13640
rect 19476 13455 19505 13595
rect 19551 13455 19564 13595
rect 19476 13396 19564 13455
rect 19636 13595 19724 13640
rect 19636 13455 19649 13595
rect 19695 13455 19724 13595
rect 19636 13396 19724 13455
rect 19924 13595 20012 13640
rect 19924 13455 19953 13595
rect 19999 13455 20012 13595
rect 19924 13396 20012 13455
rect 20084 13595 20172 13640
rect 20084 13455 20097 13595
rect 20143 13455 20172 13595
rect 20084 13396 20172 13455
rect 20372 13595 20460 13640
rect 20372 13455 20401 13595
rect 20447 13455 20460 13595
rect 20372 13396 20460 13455
rect 20532 13595 20620 13640
rect 20532 13455 20545 13595
rect 20591 13455 20620 13595
rect 20532 13396 20620 13455
rect 20820 13595 20908 13640
rect 20820 13455 20849 13595
rect 20895 13455 20908 13595
rect 20820 13396 20908 13455
rect 20980 13595 21068 13640
rect 20980 13455 20993 13595
rect 21039 13455 21068 13595
rect 20980 13396 21068 13455
rect 21268 13595 21356 13640
rect 21268 13455 21297 13595
rect 21343 13455 21356 13595
rect 21268 13396 21356 13455
rect 21428 13595 21516 13640
rect 21428 13455 21441 13595
rect 21487 13455 21516 13595
rect 21428 13396 21516 13455
rect 21716 13595 21804 13640
rect 21716 13455 21745 13595
rect 21791 13455 21804 13595
rect 21716 13396 21804 13455
rect 21876 13595 21964 13640
rect 21876 13455 21889 13595
rect 21935 13455 21964 13595
rect 21876 13396 21964 13455
rect 22164 13595 22252 13640
rect 22164 13455 22193 13595
rect 22239 13455 22252 13595
rect 22164 13396 22252 13455
rect 1604 13201 1692 13260
rect 1604 13061 1617 13201
rect 1663 13061 1692 13201
rect 1604 13016 1692 13061
rect 1892 13201 1980 13260
rect 1892 13061 1921 13201
rect 1967 13061 1980 13201
rect 1892 13016 1980 13061
rect 2052 13201 2140 13260
rect 2052 13061 2065 13201
rect 2111 13061 2140 13201
rect 2052 13016 2140 13061
rect 2340 13201 2428 13260
rect 2340 13061 2369 13201
rect 2415 13061 2428 13201
rect 2340 13016 2428 13061
rect 2500 13201 2588 13260
rect 2500 13061 2513 13201
rect 2559 13061 2588 13201
rect 2500 13016 2588 13061
rect 2788 13201 2876 13260
rect 2788 13061 2817 13201
rect 2863 13061 2876 13201
rect 2788 13016 2876 13061
rect 2948 13201 3036 13260
rect 2948 13061 2961 13201
rect 3007 13061 3036 13201
rect 2948 13016 3036 13061
rect 3236 13201 3324 13260
rect 3236 13061 3265 13201
rect 3311 13061 3324 13201
rect 3236 13016 3324 13061
rect 3396 13201 3484 13260
rect 3396 13061 3409 13201
rect 3455 13061 3484 13201
rect 3396 13016 3484 13061
rect 3684 13201 3772 13260
rect 3684 13061 3713 13201
rect 3759 13061 3772 13201
rect 3684 13016 3772 13061
rect 3844 13201 3932 13260
rect 3844 13061 3857 13201
rect 3903 13061 3932 13201
rect 3844 13016 3932 13061
rect 4132 13201 4220 13260
rect 4132 13061 4161 13201
rect 4207 13061 4220 13201
rect 4132 13016 4220 13061
rect 4292 13201 4380 13260
rect 4292 13061 4305 13201
rect 4351 13061 4380 13201
rect 4292 13016 4380 13061
rect 4580 13201 4668 13260
rect 4580 13061 4609 13201
rect 4655 13061 4668 13201
rect 4580 13016 4668 13061
rect 4740 13201 4828 13260
rect 4740 13061 4753 13201
rect 4799 13061 4828 13201
rect 4740 13016 4828 13061
rect 5028 13201 5116 13260
rect 5028 13061 5057 13201
rect 5103 13061 5116 13201
rect 5028 13016 5116 13061
rect 5524 13201 5612 13260
rect 5524 13061 5537 13201
rect 5583 13061 5612 13201
rect 5524 13016 5612 13061
rect 5812 13201 5900 13260
rect 5812 13061 5841 13201
rect 5887 13061 5900 13201
rect 5812 13016 5900 13061
rect 5972 13201 6060 13260
rect 5972 13061 5985 13201
rect 6031 13061 6060 13201
rect 5972 13016 6060 13061
rect 6260 13201 6348 13260
rect 6260 13061 6289 13201
rect 6335 13061 6348 13201
rect 6260 13016 6348 13061
rect 6420 13201 6508 13260
rect 6420 13061 6433 13201
rect 6479 13061 6508 13201
rect 6420 13016 6508 13061
rect 6708 13201 6796 13260
rect 6708 13061 6737 13201
rect 6783 13061 6796 13201
rect 6708 13016 6796 13061
rect 6868 13201 6956 13260
rect 6868 13061 6881 13201
rect 6927 13061 6956 13201
rect 6868 13016 6956 13061
rect 7156 13201 7244 13260
rect 7156 13061 7185 13201
rect 7231 13061 7244 13201
rect 7156 13016 7244 13061
rect 7316 13201 7404 13260
rect 7316 13061 7329 13201
rect 7375 13061 7404 13201
rect 7316 13016 7404 13061
rect 7604 13201 7692 13260
rect 7604 13061 7633 13201
rect 7679 13061 7692 13201
rect 7604 13016 7692 13061
rect 7764 13201 7852 13260
rect 7764 13061 7777 13201
rect 7823 13061 7852 13201
rect 7764 13016 7852 13061
rect 8052 13201 8140 13260
rect 8052 13061 8081 13201
rect 8127 13061 8140 13201
rect 8052 13016 8140 13061
rect 8212 13201 8300 13260
rect 8212 13061 8225 13201
rect 8271 13061 8300 13201
rect 8212 13016 8300 13061
rect 8500 13201 8588 13260
rect 8500 13061 8529 13201
rect 8575 13061 8588 13201
rect 8500 13016 8588 13061
rect 8660 13201 8748 13260
rect 8660 13061 8673 13201
rect 8719 13061 8748 13201
rect 8660 13016 8748 13061
rect 8948 13201 9036 13260
rect 8948 13061 8977 13201
rect 9023 13061 9036 13201
rect 8948 13016 9036 13061
rect 9108 13201 9196 13260
rect 9108 13061 9121 13201
rect 9167 13061 9196 13201
rect 9108 13016 9196 13061
rect 9396 13201 9484 13260
rect 9396 13061 9425 13201
rect 9471 13061 9484 13201
rect 9396 13016 9484 13061
rect 9556 13201 9644 13260
rect 9556 13061 9569 13201
rect 9615 13061 9644 13201
rect 9556 13016 9644 13061
rect 9844 13201 9932 13260
rect 9844 13061 9873 13201
rect 9919 13061 9932 13201
rect 9844 13016 9932 13061
rect 10004 13201 10092 13260
rect 10004 13061 10017 13201
rect 10063 13061 10092 13201
rect 10004 13016 10092 13061
rect 10292 13201 10380 13260
rect 10292 13061 10321 13201
rect 10367 13061 10380 13201
rect 10292 13016 10380 13061
rect 10452 13201 10540 13260
rect 10452 13061 10465 13201
rect 10511 13061 10540 13201
rect 10452 13016 10540 13061
rect 10740 13201 10828 13260
rect 10740 13061 10769 13201
rect 10815 13061 10828 13201
rect 10740 13016 10828 13061
rect 10900 13201 10988 13260
rect 10900 13061 10913 13201
rect 10959 13061 10988 13201
rect 10900 13016 10988 13061
rect 11188 13201 11276 13260
rect 11188 13061 11217 13201
rect 11263 13061 11276 13201
rect 11188 13016 11276 13061
rect 11348 13201 11436 13260
rect 11348 13061 11361 13201
rect 11407 13061 11436 13201
rect 11348 13016 11436 13061
rect 11636 13201 11724 13260
rect 11636 13061 11665 13201
rect 11711 13061 11724 13201
rect 11636 13016 11724 13061
rect 11796 13201 11884 13260
rect 11796 13061 11809 13201
rect 11855 13061 11884 13201
rect 11796 13016 11884 13061
rect 12084 13201 12172 13260
rect 12084 13061 12113 13201
rect 12159 13061 12172 13201
rect 12084 13016 12172 13061
rect 12244 13201 12332 13260
rect 12244 13061 12257 13201
rect 12303 13061 12332 13201
rect 12244 13016 12332 13061
rect 12532 13201 12620 13260
rect 12532 13061 12561 13201
rect 12607 13061 12620 13201
rect 12532 13016 12620 13061
rect 12692 13201 12780 13260
rect 12692 13061 12705 13201
rect 12751 13061 12780 13201
rect 12692 13016 12780 13061
rect 12980 13201 13068 13260
rect 12980 13061 13009 13201
rect 13055 13061 13068 13201
rect 12980 13016 13068 13061
rect 13476 13201 13564 13260
rect 13476 13061 13489 13201
rect 13535 13061 13564 13201
rect 13476 13016 13564 13061
rect 13764 13201 13852 13260
rect 13764 13061 13793 13201
rect 13839 13061 13852 13201
rect 13764 13016 13852 13061
rect 13924 13201 14012 13260
rect 13924 13061 13937 13201
rect 13983 13061 14012 13201
rect 13924 13016 14012 13061
rect 14212 13201 14300 13260
rect 14212 13061 14241 13201
rect 14287 13061 14300 13201
rect 14212 13016 14300 13061
rect 14728 13209 14816 13260
rect 14728 13069 14741 13209
rect 14787 13069 14816 13209
rect 14728 13016 14816 13069
rect 14916 13209 15004 13260
rect 14916 13069 14945 13209
rect 14991 13069 15004 13209
rect 14916 13016 15004 13069
rect 15400 13209 15488 13260
rect 15400 13069 15413 13209
rect 15459 13069 15488 13209
rect 15400 13016 15488 13069
rect 15588 13209 15676 13260
rect 15588 13069 15617 13209
rect 15663 13069 15676 13209
rect 15588 13016 15676 13069
rect 16072 13209 16160 13260
rect 16072 13069 16085 13209
rect 16131 13069 16160 13209
rect 16072 13016 16160 13069
rect 16260 13209 16348 13260
rect 16260 13069 16289 13209
rect 16335 13069 16348 13209
rect 16260 13016 16348 13069
rect 16744 13209 16832 13260
rect 16744 13069 16757 13209
rect 16803 13069 16832 13209
rect 16744 13016 16832 13069
rect 16932 13209 17020 13260
rect 16932 13069 16961 13209
rect 17007 13069 17020 13209
rect 16932 13016 17020 13069
rect 17416 13209 17504 13260
rect 17416 13069 17429 13209
rect 17475 13069 17504 13209
rect 17416 13016 17504 13069
rect 17604 13209 17692 13260
rect 17604 13069 17633 13209
rect 17679 13069 17692 13209
rect 17604 13016 17692 13069
rect 18088 13209 18176 13260
rect 18088 13069 18101 13209
rect 18147 13069 18176 13209
rect 18088 13016 18176 13069
rect 18276 13209 18364 13260
rect 18276 13069 18305 13209
rect 18351 13069 18364 13209
rect 18276 13016 18364 13069
rect 18760 13209 18848 13260
rect 18760 13069 18773 13209
rect 18819 13069 18848 13209
rect 18760 13016 18848 13069
rect 18948 13209 19036 13260
rect 18948 13069 18977 13209
rect 19023 13069 19036 13209
rect 18948 13016 19036 13069
rect 19432 13209 19520 13260
rect 19432 13069 19445 13209
rect 19491 13069 19520 13209
rect 19432 13016 19520 13069
rect 19620 13209 19708 13260
rect 19620 13069 19649 13209
rect 19695 13069 19708 13209
rect 19620 13016 19708 13069
rect 19860 13201 19948 13260
rect 19860 13061 19873 13201
rect 19919 13061 19948 13201
rect 19860 13016 19948 13061
rect 20148 13201 20236 13260
rect 20148 13061 20177 13201
rect 20223 13061 20236 13201
rect 20148 13016 20236 13061
rect 20308 13201 20396 13260
rect 20308 13061 20321 13201
rect 20367 13061 20396 13201
rect 20308 13016 20396 13061
rect 20596 13201 20684 13260
rect 20596 13061 20625 13201
rect 20671 13061 20684 13201
rect 20596 13016 20684 13061
rect 20756 13201 20844 13260
rect 20756 13061 20769 13201
rect 20815 13061 20844 13201
rect 20756 13016 20844 13061
rect 21044 13201 21132 13260
rect 21044 13061 21073 13201
rect 21119 13061 21132 13201
rect 21044 13016 21132 13061
rect 21428 13201 21516 13260
rect 21428 13061 21441 13201
rect 21487 13061 21516 13201
rect 21428 13016 21516 13061
rect 21716 13201 21804 13260
rect 21716 13061 21745 13201
rect 21791 13061 21804 13201
rect 21716 13016 21804 13061
rect 21876 13201 21964 13260
rect 21876 13061 21889 13201
rect 21935 13061 21964 13201
rect 21876 13016 21964 13061
rect 22164 13201 22252 13260
rect 22164 13061 22193 13201
rect 22239 13061 22252 13201
rect 22164 13016 22252 13061
rect 1604 12027 1692 12072
rect 1604 11887 1617 12027
rect 1663 11887 1692 12027
rect 1604 11828 1692 11887
rect 1892 12027 1980 12072
rect 1892 11887 1921 12027
rect 1967 11887 1980 12027
rect 1892 11828 1980 11887
rect 2052 12027 2140 12072
rect 2052 11887 2065 12027
rect 2111 11887 2140 12027
rect 2052 11828 2140 11887
rect 2340 12027 2428 12072
rect 2340 11887 2369 12027
rect 2415 11887 2428 12027
rect 2340 11828 2428 11887
rect 2500 12027 2588 12072
rect 2500 11887 2513 12027
rect 2559 11887 2588 12027
rect 2500 11828 2588 11887
rect 2788 12027 2876 12072
rect 2788 11887 2817 12027
rect 2863 11887 2876 12027
rect 2788 11828 2876 11887
rect 2948 12027 3036 12072
rect 2948 11887 2961 12027
rect 3007 11887 3036 12027
rect 2948 11828 3036 11887
rect 3236 12027 3324 12072
rect 3236 11887 3265 12027
rect 3311 11887 3324 12027
rect 3236 11828 3324 11887
rect 3396 12027 3484 12072
rect 3396 11887 3409 12027
rect 3455 11887 3484 12027
rect 3396 11828 3484 11887
rect 3684 12027 3772 12072
rect 3684 11887 3713 12027
rect 3759 11887 3772 12027
rect 3684 11828 3772 11887
rect 3844 12027 3932 12072
rect 3844 11887 3857 12027
rect 3903 11887 3932 12027
rect 3844 11828 3932 11887
rect 4132 12027 4220 12072
rect 4132 11887 4161 12027
rect 4207 11887 4220 12027
rect 4132 11828 4220 11887
rect 4292 12027 4380 12072
rect 4292 11887 4305 12027
rect 4351 11887 4380 12027
rect 4292 11828 4380 11887
rect 4580 12027 4668 12072
rect 4580 11887 4609 12027
rect 4655 11887 4668 12027
rect 4580 11828 4668 11887
rect 4740 12027 4828 12072
rect 4740 11887 4753 12027
rect 4799 11887 4828 12027
rect 4740 11828 4828 11887
rect 5028 12027 5116 12072
rect 5028 11887 5057 12027
rect 5103 11887 5116 12027
rect 5028 11828 5116 11887
rect 5188 12027 5276 12072
rect 5188 11887 5201 12027
rect 5247 11887 5276 12027
rect 5188 11828 5276 11887
rect 5476 12027 5564 12072
rect 5476 11887 5505 12027
rect 5551 11887 5564 12027
rect 5476 11828 5564 11887
rect 5636 12027 5724 12072
rect 5636 11887 5649 12027
rect 5695 11887 5724 12027
rect 5636 11828 5724 11887
rect 5924 12027 6012 12072
rect 5924 11887 5953 12027
rect 5999 11887 6012 12027
rect 5924 11828 6012 11887
rect 6084 12027 6172 12072
rect 6084 11887 6097 12027
rect 6143 11887 6172 12027
rect 6084 11828 6172 11887
rect 6372 12027 6460 12072
rect 6372 11887 6401 12027
rect 6447 11887 6460 12027
rect 6372 11828 6460 11887
rect 6532 12027 6620 12072
rect 6532 11887 6545 12027
rect 6591 11887 6620 12027
rect 6532 11828 6620 11887
rect 6820 12027 6908 12072
rect 6820 11887 6849 12027
rect 6895 11887 6908 12027
rect 6820 11828 6908 11887
rect 6980 12027 7068 12072
rect 6980 11887 6993 12027
rect 7039 11887 7068 12027
rect 6980 11828 7068 11887
rect 7268 12027 7356 12072
rect 7268 11887 7297 12027
rect 7343 11887 7356 12027
rect 7268 11828 7356 11887
rect 7428 12027 7516 12072
rect 7428 11887 7441 12027
rect 7487 11887 7516 12027
rect 7428 11828 7516 11887
rect 7716 12027 7804 12072
rect 7716 11887 7745 12027
rect 7791 11887 7804 12027
rect 7716 11828 7804 11887
rect 7876 12027 7964 12072
rect 7876 11887 7889 12027
rect 7935 11887 7964 12027
rect 7876 11828 7964 11887
rect 8164 12027 8252 12072
rect 8164 11887 8193 12027
rect 8239 11887 8252 12027
rect 8164 11828 8252 11887
rect 8324 12027 8412 12072
rect 8324 11887 8337 12027
rect 8383 11887 8412 12027
rect 8324 11828 8412 11887
rect 8612 12027 8700 12072
rect 8612 11887 8641 12027
rect 8687 11887 8700 12027
rect 8612 11828 8700 11887
rect 8772 12027 8860 12072
rect 8772 11887 8785 12027
rect 8831 11887 8860 12027
rect 8772 11828 8860 11887
rect 9060 12027 9148 12072
rect 9060 11887 9089 12027
rect 9135 11887 9148 12027
rect 9060 11828 9148 11887
rect 9556 12027 9644 12072
rect 9556 11887 9569 12027
rect 9615 11887 9644 12027
rect 9556 11828 9644 11887
rect 9844 12027 9932 12072
rect 9844 11887 9873 12027
rect 9919 11887 9932 12027
rect 9844 11828 9932 11887
rect 10004 12027 10092 12072
rect 10004 11887 10017 12027
rect 10063 11887 10092 12027
rect 10004 11828 10092 11887
rect 10292 12027 10380 12072
rect 10292 11887 10321 12027
rect 10367 11887 10380 12027
rect 10292 11828 10380 11887
rect 10452 12027 10540 12072
rect 10452 11887 10465 12027
rect 10511 11887 10540 12027
rect 10452 11828 10540 11887
rect 10740 12027 10828 12072
rect 10740 11887 10769 12027
rect 10815 11887 10828 12027
rect 10740 11828 10828 11887
rect 10900 12027 10988 12072
rect 10900 11887 10913 12027
rect 10959 11887 10988 12027
rect 10900 11828 10988 11887
rect 11188 12027 11276 12072
rect 11188 11887 11217 12027
rect 11263 11887 11276 12027
rect 11188 11828 11276 11887
rect 11348 12027 11436 12072
rect 11348 11887 11361 12027
rect 11407 11887 11436 12027
rect 11348 11828 11436 11887
rect 11636 12027 11724 12072
rect 11636 11887 11665 12027
rect 11711 11887 11724 12027
rect 11636 11828 11724 11887
rect 11796 12027 11884 12072
rect 11796 11887 11809 12027
rect 11855 11887 11884 12027
rect 11796 11828 11884 11887
rect 12084 12027 12172 12072
rect 12084 11887 12113 12027
rect 12159 11887 12172 12027
rect 12084 11828 12172 11887
rect 12244 12027 12332 12072
rect 12244 11887 12257 12027
rect 12303 11887 12332 12027
rect 12244 11828 12332 11887
rect 12532 12027 12620 12072
rect 12532 11887 12561 12027
rect 12607 11887 12620 12027
rect 12532 11828 12620 11887
rect 12692 12027 12780 12072
rect 12692 11887 12705 12027
rect 12751 11887 12780 12027
rect 12692 11828 12780 11887
rect 12980 12027 13068 12072
rect 12980 11887 13009 12027
rect 13055 11887 13068 12027
rect 12980 11828 13068 11887
rect 13140 12027 13228 12072
rect 13140 11887 13153 12027
rect 13199 11887 13228 12027
rect 13140 11828 13228 11887
rect 13428 12027 13516 12072
rect 13428 11887 13457 12027
rect 13503 11887 13516 12027
rect 13428 11828 13516 11887
rect 13588 12027 13676 12072
rect 13588 11887 13601 12027
rect 13647 11887 13676 12027
rect 13588 11828 13676 11887
rect 13876 12027 13964 12072
rect 13876 11887 13905 12027
rect 13951 11887 13964 12027
rect 13876 11828 13964 11887
rect 14056 12019 14144 12072
rect 14056 11879 14069 12019
rect 14115 11879 14144 12019
rect 14056 11828 14144 11879
rect 14244 12019 14332 12072
rect 14244 11879 14273 12019
rect 14319 11879 14332 12019
rect 14244 11828 14332 11879
rect 14728 12019 14816 12072
rect 14728 11879 14741 12019
rect 14787 11879 14816 12019
rect 14728 11828 14816 11879
rect 14916 12019 15004 12072
rect 14916 11879 14945 12019
rect 14991 11879 15004 12019
rect 14916 11828 15004 11879
rect 15400 12019 15488 12072
rect 15400 11879 15413 12019
rect 15459 11879 15488 12019
rect 15400 11828 15488 11879
rect 15588 12019 15676 12072
rect 15588 11879 15617 12019
rect 15663 11879 15676 12019
rect 15588 11828 15676 11879
rect 16072 12019 16160 12072
rect 16072 11879 16085 12019
rect 16131 11879 16160 12019
rect 16072 11828 16160 11879
rect 16260 12019 16348 12072
rect 16260 11879 16289 12019
rect 16335 11879 16348 12019
rect 16260 11828 16348 11879
rect 16744 12019 16832 12072
rect 16744 11879 16757 12019
rect 16803 11879 16832 12019
rect 16744 11828 16832 11879
rect 16932 12019 17020 12072
rect 16932 11879 16961 12019
rect 17007 11879 17020 12019
rect 16932 11828 17020 11879
rect 17640 12019 17728 12072
rect 17640 11879 17653 12019
rect 17699 11879 17728 12019
rect 17640 11828 17728 11879
rect 17828 12019 17916 12072
rect 17828 11879 17857 12019
rect 17903 11879 17916 12019
rect 17828 11828 17916 11879
rect 18312 12019 18400 12072
rect 18312 11879 18325 12019
rect 18371 11879 18400 12019
rect 18312 11828 18400 11879
rect 18500 12019 18588 12072
rect 18500 11879 18529 12019
rect 18575 11879 18588 12019
rect 18500 11828 18588 11879
rect 18984 12019 19072 12072
rect 18984 11879 18997 12019
rect 19043 11879 19072 12019
rect 18984 11828 19072 11879
rect 19172 12019 19260 12072
rect 19172 11879 19201 12019
rect 19247 11879 19260 12019
rect 19172 11828 19260 11879
rect 19656 12019 19744 12072
rect 19656 11879 19669 12019
rect 19715 11879 19744 12019
rect 19656 11828 19744 11879
rect 19844 12019 19932 12072
rect 19844 11879 19873 12019
rect 19919 11879 19932 12019
rect 19844 11828 19932 11879
rect 20328 12019 20416 12072
rect 20328 11879 20341 12019
rect 20387 11879 20416 12019
rect 20328 11828 20416 11879
rect 20516 12019 20604 12072
rect 20516 11879 20545 12019
rect 20591 11879 20604 12019
rect 20516 11828 20604 11879
rect 20756 12027 20844 12072
rect 20756 11887 20769 12027
rect 20815 11887 20844 12027
rect 20756 11828 20844 11887
rect 21044 12027 21132 12072
rect 21044 11887 21073 12027
rect 21119 11887 21132 12027
rect 21044 11828 21132 11887
rect 21204 12027 21292 12072
rect 21204 11887 21217 12027
rect 21263 11887 21292 12027
rect 21204 11828 21292 11887
rect 21492 12027 21580 12072
rect 21492 11887 21521 12027
rect 21567 11887 21580 12027
rect 21492 11828 21580 11887
rect 21652 12027 21740 12072
rect 21652 11887 21665 12027
rect 21711 11887 21740 12027
rect 21652 11828 21740 11887
rect 21940 12027 22028 12072
rect 21940 11887 21969 12027
rect 22015 11887 22028 12027
rect 21940 11828 22028 11887
rect 1604 11633 1692 11692
rect 1604 11493 1617 11633
rect 1663 11493 1692 11633
rect 1604 11448 1692 11493
rect 1892 11633 1980 11692
rect 1892 11493 1921 11633
rect 1967 11493 1980 11633
rect 1892 11448 1980 11493
rect 2052 11633 2140 11692
rect 2052 11493 2065 11633
rect 2111 11493 2140 11633
rect 2052 11448 2140 11493
rect 2340 11633 2428 11692
rect 2340 11493 2369 11633
rect 2415 11493 2428 11633
rect 2340 11448 2428 11493
rect 2500 11633 2588 11692
rect 2500 11493 2513 11633
rect 2559 11493 2588 11633
rect 2500 11448 2588 11493
rect 2788 11633 2876 11692
rect 2788 11493 2817 11633
rect 2863 11493 2876 11633
rect 2788 11448 2876 11493
rect 2948 11633 3036 11692
rect 2948 11493 2961 11633
rect 3007 11493 3036 11633
rect 2948 11448 3036 11493
rect 3236 11633 3324 11692
rect 3236 11493 3265 11633
rect 3311 11493 3324 11633
rect 3236 11448 3324 11493
rect 3396 11633 3484 11692
rect 3396 11493 3409 11633
rect 3455 11493 3484 11633
rect 3396 11448 3484 11493
rect 3684 11633 3772 11692
rect 3684 11493 3713 11633
rect 3759 11493 3772 11633
rect 3684 11448 3772 11493
rect 3844 11633 3932 11692
rect 3844 11493 3857 11633
rect 3903 11493 3932 11633
rect 3844 11448 3932 11493
rect 4132 11633 4220 11692
rect 4132 11493 4161 11633
rect 4207 11493 4220 11633
rect 4132 11448 4220 11493
rect 4292 11633 4380 11692
rect 4292 11493 4305 11633
rect 4351 11493 4380 11633
rect 4292 11448 4380 11493
rect 4580 11633 4668 11692
rect 4580 11493 4609 11633
rect 4655 11493 4668 11633
rect 4580 11448 4668 11493
rect 4740 11633 4828 11692
rect 4740 11493 4753 11633
rect 4799 11493 4828 11633
rect 4740 11448 4828 11493
rect 5028 11633 5116 11692
rect 5028 11493 5057 11633
rect 5103 11493 5116 11633
rect 5028 11448 5116 11493
rect 5524 11633 5612 11692
rect 5524 11493 5537 11633
rect 5583 11493 5612 11633
rect 5524 11448 5612 11493
rect 5812 11633 5900 11692
rect 5812 11493 5841 11633
rect 5887 11493 5900 11633
rect 5812 11448 5900 11493
rect 6052 11641 6140 11692
rect 6052 11501 6065 11641
rect 6111 11501 6140 11641
rect 6052 11448 6140 11501
rect 6240 11641 6328 11692
rect 6240 11501 6269 11641
rect 6315 11501 6328 11641
rect 6240 11448 6328 11501
rect 6836 11641 6924 11692
rect 6836 11501 6849 11641
rect 6895 11501 6924 11641
rect 6836 11448 6924 11501
rect 7024 11641 7112 11692
rect 7024 11501 7053 11641
rect 7099 11501 7112 11641
rect 7024 11448 7112 11501
rect 7508 11641 7596 11692
rect 7508 11501 7521 11641
rect 7567 11501 7596 11641
rect 7508 11448 7596 11501
rect 7696 11641 7784 11692
rect 7696 11501 7725 11641
rect 7771 11501 7784 11641
rect 7696 11448 7784 11501
rect 8180 11641 8268 11692
rect 8180 11501 8193 11641
rect 8239 11501 8268 11641
rect 8180 11448 8268 11501
rect 8368 11641 8456 11692
rect 8368 11501 8397 11641
rect 8443 11501 8456 11641
rect 8368 11448 8456 11501
rect 8548 11633 8636 11692
rect 8548 11493 8561 11633
rect 8607 11493 8636 11633
rect 8548 11448 8636 11493
rect 8836 11633 8924 11692
rect 8836 11493 8865 11633
rect 8911 11493 8924 11633
rect 8836 11448 8924 11493
rect 9128 11641 9216 11692
rect 9128 11501 9141 11641
rect 9187 11501 9216 11641
rect 9128 11448 9216 11501
rect 9316 11641 9404 11692
rect 9316 11501 9345 11641
rect 9391 11501 9404 11641
rect 9316 11448 9404 11501
rect 9800 11641 9888 11692
rect 9800 11501 9813 11641
rect 9859 11501 9888 11641
rect 9800 11448 9888 11501
rect 9988 11641 10076 11692
rect 9988 11501 10017 11641
rect 10063 11501 10076 11641
rect 9988 11448 10076 11501
rect 10472 11641 10560 11692
rect 10472 11501 10485 11641
rect 10531 11501 10560 11641
rect 10472 11448 10560 11501
rect 10660 11641 10748 11692
rect 10660 11501 10689 11641
rect 10735 11501 10748 11641
rect 10660 11448 10748 11501
rect 10900 11633 10988 11692
rect 10900 11493 10913 11633
rect 10959 11493 10988 11633
rect 10900 11448 10988 11493
rect 11188 11633 11276 11692
rect 11188 11493 11217 11633
rect 11263 11493 11276 11633
rect 11188 11448 11276 11493
rect 11348 11633 11436 11692
rect 11348 11493 11361 11633
rect 11407 11493 11436 11633
rect 11348 11448 11436 11493
rect 11636 11633 11724 11692
rect 11636 11493 11665 11633
rect 11711 11493 11724 11633
rect 11636 11448 11724 11493
rect 12040 11641 12128 11692
rect 12040 11501 12053 11641
rect 12099 11501 12128 11641
rect 12040 11448 12128 11501
rect 12228 11641 12316 11692
rect 12228 11501 12257 11641
rect 12303 11501 12316 11641
rect 12228 11448 12316 11501
rect 12712 11641 12800 11692
rect 12712 11501 12725 11641
rect 12771 11501 12800 11641
rect 12712 11448 12800 11501
rect 12900 11641 12988 11692
rect 12900 11501 12929 11641
rect 12975 11501 12988 11641
rect 12900 11448 12988 11501
rect 13608 11641 13696 11692
rect 13608 11501 13621 11641
rect 13667 11501 13696 11641
rect 13608 11448 13696 11501
rect 13796 11641 13884 11692
rect 13796 11501 13825 11641
rect 13871 11501 13884 11641
rect 13796 11448 13884 11501
rect 14036 11633 14124 11692
rect 14036 11493 14049 11633
rect 14095 11493 14124 11633
rect 14036 11448 14124 11493
rect 14324 11633 14412 11692
rect 14324 11493 14353 11633
rect 14399 11493 14412 11633
rect 14324 11448 14412 11493
rect 14728 11641 14816 11692
rect 14728 11501 14741 11641
rect 14787 11501 14816 11641
rect 14728 11448 14816 11501
rect 14916 11641 15004 11692
rect 14916 11501 14945 11641
rect 14991 11501 15004 11641
rect 14916 11448 15004 11501
rect 15400 11641 15488 11692
rect 15400 11501 15413 11641
rect 15459 11501 15488 11641
rect 15400 11448 15488 11501
rect 15588 11641 15676 11692
rect 15588 11501 15617 11641
rect 15663 11501 15676 11641
rect 15588 11448 15676 11501
rect 16072 11641 16160 11692
rect 16072 11501 16085 11641
rect 16131 11501 16160 11641
rect 16072 11448 16160 11501
rect 16260 11641 16348 11692
rect 16260 11501 16289 11641
rect 16335 11501 16348 11641
rect 16260 11448 16348 11501
rect 16744 11641 16832 11692
rect 16744 11501 16757 11641
rect 16803 11501 16832 11641
rect 16744 11448 16832 11501
rect 16932 11641 17020 11692
rect 16932 11501 16961 11641
rect 17007 11501 17020 11641
rect 16932 11448 17020 11501
rect 17416 11641 17504 11692
rect 17416 11501 17429 11641
rect 17475 11501 17504 11641
rect 17416 11448 17504 11501
rect 17604 11641 17692 11692
rect 17604 11501 17633 11641
rect 17679 11501 17692 11641
rect 17604 11448 17692 11501
rect 18088 11641 18176 11692
rect 18088 11501 18101 11641
rect 18147 11501 18176 11641
rect 18088 11448 18176 11501
rect 18276 11641 18364 11692
rect 18276 11501 18305 11641
rect 18351 11501 18364 11641
rect 18276 11448 18364 11501
rect 18760 11641 18848 11692
rect 18760 11501 18773 11641
rect 18819 11501 18848 11641
rect 18760 11448 18848 11501
rect 18948 11641 19036 11692
rect 18948 11501 18977 11641
rect 19023 11501 19036 11641
rect 18948 11448 19036 11501
rect 19432 11641 19520 11692
rect 19432 11501 19445 11641
rect 19491 11501 19520 11641
rect 19432 11448 19520 11501
rect 19620 11641 19708 11692
rect 19620 11501 19649 11641
rect 19695 11501 19708 11641
rect 19620 11448 19708 11501
rect 20104 11641 20192 11692
rect 20104 11501 20117 11641
rect 20163 11501 20192 11641
rect 20104 11448 20192 11501
rect 20292 11641 20380 11692
rect 20292 11501 20321 11641
rect 20367 11501 20380 11641
rect 20292 11448 20380 11501
rect 20532 11633 20620 11692
rect 20532 11493 20545 11633
rect 20591 11493 20620 11633
rect 20532 11448 20620 11493
rect 20820 11633 20908 11692
rect 20820 11493 20849 11633
rect 20895 11493 20908 11633
rect 20820 11448 20908 11493
rect 21428 11633 21516 11692
rect 21428 11493 21441 11633
rect 21487 11493 21516 11633
rect 21428 11448 21516 11493
rect 21716 11633 21804 11692
rect 21716 11493 21745 11633
rect 21791 11493 21804 11633
rect 21716 11448 21804 11493
rect 21876 11633 21964 11692
rect 21876 11493 21889 11633
rect 21935 11493 21964 11633
rect 21876 11448 21964 11493
rect 22164 11633 22252 11692
rect 22164 11493 22193 11633
rect 22239 11493 22252 11633
rect 22164 11448 22252 11493
rect 1604 10459 1692 10504
rect 1604 10319 1617 10459
rect 1663 10319 1692 10459
rect 1604 10260 1692 10319
rect 1892 10459 1980 10504
rect 1892 10319 1921 10459
rect 1967 10319 1980 10459
rect 1892 10260 1980 10319
rect 2052 10459 2140 10504
rect 2052 10319 2065 10459
rect 2111 10319 2140 10459
rect 2052 10260 2140 10319
rect 2340 10459 2428 10504
rect 2340 10319 2369 10459
rect 2415 10319 2428 10459
rect 2340 10260 2428 10319
rect 2500 10459 2588 10504
rect 2500 10319 2513 10459
rect 2559 10319 2588 10459
rect 2500 10260 2588 10319
rect 2788 10459 2876 10504
rect 2788 10319 2817 10459
rect 2863 10319 2876 10459
rect 2788 10260 2876 10319
rect 2948 10459 3036 10504
rect 2948 10319 2961 10459
rect 3007 10319 3036 10459
rect 2948 10260 3036 10319
rect 3236 10459 3324 10504
rect 3236 10319 3265 10459
rect 3311 10319 3324 10459
rect 3236 10260 3324 10319
rect 3396 10459 3484 10504
rect 3396 10319 3409 10459
rect 3455 10319 3484 10459
rect 3396 10260 3484 10319
rect 3684 10459 3772 10504
rect 3684 10319 3713 10459
rect 3759 10319 3772 10459
rect 3684 10260 3772 10319
rect 3844 10459 3932 10504
rect 3844 10319 3857 10459
rect 3903 10319 3932 10459
rect 3844 10260 3932 10319
rect 4132 10459 4220 10504
rect 4132 10319 4161 10459
rect 4207 10319 4220 10459
rect 4132 10260 4220 10319
rect 4292 10459 4380 10504
rect 4292 10319 4305 10459
rect 4351 10319 4380 10459
rect 4292 10260 4380 10319
rect 4580 10459 4668 10504
rect 4580 10319 4609 10459
rect 4655 10319 4668 10459
rect 4580 10260 4668 10319
rect 4740 10459 4828 10504
rect 4740 10319 4753 10459
rect 4799 10319 4828 10459
rect 4740 10260 4828 10319
rect 5028 10459 5116 10504
rect 5028 10319 5057 10459
rect 5103 10319 5116 10459
rect 5028 10260 5116 10319
rect 5320 10451 5408 10504
rect 5320 10311 5333 10451
rect 5379 10311 5408 10451
rect 5320 10260 5408 10311
rect 5508 10451 5596 10504
rect 5508 10311 5537 10451
rect 5583 10311 5596 10451
rect 5508 10260 5596 10311
rect 5992 10451 6080 10504
rect 5992 10311 6005 10451
rect 6051 10311 6080 10451
rect 5992 10260 6080 10311
rect 6180 10451 6268 10504
rect 6180 10311 6209 10451
rect 6255 10311 6268 10451
rect 6180 10260 6268 10311
rect 6664 10451 6752 10504
rect 6664 10311 6677 10451
rect 6723 10311 6752 10451
rect 6664 10260 6752 10311
rect 6852 10451 6940 10504
rect 6852 10311 6881 10451
rect 6927 10311 6940 10451
rect 6852 10260 6940 10311
rect 7336 10451 7424 10504
rect 7336 10311 7349 10451
rect 7395 10311 7424 10451
rect 7336 10260 7424 10311
rect 7524 10451 7612 10504
rect 7524 10311 7553 10451
rect 7599 10311 7612 10451
rect 7524 10260 7612 10311
rect 8008 10451 8096 10504
rect 8008 10311 8021 10451
rect 8067 10311 8096 10451
rect 8008 10260 8096 10311
rect 8196 10451 8284 10504
rect 8196 10311 8225 10451
rect 8271 10311 8284 10451
rect 8196 10260 8284 10311
rect 8792 10451 8880 10504
rect 8792 10311 8805 10451
rect 8851 10311 8880 10451
rect 8792 10260 8880 10311
rect 8980 10451 9068 10504
rect 8980 10311 9009 10451
rect 9055 10311 9068 10451
rect 8980 10260 9068 10311
rect 9800 10451 9888 10504
rect 9800 10311 9813 10451
rect 9859 10311 9888 10451
rect 9800 10260 9888 10311
rect 9988 10451 10076 10504
rect 9988 10311 10017 10451
rect 10063 10311 10076 10451
rect 9988 10260 10076 10311
rect 10472 10451 10560 10504
rect 10472 10311 10485 10451
rect 10531 10311 10560 10451
rect 10472 10260 10560 10311
rect 10660 10451 10748 10504
rect 10660 10311 10689 10451
rect 10735 10311 10748 10451
rect 10660 10260 10748 10311
rect 11144 10451 11232 10504
rect 11144 10311 11157 10451
rect 11203 10311 11232 10451
rect 11144 10260 11232 10311
rect 11332 10451 11420 10504
rect 11332 10311 11361 10451
rect 11407 10311 11420 10451
rect 11332 10260 11420 10311
rect 11928 10451 12016 10504
rect 11928 10311 11941 10451
rect 11987 10311 12016 10451
rect 11928 10260 12016 10311
rect 12116 10451 12204 10504
rect 12116 10311 12145 10451
rect 12191 10311 12204 10451
rect 12116 10260 12204 10311
rect 12600 10451 12688 10504
rect 12600 10311 12613 10451
rect 12659 10311 12688 10451
rect 12600 10260 12688 10311
rect 12788 10451 12876 10504
rect 12788 10311 12817 10451
rect 12863 10311 12876 10451
rect 12788 10260 12876 10311
rect 13272 10451 13360 10504
rect 13272 10311 13285 10451
rect 13331 10311 13360 10451
rect 13272 10260 13360 10311
rect 13460 10451 13548 10504
rect 13460 10311 13489 10451
rect 13535 10311 13548 10451
rect 13460 10260 13548 10311
rect 13944 10451 14032 10504
rect 13944 10311 13957 10451
rect 14003 10311 14032 10451
rect 13944 10260 14032 10311
rect 14132 10451 14220 10504
rect 14132 10311 14161 10451
rect 14207 10311 14220 10451
rect 14132 10260 14220 10311
rect 14616 10451 14704 10504
rect 14616 10311 14629 10451
rect 14675 10311 14704 10451
rect 14616 10260 14704 10311
rect 14804 10451 14892 10504
rect 14804 10311 14833 10451
rect 14879 10311 14892 10451
rect 14804 10260 14892 10311
rect 15288 10451 15376 10504
rect 15288 10311 15301 10451
rect 15347 10311 15376 10451
rect 15288 10260 15376 10311
rect 15476 10451 15564 10504
rect 15476 10311 15505 10451
rect 15551 10311 15564 10451
rect 15476 10260 15564 10311
rect 15960 10451 16048 10504
rect 15960 10311 15973 10451
rect 16019 10311 16048 10451
rect 15960 10260 16048 10311
rect 16148 10451 16236 10504
rect 16148 10311 16177 10451
rect 16223 10311 16236 10451
rect 16148 10260 16236 10311
rect 16632 10451 16720 10504
rect 16632 10311 16645 10451
rect 16691 10311 16720 10451
rect 16632 10260 16720 10311
rect 16820 10451 16908 10504
rect 16820 10311 16849 10451
rect 16895 10311 16908 10451
rect 16820 10260 16908 10311
rect 17640 10451 17728 10504
rect 17640 10311 17653 10451
rect 17699 10311 17728 10451
rect 17640 10260 17728 10311
rect 17828 10451 17916 10504
rect 17828 10311 17857 10451
rect 17903 10311 17916 10451
rect 17828 10260 17916 10311
rect 18312 10451 18400 10504
rect 18312 10311 18325 10451
rect 18371 10311 18400 10451
rect 18312 10260 18400 10311
rect 18500 10451 18588 10504
rect 18500 10311 18529 10451
rect 18575 10311 18588 10451
rect 18500 10260 18588 10311
rect 18984 10451 19072 10504
rect 18984 10311 18997 10451
rect 19043 10311 19072 10451
rect 18984 10260 19072 10311
rect 19172 10451 19260 10504
rect 19172 10311 19201 10451
rect 19247 10311 19260 10451
rect 19172 10260 19260 10311
rect 19656 10451 19744 10504
rect 19656 10311 19669 10451
rect 19715 10311 19744 10451
rect 19656 10260 19744 10311
rect 19844 10451 19932 10504
rect 19844 10311 19873 10451
rect 19919 10311 19932 10451
rect 19844 10260 19932 10311
rect 20328 10451 20416 10504
rect 20328 10311 20341 10451
rect 20387 10311 20416 10451
rect 20328 10260 20416 10311
rect 20516 10451 20604 10504
rect 20516 10311 20545 10451
rect 20591 10311 20604 10451
rect 20516 10260 20604 10311
rect 21000 10451 21088 10504
rect 21000 10311 21013 10451
rect 21059 10311 21088 10451
rect 21000 10260 21088 10311
rect 21188 10451 21276 10504
rect 21188 10311 21217 10451
rect 21263 10311 21276 10451
rect 21188 10260 21276 10311
rect 21672 10451 21760 10504
rect 21672 10311 21685 10451
rect 21731 10311 21760 10451
rect 21672 10260 21760 10311
rect 21860 10451 21948 10504
rect 21860 10311 21889 10451
rect 21935 10311 21948 10451
rect 21860 10260 21948 10311
rect 1604 10065 1692 10124
rect 1604 9925 1617 10065
rect 1663 9925 1692 10065
rect 1604 9880 1692 9925
rect 1892 10065 1980 10124
rect 1892 9925 1921 10065
rect 1967 9925 1980 10065
rect 1892 9880 1980 9925
rect 2052 10065 2140 10124
rect 2052 9925 2065 10065
rect 2111 9925 2140 10065
rect 2052 9880 2140 9925
rect 2340 10065 2428 10124
rect 2340 9925 2369 10065
rect 2415 9925 2428 10065
rect 2340 9880 2428 9925
rect 2500 10065 2588 10124
rect 2500 9925 2513 10065
rect 2559 9925 2588 10065
rect 2500 9880 2588 9925
rect 2788 10065 2876 10124
rect 2788 9925 2817 10065
rect 2863 9925 2876 10065
rect 2788 9880 2876 9925
rect 2948 10065 3036 10124
rect 2948 9925 2961 10065
rect 3007 9925 3036 10065
rect 2948 9880 3036 9925
rect 3236 10065 3324 10124
rect 3236 9925 3265 10065
rect 3311 9925 3324 10065
rect 3236 9880 3324 9925
rect 3396 10065 3484 10124
rect 3396 9925 3409 10065
rect 3455 9925 3484 10065
rect 3396 9880 3484 9925
rect 3684 10065 3772 10124
rect 3684 9925 3713 10065
rect 3759 9925 3772 10065
rect 3684 9880 3772 9925
rect 4088 10073 4176 10124
rect 4088 9933 4101 10073
rect 4147 9933 4176 10073
rect 4088 9880 4176 9933
rect 4276 10073 4364 10124
rect 4276 9933 4305 10073
rect 4351 9933 4364 10073
rect 4276 9880 4364 9933
rect 4760 10073 4848 10124
rect 4760 9933 4773 10073
rect 4819 9933 4848 10073
rect 4760 9880 4848 9933
rect 4948 10073 5036 10124
rect 4948 9933 4977 10073
rect 5023 9933 5036 10073
rect 4948 9880 5036 9933
rect 5768 10073 5856 10124
rect 5768 9933 5781 10073
rect 5827 9933 5856 10073
rect 5768 9880 5856 9933
rect 5956 10073 6044 10124
rect 5956 9933 5985 10073
rect 6031 9933 6044 10073
rect 5956 9880 6044 9933
rect 6440 10073 6528 10124
rect 6440 9933 6453 10073
rect 6499 9933 6528 10073
rect 6440 9880 6528 9933
rect 6628 10073 6716 10124
rect 6628 9933 6657 10073
rect 6703 9933 6716 10073
rect 6628 9880 6716 9933
rect 7112 10073 7200 10124
rect 7112 9933 7125 10073
rect 7171 9933 7200 10073
rect 7112 9880 7200 9933
rect 7300 10073 7388 10124
rect 7300 9933 7329 10073
rect 7375 9933 7388 10073
rect 7300 9880 7388 9933
rect 7784 10073 7872 10124
rect 7784 9933 7797 10073
rect 7843 9933 7872 10073
rect 7784 9880 7872 9933
rect 7972 10073 8060 10124
rect 7972 9933 8001 10073
rect 8047 9933 8060 10073
rect 7972 9880 8060 9933
rect 8456 10073 8544 10124
rect 8456 9933 8469 10073
rect 8515 9933 8544 10073
rect 8456 9880 8544 9933
rect 8644 10073 8732 10124
rect 8644 9933 8673 10073
rect 8719 9933 8732 10073
rect 8644 9880 8732 9933
rect 9128 10073 9216 10124
rect 9128 9933 9141 10073
rect 9187 9933 9216 10073
rect 9128 9880 9216 9933
rect 9316 10073 9404 10124
rect 9316 9933 9345 10073
rect 9391 9933 9404 10073
rect 9316 9880 9404 9933
rect 9800 10073 9888 10124
rect 9800 9933 9813 10073
rect 9859 9933 9888 10073
rect 9800 9880 9888 9933
rect 9988 10073 10076 10124
rect 9988 9933 10017 10073
rect 10063 9933 10076 10073
rect 9988 9880 10076 9933
rect 10472 10073 10560 10124
rect 10472 9933 10485 10073
rect 10531 9933 10560 10073
rect 10472 9880 10560 9933
rect 10660 10073 10748 10124
rect 10660 9933 10689 10073
rect 10735 9933 10748 10073
rect 10660 9880 10748 9933
rect 10900 10065 10988 10124
rect 10900 9925 10913 10065
rect 10959 9925 10988 10065
rect 10900 9880 10988 9925
rect 11188 10065 11276 10124
rect 11188 9925 11217 10065
rect 11263 9925 11276 10065
rect 11188 9880 11276 9925
rect 11368 10073 11456 10124
rect 11368 9933 11381 10073
rect 11427 9933 11456 10073
rect 11368 9880 11456 9933
rect 11556 10073 11644 10124
rect 11556 9933 11585 10073
rect 11631 9933 11644 10073
rect 11556 9880 11644 9933
rect 12040 10073 12128 10124
rect 12040 9933 12053 10073
rect 12099 9933 12128 10073
rect 12040 9880 12128 9933
rect 12228 10073 12316 10124
rect 12228 9933 12257 10073
rect 12303 9933 12316 10073
rect 12228 9880 12316 9933
rect 12712 10073 12800 10124
rect 12712 9933 12725 10073
rect 12771 9933 12800 10073
rect 12712 9880 12800 9933
rect 12900 10073 12988 10124
rect 12900 9933 12929 10073
rect 12975 9933 12988 10073
rect 12900 9880 12988 9933
rect 13608 10073 13696 10124
rect 13608 9933 13621 10073
rect 13667 9933 13696 10073
rect 13608 9880 13696 9933
rect 13796 10073 13884 10124
rect 13796 9933 13825 10073
rect 13871 9933 13884 10073
rect 13796 9880 13884 9933
rect 14280 10073 14368 10124
rect 14280 9933 14293 10073
rect 14339 9933 14368 10073
rect 14280 9880 14368 9933
rect 14468 10073 14556 10124
rect 14468 9933 14497 10073
rect 14543 9933 14556 10073
rect 14468 9880 14556 9933
rect 14952 10073 15040 10124
rect 14952 9933 14965 10073
rect 15011 9933 15040 10073
rect 14952 9880 15040 9933
rect 15140 10073 15228 10124
rect 15140 9933 15169 10073
rect 15215 9933 15228 10073
rect 15140 9880 15228 9933
rect 15624 10073 15712 10124
rect 15624 9933 15637 10073
rect 15683 9933 15712 10073
rect 15624 9880 15712 9933
rect 15812 10073 15900 10124
rect 15812 9933 15841 10073
rect 15887 9933 15900 10073
rect 15812 9880 15900 9933
rect 16296 10073 16384 10124
rect 16296 9933 16309 10073
rect 16355 9933 16384 10073
rect 16296 9880 16384 9933
rect 16484 10073 16572 10124
rect 16484 9933 16513 10073
rect 16559 9933 16572 10073
rect 16484 9880 16572 9933
rect 16968 10073 17056 10124
rect 16968 9933 16981 10073
rect 17027 9933 17056 10073
rect 16968 9880 17056 9933
rect 17156 10073 17244 10124
rect 17156 9933 17185 10073
rect 17231 9933 17244 10073
rect 17156 9880 17244 9933
rect 17700 10073 17788 10124
rect 17700 9933 17713 10073
rect 17759 9933 17788 10073
rect 17700 9880 17788 9933
rect 17888 10073 17976 10124
rect 17888 9933 17917 10073
rect 17963 9933 17976 10073
rect 17888 9880 17976 9933
rect 18312 10073 18400 10124
rect 18312 9933 18325 10073
rect 18371 9933 18400 10073
rect 18312 9880 18400 9933
rect 18500 10073 18588 10124
rect 18500 9933 18529 10073
rect 18575 9933 18588 10073
rect 18500 9880 18588 9933
rect 18984 10073 19072 10124
rect 18984 9933 18997 10073
rect 19043 9933 19072 10073
rect 18984 9880 19072 9933
rect 19172 10073 19260 10124
rect 19172 9933 19201 10073
rect 19247 9933 19260 10073
rect 19172 9880 19260 9933
rect 19656 10073 19744 10124
rect 19656 9933 19669 10073
rect 19715 9933 19744 10073
rect 19656 9880 19744 9933
rect 19844 10073 19932 10124
rect 19844 9933 19873 10073
rect 19919 9933 19932 10073
rect 19844 9880 19932 9933
rect 20328 10073 20416 10124
rect 20328 9933 20341 10073
rect 20387 9933 20416 10073
rect 20328 9880 20416 9933
rect 20516 10073 20604 10124
rect 20516 9933 20545 10073
rect 20591 9933 20604 10073
rect 20516 9880 20604 9933
rect 20756 10065 20844 10124
rect 20756 9925 20769 10065
rect 20815 9925 20844 10065
rect 20756 9880 20844 9925
rect 21044 10065 21132 10124
rect 21044 9925 21073 10065
rect 21119 9925 21132 10065
rect 21044 9880 21132 9925
rect 21560 10073 21648 10124
rect 21560 9933 21573 10073
rect 21619 9933 21648 10073
rect 21560 9880 21648 9933
rect 21748 10073 21836 10124
rect 21748 9933 21777 10073
rect 21823 9933 21836 10073
rect 21748 9880 21836 9933
rect 21988 10065 22076 10124
rect 21988 9925 22001 10065
rect 22047 9925 22076 10065
rect 21988 9880 22076 9925
rect 22276 10065 22364 10124
rect 22276 9925 22305 10065
rect 22351 9925 22364 10065
rect 22276 9880 22364 9925
rect 1604 8891 1692 8936
rect 1604 8751 1617 8891
rect 1663 8751 1692 8891
rect 1604 8692 1692 8751
rect 1892 8891 1980 8936
rect 1892 8751 1921 8891
rect 1967 8751 1980 8891
rect 1892 8692 1980 8751
rect 2052 8891 2140 8936
rect 2052 8751 2065 8891
rect 2111 8751 2140 8891
rect 2052 8692 2140 8751
rect 2340 8891 2428 8936
rect 2340 8751 2369 8891
rect 2415 8751 2428 8891
rect 2340 8692 2428 8751
rect 2500 8891 2588 8936
rect 2500 8751 2513 8891
rect 2559 8751 2588 8891
rect 2500 8692 2588 8751
rect 2788 8891 2876 8936
rect 2788 8751 2817 8891
rect 2863 8751 2876 8891
rect 2788 8692 2876 8751
rect 3304 8883 3392 8936
rect 3304 8743 3317 8883
rect 3363 8743 3392 8883
rect 3304 8692 3392 8743
rect 3492 8883 3580 8936
rect 3492 8743 3521 8883
rect 3567 8743 3580 8883
rect 3492 8692 3580 8743
rect 3976 8883 4064 8936
rect 3976 8743 3989 8883
rect 4035 8743 4064 8883
rect 3976 8692 4064 8743
rect 4164 8883 4252 8936
rect 4164 8743 4193 8883
rect 4239 8743 4252 8883
rect 4164 8692 4252 8743
rect 4648 8883 4736 8936
rect 4648 8743 4661 8883
rect 4707 8743 4736 8883
rect 4648 8692 4736 8743
rect 4836 8883 4924 8936
rect 4836 8743 4865 8883
rect 4911 8743 4924 8883
rect 4836 8692 4924 8743
rect 5320 8883 5408 8936
rect 5320 8743 5333 8883
rect 5379 8743 5408 8883
rect 5320 8692 5408 8743
rect 5508 8883 5596 8936
rect 5508 8743 5537 8883
rect 5583 8743 5596 8883
rect 5508 8692 5596 8743
rect 5992 8883 6080 8936
rect 5992 8743 6005 8883
rect 6051 8743 6080 8883
rect 5992 8692 6080 8743
rect 6180 8883 6268 8936
rect 6180 8743 6209 8883
rect 6255 8743 6268 8883
rect 6180 8692 6268 8743
rect 6664 8883 6752 8936
rect 6664 8743 6677 8883
rect 6723 8743 6752 8883
rect 6664 8692 6752 8743
rect 6852 8883 6940 8936
rect 6852 8743 6881 8883
rect 6927 8743 6940 8883
rect 6852 8692 6940 8743
rect 7336 8883 7424 8936
rect 7336 8743 7349 8883
rect 7395 8743 7424 8883
rect 7336 8692 7424 8743
rect 7524 8883 7612 8936
rect 7524 8743 7553 8883
rect 7599 8743 7612 8883
rect 7524 8692 7612 8743
rect 8120 8883 8208 8936
rect 8120 8743 8133 8883
rect 8179 8743 8208 8883
rect 8120 8692 8208 8743
rect 8308 8883 8396 8936
rect 8308 8743 8337 8883
rect 8383 8743 8396 8883
rect 8308 8692 8396 8743
rect 8792 8883 8880 8936
rect 8792 8743 8805 8883
rect 8851 8743 8880 8883
rect 8792 8692 8880 8743
rect 8980 8883 9068 8936
rect 8980 8743 9009 8883
rect 9055 8743 9068 8883
rect 8980 8692 9068 8743
rect 9556 8891 9644 8936
rect 9556 8751 9569 8891
rect 9615 8751 9644 8891
rect 9556 8692 9644 8751
rect 9844 8891 9932 8936
rect 9844 8751 9873 8891
rect 9919 8751 9932 8891
rect 9844 8692 9932 8751
rect 10248 8883 10336 8936
rect 10248 8743 10261 8883
rect 10307 8743 10336 8883
rect 10248 8692 10336 8743
rect 10436 8883 10524 8936
rect 10436 8743 10465 8883
rect 10511 8743 10524 8883
rect 10436 8692 10524 8743
rect 10920 8883 11008 8936
rect 10920 8743 10933 8883
rect 10979 8743 11008 8883
rect 10920 8692 11008 8743
rect 11108 8883 11196 8936
rect 11108 8743 11137 8883
rect 11183 8743 11196 8883
rect 11108 8692 11196 8743
rect 11592 8883 11680 8936
rect 11592 8743 11605 8883
rect 11651 8743 11680 8883
rect 11592 8692 11680 8743
rect 11780 8883 11868 8936
rect 11780 8743 11809 8883
rect 11855 8743 11868 8883
rect 11780 8692 11868 8743
rect 12264 8883 12352 8936
rect 12264 8743 12277 8883
rect 12323 8743 12352 8883
rect 12264 8692 12352 8743
rect 12452 8883 12540 8936
rect 12452 8743 12481 8883
rect 12527 8743 12540 8883
rect 12452 8692 12540 8743
rect 12936 8883 13024 8936
rect 12936 8743 12949 8883
rect 12995 8743 13024 8883
rect 12936 8692 13024 8743
rect 13124 8883 13212 8936
rect 13124 8743 13153 8883
rect 13199 8743 13212 8883
rect 13124 8692 13212 8743
rect 13608 8883 13696 8936
rect 13608 8743 13621 8883
rect 13667 8743 13696 8883
rect 13608 8692 13696 8743
rect 13796 8883 13884 8936
rect 13796 8743 13825 8883
rect 13871 8743 13884 8883
rect 13796 8692 13884 8743
rect 14280 8883 14368 8936
rect 14280 8743 14293 8883
rect 14339 8743 14368 8883
rect 14280 8692 14368 8743
rect 14468 8883 14556 8936
rect 14468 8743 14497 8883
rect 14543 8743 14556 8883
rect 14468 8692 14556 8743
rect 14952 8883 15040 8936
rect 14952 8743 14965 8883
rect 15011 8743 15040 8883
rect 14952 8692 15040 8743
rect 15140 8883 15228 8936
rect 15140 8743 15169 8883
rect 15215 8743 15228 8883
rect 15140 8692 15228 8743
rect 15624 8883 15712 8936
rect 15624 8743 15637 8883
rect 15683 8743 15712 8883
rect 15624 8692 15712 8743
rect 15812 8883 15900 8936
rect 15812 8743 15841 8883
rect 15887 8743 15900 8883
rect 15812 8692 15900 8743
rect 16296 8883 16384 8936
rect 16296 8743 16309 8883
rect 16355 8743 16384 8883
rect 16296 8692 16384 8743
rect 16484 8883 16572 8936
rect 16484 8743 16513 8883
rect 16559 8743 16572 8883
rect 16484 8692 16572 8743
rect 16724 8891 16812 8936
rect 16724 8751 16737 8891
rect 16783 8751 16812 8891
rect 16724 8692 16812 8751
rect 17012 8891 17100 8936
rect 17012 8751 17041 8891
rect 17087 8751 17100 8891
rect 17012 8692 17100 8751
rect 17640 8883 17728 8936
rect 17640 8743 17653 8883
rect 17699 8743 17728 8883
rect 17640 8692 17728 8743
rect 17828 8883 17916 8936
rect 17828 8743 17857 8883
rect 17903 8743 17916 8883
rect 17828 8692 17916 8743
rect 18312 8883 18400 8936
rect 18312 8743 18325 8883
rect 18371 8743 18400 8883
rect 18312 8692 18400 8743
rect 18500 8883 18588 8936
rect 18500 8743 18529 8883
rect 18575 8743 18588 8883
rect 18500 8692 18588 8743
rect 18984 8883 19072 8936
rect 18984 8743 18997 8883
rect 19043 8743 19072 8883
rect 18984 8692 19072 8743
rect 19172 8883 19260 8936
rect 19172 8743 19201 8883
rect 19247 8743 19260 8883
rect 19172 8692 19260 8743
rect 19656 8883 19744 8936
rect 19656 8743 19669 8883
rect 19715 8743 19744 8883
rect 19656 8692 19744 8743
rect 19844 8883 19932 8936
rect 19844 8743 19873 8883
rect 19919 8743 19932 8883
rect 19844 8692 19932 8743
rect 20328 8883 20416 8936
rect 20328 8743 20341 8883
rect 20387 8743 20416 8883
rect 20328 8692 20416 8743
rect 20516 8883 20604 8936
rect 20516 8743 20545 8883
rect 20591 8743 20604 8883
rect 20516 8692 20604 8743
rect 20756 8891 20844 8936
rect 20756 8751 20769 8891
rect 20815 8751 20844 8891
rect 20756 8692 20844 8751
rect 21044 8891 21132 8936
rect 21044 8751 21073 8891
rect 21119 8751 21132 8891
rect 21044 8692 21132 8751
rect 21204 8891 21292 8936
rect 21204 8751 21217 8891
rect 21263 8751 21292 8891
rect 21204 8692 21292 8751
rect 21492 8891 21580 8936
rect 21492 8751 21521 8891
rect 21567 8751 21580 8891
rect 21492 8692 21580 8751
rect 21652 8891 21740 8936
rect 21652 8751 21665 8891
rect 21711 8751 21740 8891
rect 21652 8692 21740 8751
rect 21940 8891 22028 8936
rect 21940 8751 21969 8891
rect 22015 8751 22028 8891
rect 21940 8692 22028 8751
rect 1604 8497 1692 8556
rect 1604 8357 1617 8497
rect 1663 8357 1692 8497
rect 1604 8312 1692 8357
rect 1892 8497 1980 8556
rect 1892 8357 1921 8497
rect 1967 8357 1980 8497
rect 1892 8312 1980 8357
rect 2052 8497 2140 8556
rect 2052 8357 2065 8497
rect 2111 8357 2140 8497
rect 2052 8312 2140 8357
rect 2340 8497 2428 8556
rect 2340 8357 2369 8497
rect 2415 8357 2428 8497
rect 2340 8312 2428 8357
rect 2804 8505 2892 8556
rect 2804 8365 2817 8505
rect 2863 8365 2892 8505
rect 2804 8312 2892 8365
rect 2992 8505 3080 8556
rect 2992 8365 3021 8505
rect 3067 8365 3080 8505
rect 2992 8312 3080 8365
rect 3416 8505 3504 8556
rect 3416 8365 3429 8505
rect 3475 8365 3504 8505
rect 3416 8312 3504 8365
rect 3604 8505 3692 8556
rect 3604 8365 3633 8505
rect 3679 8365 3692 8505
rect 3604 8312 3692 8365
rect 4088 8505 4176 8556
rect 4088 8365 4101 8505
rect 4147 8365 4176 8505
rect 4088 8312 4176 8365
rect 4276 8505 4364 8556
rect 4276 8365 4305 8505
rect 4351 8365 4364 8505
rect 4276 8312 4364 8365
rect 4760 8505 4848 8556
rect 4760 8365 4773 8505
rect 4819 8365 4848 8505
rect 4760 8312 4848 8365
rect 4948 8505 5036 8556
rect 4948 8365 4977 8505
rect 5023 8365 5036 8505
rect 4948 8312 5036 8365
rect 5768 8505 5856 8556
rect 5768 8365 5781 8505
rect 5827 8365 5856 8505
rect 5768 8312 5856 8365
rect 5956 8505 6044 8556
rect 5956 8365 5985 8505
rect 6031 8365 6044 8505
rect 5956 8312 6044 8365
rect 6440 8505 6528 8556
rect 6440 8365 6453 8505
rect 6499 8365 6528 8505
rect 6440 8312 6528 8365
rect 6628 8505 6716 8556
rect 6628 8365 6657 8505
rect 6703 8365 6716 8505
rect 6628 8312 6716 8365
rect 7112 8505 7200 8556
rect 7112 8365 7125 8505
rect 7171 8365 7200 8505
rect 7112 8312 7200 8365
rect 7300 8505 7388 8556
rect 7300 8365 7329 8505
rect 7375 8365 7388 8505
rect 7300 8312 7388 8365
rect 7784 8505 7872 8556
rect 7784 8365 7797 8505
rect 7843 8365 7872 8505
rect 7784 8312 7872 8365
rect 7972 8505 8060 8556
rect 7972 8365 8001 8505
rect 8047 8365 8060 8505
rect 7972 8312 8060 8365
rect 8456 8505 8544 8556
rect 8456 8365 8469 8505
rect 8515 8365 8544 8505
rect 8456 8312 8544 8365
rect 8644 8505 8732 8556
rect 8644 8365 8673 8505
rect 8719 8365 8732 8505
rect 8644 8312 8732 8365
rect 9128 8505 9216 8556
rect 9128 8365 9141 8505
rect 9187 8365 9216 8505
rect 9128 8312 9216 8365
rect 9316 8505 9404 8556
rect 9316 8365 9345 8505
rect 9391 8365 9404 8505
rect 9316 8312 9404 8365
rect 9800 8505 9888 8556
rect 9800 8365 9813 8505
rect 9859 8365 9888 8505
rect 9800 8312 9888 8365
rect 9988 8505 10076 8556
rect 9988 8365 10017 8505
rect 10063 8365 10076 8505
rect 9988 8312 10076 8365
rect 10472 8505 10560 8556
rect 10472 8365 10485 8505
rect 10531 8365 10560 8505
rect 10472 8312 10560 8365
rect 10660 8505 10748 8556
rect 10660 8365 10689 8505
rect 10735 8365 10748 8505
rect 10660 8312 10748 8365
rect 11204 8505 11292 8556
rect 11204 8365 11217 8505
rect 11263 8365 11292 8505
rect 11204 8312 11292 8365
rect 11392 8505 11480 8556
rect 11392 8365 11421 8505
rect 11467 8365 11480 8505
rect 11392 8312 11480 8365
rect 11572 8497 11660 8556
rect 11572 8357 11585 8497
rect 11631 8357 11660 8497
rect 11572 8312 11660 8357
rect 11860 8497 11948 8556
rect 11860 8357 11889 8497
rect 11935 8357 11948 8497
rect 11860 8312 11948 8357
rect 12040 8505 12128 8556
rect 12040 8365 12053 8505
rect 12099 8365 12128 8505
rect 12040 8312 12128 8365
rect 12228 8505 12316 8556
rect 12228 8365 12257 8505
rect 12303 8365 12316 8505
rect 12228 8312 12316 8365
rect 12712 8505 12800 8556
rect 12712 8365 12725 8505
rect 12771 8365 12800 8505
rect 12712 8312 12800 8365
rect 12900 8505 12988 8556
rect 12900 8365 12929 8505
rect 12975 8365 12988 8505
rect 12900 8312 12988 8365
rect 13608 8505 13696 8556
rect 13608 8365 13621 8505
rect 13667 8365 13696 8505
rect 13608 8312 13696 8365
rect 13796 8505 13884 8556
rect 13796 8365 13825 8505
rect 13871 8365 13884 8505
rect 13796 8312 13884 8365
rect 14280 8505 14368 8556
rect 14280 8365 14293 8505
rect 14339 8365 14368 8505
rect 14280 8312 14368 8365
rect 14468 8505 14556 8556
rect 14468 8365 14497 8505
rect 14543 8365 14556 8505
rect 14468 8312 14556 8365
rect 14952 8505 15040 8556
rect 14952 8365 14965 8505
rect 15011 8365 15040 8505
rect 14952 8312 15040 8365
rect 15140 8505 15228 8556
rect 15140 8365 15169 8505
rect 15215 8365 15228 8505
rect 15140 8312 15228 8365
rect 15624 8505 15712 8556
rect 15624 8365 15637 8505
rect 15683 8365 15712 8505
rect 15624 8312 15712 8365
rect 15812 8505 15900 8556
rect 15812 8365 15841 8505
rect 15887 8365 15900 8505
rect 15812 8312 15900 8365
rect 16296 8505 16384 8556
rect 16296 8365 16309 8505
rect 16355 8365 16384 8505
rect 16296 8312 16384 8365
rect 16484 8505 16572 8556
rect 16484 8365 16513 8505
rect 16559 8365 16572 8505
rect 16484 8312 16572 8365
rect 16968 8505 17056 8556
rect 16968 8365 16981 8505
rect 17027 8365 17056 8505
rect 16968 8312 17056 8365
rect 17156 8505 17244 8556
rect 17156 8365 17185 8505
rect 17231 8365 17244 8505
rect 17156 8312 17244 8365
rect 17640 8505 17728 8556
rect 17640 8365 17653 8505
rect 17699 8365 17728 8505
rect 17640 8312 17728 8365
rect 17828 8505 17916 8556
rect 17828 8365 17857 8505
rect 17903 8365 17916 8505
rect 17828 8312 17916 8365
rect 18312 8505 18400 8556
rect 18312 8365 18325 8505
rect 18371 8365 18400 8505
rect 18312 8312 18400 8365
rect 18500 8505 18588 8556
rect 18500 8365 18529 8505
rect 18575 8365 18588 8505
rect 18500 8312 18588 8365
rect 18984 8505 19072 8556
rect 18984 8365 18997 8505
rect 19043 8365 19072 8505
rect 18984 8312 19072 8365
rect 19172 8505 19260 8556
rect 19172 8365 19201 8505
rect 19247 8365 19260 8505
rect 19172 8312 19260 8365
rect 19656 8505 19744 8556
rect 19656 8365 19669 8505
rect 19715 8365 19744 8505
rect 19656 8312 19744 8365
rect 19844 8505 19932 8556
rect 19844 8365 19873 8505
rect 19919 8365 19932 8505
rect 19844 8312 19932 8365
rect 20388 8505 20476 8556
rect 20388 8365 20401 8505
rect 20447 8365 20476 8505
rect 20388 8312 20476 8365
rect 20576 8505 20664 8556
rect 20576 8365 20605 8505
rect 20651 8365 20664 8505
rect 20576 8312 20664 8365
rect 20756 8497 20844 8556
rect 20756 8357 20769 8497
rect 20815 8357 20844 8497
rect 20756 8312 20844 8357
rect 21044 8497 21132 8556
rect 21044 8357 21073 8497
rect 21119 8357 21132 8497
rect 21044 8312 21132 8357
rect 21428 8497 21516 8556
rect 21428 8357 21441 8497
rect 21487 8357 21516 8497
rect 21428 8312 21516 8357
rect 21716 8497 21804 8556
rect 21716 8357 21745 8497
rect 21791 8357 21804 8497
rect 21716 8312 21804 8357
rect 21876 8497 21964 8556
rect 21876 8357 21889 8497
rect 21935 8357 21964 8497
rect 21876 8312 21964 8357
rect 22164 8497 22252 8556
rect 22164 8357 22193 8497
rect 22239 8357 22252 8497
rect 22164 8312 22252 8357
rect 2020 7315 2108 7368
rect 2020 7175 2033 7315
rect 2079 7175 2108 7315
rect 2020 7124 2108 7175
rect 2208 7315 2296 7368
rect 2208 7175 2237 7315
rect 2283 7175 2296 7315
rect 2208 7124 2296 7175
rect 2632 7315 2720 7368
rect 2632 7175 2645 7315
rect 2691 7175 2720 7315
rect 2632 7124 2720 7175
rect 2820 7315 2908 7368
rect 2820 7175 2849 7315
rect 2895 7175 2908 7315
rect 2820 7124 2908 7175
rect 3304 7315 3392 7368
rect 3304 7175 3317 7315
rect 3363 7175 3392 7315
rect 3304 7124 3392 7175
rect 3492 7315 3580 7368
rect 3492 7175 3521 7315
rect 3567 7175 3580 7315
rect 3492 7124 3580 7175
rect 3976 7315 4064 7368
rect 3976 7175 3989 7315
rect 4035 7175 4064 7315
rect 3976 7124 4064 7175
rect 4164 7315 4252 7368
rect 4164 7175 4193 7315
rect 4239 7175 4252 7315
rect 4164 7124 4252 7175
rect 4648 7315 4736 7368
rect 4648 7175 4661 7315
rect 4707 7175 4736 7315
rect 4648 7124 4736 7175
rect 4836 7315 4924 7368
rect 4836 7175 4865 7315
rect 4911 7175 4924 7315
rect 4836 7124 4924 7175
rect 5320 7315 5408 7368
rect 5320 7175 5333 7315
rect 5379 7175 5408 7315
rect 5320 7124 5408 7175
rect 5508 7315 5596 7368
rect 5508 7175 5537 7315
rect 5583 7175 5596 7315
rect 5508 7124 5596 7175
rect 5992 7315 6080 7368
rect 5992 7175 6005 7315
rect 6051 7175 6080 7315
rect 5992 7124 6080 7175
rect 6180 7315 6268 7368
rect 6180 7175 6209 7315
rect 6255 7175 6268 7315
rect 6180 7124 6268 7175
rect 6664 7315 6752 7368
rect 6664 7175 6677 7315
rect 6723 7175 6752 7315
rect 6664 7124 6752 7175
rect 6852 7315 6940 7368
rect 6852 7175 6881 7315
rect 6927 7175 6940 7315
rect 6852 7124 6940 7175
rect 7336 7315 7424 7368
rect 7336 7175 7349 7315
rect 7395 7175 7424 7315
rect 7336 7124 7424 7175
rect 7524 7315 7612 7368
rect 7524 7175 7553 7315
rect 7599 7175 7612 7315
rect 7524 7124 7612 7175
rect 8120 7315 8208 7368
rect 8120 7175 8133 7315
rect 8179 7175 8208 7315
rect 8120 7124 8208 7175
rect 8308 7315 8396 7368
rect 8308 7175 8337 7315
rect 8383 7175 8396 7315
rect 8308 7124 8396 7175
rect 8792 7315 8880 7368
rect 8792 7175 8805 7315
rect 8851 7175 8880 7315
rect 8792 7124 8880 7175
rect 8980 7315 9068 7368
rect 8980 7175 9009 7315
rect 9055 7175 9068 7315
rect 8980 7124 9068 7175
rect 9800 7315 9888 7368
rect 9800 7175 9813 7315
rect 9859 7175 9888 7315
rect 9800 7124 9888 7175
rect 9988 7315 10076 7368
rect 9988 7175 10017 7315
rect 10063 7175 10076 7315
rect 9988 7124 10076 7175
rect 10472 7315 10560 7368
rect 10472 7175 10485 7315
rect 10531 7175 10560 7315
rect 10472 7124 10560 7175
rect 10660 7315 10748 7368
rect 10660 7175 10689 7315
rect 10735 7175 10748 7315
rect 10660 7124 10748 7175
rect 11204 7315 11292 7368
rect 11204 7175 11217 7315
rect 11263 7175 11292 7315
rect 11204 7124 11292 7175
rect 11392 7315 11480 7368
rect 11392 7175 11421 7315
rect 11467 7175 11480 7315
rect 11392 7124 11480 7175
rect 11816 7315 11904 7368
rect 11816 7175 11829 7315
rect 11875 7175 11904 7315
rect 11816 7124 11904 7175
rect 12004 7315 12092 7368
rect 12004 7175 12033 7315
rect 12079 7175 12092 7315
rect 12004 7124 12092 7175
rect 12488 7315 12576 7368
rect 12488 7175 12501 7315
rect 12547 7175 12576 7315
rect 12488 7124 12576 7175
rect 12676 7315 12764 7368
rect 12676 7175 12705 7315
rect 12751 7175 12764 7315
rect 12676 7124 12764 7175
rect 13160 7315 13248 7368
rect 13160 7175 13173 7315
rect 13219 7175 13248 7315
rect 13160 7124 13248 7175
rect 13348 7315 13436 7368
rect 13348 7175 13377 7315
rect 13423 7175 13436 7315
rect 13348 7124 13436 7175
rect 13832 7315 13920 7368
rect 13832 7175 13845 7315
rect 13891 7175 13920 7315
rect 13832 7124 13920 7175
rect 14020 7315 14108 7368
rect 14020 7175 14049 7315
rect 14095 7175 14108 7315
rect 14020 7124 14108 7175
rect 14504 7315 14592 7368
rect 14504 7175 14517 7315
rect 14563 7175 14592 7315
rect 14504 7124 14592 7175
rect 14692 7315 14780 7368
rect 14692 7175 14721 7315
rect 14767 7175 14780 7315
rect 14692 7124 14780 7175
rect 15176 7315 15264 7368
rect 15176 7175 15189 7315
rect 15235 7175 15264 7315
rect 15176 7124 15264 7175
rect 15364 7315 15452 7368
rect 15364 7175 15393 7315
rect 15439 7175 15452 7315
rect 15364 7124 15452 7175
rect 15848 7315 15936 7368
rect 15848 7175 15861 7315
rect 15907 7175 15936 7315
rect 15848 7124 15936 7175
rect 16036 7315 16124 7368
rect 16036 7175 16065 7315
rect 16111 7175 16124 7315
rect 16036 7124 16124 7175
rect 16520 7315 16608 7368
rect 16520 7175 16533 7315
rect 16579 7175 16608 7315
rect 16520 7124 16608 7175
rect 16708 7315 16796 7368
rect 16708 7175 16737 7315
rect 16783 7175 16796 7315
rect 16708 7124 16796 7175
rect 17640 7315 17728 7368
rect 17640 7175 17653 7315
rect 17699 7175 17728 7315
rect 17640 7124 17728 7175
rect 17828 7315 17916 7368
rect 17828 7175 17857 7315
rect 17903 7175 17916 7315
rect 17828 7124 17916 7175
rect 18312 7315 18400 7368
rect 18312 7175 18325 7315
rect 18371 7175 18400 7315
rect 18312 7124 18400 7175
rect 18500 7315 18588 7368
rect 18500 7175 18529 7315
rect 18575 7175 18588 7315
rect 18500 7124 18588 7175
rect 18984 7315 19072 7368
rect 18984 7175 18997 7315
rect 19043 7175 19072 7315
rect 18984 7124 19072 7175
rect 19172 7315 19260 7368
rect 19172 7175 19201 7315
rect 19247 7175 19260 7315
rect 19172 7124 19260 7175
rect 19656 7315 19744 7368
rect 19656 7175 19669 7315
rect 19715 7175 19744 7315
rect 19656 7124 19744 7175
rect 19844 7315 19932 7368
rect 19844 7175 19873 7315
rect 19919 7175 19932 7315
rect 19844 7124 19932 7175
rect 20328 7315 20416 7368
rect 20328 7175 20341 7315
rect 20387 7175 20416 7315
rect 20328 7124 20416 7175
rect 20516 7315 20604 7368
rect 20516 7175 20545 7315
rect 20591 7175 20604 7315
rect 20516 7124 20604 7175
rect 21000 7315 21088 7368
rect 21000 7175 21013 7315
rect 21059 7175 21088 7315
rect 21000 7124 21088 7175
rect 21188 7315 21276 7368
rect 21188 7175 21217 7315
rect 21263 7175 21276 7315
rect 21188 7124 21276 7175
rect 21428 7323 21516 7368
rect 21428 7183 21441 7323
rect 21487 7183 21516 7323
rect 21428 7124 21516 7183
rect 21716 7323 21804 7368
rect 21716 7183 21745 7323
rect 21791 7183 21804 7323
rect 21716 7124 21804 7183
rect 21876 7323 21964 7368
rect 21876 7183 21889 7323
rect 21935 7183 21964 7323
rect 21876 7124 21964 7183
rect 22164 7323 22252 7368
rect 22164 7183 22193 7323
rect 22239 7183 22252 7323
rect 22164 7124 22252 7183
rect 1604 6929 1692 6988
rect 1604 6789 1617 6929
rect 1663 6789 1692 6929
rect 1604 6744 1692 6789
rect 1892 6929 1980 6988
rect 1892 6789 1921 6929
rect 1967 6789 1980 6929
rect 1892 6744 1980 6789
rect 2072 6937 2160 6988
rect 2072 6797 2085 6937
rect 2131 6797 2160 6937
rect 2072 6744 2160 6797
rect 2260 6937 2348 6988
rect 2260 6797 2289 6937
rect 2335 6797 2348 6937
rect 2260 6744 2348 6797
rect 2744 6937 2832 6988
rect 2744 6797 2757 6937
rect 2803 6797 2832 6937
rect 2744 6744 2832 6797
rect 2932 6937 3020 6988
rect 2932 6797 2961 6937
rect 3007 6797 3020 6937
rect 2932 6744 3020 6797
rect 3416 6937 3504 6988
rect 3416 6797 3429 6937
rect 3475 6797 3504 6937
rect 3416 6744 3504 6797
rect 3604 6937 3692 6988
rect 3604 6797 3633 6937
rect 3679 6797 3692 6937
rect 3604 6744 3692 6797
rect 4088 6937 4176 6988
rect 4088 6797 4101 6937
rect 4147 6797 4176 6937
rect 4088 6744 4176 6797
rect 4276 6937 4364 6988
rect 4276 6797 4305 6937
rect 4351 6797 4364 6937
rect 4276 6744 4364 6797
rect 4760 6937 4848 6988
rect 4760 6797 4773 6937
rect 4819 6797 4848 6937
rect 4760 6744 4848 6797
rect 4948 6937 5036 6988
rect 4948 6797 4977 6937
rect 5023 6797 5036 6937
rect 4948 6744 5036 6797
rect 5656 6937 5744 6988
rect 5656 6797 5669 6937
rect 5715 6797 5744 6937
rect 5656 6744 5744 6797
rect 5844 6937 5932 6988
rect 5844 6797 5873 6937
rect 5919 6797 5932 6937
rect 5844 6744 5932 6797
rect 6328 6937 6416 6988
rect 6328 6797 6341 6937
rect 6387 6797 6416 6937
rect 6328 6744 6416 6797
rect 6516 6937 6604 6988
rect 6516 6797 6545 6937
rect 6591 6797 6604 6937
rect 6516 6744 6604 6797
rect 7000 6937 7088 6988
rect 7000 6797 7013 6937
rect 7059 6797 7088 6937
rect 7000 6744 7088 6797
rect 7188 6937 7276 6988
rect 7188 6797 7217 6937
rect 7263 6797 7276 6937
rect 7188 6744 7276 6797
rect 7672 6937 7760 6988
rect 7672 6797 7685 6937
rect 7731 6797 7760 6937
rect 7672 6744 7760 6797
rect 7860 6937 7948 6988
rect 7860 6797 7889 6937
rect 7935 6797 7948 6937
rect 7860 6744 7948 6797
rect 8344 6937 8432 6988
rect 8344 6797 8357 6937
rect 8403 6797 8432 6937
rect 8344 6744 8432 6797
rect 8532 6937 8620 6988
rect 8532 6797 8561 6937
rect 8607 6797 8620 6937
rect 8532 6744 8620 6797
rect 9016 6937 9104 6988
rect 9016 6797 9029 6937
rect 9075 6797 9104 6937
rect 9016 6744 9104 6797
rect 9204 6937 9292 6988
rect 9204 6797 9233 6937
rect 9279 6797 9292 6937
rect 9204 6744 9292 6797
rect 9688 6937 9776 6988
rect 9688 6797 9701 6937
rect 9747 6797 9776 6937
rect 9688 6744 9776 6797
rect 9876 6937 9964 6988
rect 9876 6797 9905 6937
rect 9951 6797 9964 6937
rect 9876 6744 9964 6797
rect 10360 6937 10448 6988
rect 10360 6797 10373 6937
rect 10419 6797 10448 6937
rect 10360 6744 10448 6797
rect 10548 6937 10636 6988
rect 10548 6797 10577 6937
rect 10623 6797 10636 6937
rect 10548 6744 10636 6797
rect 11032 6937 11120 6988
rect 11032 6797 11045 6937
rect 11091 6797 11120 6937
rect 11032 6744 11120 6797
rect 11220 6937 11308 6988
rect 11220 6797 11249 6937
rect 11295 6797 11308 6937
rect 11220 6744 11308 6797
rect 11704 6937 11792 6988
rect 11704 6797 11717 6937
rect 11763 6797 11792 6937
rect 11704 6744 11792 6797
rect 11892 6937 11980 6988
rect 11892 6797 11921 6937
rect 11967 6797 11980 6937
rect 11892 6744 11980 6797
rect 12376 6937 12464 6988
rect 12376 6797 12389 6937
rect 12435 6797 12464 6937
rect 12376 6744 12464 6797
rect 12564 6937 12652 6988
rect 12564 6797 12593 6937
rect 12639 6797 12652 6937
rect 12564 6744 12652 6797
rect 12804 6929 12892 6988
rect 12804 6789 12817 6929
rect 12863 6789 12892 6929
rect 12804 6744 12892 6789
rect 13092 6929 13180 6988
rect 13092 6789 13121 6929
rect 13167 6789 13180 6929
rect 13092 6744 13180 6789
rect 13476 6929 13564 6988
rect 13476 6789 13489 6929
rect 13535 6789 13564 6929
rect 13476 6744 13564 6789
rect 13764 6929 13852 6988
rect 13764 6789 13793 6929
rect 13839 6789 13852 6929
rect 13764 6744 13852 6789
rect 14056 6937 14144 6988
rect 14056 6797 14069 6937
rect 14115 6797 14144 6937
rect 14056 6744 14144 6797
rect 14244 6937 14332 6988
rect 14244 6797 14273 6937
rect 14319 6797 14332 6937
rect 14244 6744 14332 6797
rect 14728 6937 14816 6988
rect 14728 6797 14741 6937
rect 14787 6797 14816 6937
rect 14728 6744 14816 6797
rect 14916 6937 15004 6988
rect 14916 6797 14945 6937
rect 14991 6797 15004 6937
rect 14916 6744 15004 6797
rect 15400 6937 15488 6988
rect 15400 6797 15413 6937
rect 15459 6797 15488 6937
rect 15400 6744 15488 6797
rect 15588 6937 15676 6988
rect 15588 6797 15617 6937
rect 15663 6797 15676 6937
rect 15588 6744 15676 6797
rect 16072 6937 16160 6988
rect 16072 6797 16085 6937
rect 16131 6797 16160 6937
rect 16072 6744 16160 6797
rect 16260 6937 16348 6988
rect 16260 6797 16289 6937
rect 16335 6797 16348 6937
rect 16260 6744 16348 6797
rect 16744 6937 16832 6988
rect 16744 6797 16757 6937
rect 16803 6797 16832 6937
rect 16744 6744 16832 6797
rect 16932 6937 17020 6988
rect 16932 6797 16961 6937
rect 17007 6797 17020 6937
rect 16932 6744 17020 6797
rect 17416 6937 17504 6988
rect 17416 6797 17429 6937
rect 17475 6797 17504 6937
rect 17416 6744 17504 6797
rect 17604 6937 17692 6988
rect 17604 6797 17633 6937
rect 17679 6797 17692 6937
rect 17604 6744 17692 6797
rect 18088 6937 18176 6988
rect 18088 6797 18101 6937
rect 18147 6797 18176 6937
rect 18088 6744 18176 6797
rect 18276 6937 18364 6988
rect 18276 6797 18305 6937
rect 18351 6797 18364 6937
rect 18276 6744 18364 6797
rect 18760 6937 18848 6988
rect 18760 6797 18773 6937
rect 18819 6797 18848 6937
rect 18760 6744 18848 6797
rect 18948 6937 19036 6988
rect 18948 6797 18977 6937
rect 19023 6797 19036 6937
rect 18948 6744 19036 6797
rect 19432 6937 19520 6988
rect 19432 6797 19445 6937
rect 19491 6797 19520 6937
rect 19432 6744 19520 6797
rect 19620 6937 19708 6988
rect 19620 6797 19649 6937
rect 19695 6797 19708 6937
rect 19620 6744 19708 6797
rect 20164 6937 20252 6988
rect 20164 6797 20177 6937
rect 20223 6797 20252 6937
rect 20164 6744 20252 6797
rect 20352 6937 20440 6988
rect 20352 6797 20381 6937
rect 20427 6797 20440 6937
rect 20352 6744 20440 6797
rect 20532 6929 20620 6988
rect 20532 6789 20545 6929
rect 20591 6789 20620 6929
rect 20532 6744 20620 6789
rect 20820 6929 20908 6988
rect 20820 6789 20849 6929
rect 20895 6789 20908 6929
rect 20820 6744 20908 6789
rect 21560 6937 21648 6988
rect 21560 6797 21573 6937
rect 21619 6797 21648 6937
rect 21560 6744 21648 6797
rect 21748 6937 21836 6988
rect 21748 6797 21777 6937
rect 21823 6797 21836 6937
rect 21748 6744 21836 6797
rect 21988 6929 22076 6988
rect 21988 6789 22001 6929
rect 22047 6789 22076 6929
rect 21988 6744 22076 6789
rect 22276 6929 22364 6988
rect 22276 6789 22305 6929
rect 22351 6789 22364 6929
rect 22276 6744 22364 6789
rect 1960 5747 2048 5800
rect 1960 5607 1973 5747
rect 2019 5607 2048 5747
rect 1960 5556 2048 5607
rect 2148 5747 2236 5800
rect 2148 5607 2177 5747
rect 2223 5607 2236 5747
rect 2148 5556 2236 5607
rect 2632 5747 2720 5800
rect 2632 5607 2645 5747
rect 2691 5607 2720 5747
rect 2632 5556 2720 5607
rect 2820 5747 2908 5800
rect 2820 5607 2849 5747
rect 2895 5607 2908 5747
rect 2820 5556 2908 5607
rect 3304 5747 3392 5800
rect 3304 5607 3317 5747
rect 3363 5607 3392 5747
rect 3304 5556 3392 5607
rect 3492 5747 3580 5800
rect 3492 5607 3521 5747
rect 3567 5607 3580 5747
rect 3492 5556 3580 5607
rect 3976 5747 4064 5800
rect 3976 5607 3989 5747
rect 4035 5607 4064 5747
rect 3976 5556 4064 5607
rect 4164 5747 4252 5800
rect 4164 5607 4193 5747
rect 4239 5607 4252 5747
rect 4164 5556 4252 5607
rect 4648 5747 4736 5800
rect 4648 5607 4661 5747
rect 4707 5607 4736 5747
rect 4648 5556 4736 5607
rect 4836 5747 4924 5800
rect 4836 5607 4865 5747
rect 4911 5607 4924 5747
rect 4836 5556 4924 5607
rect 5320 5747 5408 5800
rect 5320 5607 5333 5747
rect 5379 5607 5408 5747
rect 5320 5556 5408 5607
rect 5508 5747 5596 5800
rect 5508 5607 5537 5747
rect 5583 5607 5596 5747
rect 5508 5556 5596 5607
rect 5992 5747 6080 5800
rect 5992 5607 6005 5747
rect 6051 5607 6080 5747
rect 5992 5556 6080 5607
rect 6180 5747 6268 5800
rect 6180 5607 6209 5747
rect 6255 5607 6268 5747
rect 6180 5556 6268 5607
rect 6664 5747 6752 5800
rect 6664 5607 6677 5747
rect 6723 5607 6752 5747
rect 6664 5556 6752 5607
rect 6852 5747 6940 5800
rect 6852 5607 6881 5747
rect 6927 5607 6940 5747
rect 6852 5556 6940 5607
rect 7336 5747 7424 5800
rect 7336 5607 7349 5747
rect 7395 5607 7424 5747
rect 7336 5556 7424 5607
rect 7524 5747 7612 5800
rect 7524 5607 7553 5747
rect 7599 5607 7612 5747
rect 7524 5556 7612 5607
rect 8008 5747 8096 5800
rect 8008 5607 8021 5747
rect 8067 5607 8096 5747
rect 8008 5556 8096 5607
rect 8196 5747 8284 5800
rect 8196 5607 8225 5747
rect 8271 5607 8284 5747
rect 8196 5556 8284 5607
rect 8680 5747 8768 5800
rect 8680 5607 8693 5747
rect 8739 5607 8768 5747
rect 8680 5556 8768 5607
rect 8868 5747 8956 5800
rect 8868 5607 8897 5747
rect 8943 5607 8956 5747
rect 8868 5556 8956 5607
rect 9688 5747 9776 5800
rect 9688 5607 9701 5747
rect 9747 5607 9776 5747
rect 9688 5556 9776 5607
rect 9876 5747 9964 5800
rect 9876 5607 9905 5747
rect 9951 5607 9964 5747
rect 9876 5556 9964 5607
rect 10360 5747 10448 5800
rect 10360 5607 10373 5747
rect 10419 5607 10448 5747
rect 10360 5556 10448 5607
rect 10548 5747 10636 5800
rect 10548 5607 10577 5747
rect 10623 5607 10636 5747
rect 10548 5556 10636 5607
rect 11032 5747 11120 5800
rect 11032 5607 11045 5747
rect 11091 5607 11120 5747
rect 11032 5556 11120 5607
rect 11220 5747 11308 5800
rect 11220 5607 11249 5747
rect 11295 5607 11308 5747
rect 11220 5556 11308 5607
rect 11704 5747 11792 5800
rect 11704 5607 11717 5747
rect 11763 5607 11792 5747
rect 11704 5556 11792 5607
rect 11892 5747 11980 5800
rect 11892 5607 11921 5747
rect 11967 5607 11980 5747
rect 11892 5556 11980 5607
rect 12488 5747 12576 5800
rect 12488 5607 12501 5747
rect 12547 5607 12576 5747
rect 12488 5556 12576 5607
rect 12676 5747 12764 5800
rect 12676 5607 12705 5747
rect 12751 5607 12764 5747
rect 12676 5556 12764 5607
rect 13160 5747 13248 5800
rect 13160 5607 13173 5747
rect 13219 5607 13248 5747
rect 13160 5556 13248 5607
rect 13348 5747 13436 5800
rect 13348 5607 13377 5747
rect 13423 5607 13436 5747
rect 13348 5556 13436 5607
rect 13832 5747 13920 5800
rect 13832 5607 13845 5747
rect 13891 5607 13920 5747
rect 13832 5556 13920 5607
rect 14020 5747 14108 5800
rect 14020 5607 14049 5747
rect 14095 5607 14108 5747
rect 14020 5556 14108 5607
rect 14504 5747 14592 5800
rect 14504 5607 14517 5747
rect 14563 5607 14592 5747
rect 14504 5556 14592 5607
rect 14692 5747 14780 5800
rect 14692 5607 14721 5747
rect 14767 5607 14780 5747
rect 14692 5556 14780 5607
rect 15176 5747 15264 5800
rect 15176 5607 15189 5747
rect 15235 5607 15264 5747
rect 15176 5556 15264 5607
rect 15364 5747 15452 5800
rect 15364 5607 15393 5747
rect 15439 5607 15452 5747
rect 15364 5556 15452 5607
rect 15848 5747 15936 5800
rect 15848 5607 15861 5747
rect 15907 5607 15936 5747
rect 15848 5556 15936 5607
rect 16036 5747 16124 5800
rect 16036 5607 16065 5747
rect 16111 5607 16124 5747
rect 16036 5556 16124 5607
rect 16520 5747 16608 5800
rect 16520 5607 16533 5747
rect 16579 5607 16608 5747
rect 16520 5556 16608 5607
rect 16708 5747 16796 5800
rect 16708 5607 16737 5747
rect 16783 5607 16796 5747
rect 16708 5556 16796 5607
rect 17640 5747 17728 5800
rect 17640 5607 17653 5747
rect 17699 5607 17728 5747
rect 17640 5556 17728 5607
rect 17828 5747 17916 5800
rect 17828 5607 17857 5747
rect 17903 5607 17916 5747
rect 17828 5556 17916 5607
rect 18312 5747 18400 5800
rect 18312 5607 18325 5747
rect 18371 5607 18400 5747
rect 18312 5556 18400 5607
rect 18500 5747 18588 5800
rect 18500 5607 18529 5747
rect 18575 5607 18588 5747
rect 18500 5556 18588 5607
rect 18984 5747 19072 5800
rect 18984 5607 18997 5747
rect 19043 5607 19072 5747
rect 18984 5556 19072 5607
rect 19172 5747 19260 5800
rect 19172 5607 19201 5747
rect 19247 5607 19260 5747
rect 19172 5556 19260 5607
rect 19656 5747 19744 5800
rect 19656 5607 19669 5747
rect 19715 5607 19744 5747
rect 19656 5556 19744 5607
rect 19844 5747 19932 5800
rect 19844 5607 19873 5747
rect 19919 5607 19932 5747
rect 19844 5556 19932 5607
rect 20328 5747 20416 5800
rect 20328 5607 20341 5747
rect 20387 5607 20416 5747
rect 20328 5556 20416 5607
rect 20516 5747 20604 5800
rect 20516 5607 20545 5747
rect 20591 5607 20604 5747
rect 20516 5556 20604 5607
rect 21000 5747 21088 5800
rect 21000 5607 21013 5747
rect 21059 5607 21088 5747
rect 21000 5556 21088 5607
rect 21188 5747 21276 5800
rect 21188 5607 21217 5747
rect 21263 5607 21276 5747
rect 21188 5556 21276 5607
rect 21732 5747 21820 5800
rect 21732 5607 21745 5747
rect 21791 5607 21820 5747
rect 21732 5556 21820 5607
rect 21920 5747 22008 5800
rect 21920 5607 21949 5747
rect 21995 5607 22008 5747
rect 21920 5556 22008 5607
rect 1604 5361 1692 5420
rect 1604 5221 1617 5361
rect 1663 5221 1692 5361
rect 1604 5176 1692 5221
rect 1892 5361 1980 5420
rect 1892 5221 1921 5361
rect 1967 5221 1980 5361
rect 1892 5176 1980 5221
rect 2072 5369 2160 5420
rect 2072 5229 2085 5369
rect 2131 5229 2160 5369
rect 2072 5176 2160 5229
rect 2260 5369 2348 5420
rect 2260 5229 2289 5369
rect 2335 5229 2348 5369
rect 2260 5176 2348 5229
rect 2744 5369 2832 5420
rect 2744 5229 2757 5369
rect 2803 5229 2832 5369
rect 2744 5176 2832 5229
rect 2932 5369 3020 5420
rect 2932 5229 2961 5369
rect 3007 5229 3020 5369
rect 2932 5176 3020 5229
rect 3416 5369 3504 5420
rect 3416 5229 3429 5369
rect 3475 5229 3504 5369
rect 3416 5176 3504 5229
rect 3604 5369 3692 5420
rect 3604 5229 3633 5369
rect 3679 5229 3692 5369
rect 3604 5176 3692 5229
rect 4088 5369 4176 5420
rect 4088 5229 4101 5369
rect 4147 5229 4176 5369
rect 4088 5176 4176 5229
rect 4276 5369 4364 5420
rect 4276 5229 4305 5369
rect 4351 5229 4364 5369
rect 4276 5176 4364 5229
rect 4760 5369 4848 5420
rect 4760 5229 4773 5369
rect 4819 5229 4848 5369
rect 4760 5176 4848 5229
rect 4948 5369 5036 5420
rect 4948 5229 4977 5369
rect 5023 5229 5036 5369
rect 4948 5176 5036 5229
rect 5656 5369 5744 5420
rect 5656 5229 5669 5369
rect 5715 5229 5744 5369
rect 5656 5176 5744 5229
rect 5844 5369 5932 5420
rect 5844 5229 5873 5369
rect 5919 5229 5932 5369
rect 5844 5176 5932 5229
rect 6328 5369 6416 5420
rect 6328 5229 6341 5369
rect 6387 5229 6416 5369
rect 6328 5176 6416 5229
rect 6516 5369 6604 5420
rect 6516 5229 6545 5369
rect 6591 5229 6604 5369
rect 6516 5176 6604 5229
rect 7000 5369 7088 5420
rect 7000 5229 7013 5369
rect 7059 5229 7088 5369
rect 7000 5176 7088 5229
rect 7188 5369 7276 5420
rect 7188 5229 7217 5369
rect 7263 5229 7276 5369
rect 7188 5176 7276 5229
rect 7672 5369 7760 5420
rect 7672 5229 7685 5369
rect 7731 5229 7760 5369
rect 7672 5176 7760 5229
rect 7860 5369 7948 5420
rect 7860 5229 7889 5369
rect 7935 5229 7948 5369
rect 7860 5176 7948 5229
rect 8344 5369 8432 5420
rect 8344 5229 8357 5369
rect 8403 5229 8432 5369
rect 8344 5176 8432 5229
rect 8532 5369 8620 5420
rect 8532 5229 8561 5369
rect 8607 5229 8620 5369
rect 8532 5176 8620 5229
rect 9016 5369 9104 5420
rect 9016 5229 9029 5369
rect 9075 5229 9104 5369
rect 9016 5176 9104 5229
rect 9204 5369 9292 5420
rect 9204 5229 9233 5369
rect 9279 5229 9292 5369
rect 9204 5176 9292 5229
rect 9688 5369 9776 5420
rect 9688 5229 9701 5369
rect 9747 5229 9776 5369
rect 9688 5176 9776 5229
rect 9876 5369 9964 5420
rect 9876 5229 9905 5369
rect 9951 5229 9964 5369
rect 9876 5176 9964 5229
rect 10360 5369 10448 5420
rect 10360 5229 10373 5369
rect 10419 5229 10448 5369
rect 10360 5176 10448 5229
rect 10548 5369 10636 5420
rect 10548 5229 10577 5369
rect 10623 5229 10636 5369
rect 10548 5176 10636 5229
rect 10788 5361 10876 5420
rect 10788 5221 10801 5361
rect 10847 5221 10876 5361
rect 10788 5176 10876 5221
rect 11076 5361 11164 5420
rect 11076 5221 11105 5361
rect 11151 5221 11164 5361
rect 11076 5176 11164 5221
rect 11368 5369 11456 5420
rect 11368 5229 11381 5369
rect 11427 5229 11456 5369
rect 11368 5176 11456 5229
rect 11556 5369 11644 5420
rect 11556 5229 11585 5369
rect 11631 5229 11644 5369
rect 11556 5176 11644 5229
rect 12040 5369 12128 5420
rect 12040 5229 12053 5369
rect 12099 5229 12128 5369
rect 12040 5176 12128 5229
rect 12228 5369 12316 5420
rect 12228 5229 12257 5369
rect 12303 5229 12316 5369
rect 12228 5176 12316 5229
rect 12712 5369 12800 5420
rect 12712 5229 12725 5369
rect 12771 5229 12800 5369
rect 12712 5176 12800 5229
rect 12900 5369 12988 5420
rect 12900 5229 12929 5369
rect 12975 5229 12988 5369
rect 12900 5176 12988 5229
rect 13476 5361 13564 5420
rect 13476 5221 13489 5361
rect 13535 5221 13564 5361
rect 13476 5176 13564 5221
rect 13764 5361 13852 5420
rect 13764 5221 13793 5361
rect 13839 5221 13852 5361
rect 13764 5176 13852 5221
rect 13944 5369 14032 5420
rect 13944 5229 13957 5369
rect 14003 5229 14032 5369
rect 13944 5176 14032 5229
rect 14132 5369 14220 5420
rect 14132 5229 14161 5369
rect 14207 5229 14220 5369
rect 14132 5176 14220 5229
rect 14616 5369 14704 5420
rect 14616 5229 14629 5369
rect 14675 5229 14704 5369
rect 14616 5176 14704 5229
rect 14804 5369 14892 5420
rect 14804 5229 14833 5369
rect 14879 5229 14892 5369
rect 14804 5176 14892 5229
rect 15288 5369 15376 5420
rect 15288 5229 15301 5369
rect 15347 5229 15376 5369
rect 15288 5176 15376 5229
rect 15476 5369 15564 5420
rect 15476 5229 15505 5369
rect 15551 5229 15564 5369
rect 15476 5176 15564 5229
rect 15960 5369 16048 5420
rect 15960 5229 15973 5369
rect 16019 5229 16048 5369
rect 15960 5176 16048 5229
rect 16148 5369 16236 5420
rect 16148 5229 16177 5369
rect 16223 5229 16236 5369
rect 16148 5176 16236 5229
rect 16632 5369 16720 5420
rect 16632 5229 16645 5369
rect 16691 5229 16720 5369
rect 16632 5176 16720 5229
rect 16820 5369 16908 5420
rect 16820 5229 16849 5369
rect 16895 5229 16908 5369
rect 16820 5176 16908 5229
rect 17304 5369 17392 5420
rect 17304 5229 17317 5369
rect 17363 5229 17392 5369
rect 17304 5176 17392 5229
rect 17492 5369 17580 5420
rect 17492 5229 17521 5369
rect 17567 5229 17580 5369
rect 17492 5176 17580 5229
rect 17976 5369 18064 5420
rect 17976 5229 17989 5369
rect 18035 5229 18064 5369
rect 17976 5176 18064 5229
rect 18164 5369 18252 5420
rect 18164 5229 18193 5369
rect 18239 5229 18252 5369
rect 18164 5176 18252 5229
rect 18648 5369 18736 5420
rect 18648 5229 18661 5369
rect 18707 5229 18736 5369
rect 18648 5176 18736 5229
rect 18836 5369 18924 5420
rect 18836 5229 18865 5369
rect 18911 5229 18924 5369
rect 18836 5176 18924 5229
rect 19320 5369 19408 5420
rect 19320 5229 19333 5369
rect 19379 5229 19408 5369
rect 19320 5176 19408 5229
rect 19508 5369 19596 5420
rect 19508 5229 19537 5369
rect 19583 5229 19596 5369
rect 19508 5176 19596 5229
rect 19992 5369 20080 5420
rect 19992 5229 20005 5369
rect 20051 5229 20080 5369
rect 19992 5176 20080 5229
rect 20180 5369 20268 5420
rect 20180 5229 20209 5369
rect 20255 5229 20268 5369
rect 20180 5176 20268 5229
rect 20664 5369 20752 5420
rect 20664 5229 20677 5369
rect 20723 5229 20752 5369
rect 20664 5176 20752 5229
rect 20852 5369 20940 5420
rect 20852 5229 20881 5369
rect 20927 5229 20940 5369
rect 20852 5176 20940 5229
rect 21560 5369 21648 5420
rect 21560 5229 21573 5369
rect 21619 5229 21648 5369
rect 21560 5176 21648 5229
rect 21748 5369 21836 5420
rect 21748 5229 21777 5369
rect 21823 5229 21836 5369
rect 21748 5176 21836 5229
rect 21988 5361 22076 5420
rect 21988 5221 22001 5361
rect 22047 5221 22076 5361
rect 21988 5176 22076 5221
rect 22276 5361 22364 5420
rect 22276 5221 22305 5361
rect 22351 5221 22364 5361
rect 22276 5176 22364 5221
rect 1604 4187 1692 4232
rect 1604 4047 1617 4187
rect 1663 4047 1692 4187
rect 1604 3988 1692 4047
rect 1892 4187 1980 4232
rect 1892 4047 1921 4187
rect 1967 4047 1980 4187
rect 1892 3988 1980 4047
rect 2296 4179 2384 4232
rect 2296 4039 2309 4179
rect 2355 4039 2384 4179
rect 2296 3988 2384 4039
rect 2484 4179 2572 4232
rect 2484 4039 2513 4179
rect 2559 4039 2572 4179
rect 2484 3988 2572 4039
rect 2968 4179 3056 4232
rect 2968 4039 2981 4179
rect 3027 4039 3056 4179
rect 2968 3988 3056 4039
rect 3156 4179 3244 4232
rect 3156 4039 3185 4179
rect 3231 4039 3244 4179
rect 3156 3988 3244 4039
rect 3640 4179 3728 4232
rect 3640 4039 3653 4179
rect 3699 4039 3728 4179
rect 3640 3988 3728 4039
rect 3828 4179 3916 4232
rect 3828 4039 3857 4179
rect 3903 4039 3916 4179
rect 3828 3988 3916 4039
rect 4312 4179 4400 4232
rect 4312 4039 4325 4179
rect 4371 4039 4400 4179
rect 4312 3988 4400 4039
rect 4500 4179 4588 4232
rect 4500 4039 4529 4179
rect 4575 4039 4588 4179
rect 4500 3988 4588 4039
rect 4984 4179 5072 4232
rect 4984 4039 4997 4179
rect 5043 4039 5072 4179
rect 4984 3988 5072 4039
rect 5172 4179 5260 4232
rect 5172 4039 5201 4179
rect 5247 4039 5260 4179
rect 5172 3988 5260 4039
rect 5656 4179 5744 4232
rect 5656 4039 5669 4179
rect 5715 4039 5744 4179
rect 5656 3988 5744 4039
rect 5844 4179 5932 4232
rect 5844 4039 5873 4179
rect 5919 4039 5932 4179
rect 5844 3988 5932 4039
rect 6328 4179 6416 4232
rect 6328 4039 6341 4179
rect 6387 4039 6416 4179
rect 6328 3988 6416 4039
rect 6516 4179 6604 4232
rect 6516 4039 6545 4179
rect 6591 4039 6604 4179
rect 6516 3988 6604 4039
rect 7000 4179 7088 4232
rect 7000 4039 7013 4179
rect 7059 4039 7088 4179
rect 7000 3988 7088 4039
rect 7188 4179 7276 4232
rect 7188 4039 7217 4179
rect 7263 4039 7276 4179
rect 7188 3988 7276 4039
rect 7672 4179 7760 4232
rect 7672 4039 7685 4179
rect 7731 4039 7760 4179
rect 7672 3988 7760 4039
rect 7860 4179 7948 4232
rect 7860 4039 7889 4179
rect 7935 4039 7948 4179
rect 7860 3988 7948 4039
rect 8344 4179 8432 4232
rect 8344 4039 8357 4179
rect 8403 4039 8432 4179
rect 8344 3988 8432 4039
rect 8532 4179 8620 4232
rect 8532 4039 8561 4179
rect 8607 4039 8620 4179
rect 8532 3988 8620 4039
rect 8772 4187 8860 4232
rect 8772 4047 8785 4187
rect 8831 4047 8860 4187
rect 8772 3988 8860 4047
rect 9060 4187 9148 4232
rect 9060 4047 9089 4187
rect 9135 4047 9148 4187
rect 9060 3988 9148 4047
rect 9688 4179 9776 4232
rect 9688 4039 9701 4179
rect 9747 4039 9776 4179
rect 9688 3988 9776 4039
rect 9876 4179 9964 4232
rect 9876 4039 9905 4179
rect 9951 4039 9964 4179
rect 9876 3988 9964 4039
rect 10360 4179 10448 4232
rect 10360 4039 10373 4179
rect 10419 4039 10448 4179
rect 10360 3988 10448 4039
rect 10548 4179 10636 4232
rect 10548 4039 10577 4179
rect 10623 4039 10636 4179
rect 10548 3988 10636 4039
rect 11032 4179 11120 4232
rect 11032 4039 11045 4179
rect 11091 4039 11120 4179
rect 11032 3988 11120 4039
rect 11220 4179 11308 4232
rect 11220 4039 11249 4179
rect 11295 4039 11308 4179
rect 11220 3988 11308 4039
rect 11460 4187 11548 4232
rect 11460 4047 11473 4187
rect 11519 4047 11548 4187
rect 11460 3988 11548 4047
rect 11748 4187 11836 4232
rect 11748 4047 11777 4187
rect 11823 4047 11836 4187
rect 11748 3988 11836 4047
rect 12264 4179 12352 4232
rect 12264 4039 12277 4179
rect 12323 4039 12352 4179
rect 12264 3988 12352 4039
rect 12452 4179 12540 4232
rect 12452 4039 12481 4179
rect 12527 4039 12540 4179
rect 12452 3988 12540 4039
rect 12936 4179 13024 4232
rect 12936 4039 12949 4179
rect 12995 4039 13024 4179
rect 12936 3988 13024 4039
rect 13124 4179 13212 4232
rect 13124 4039 13153 4179
rect 13199 4039 13212 4179
rect 13124 3988 13212 4039
rect 13608 4179 13696 4232
rect 13608 4039 13621 4179
rect 13667 4039 13696 4179
rect 13608 3988 13696 4039
rect 13796 4179 13884 4232
rect 13796 4039 13825 4179
rect 13871 4039 13884 4179
rect 13796 3988 13884 4039
rect 14280 4179 14368 4232
rect 14280 4039 14293 4179
rect 14339 4039 14368 4179
rect 14280 3988 14368 4039
rect 14468 4179 14556 4232
rect 14468 4039 14497 4179
rect 14543 4039 14556 4179
rect 14468 3988 14556 4039
rect 14952 4179 15040 4232
rect 14952 4039 14965 4179
rect 15011 4039 15040 4179
rect 14952 3988 15040 4039
rect 15140 4179 15228 4232
rect 15140 4039 15169 4179
rect 15215 4039 15228 4179
rect 15140 3988 15228 4039
rect 15624 4179 15712 4232
rect 15624 4039 15637 4179
rect 15683 4039 15712 4179
rect 15624 3988 15712 4039
rect 15812 4179 15900 4232
rect 15812 4039 15841 4179
rect 15887 4039 15900 4179
rect 15812 3988 15900 4039
rect 16296 4179 16384 4232
rect 16296 4039 16309 4179
rect 16355 4039 16384 4179
rect 16296 3988 16384 4039
rect 16484 4179 16572 4232
rect 16484 4039 16513 4179
rect 16559 4039 16572 4179
rect 16484 3988 16572 4039
rect 16724 4187 16812 4232
rect 16724 4047 16737 4187
rect 16783 4047 16812 4187
rect 16724 3988 16812 4047
rect 17012 4187 17100 4232
rect 17012 4047 17041 4187
rect 17087 4047 17100 4187
rect 17012 3988 17100 4047
rect 17640 4179 17728 4232
rect 17640 4039 17653 4179
rect 17699 4039 17728 4179
rect 17640 3988 17728 4039
rect 17828 4179 17916 4232
rect 17828 4039 17857 4179
rect 17903 4039 17916 4179
rect 17828 3988 17916 4039
rect 18312 4179 18400 4232
rect 18312 4039 18325 4179
rect 18371 4039 18400 4179
rect 18312 3988 18400 4039
rect 18500 4179 18588 4232
rect 18500 4039 18529 4179
rect 18575 4039 18588 4179
rect 18500 3988 18588 4039
rect 18984 4179 19072 4232
rect 18984 4039 18997 4179
rect 19043 4039 19072 4179
rect 18984 3988 19072 4039
rect 19172 4179 19260 4232
rect 19172 4039 19201 4179
rect 19247 4039 19260 4179
rect 19172 3988 19260 4039
rect 19656 4179 19744 4232
rect 19656 4039 19669 4179
rect 19715 4039 19744 4179
rect 19656 3988 19744 4039
rect 19844 4179 19932 4232
rect 19844 4039 19873 4179
rect 19919 4039 19932 4179
rect 19844 3988 19932 4039
rect 20328 4179 20416 4232
rect 20328 4039 20341 4179
rect 20387 4039 20416 4179
rect 20328 3988 20416 4039
rect 20516 4179 20604 4232
rect 20516 4039 20545 4179
rect 20591 4039 20604 4179
rect 20516 3988 20604 4039
rect 21000 4179 21088 4232
rect 21000 4039 21013 4179
rect 21059 4039 21088 4179
rect 21000 3988 21088 4039
rect 21188 4179 21276 4232
rect 21188 4039 21217 4179
rect 21263 4039 21276 4179
rect 21188 3988 21276 4039
rect 21732 4179 21820 4232
rect 21732 4039 21745 4179
rect 21791 4039 21820 4179
rect 21732 3988 21820 4039
rect 21920 4179 22008 4232
rect 21920 4039 21949 4179
rect 21995 4039 22008 4179
rect 21920 3988 22008 4039
rect 1604 3793 1692 3852
rect 1604 3653 1617 3793
rect 1663 3653 1692 3793
rect 1604 3608 1692 3653
rect 1892 3793 1980 3852
rect 1892 3653 1921 3793
rect 1967 3653 1980 3793
rect 1892 3608 1980 3653
rect 2052 3793 2140 3852
rect 2052 3653 2065 3793
rect 2111 3653 2140 3793
rect 2052 3608 2140 3653
rect 2340 3793 2428 3852
rect 2340 3653 2369 3793
rect 2415 3653 2428 3793
rect 2340 3608 2428 3653
rect 2744 3801 2832 3852
rect 2744 3661 2757 3801
rect 2803 3661 2832 3801
rect 2744 3608 2832 3661
rect 2932 3801 3020 3852
rect 2932 3661 2961 3801
rect 3007 3661 3020 3801
rect 2932 3608 3020 3661
rect 3416 3801 3504 3852
rect 3416 3661 3429 3801
rect 3475 3661 3504 3801
rect 3416 3608 3504 3661
rect 3604 3801 3692 3852
rect 3604 3661 3633 3801
rect 3679 3661 3692 3801
rect 3604 3608 3692 3661
rect 4088 3801 4176 3852
rect 4088 3661 4101 3801
rect 4147 3661 4176 3801
rect 4088 3608 4176 3661
rect 4276 3801 4364 3852
rect 4276 3661 4305 3801
rect 4351 3661 4364 3801
rect 4276 3608 4364 3661
rect 4760 3801 4848 3852
rect 4760 3661 4773 3801
rect 4819 3661 4848 3801
rect 4760 3608 4848 3661
rect 4948 3801 5036 3852
rect 4948 3661 4977 3801
rect 5023 3661 5036 3801
rect 4948 3608 5036 3661
rect 5716 3801 5804 3852
rect 5716 3661 5729 3801
rect 5775 3661 5804 3801
rect 5716 3608 5804 3661
rect 5904 3801 5992 3852
rect 5904 3661 5933 3801
rect 5979 3661 5992 3801
rect 5904 3608 5992 3661
rect 6388 3801 6476 3852
rect 6388 3661 6401 3801
rect 6447 3661 6476 3801
rect 6388 3608 6476 3661
rect 6576 3801 6664 3852
rect 6576 3661 6605 3801
rect 6651 3661 6664 3801
rect 6576 3608 6664 3661
rect 7060 3801 7148 3852
rect 7060 3661 7073 3801
rect 7119 3661 7148 3801
rect 7060 3608 7148 3661
rect 7248 3801 7336 3852
rect 7248 3661 7277 3801
rect 7323 3661 7336 3801
rect 7248 3608 7336 3661
rect 7672 3801 7760 3852
rect 7672 3661 7685 3801
rect 7731 3661 7760 3801
rect 7672 3608 7760 3661
rect 7860 3801 7948 3852
rect 7860 3661 7889 3801
rect 7935 3661 7948 3801
rect 7860 3608 7948 3661
rect 8404 3801 8492 3852
rect 8404 3661 8417 3801
rect 8463 3661 8492 3801
rect 8404 3608 8492 3661
rect 8592 3801 8680 3852
rect 8592 3661 8621 3801
rect 8667 3661 8680 3801
rect 8592 3608 8680 3661
rect 8772 3793 8860 3852
rect 8772 3653 8785 3793
rect 8831 3653 8860 3793
rect 8772 3608 8860 3653
rect 9060 3793 9148 3852
rect 9060 3653 9089 3793
rect 9135 3653 9148 3793
rect 9060 3608 9148 3653
rect 9636 3801 9724 3852
rect 9636 3661 9649 3801
rect 9695 3661 9724 3801
rect 9636 3608 9724 3661
rect 9824 3801 9912 3852
rect 9824 3661 9853 3801
rect 9899 3661 9912 3801
rect 9824 3608 9912 3661
rect 10248 3801 10336 3852
rect 10248 3661 10261 3801
rect 10307 3661 10336 3801
rect 10248 3608 10336 3661
rect 10436 3801 10524 3852
rect 10436 3661 10465 3801
rect 10511 3661 10524 3801
rect 10436 3608 10524 3661
rect 10920 3801 11008 3852
rect 10920 3661 10933 3801
rect 10979 3661 11008 3801
rect 10920 3608 11008 3661
rect 11108 3801 11196 3852
rect 11108 3661 11137 3801
rect 11183 3661 11196 3801
rect 11108 3608 11196 3661
rect 11652 3801 11740 3852
rect 11652 3661 11665 3801
rect 11711 3661 11740 3801
rect 11652 3608 11740 3661
rect 11840 3801 11928 3852
rect 11840 3661 11869 3801
rect 11915 3661 11928 3801
rect 11840 3608 11928 3661
rect 12020 3793 12108 3852
rect 12020 3653 12033 3793
rect 12079 3653 12108 3793
rect 12020 3608 12108 3653
rect 12308 3793 12396 3852
rect 12308 3653 12337 3793
rect 12383 3653 12396 3793
rect 12308 3608 12396 3653
rect 12468 3793 12556 3852
rect 12468 3653 12481 3793
rect 12527 3653 12556 3793
rect 12468 3608 12556 3653
rect 12756 3793 12844 3852
rect 12756 3653 12785 3793
rect 12831 3653 12844 3793
rect 12756 3608 12844 3653
rect 13364 3793 13452 3852
rect 13364 3653 13377 3793
rect 13423 3653 13452 3793
rect 13364 3608 13452 3653
rect 13652 3793 13740 3852
rect 13652 3653 13681 3793
rect 13727 3653 13740 3793
rect 13652 3608 13740 3653
rect 13832 3801 13920 3852
rect 13832 3661 13845 3801
rect 13891 3661 13920 3801
rect 13832 3608 13920 3661
rect 14020 3801 14108 3852
rect 14020 3661 14049 3801
rect 14095 3661 14108 3801
rect 14020 3608 14108 3661
rect 14504 3801 14592 3852
rect 14504 3661 14517 3801
rect 14563 3661 14592 3801
rect 14504 3608 14592 3661
rect 14692 3801 14780 3852
rect 14692 3661 14721 3801
rect 14767 3661 14780 3801
rect 14692 3608 14780 3661
rect 15176 3801 15264 3852
rect 15176 3661 15189 3801
rect 15235 3661 15264 3801
rect 15176 3608 15264 3661
rect 15364 3801 15452 3852
rect 15364 3661 15393 3801
rect 15439 3661 15452 3801
rect 15364 3608 15452 3661
rect 15848 3801 15936 3852
rect 15848 3661 15861 3801
rect 15907 3661 15936 3801
rect 15848 3608 15936 3661
rect 16036 3801 16124 3852
rect 16036 3661 16065 3801
rect 16111 3661 16124 3801
rect 16036 3608 16124 3661
rect 16520 3801 16608 3852
rect 16520 3661 16533 3801
rect 16579 3661 16608 3801
rect 16520 3608 16608 3661
rect 16708 3801 16796 3852
rect 16708 3661 16737 3801
rect 16783 3661 16796 3801
rect 16708 3608 16796 3661
rect 17416 3801 17504 3852
rect 17416 3661 17429 3801
rect 17475 3661 17504 3801
rect 17416 3608 17504 3661
rect 17604 3801 17692 3852
rect 17604 3661 17633 3801
rect 17679 3661 17692 3801
rect 17604 3608 17692 3661
rect 18088 3801 18176 3852
rect 18088 3661 18101 3801
rect 18147 3661 18176 3801
rect 18088 3608 18176 3661
rect 18276 3801 18364 3852
rect 18276 3661 18305 3801
rect 18351 3661 18364 3801
rect 18276 3608 18364 3661
rect 18760 3801 18848 3852
rect 18760 3661 18773 3801
rect 18819 3661 18848 3801
rect 18760 3608 18848 3661
rect 18948 3801 19036 3852
rect 18948 3661 18977 3801
rect 19023 3661 19036 3801
rect 18948 3608 19036 3661
rect 19432 3801 19520 3852
rect 19432 3661 19445 3801
rect 19491 3661 19520 3801
rect 19432 3608 19520 3661
rect 19620 3801 19708 3852
rect 19620 3661 19649 3801
rect 19695 3661 19708 3801
rect 19620 3608 19708 3661
rect 20104 3801 20192 3852
rect 20104 3661 20117 3801
rect 20163 3661 20192 3801
rect 20104 3608 20192 3661
rect 20292 3801 20380 3852
rect 20292 3661 20321 3801
rect 20367 3661 20380 3801
rect 20292 3608 20380 3661
rect 20532 3793 20620 3852
rect 20532 3653 20545 3793
rect 20591 3653 20620 3793
rect 20532 3608 20620 3653
rect 20820 3793 20908 3852
rect 20820 3653 20849 3793
rect 20895 3653 20908 3793
rect 20820 3608 20908 3653
rect 21204 3793 21292 3852
rect 21204 3653 21217 3793
rect 21263 3653 21292 3793
rect 21204 3608 21292 3653
rect 21492 3793 21580 3852
rect 21492 3653 21521 3793
rect 21567 3653 21580 3793
rect 21492 3608 21580 3653
rect 21652 3793 21740 3852
rect 21652 3653 21665 3793
rect 21711 3653 21740 3793
rect 21652 3608 21740 3653
rect 21940 3793 22028 3852
rect 21940 3653 21969 3793
rect 22015 3653 22028 3793
rect 21940 3608 22028 3653
<< mvndiffc >>
rect 1617 15826 1663 15872
rect 1921 15826 1967 15872
rect 2065 15826 2111 15872
rect 2369 15826 2415 15872
rect 2513 15826 2559 15872
rect 2817 15826 2863 15872
rect 2961 15826 3007 15872
rect 3265 15826 3311 15872
rect 3409 15826 3455 15872
rect 3713 15826 3759 15872
rect 3857 15826 3903 15872
rect 4161 15826 4207 15872
rect 4305 15826 4351 15872
rect 4609 15826 4655 15872
rect 4753 15826 4799 15872
rect 5057 15826 5103 15872
rect 5537 15826 5583 15872
rect 5841 15826 5887 15872
rect 5985 15826 6031 15872
rect 6289 15826 6335 15872
rect 6433 15826 6479 15872
rect 6737 15826 6783 15872
rect 6881 15826 6927 15872
rect 7185 15826 7231 15872
rect 7329 15826 7375 15872
rect 7633 15826 7679 15872
rect 7777 15826 7823 15872
rect 8081 15826 8127 15872
rect 8225 15826 8271 15872
rect 8529 15826 8575 15872
rect 8673 15826 8719 15872
rect 8977 15826 9023 15872
rect 9457 15826 9503 15872
rect 9761 15826 9807 15872
rect 9905 15826 9951 15872
rect 10209 15826 10255 15872
rect 10353 15826 10399 15872
rect 10657 15826 10703 15872
rect 10801 15826 10847 15872
rect 11105 15826 11151 15872
rect 11249 15826 11295 15872
rect 11553 15826 11599 15872
rect 11697 15826 11743 15872
rect 12001 15826 12047 15872
rect 12145 15826 12191 15872
rect 12449 15826 12495 15872
rect 12593 15826 12639 15872
rect 12897 15826 12943 15872
rect 13377 15826 13423 15872
rect 13681 15826 13727 15872
rect 13825 15826 13871 15872
rect 14129 15826 14175 15872
rect 14273 15826 14319 15872
rect 14577 15826 14623 15872
rect 14721 15826 14767 15872
rect 15025 15826 15071 15872
rect 15169 15826 15215 15872
rect 15473 15826 15519 15872
rect 15617 15826 15663 15872
rect 15921 15826 15967 15872
rect 16065 15826 16111 15872
rect 16369 15826 16415 15872
rect 16513 15826 16559 15872
rect 16817 15826 16863 15872
rect 17297 15826 17343 15872
rect 17601 15826 17647 15872
rect 17745 15826 17791 15872
rect 18049 15826 18095 15872
rect 18193 15826 18239 15872
rect 18497 15826 18543 15872
rect 18641 15826 18687 15872
rect 18945 15826 18991 15872
rect 19089 15826 19135 15872
rect 19393 15826 19439 15872
rect 19537 15826 19583 15872
rect 19841 15826 19887 15872
rect 19985 15826 20031 15872
rect 20289 15826 20335 15872
rect 20433 15826 20479 15872
rect 20737 15826 20783 15872
rect 21217 15826 21263 15872
rect 21521 15826 21567 15872
rect 21665 15826 21711 15872
rect 21969 15826 22015 15872
rect 1617 15488 1663 15534
rect 1921 15488 1967 15534
rect 2065 15488 2111 15534
rect 2369 15488 2415 15534
rect 2513 15488 2559 15534
rect 2817 15488 2863 15534
rect 2961 15488 3007 15534
rect 3265 15488 3311 15534
rect 3409 15488 3455 15534
rect 3713 15488 3759 15534
rect 3857 15488 3903 15534
rect 4161 15488 4207 15534
rect 4305 15488 4351 15534
rect 4609 15488 4655 15534
rect 4753 15488 4799 15534
rect 5057 15488 5103 15534
rect 5201 15488 5247 15534
rect 5505 15488 5551 15534
rect 5649 15488 5695 15534
rect 5953 15488 5999 15534
rect 6097 15488 6143 15534
rect 6401 15488 6447 15534
rect 6545 15488 6591 15534
rect 6849 15488 6895 15534
rect 6993 15488 7039 15534
rect 7297 15488 7343 15534
rect 7441 15488 7487 15534
rect 7745 15488 7791 15534
rect 7889 15488 7935 15534
rect 8193 15488 8239 15534
rect 8337 15488 8383 15534
rect 8641 15488 8687 15534
rect 8785 15488 8831 15534
rect 9089 15488 9135 15534
rect 9569 15488 9615 15534
rect 9873 15488 9919 15534
rect 10017 15488 10063 15534
rect 10321 15488 10367 15534
rect 10465 15488 10511 15534
rect 10769 15488 10815 15534
rect 10913 15488 10959 15534
rect 11217 15488 11263 15534
rect 11361 15488 11407 15534
rect 11665 15488 11711 15534
rect 11809 15488 11855 15534
rect 12113 15488 12159 15534
rect 12257 15488 12303 15534
rect 12561 15488 12607 15534
rect 12705 15488 12751 15534
rect 13009 15488 13055 15534
rect 13153 15488 13199 15534
rect 13457 15488 13503 15534
rect 13601 15488 13647 15534
rect 13905 15488 13951 15534
rect 14049 15488 14095 15534
rect 14353 15488 14399 15534
rect 14497 15488 14543 15534
rect 14801 15488 14847 15534
rect 14945 15488 14991 15534
rect 15249 15488 15295 15534
rect 15393 15488 15439 15534
rect 15697 15488 15743 15534
rect 15841 15488 15887 15534
rect 16145 15488 16191 15534
rect 16289 15488 16335 15534
rect 16593 15488 16639 15534
rect 16737 15488 16783 15534
rect 17041 15488 17087 15534
rect 17521 15488 17567 15534
rect 17825 15488 17871 15534
rect 17969 15488 18015 15534
rect 18273 15488 18319 15534
rect 18417 15488 18463 15534
rect 18721 15488 18767 15534
rect 18865 15488 18911 15534
rect 19169 15488 19215 15534
rect 19313 15488 19359 15534
rect 19617 15488 19663 15534
rect 19761 15488 19807 15534
rect 20065 15488 20111 15534
rect 20209 15488 20255 15534
rect 20513 15488 20559 15534
rect 20657 15488 20703 15534
rect 20961 15488 21007 15534
rect 21105 15488 21151 15534
rect 21409 15488 21455 15534
rect 21553 15488 21599 15534
rect 21857 15488 21903 15534
rect 22001 15488 22047 15534
rect 22305 15488 22351 15534
rect 1617 14258 1663 14304
rect 1921 14258 1967 14304
rect 2065 14258 2111 14304
rect 2369 14258 2415 14304
rect 2513 14258 2559 14304
rect 2817 14258 2863 14304
rect 2961 14258 3007 14304
rect 3265 14258 3311 14304
rect 3409 14258 3455 14304
rect 3713 14258 3759 14304
rect 3857 14258 3903 14304
rect 4161 14258 4207 14304
rect 4305 14258 4351 14304
rect 4609 14258 4655 14304
rect 4753 14258 4799 14304
rect 5057 14258 5103 14304
rect 5537 14258 5583 14304
rect 5841 14258 5887 14304
rect 5985 14258 6031 14304
rect 6289 14258 6335 14304
rect 6433 14258 6479 14304
rect 6737 14258 6783 14304
rect 6881 14258 6927 14304
rect 7185 14258 7231 14304
rect 7329 14258 7375 14304
rect 7633 14258 7679 14304
rect 7777 14258 7823 14304
rect 8081 14258 8127 14304
rect 8225 14258 8271 14304
rect 8529 14258 8575 14304
rect 8673 14258 8719 14304
rect 8977 14258 9023 14304
rect 9121 14258 9167 14304
rect 9425 14258 9471 14304
rect 9569 14258 9615 14304
rect 9873 14258 9919 14304
rect 10017 14258 10063 14304
rect 10321 14258 10367 14304
rect 10465 14258 10511 14304
rect 10769 14258 10815 14304
rect 10913 14258 10959 14304
rect 11217 14258 11263 14304
rect 11361 14258 11407 14304
rect 11665 14258 11711 14304
rect 11809 14258 11855 14304
rect 12113 14258 12159 14304
rect 12257 14258 12303 14304
rect 12561 14258 12607 14304
rect 12705 14258 12751 14304
rect 13009 14258 13055 14304
rect 13489 14258 13535 14304
rect 13793 14258 13839 14304
rect 13937 14258 13983 14304
rect 14241 14258 14287 14304
rect 14385 14258 14431 14304
rect 14689 14258 14735 14304
rect 14833 14258 14879 14304
rect 15137 14258 15183 14304
rect 15281 14258 15327 14304
rect 15585 14258 15631 14304
rect 15729 14258 15775 14304
rect 16033 14258 16079 14304
rect 16177 14258 16223 14304
rect 16481 14258 16527 14304
rect 16817 14258 16863 14304
rect 17041 14258 17087 14304
rect 17489 14258 17535 14304
rect 17713 14258 17759 14304
rect 17857 14258 17903 14304
rect 18161 14258 18207 14304
rect 18305 14258 18351 14304
rect 18609 14258 18655 14304
rect 18753 14258 18799 14304
rect 19057 14258 19103 14304
rect 19201 14258 19247 14304
rect 19505 14258 19551 14304
rect 19649 14258 19695 14304
rect 19953 14258 19999 14304
rect 20097 14258 20143 14304
rect 20401 14258 20447 14304
rect 20545 14258 20591 14304
rect 20849 14258 20895 14304
rect 21441 14258 21487 14304
rect 21745 14258 21791 14304
rect 21889 14258 21935 14304
rect 22193 14258 22239 14304
rect 1617 13920 1663 13966
rect 1921 13920 1967 13966
rect 2065 13920 2111 13966
rect 2369 13920 2415 13966
rect 2513 13920 2559 13966
rect 2817 13920 2863 13966
rect 2961 13920 3007 13966
rect 3265 13920 3311 13966
rect 3409 13920 3455 13966
rect 3713 13920 3759 13966
rect 3857 13920 3903 13966
rect 4161 13920 4207 13966
rect 4305 13920 4351 13966
rect 4609 13920 4655 13966
rect 4753 13920 4799 13966
rect 5057 13920 5103 13966
rect 5201 13920 5247 13966
rect 5505 13920 5551 13966
rect 5649 13920 5695 13966
rect 5953 13920 5999 13966
rect 6097 13920 6143 13966
rect 6401 13920 6447 13966
rect 6545 13920 6591 13966
rect 6849 13920 6895 13966
rect 6993 13920 7039 13966
rect 7297 13920 7343 13966
rect 7441 13920 7487 13966
rect 7745 13920 7791 13966
rect 7889 13920 7935 13966
rect 8193 13920 8239 13966
rect 8337 13920 8383 13966
rect 8641 13920 8687 13966
rect 8785 13920 8831 13966
rect 9089 13920 9135 13966
rect 9569 13920 9615 13966
rect 9873 13920 9919 13966
rect 10017 13920 10063 13966
rect 10321 13920 10367 13966
rect 10465 13920 10511 13966
rect 10769 13920 10815 13966
rect 10913 13920 10959 13966
rect 11217 13920 11263 13966
rect 11361 13920 11407 13966
rect 11665 13920 11711 13966
rect 11809 13920 11855 13966
rect 12113 13920 12159 13966
rect 12257 13920 12303 13966
rect 12561 13920 12607 13966
rect 12705 13920 12751 13966
rect 13009 13920 13055 13966
rect 13153 13920 13199 13966
rect 13457 13920 13503 13966
rect 13601 13920 13647 13966
rect 13905 13920 13951 13966
rect 14049 13920 14095 13966
rect 14353 13920 14399 13966
rect 14497 13920 14543 13966
rect 14801 13920 14847 13966
rect 14945 13920 14991 13966
rect 15249 13920 15295 13966
rect 15393 13920 15439 13966
rect 15697 13920 15743 13966
rect 16065 13920 16111 13966
rect 16289 13920 16335 13966
rect 16737 13920 16783 13966
rect 16961 13920 17007 13966
rect 17633 13920 17679 13966
rect 17857 13920 17903 13966
rect 18305 13920 18351 13966
rect 18529 13920 18575 13966
rect 18753 13920 18799 13966
rect 19057 13920 19103 13966
rect 19201 13920 19247 13966
rect 19505 13920 19551 13966
rect 19649 13920 19695 13966
rect 19953 13920 19999 13966
rect 20097 13920 20143 13966
rect 20401 13920 20447 13966
rect 20545 13920 20591 13966
rect 20849 13920 20895 13966
rect 20993 13920 21039 13966
rect 21297 13920 21343 13966
rect 21441 13920 21487 13966
rect 21745 13920 21791 13966
rect 21889 13920 21935 13966
rect 22193 13920 22239 13966
rect 1617 12690 1663 12736
rect 1921 12690 1967 12736
rect 2065 12690 2111 12736
rect 2369 12690 2415 12736
rect 2513 12690 2559 12736
rect 2817 12690 2863 12736
rect 2961 12690 3007 12736
rect 3265 12690 3311 12736
rect 3409 12690 3455 12736
rect 3713 12690 3759 12736
rect 3857 12690 3903 12736
rect 4161 12690 4207 12736
rect 4305 12690 4351 12736
rect 4609 12690 4655 12736
rect 4753 12690 4799 12736
rect 5057 12690 5103 12736
rect 5537 12690 5583 12736
rect 5841 12690 5887 12736
rect 5985 12690 6031 12736
rect 6289 12690 6335 12736
rect 6433 12690 6479 12736
rect 6737 12690 6783 12736
rect 6881 12690 6927 12736
rect 7185 12690 7231 12736
rect 7329 12690 7375 12736
rect 7633 12690 7679 12736
rect 7777 12690 7823 12736
rect 8081 12690 8127 12736
rect 8225 12690 8271 12736
rect 8529 12690 8575 12736
rect 8673 12690 8719 12736
rect 8977 12690 9023 12736
rect 9121 12690 9167 12736
rect 9425 12690 9471 12736
rect 9569 12690 9615 12736
rect 9873 12690 9919 12736
rect 10017 12690 10063 12736
rect 10321 12690 10367 12736
rect 10465 12690 10511 12736
rect 10769 12690 10815 12736
rect 10913 12690 10959 12736
rect 11217 12690 11263 12736
rect 11361 12690 11407 12736
rect 11665 12690 11711 12736
rect 11809 12690 11855 12736
rect 12113 12690 12159 12736
rect 12257 12690 12303 12736
rect 12561 12690 12607 12736
rect 12705 12690 12751 12736
rect 13009 12690 13055 12736
rect 13489 12690 13535 12736
rect 13793 12690 13839 12736
rect 13937 12690 13983 12736
rect 14241 12690 14287 12736
rect 14721 12690 14767 12736
rect 14945 12690 14991 12736
rect 15393 12690 15439 12736
rect 15617 12690 15663 12736
rect 16065 12690 16111 12736
rect 16289 12690 16335 12736
rect 16737 12690 16783 12736
rect 16961 12690 17007 12736
rect 17409 12690 17455 12736
rect 17633 12690 17679 12736
rect 18081 12690 18127 12736
rect 18305 12690 18351 12736
rect 18753 12690 18799 12736
rect 18977 12690 19023 12736
rect 19425 12690 19471 12736
rect 19649 12690 19695 12736
rect 19873 12690 19919 12736
rect 20177 12690 20223 12736
rect 20321 12690 20367 12736
rect 20625 12690 20671 12736
rect 20769 12690 20815 12736
rect 21073 12690 21119 12736
rect 21441 12690 21487 12736
rect 21745 12690 21791 12736
rect 21889 12690 21935 12736
rect 22193 12690 22239 12736
rect 1617 12352 1663 12398
rect 1921 12352 1967 12398
rect 2065 12352 2111 12398
rect 2369 12352 2415 12398
rect 2513 12352 2559 12398
rect 2817 12352 2863 12398
rect 2961 12352 3007 12398
rect 3265 12352 3311 12398
rect 3409 12352 3455 12398
rect 3713 12352 3759 12398
rect 3857 12352 3903 12398
rect 4161 12352 4207 12398
rect 4305 12352 4351 12398
rect 4609 12352 4655 12398
rect 4753 12352 4799 12398
rect 5057 12352 5103 12398
rect 5201 12352 5247 12398
rect 5505 12352 5551 12398
rect 5649 12352 5695 12398
rect 5953 12352 5999 12398
rect 6097 12352 6143 12398
rect 6401 12352 6447 12398
rect 6545 12352 6591 12398
rect 6849 12352 6895 12398
rect 6993 12352 7039 12398
rect 7297 12352 7343 12398
rect 7441 12352 7487 12398
rect 7745 12352 7791 12398
rect 7889 12352 7935 12398
rect 8193 12352 8239 12398
rect 8337 12352 8383 12398
rect 8641 12352 8687 12398
rect 8785 12352 8831 12398
rect 9089 12352 9135 12398
rect 9569 12352 9615 12398
rect 9873 12352 9919 12398
rect 10017 12352 10063 12398
rect 10321 12352 10367 12398
rect 10465 12352 10511 12398
rect 10769 12352 10815 12398
rect 10913 12352 10959 12398
rect 11217 12352 11263 12398
rect 11361 12352 11407 12398
rect 11665 12352 11711 12398
rect 11809 12352 11855 12398
rect 12113 12352 12159 12398
rect 12257 12352 12303 12398
rect 12561 12352 12607 12398
rect 12705 12352 12751 12398
rect 13009 12352 13055 12398
rect 13153 12352 13199 12398
rect 13457 12352 13503 12398
rect 13601 12352 13647 12398
rect 13905 12352 13951 12398
rect 14049 12352 14095 12398
rect 14273 12352 14319 12398
rect 14721 12352 14767 12398
rect 14945 12352 14991 12398
rect 15393 12352 15439 12398
rect 15617 12352 15663 12398
rect 16065 12352 16111 12398
rect 16289 12352 16335 12398
rect 16737 12352 16783 12398
rect 16961 12352 17007 12398
rect 17633 12352 17679 12398
rect 17857 12352 17903 12398
rect 18305 12352 18351 12398
rect 18529 12352 18575 12398
rect 18977 12352 19023 12398
rect 19201 12352 19247 12398
rect 19649 12352 19695 12398
rect 19873 12352 19919 12398
rect 20321 12352 20367 12398
rect 20545 12352 20591 12398
rect 20769 12352 20815 12398
rect 21073 12352 21119 12398
rect 21217 12352 21263 12398
rect 21521 12352 21567 12398
rect 21665 12352 21711 12398
rect 21969 12352 22015 12398
rect 1617 11122 1663 11168
rect 1921 11122 1967 11168
rect 2065 11122 2111 11168
rect 2369 11122 2415 11168
rect 2513 11122 2559 11168
rect 2817 11122 2863 11168
rect 2961 11122 3007 11168
rect 3265 11122 3311 11168
rect 3409 11122 3455 11168
rect 3713 11122 3759 11168
rect 3857 11122 3903 11168
rect 4161 11122 4207 11168
rect 4305 11122 4351 11168
rect 4609 11122 4655 11168
rect 4753 11122 4799 11168
rect 5057 11122 5103 11168
rect 5537 11122 5583 11168
rect 5841 11122 5887 11168
rect 6065 11122 6111 11168
rect 6289 11122 6335 11168
rect 6849 11122 6895 11168
rect 7073 11122 7119 11168
rect 7521 11122 7567 11168
rect 7745 11122 7791 11168
rect 8193 11122 8239 11168
rect 8417 11122 8463 11168
rect 8561 11122 8607 11168
rect 8865 11122 8911 11168
rect 9121 11122 9167 11168
rect 9345 11122 9391 11168
rect 9793 11122 9839 11168
rect 10017 11122 10063 11168
rect 10465 11122 10511 11168
rect 10689 11122 10735 11168
rect 10913 11122 10959 11168
rect 11217 11122 11263 11168
rect 11361 11122 11407 11168
rect 11665 11122 11711 11168
rect 12033 11122 12079 11168
rect 12257 11122 12303 11168
rect 12705 11122 12751 11168
rect 12929 11122 12975 11168
rect 13601 11122 13647 11168
rect 13825 11122 13871 11168
rect 14049 11122 14095 11168
rect 14353 11122 14399 11168
rect 14721 11122 14767 11168
rect 14945 11122 14991 11168
rect 15393 11122 15439 11168
rect 15617 11122 15663 11168
rect 16065 11122 16111 11168
rect 16289 11122 16335 11168
rect 16737 11122 16783 11168
rect 16961 11122 17007 11168
rect 17409 11122 17455 11168
rect 17633 11122 17679 11168
rect 18081 11122 18127 11168
rect 18305 11122 18351 11168
rect 18753 11122 18799 11168
rect 18977 11122 19023 11168
rect 19425 11122 19471 11168
rect 19649 11122 19695 11168
rect 20097 11122 20143 11168
rect 20321 11122 20367 11168
rect 20545 11122 20591 11168
rect 20849 11122 20895 11168
rect 21441 11122 21487 11168
rect 21745 11122 21791 11168
rect 21889 11122 21935 11168
rect 22193 11122 22239 11168
rect 1617 10784 1663 10830
rect 1921 10784 1967 10830
rect 2065 10784 2111 10830
rect 2369 10784 2415 10830
rect 2513 10784 2559 10830
rect 2817 10784 2863 10830
rect 2961 10784 3007 10830
rect 3265 10784 3311 10830
rect 3409 10784 3455 10830
rect 3713 10784 3759 10830
rect 3857 10784 3903 10830
rect 4161 10784 4207 10830
rect 4305 10784 4351 10830
rect 4609 10784 4655 10830
rect 4753 10784 4799 10830
rect 5057 10784 5103 10830
rect 5313 10784 5359 10830
rect 5537 10784 5583 10830
rect 5985 10784 6031 10830
rect 6209 10784 6255 10830
rect 6657 10784 6703 10830
rect 6881 10784 6927 10830
rect 7329 10784 7375 10830
rect 7553 10784 7599 10830
rect 8001 10784 8047 10830
rect 8225 10784 8271 10830
rect 8785 10784 8831 10830
rect 9009 10784 9055 10830
rect 9793 10784 9839 10830
rect 10017 10784 10063 10830
rect 10465 10784 10511 10830
rect 10689 10784 10735 10830
rect 11137 10784 11183 10830
rect 11361 10784 11407 10830
rect 11921 10784 11967 10830
rect 12145 10784 12191 10830
rect 12593 10784 12639 10830
rect 12817 10784 12863 10830
rect 13265 10784 13311 10830
rect 13489 10784 13535 10830
rect 13937 10784 13983 10830
rect 14161 10784 14207 10830
rect 14609 10784 14655 10830
rect 14833 10784 14879 10830
rect 15281 10784 15327 10830
rect 15505 10784 15551 10830
rect 15953 10784 15999 10830
rect 16177 10784 16223 10830
rect 16625 10784 16671 10830
rect 16849 10784 16895 10830
rect 17633 10784 17679 10830
rect 17857 10784 17903 10830
rect 18305 10784 18351 10830
rect 18529 10784 18575 10830
rect 18977 10784 19023 10830
rect 19201 10784 19247 10830
rect 19649 10784 19695 10830
rect 19873 10784 19919 10830
rect 20321 10784 20367 10830
rect 20545 10784 20591 10830
rect 20993 10784 21039 10830
rect 21217 10784 21263 10830
rect 21665 10784 21711 10830
rect 21889 10784 21935 10830
rect 1617 9554 1663 9600
rect 1921 9554 1967 9600
rect 2065 9554 2111 9600
rect 2369 9554 2415 9600
rect 2513 9554 2559 9600
rect 2817 9554 2863 9600
rect 2961 9554 3007 9600
rect 3265 9554 3311 9600
rect 3409 9554 3455 9600
rect 3713 9554 3759 9600
rect 4081 9554 4127 9600
rect 4305 9554 4351 9600
rect 4753 9554 4799 9600
rect 4977 9554 5023 9600
rect 5761 9554 5807 9600
rect 5985 9554 6031 9600
rect 6433 9554 6479 9600
rect 6657 9554 6703 9600
rect 7105 9554 7151 9600
rect 7329 9554 7375 9600
rect 7777 9554 7823 9600
rect 8001 9554 8047 9600
rect 8449 9554 8495 9600
rect 8673 9554 8719 9600
rect 9121 9554 9167 9600
rect 9345 9554 9391 9600
rect 9793 9554 9839 9600
rect 10017 9554 10063 9600
rect 10465 9554 10511 9600
rect 10689 9554 10735 9600
rect 10913 9554 10959 9600
rect 11217 9554 11263 9600
rect 11361 9554 11407 9600
rect 11585 9554 11631 9600
rect 12033 9554 12079 9600
rect 12257 9554 12303 9600
rect 12705 9554 12751 9600
rect 12929 9554 12975 9600
rect 13601 9554 13647 9600
rect 13825 9554 13871 9600
rect 14273 9554 14319 9600
rect 14497 9554 14543 9600
rect 14945 9554 14991 9600
rect 15169 9554 15215 9600
rect 15617 9554 15663 9600
rect 15841 9554 15887 9600
rect 16289 9554 16335 9600
rect 16513 9554 16559 9600
rect 16961 9554 17007 9600
rect 17185 9554 17231 9600
rect 17713 9554 17759 9600
rect 17937 9554 17983 9600
rect 18305 9554 18351 9600
rect 18529 9554 18575 9600
rect 18977 9554 19023 9600
rect 19201 9554 19247 9600
rect 19649 9554 19695 9600
rect 19873 9554 19919 9600
rect 20321 9554 20367 9600
rect 20545 9554 20591 9600
rect 20769 9554 20815 9600
rect 21073 9554 21119 9600
rect 21553 9554 21599 9600
rect 21777 9554 21823 9600
rect 22001 9554 22047 9600
rect 22305 9554 22351 9600
rect 1617 9216 1663 9262
rect 1921 9216 1967 9262
rect 2065 9216 2111 9262
rect 2369 9216 2415 9262
rect 2513 9216 2559 9262
rect 2817 9216 2863 9262
rect 3297 9216 3343 9262
rect 3521 9216 3567 9262
rect 3969 9216 4015 9262
rect 4193 9216 4239 9262
rect 4641 9216 4687 9262
rect 4865 9216 4911 9262
rect 5313 9216 5359 9262
rect 5537 9216 5583 9262
rect 5985 9216 6031 9262
rect 6209 9216 6255 9262
rect 6657 9216 6703 9262
rect 6881 9216 6927 9262
rect 7329 9216 7375 9262
rect 7553 9216 7599 9262
rect 8113 9216 8159 9262
rect 8337 9216 8383 9262
rect 8785 9216 8831 9262
rect 9009 9216 9055 9262
rect 9569 9216 9615 9262
rect 9873 9216 9919 9262
rect 10241 9216 10287 9262
rect 10465 9216 10511 9262
rect 10913 9216 10959 9262
rect 11137 9216 11183 9262
rect 11585 9216 11631 9262
rect 11809 9216 11855 9262
rect 12257 9216 12303 9262
rect 12481 9216 12527 9262
rect 12929 9216 12975 9262
rect 13153 9216 13199 9262
rect 13601 9216 13647 9262
rect 13825 9216 13871 9262
rect 14273 9216 14319 9262
rect 14497 9216 14543 9262
rect 14945 9216 14991 9262
rect 15169 9216 15215 9262
rect 15617 9216 15663 9262
rect 15841 9216 15887 9262
rect 16289 9216 16335 9262
rect 16513 9216 16559 9262
rect 16737 9216 16783 9262
rect 17041 9216 17087 9262
rect 17633 9216 17679 9262
rect 17857 9216 17903 9262
rect 18305 9216 18351 9262
rect 18529 9216 18575 9262
rect 18977 9216 19023 9262
rect 19201 9216 19247 9262
rect 19649 9216 19695 9262
rect 19873 9216 19919 9262
rect 20321 9216 20367 9262
rect 20545 9216 20591 9262
rect 20769 9216 20815 9262
rect 21073 9216 21119 9262
rect 21217 9216 21263 9262
rect 21521 9216 21567 9262
rect 21665 9216 21711 9262
rect 21969 9216 22015 9262
rect 1617 7986 1663 8032
rect 1921 7986 1967 8032
rect 2065 7986 2111 8032
rect 2369 7986 2415 8032
rect 2817 7986 2863 8032
rect 3041 7986 3087 8032
rect 3409 7986 3455 8032
rect 3633 7986 3679 8032
rect 4081 7986 4127 8032
rect 4305 7986 4351 8032
rect 4753 7986 4799 8032
rect 4977 7986 5023 8032
rect 5761 7986 5807 8032
rect 5985 7986 6031 8032
rect 6433 7986 6479 8032
rect 6657 7986 6703 8032
rect 7105 7986 7151 8032
rect 7329 7986 7375 8032
rect 7777 7986 7823 8032
rect 8001 7986 8047 8032
rect 8449 7986 8495 8032
rect 8673 7986 8719 8032
rect 9121 7986 9167 8032
rect 9345 7986 9391 8032
rect 9793 7986 9839 8032
rect 10017 7986 10063 8032
rect 10465 7986 10511 8032
rect 10689 7986 10735 8032
rect 11217 7986 11263 8032
rect 11441 7986 11487 8032
rect 11585 7986 11631 8032
rect 11889 7986 11935 8032
rect 12033 7986 12079 8032
rect 12257 7986 12303 8032
rect 12705 7986 12751 8032
rect 12929 7986 12975 8032
rect 13601 7986 13647 8032
rect 13825 7986 13871 8032
rect 14273 7986 14319 8032
rect 14497 7986 14543 8032
rect 14945 7986 14991 8032
rect 15169 7986 15215 8032
rect 15617 7986 15663 8032
rect 15841 7986 15887 8032
rect 16289 7986 16335 8032
rect 16513 7986 16559 8032
rect 16961 7986 17007 8032
rect 17185 7986 17231 8032
rect 17633 7986 17679 8032
rect 17857 7986 17903 8032
rect 18305 7986 18351 8032
rect 18529 7986 18575 8032
rect 18977 7986 19023 8032
rect 19201 7986 19247 8032
rect 19649 7986 19695 8032
rect 19873 7986 19919 8032
rect 20401 7986 20447 8032
rect 20625 7986 20671 8032
rect 20769 7986 20815 8032
rect 21073 7986 21119 8032
rect 21441 7986 21487 8032
rect 21745 7986 21791 8032
rect 21889 7986 21935 8032
rect 22193 7986 22239 8032
rect 2033 7648 2079 7694
rect 2257 7648 2303 7694
rect 2625 7648 2671 7694
rect 2849 7648 2895 7694
rect 3297 7648 3343 7694
rect 3521 7648 3567 7694
rect 3969 7648 4015 7694
rect 4193 7648 4239 7694
rect 4641 7648 4687 7694
rect 4865 7648 4911 7694
rect 5313 7648 5359 7694
rect 5537 7648 5583 7694
rect 5985 7648 6031 7694
rect 6209 7648 6255 7694
rect 6657 7648 6703 7694
rect 6881 7648 6927 7694
rect 7329 7648 7375 7694
rect 7553 7648 7599 7694
rect 8113 7648 8159 7694
rect 8337 7648 8383 7694
rect 8785 7648 8831 7694
rect 9009 7648 9055 7694
rect 9793 7648 9839 7694
rect 10017 7648 10063 7694
rect 10465 7648 10511 7694
rect 10689 7648 10735 7694
rect 11217 7648 11263 7694
rect 11441 7648 11487 7694
rect 11809 7648 11855 7694
rect 12033 7648 12079 7694
rect 12481 7648 12527 7694
rect 12705 7648 12751 7694
rect 13153 7648 13199 7694
rect 13377 7648 13423 7694
rect 13825 7648 13871 7694
rect 14049 7648 14095 7694
rect 14497 7648 14543 7694
rect 14721 7648 14767 7694
rect 15169 7648 15215 7694
rect 15393 7648 15439 7694
rect 15841 7648 15887 7694
rect 16065 7648 16111 7694
rect 16513 7648 16559 7694
rect 16737 7648 16783 7694
rect 17633 7648 17679 7694
rect 17857 7648 17903 7694
rect 18305 7648 18351 7694
rect 18529 7648 18575 7694
rect 18977 7648 19023 7694
rect 19201 7648 19247 7694
rect 19649 7648 19695 7694
rect 19873 7648 19919 7694
rect 20321 7648 20367 7694
rect 20545 7648 20591 7694
rect 20993 7648 21039 7694
rect 21217 7648 21263 7694
rect 21441 7648 21487 7694
rect 21745 7648 21791 7694
rect 21889 7648 21935 7694
rect 22193 7648 22239 7694
rect 1617 6418 1663 6464
rect 1921 6418 1967 6464
rect 2065 6418 2111 6464
rect 2289 6418 2335 6464
rect 2737 6418 2783 6464
rect 2961 6418 3007 6464
rect 3409 6418 3455 6464
rect 3633 6418 3679 6464
rect 4081 6418 4127 6464
rect 4305 6418 4351 6464
rect 4753 6418 4799 6464
rect 4977 6418 5023 6464
rect 5649 6418 5695 6464
rect 5873 6418 5919 6464
rect 6321 6418 6367 6464
rect 6545 6418 6591 6464
rect 6993 6418 7039 6464
rect 7217 6418 7263 6464
rect 7665 6418 7711 6464
rect 7889 6418 7935 6464
rect 8337 6418 8383 6464
rect 8561 6418 8607 6464
rect 9009 6418 9055 6464
rect 9233 6418 9279 6464
rect 9681 6418 9727 6464
rect 9905 6418 9951 6464
rect 10353 6418 10399 6464
rect 10577 6418 10623 6464
rect 11025 6418 11071 6464
rect 11249 6418 11295 6464
rect 11697 6418 11743 6464
rect 11921 6418 11967 6464
rect 12369 6418 12415 6464
rect 12593 6418 12639 6464
rect 12817 6418 12863 6464
rect 13121 6418 13167 6464
rect 13489 6418 13535 6464
rect 13793 6418 13839 6464
rect 14049 6418 14095 6464
rect 14273 6418 14319 6464
rect 14721 6418 14767 6464
rect 14945 6418 14991 6464
rect 15393 6418 15439 6464
rect 15617 6418 15663 6464
rect 16065 6418 16111 6464
rect 16289 6418 16335 6464
rect 16737 6418 16783 6464
rect 16961 6418 17007 6464
rect 17409 6418 17455 6464
rect 17633 6418 17679 6464
rect 18081 6418 18127 6464
rect 18305 6418 18351 6464
rect 18753 6418 18799 6464
rect 18977 6418 19023 6464
rect 19425 6418 19471 6464
rect 19649 6418 19695 6464
rect 20177 6418 20223 6464
rect 20401 6418 20447 6464
rect 20545 6418 20591 6464
rect 20849 6418 20895 6464
rect 21553 6418 21599 6464
rect 21777 6418 21823 6464
rect 22001 6418 22047 6464
rect 22305 6418 22351 6464
rect 1953 6080 1999 6126
rect 2177 6080 2223 6126
rect 2625 6080 2671 6126
rect 2849 6080 2895 6126
rect 3297 6080 3343 6126
rect 3521 6080 3567 6126
rect 3969 6080 4015 6126
rect 4193 6080 4239 6126
rect 4641 6080 4687 6126
rect 4865 6080 4911 6126
rect 5313 6080 5359 6126
rect 5537 6080 5583 6126
rect 5985 6080 6031 6126
rect 6209 6080 6255 6126
rect 6657 6080 6703 6126
rect 6881 6080 6927 6126
rect 7329 6080 7375 6126
rect 7553 6080 7599 6126
rect 8001 6080 8047 6126
rect 8225 6080 8271 6126
rect 8673 6080 8719 6126
rect 8897 6080 8943 6126
rect 9681 6080 9727 6126
rect 9905 6080 9951 6126
rect 10353 6080 10399 6126
rect 10577 6080 10623 6126
rect 11025 6080 11071 6126
rect 11249 6080 11295 6126
rect 11697 6080 11743 6126
rect 11921 6080 11967 6126
rect 12481 6080 12527 6126
rect 12705 6080 12751 6126
rect 13153 6080 13199 6126
rect 13377 6080 13423 6126
rect 13825 6080 13871 6126
rect 14049 6080 14095 6126
rect 14497 6080 14543 6126
rect 14721 6080 14767 6126
rect 15169 6080 15215 6126
rect 15393 6080 15439 6126
rect 15841 6080 15887 6126
rect 16065 6080 16111 6126
rect 16513 6080 16559 6126
rect 16737 6080 16783 6126
rect 17633 6080 17679 6126
rect 17857 6080 17903 6126
rect 18305 6080 18351 6126
rect 18529 6080 18575 6126
rect 18977 6080 19023 6126
rect 19201 6080 19247 6126
rect 19649 6080 19695 6126
rect 19873 6080 19919 6126
rect 20321 6080 20367 6126
rect 20545 6080 20591 6126
rect 20993 6080 21039 6126
rect 21217 6080 21263 6126
rect 21745 6080 21791 6126
rect 21969 6080 22015 6126
rect 1617 4850 1663 4896
rect 1921 4850 1967 4896
rect 2065 4850 2111 4896
rect 2289 4850 2335 4896
rect 2737 4850 2783 4896
rect 2961 4850 3007 4896
rect 3409 4850 3455 4896
rect 3633 4850 3679 4896
rect 4081 4850 4127 4896
rect 4305 4850 4351 4896
rect 4753 4850 4799 4896
rect 4977 4850 5023 4896
rect 5649 4850 5695 4896
rect 5873 4850 5919 4896
rect 6321 4850 6367 4896
rect 6545 4850 6591 4896
rect 6993 4850 7039 4896
rect 7217 4850 7263 4896
rect 7665 4850 7711 4896
rect 7889 4850 7935 4896
rect 8337 4850 8383 4896
rect 8561 4850 8607 4896
rect 9009 4850 9055 4896
rect 9233 4850 9279 4896
rect 9681 4850 9727 4896
rect 9905 4850 9951 4896
rect 10353 4850 10399 4896
rect 10577 4850 10623 4896
rect 10801 4850 10847 4896
rect 11105 4850 11151 4896
rect 11361 4850 11407 4896
rect 11585 4850 11631 4896
rect 12033 4850 12079 4896
rect 12257 4850 12303 4896
rect 12705 4850 12751 4896
rect 12929 4850 12975 4896
rect 13489 4850 13535 4896
rect 13793 4850 13839 4896
rect 13937 4850 13983 4896
rect 14161 4850 14207 4896
rect 14609 4850 14655 4896
rect 14833 4850 14879 4896
rect 15281 4850 15327 4896
rect 15505 4850 15551 4896
rect 15953 4850 15999 4896
rect 16177 4850 16223 4896
rect 16625 4850 16671 4896
rect 16849 4850 16895 4896
rect 17297 4850 17343 4896
rect 17521 4850 17567 4896
rect 17969 4850 18015 4896
rect 18193 4850 18239 4896
rect 18641 4850 18687 4896
rect 18865 4850 18911 4896
rect 19313 4850 19359 4896
rect 19537 4850 19583 4896
rect 19985 4850 20031 4896
rect 20209 4850 20255 4896
rect 20657 4850 20703 4896
rect 20881 4850 20927 4896
rect 21553 4850 21599 4896
rect 21777 4850 21823 4896
rect 22001 4850 22047 4896
rect 22305 4850 22351 4896
rect 1617 4512 1663 4558
rect 1921 4512 1967 4558
rect 2289 4512 2335 4558
rect 2513 4512 2559 4558
rect 2961 4512 3007 4558
rect 3185 4512 3231 4558
rect 3633 4512 3679 4558
rect 3857 4512 3903 4558
rect 4305 4512 4351 4558
rect 4529 4512 4575 4558
rect 4977 4512 5023 4558
rect 5201 4512 5247 4558
rect 5649 4512 5695 4558
rect 5873 4512 5919 4558
rect 6321 4512 6367 4558
rect 6545 4512 6591 4558
rect 6993 4512 7039 4558
rect 7217 4512 7263 4558
rect 7665 4512 7711 4558
rect 7889 4512 7935 4558
rect 8337 4512 8383 4558
rect 8561 4512 8607 4558
rect 8785 4512 8831 4558
rect 9089 4512 9135 4558
rect 9681 4512 9727 4558
rect 9905 4512 9951 4558
rect 10353 4512 10399 4558
rect 10577 4512 10623 4558
rect 11025 4512 11071 4558
rect 11249 4512 11295 4558
rect 11473 4512 11519 4558
rect 11777 4512 11823 4558
rect 12257 4512 12303 4558
rect 12481 4512 12527 4558
rect 12929 4512 12975 4558
rect 13153 4512 13199 4558
rect 13601 4512 13647 4558
rect 13825 4512 13871 4558
rect 14273 4512 14319 4558
rect 14497 4512 14543 4558
rect 14945 4512 14991 4558
rect 15169 4512 15215 4558
rect 15617 4512 15663 4558
rect 15841 4512 15887 4558
rect 16289 4512 16335 4558
rect 16513 4512 16559 4558
rect 16737 4512 16783 4558
rect 17041 4512 17087 4558
rect 17633 4512 17679 4558
rect 17857 4512 17903 4558
rect 18305 4512 18351 4558
rect 18529 4512 18575 4558
rect 18977 4512 19023 4558
rect 19201 4512 19247 4558
rect 19649 4512 19695 4558
rect 19873 4512 19919 4558
rect 20321 4512 20367 4558
rect 20545 4512 20591 4558
rect 20993 4512 21039 4558
rect 21217 4512 21263 4558
rect 21745 4512 21791 4558
rect 21969 4512 22015 4558
rect 1617 3282 1663 3328
rect 1921 3282 1967 3328
rect 2065 3282 2111 3328
rect 2369 3282 2415 3328
rect 2737 3282 2783 3328
rect 2961 3282 3007 3328
rect 3409 3282 3455 3328
rect 3633 3282 3679 3328
rect 4081 3282 4127 3328
rect 4305 3282 4351 3328
rect 4753 3282 4799 3328
rect 4977 3282 5023 3328
rect 5729 3282 5775 3328
rect 5953 3282 5999 3328
rect 6401 3282 6447 3328
rect 6625 3282 6671 3328
rect 7073 3282 7119 3328
rect 7297 3282 7343 3328
rect 7665 3282 7711 3328
rect 7889 3282 7935 3328
rect 8417 3282 8463 3328
rect 8641 3282 8687 3328
rect 8785 3282 8831 3328
rect 9089 3282 9135 3328
rect 9649 3282 9695 3328
rect 9873 3282 9919 3328
rect 10241 3282 10287 3328
rect 10465 3282 10511 3328
rect 10913 3282 10959 3328
rect 11137 3282 11183 3328
rect 11665 3282 11711 3328
rect 11889 3282 11935 3328
rect 12033 3282 12079 3328
rect 12337 3282 12383 3328
rect 12481 3282 12527 3328
rect 12785 3282 12831 3328
rect 13377 3282 13423 3328
rect 13681 3282 13727 3328
rect 13825 3282 13871 3328
rect 14049 3282 14095 3328
rect 14497 3282 14543 3328
rect 14721 3282 14767 3328
rect 15169 3282 15215 3328
rect 15393 3282 15439 3328
rect 15841 3282 15887 3328
rect 16065 3282 16111 3328
rect 16513 3282 16559 3328
rect 16737 3282 16783 3328
rect 17409 3282 17455 3328
rect 17633 3282 17679 3328
rect 18081 3282 18127 3328
rect 18305 3282 18351 3328
rect 18753 3282 18799 3328
rect 18977 3282 19023 3328
rect 19425 3282 19471 3328
rect 19649 3282 19695 3328
rect 20097 3282 20143 3328
rect 20321 3282 20367 3328
rect 20545 3282 20591 3328
rect 20849 3282 20895 3328
rect 21217 3282 21263 3328
rect 21521 3282 21567 3328
rect 21665 3282 21711 3328
rect 21969 3282 22015 3328
<< mvpdiffc >>
rect 1617 16197 1663 16337
rect 1921 16197 1967 16337
rect 2065 16197 2111 16337
rect 2369 16197 2415 16337
rect 2513 16197 2559 16337
rect 2817 16197 2863 16337
rect 2961 16197 3007 16337
rect 3265 16197 3311 16337
rect 3409 16197 3455 16337
rect 3713 16197 3759 16337
rect 3857 16197 3903 16337
rect 4161 16197 4207 16337
rect 4305 16197 4351 16337
rect 4609 16197 4655 16337
rect 4753 16197 4799 16337
rect 5057 16197 5103 16337
rect 5537 16197 5583 16337
rect 5841 16197 5887 16337
rect 5985 16197 6031 16337
rect 6289 16197 6335 16337
rect 6433 16197 6479 16337
rect 6737 16197 6783 16337
rect 6881 16197 6927 16337
rect 7185 16197 7231 16337
rect 7329 16197 7375 16337
rect 7633 16197 7679 16337
rect 7777 16197 7823 16337
rect 8081 16197 8127 16337
rect 8225 16197 8271 16337
rect 8529 16197 8575 16337
rect 8673 16197 8719 16337
rect 8977 16197 9023 16337
rect 9457 16197 9503 16337
rect 9761 16197 9807 16337
rect 9905 16197 9951 16337
rect 10209 16197 10255 16337
rect 10353 16197 10399 16337
rect 10657 16197 10703 16337
rect 10801 16197 10847 16337
rect 11105 16197 11151 16337
rect 11249 16197 11295 16337
rect 11553 16197 11599 16337
rect 11697 16197 11743 16337
rect 12001 16197 12047 16337
rect 12145 16197 12191 16337
rect 12449 16197 12495 16337
rect 12593 16197 12639 16337
rect 12897 16197 12943 16337
rect 13377 16197 13423 16337
rect 13681 16197 13727 16337
rect 13825 16197 13871 16337
rect 14129 16197 14175 16337
rect 14273 16197 14319 16337
rect 14577 16197 14623 16337
rect 14721 16197 14767 16337
rect 15025 16197 15071 16337
rect 15169 16197 15215 16337
rect 15473 16197 15519 16337
rect 15617 16197 15663 16337
rect 15921 16197 15967 16337
rect 16065 16197 16111 16337
rect 16369 16197 16415 16337
rect 16513 16197 16559 16337
rect 16817 16197 16863 16337
rect 17297 16197 17343 16337
rect 17601 16197 17647 16337
rect 17745 16197 17791 16337
rect 18049 16197 18095 16337
rect 18193 16197 18239 16337
rect 18497 16197 18543 16337
rect 18641 16197 18687 16337
rect 18945 16197 18991 16337
rect 19089 16197 19135 16337
rect 19393 16197 19439 16337
rect 19537 16197 19583 16337
rect 19841 16197 19887 16337
rect 19985 16197 20031 16337
rect 20289 16197 20335 16337
rect 20433 16197 20479 16337
rect 20737 16197 20783 16337
rect 21217 16197 21263 16337
rect 21521 16197 21567 16337
rect 21665 16197 21711 16337
rect 21969 16197 22015 16337
rect 1617 15023 1663 15163
rect 1921 15023 1967 15163
rect 2065 15023 2111 15163
rect 2369 15023 2415 15163
rect 2513 15023 2559 15163
rect 2817 15023 2863 15163
rect 2961 15023 3007 15163
rect 3265 15023 3311 15163
rect 3409 15023 3455 15163
rect 3713 15023 3759 15163
rect 3857 15023 3903 15163
rect 4161 15023 4207 15163
rect 4305 15023 4351 15163
rect 4609 15023 4655 15163
rect 4753 15023 4799 15163
rect 5057 15023 5103 15163
rect 5201 15023 5247 15163
rect 5505 15023 5551 15163
rect 5649 15023 5695 15163
rect 5953 15023 5999 15163
rect 6097 15023 6143 15163
rect 6401 15023 6447 15163
rect 6545 15023 6591 15163
rect 6849 15023 6895 15163
rect 6993 15023 7039 15163
rect 7297 15023 7343 15163
rect 7441 15023 7487 15163
rect 7745 15023 7791 15163
rect 7889 15023 7935 15163
rect 8193 15023 8239 15163
rect 8337 15023 8383 15163
rect 8641 15023 8687 15163
rect 8785 15023 8831 15163
rect 9089 15023 9135 15163
rect 9569 15023 9615 15163
rect 9873 15023 9919 15163
rect 10017 15023 10063 15163
rect 10321 15023 10367 15163
rect 10465 15023 10511 15163
rect 10769 15023 10815 15163
rect 10913 15023 10959 15163
rect 11217 15023 11263 15163
rect 11361 15023 11407 15163
rect 11665 15023 11711 15163
rect 11809 15023 11855 15163
rect 12113 15023 12159 15163
rect 12257 15023 12303 15163
rect 12561 15023 12607 15163
rect 12705 15023 12751 15163
rect 13009 15023 13055 15163
rect 13153 15023 13199 15163
rect 13457 15023 13503 15163
rect 13601 15023 13647 15163
rect 13905 15023 13951 15163
rect 14049 15023 14095 15163
rect 14353 15023 14399 15163
rect 14497 15023 14543 15163
rect 14801 15023 14847 15163
rect 14945 15023 14991 15163
rect 15249 15023 15295 15163
rect 15393 15023 15439 15163
rect 15697 15023 15743 15163
rect 15841 15023 15887 15163
rect 16145 15023 16191 15163
rect 16289 15023 16335 15163
rect 16593 15023 16639 15163
rect 16737 15023 16783 15163
rect 17041 15023 17087 15163
rect 17521 15023 17567 15163
rect 17825 15023 17871 15163
rect 17969 15023 18015 15163
rect 18273 15023 18319 15163
rect 18417 15023 18463 15163
rect 18721 15023 18767 15163
rect 18865 15023 18911 15163
rect 19169 15023 19215 15163
rect 19313 15023 19359 15163
rect 19617 15023 19663 15163
rect 19761 15023 19807 15163
rect 20065 15023 20111 15163
rect 20209 15023 20255 15163
rect 20513 15023 20559 15163
rect 20657 15023 20703 15163
rect 20961 15023 21007 15163
rect 21105 15023 21151 15163
rect 21409 15023 21455 15163
rect 21553 15023 21599 15163
rect 21857 15023 21903 15163
rect 22001 15023 22047 15163
rect 22305 15023 22351 15163
rect 1617 14629 1663 14769
rect 1921 14629 1967 14769
rect 2065 14629 2111 14769
rect 2369 14629 2415 14769
rect 2513 14629 2559 14769
rect 2817 14629 2863 14769
rect 2961 14629 3007 14769
rect 3265 14629 3311 14769
rect 3409 14629 3455 14769
rect 3713 14629 3759 14769
rect 3857 14629 3903 14769
rect 4161 14629 4207 14769
rect 4305 14629 4351 14769
rect 4609 14629 4655 14769
rect 4753 14629 4799 14769
rect 5057 14629 5103 14769
rect 5537 14629 5583 14769
rect 5841 14629 5887 14769
rect 5985 14629 6031 14769
rect 6289 14629 6335 14769
rect 6433 14629 6479 14769
rect 6737 14629 6783 14769
rect 6881 14629 6927 14769
rect 7185 14629 7231 14769
rect 7329 14629 7375 14769
rect 7633 14629 7679 14769
rect 7777 14629 7823 14769
rect 8081 14629 8127 14769
rect 8225 14629 8271 14769
rect 8529 14629 8575 14769
rect 8673 14629 8719 14769
rect 8977 14629 9023 14769
rect 9121 14629 9167 14769
rect 9425 14629 9471 14769
rect 9569 14629 9615 14769
rect 9873 14629 9919 14769
rect 10017 14629 10063 14769
rect 10321 14629 10367 14769
rect 10465 14629 10511 14769
rect 10769 14629 10815 14769
rect 10913 14629 10959 14769
rect 11217 14629 11263 14769
rect 11361 14629 11407 14769
rect 11665 14629 11711 14769
rect 11809 14629 11855 14769
rect 12113 14629 12159 14769
rect 12257 14629 12303 14769
rect 12561 14629 12607 14769
rect 12705 14629 12751 14769
rect 13009 14629 13055 14769
rect 13489 14629 13535 14769
rect 13793 14629 13839 14769
rect 13937 14629 13983 14769
rect 14241 14629 14287 14769
rect 14385 14629 14431 14769
rect 14689 14629 14735 14769
rect 14833 14629 14879 14769
rect 15137 14629 15183 14769
rect 15281 14629 15327 14769
rect 15585 14629 15631 14769
rect 15729 14629 15775 14769
rect 16033 14629 16079 14769
rect 16177 14629 16223 14769
rect 16481 14629 16527 14769
rect 16817 14637 16863 14777
rect 17021 14637 17067 14777
rect 17489 14637 17535 14777
rect 17693 14637 17739 14777
rect 17857 14629 17903 14769
rect 18161 14629 18207 14769
rect 18305 14629 18351 14769
rect 18609 14629 18655 14769
rect 18753 14629 18799 14769
rect 19057 14629 19103 14769
rect 19201 14629 19247 14769
rect 19505 14629 19551 14769
rect 19649 14629 19695 14769
rect 19953 14629 19999 14769
rect 20097 14629 20143 14769
rect 20401 14629 20447 14769
rect 20545 14629 20591 14769
rect 20849 14629 20895 14769
rect 21441 14629 21487 14769
rect 21745 14629 21791 14769
rect 21889 14629 21935 14769
rect 22193 14629 22239 14769
rect 1617 13455 1663 13595
rect 1921 13455 1967 13595
rect 2065 13455 2111 13595
rect 2369 13455 2415 13595
rect 2513 13455 2559 13595
rect 2817 13455 2863 13595
rect 2961 13455 3007 13595
rect 3265 13455 3311 13595
rect 3409 13455 3455 13595
rect 3713 13455 3759 13595
rect 3857 13455 3903 13595
rect 4161 13455 4207 13595
rect 4305 13455 4351 13595
rect 4609 13455 4655 13595
rect 4753 13455 4799 13595
rect 5057 13455 5103 13595
rect 5201 13455 5247 13595
rect 5505 13455 5551 13595
rect 5649 13455 5695 13595
rect 5953 13455 5999 13595
rect 6097 13455 6143 13595
rect 6401 13455 6447 13595
rect 6545 13455 6591 13595
rect 6849 13455 6895 13595
rect 6993 13455 7039 13595
rect 7297 13455 7343 13595
rect 7441 13455 7487 13595
rect 7745 13455 7791 13595
rect 7889 13455 7935 13595
rect 8193 13455 8239 13595
rect 8337 13455 8383 13595
rect 8641 13455 8687 13595
rect 8785 13455 8831 13595
rect 9089 13455 9135 13595
rect 9569 13455 9615 13595
rect 9873 13455 9919 13595
rect 10017 13455 10063 13595
rect 10321 13455 10367 13595
rect 10465 13455 10511 13595
rect 10769 13455 10815 13595
rect 10913 13455 10959 13595
rect 11217 13455 11263 13595
rect 11361 13455 11407 13595
rect 11665 13455 11711 13595
rect 11809 13455 11855 13595
rect 12113 13455 12159 13595
rect 12257 13455 12303 13595
rect 12561 13455 12607 13595
rect 12705 13455 12751 13595
rect 13009 13455 13055 13595
rect 13153 13455 13199 13595
rect 13457 13455 13503 13595
rect 13601 13455 13647 13595
rect 13905 13455 13951 13595
rect 14049 13455 14095 13595
rect 14353 13455 14399 13595
rect 14497 13455 14543 13595
rect 14801 13455 14847 13595
rect 14945 13455 14991 13595
rect 15249 13455 15295 13595
rect 15393 13455 15439 13595
rect 15697 13455 15743 13595
rect 16085 13447 16131 13587
rect 16289 13447 16335 13587
rect 16757 13447 16803 13587
rect 16961 13447 17007 13587
rect 17653 13447 17699 13587
rect 17857 13447 17903 13587
rect 18325 13447 18371 13587
rect 18529 13447 18575 13587
rect 18753 13455 18799 13595
rect 19057 13455 19103 13595
rect 19201 13455 19247 13595
rect 19505 13455 19551 13595
rect 19649 13455 19695 13595
rect 19953 13455 19999 13595
rect 20097 13455 20143 13595
rect 20401 13455 20447 13595
rect 20545 13455 20591 13595
rect 20849 13455 20895 13595
rect 20993 13455 21039 13595
rect 21297 13455 21343 13595
rect 21441 13455 21487 13595
rect 21745 13455 21791 13595
rect 21889 13455 21935 13595
rect 22193 13455 22239 13595
rect 1617 13061 1663 13201
rect 1921 13061 1967 13201
rect 2065 13061 2111 13201
rect 2369 13061 2415 13201
rect 2513 13061 2559 13201
rect 2817 13061 2863 13201
rect 2961 13061 3007 13201
rect 3265 13061 3311 13201
rect 3409 13061 3455 13201
rect 3713 13061 3759 13201
rect 3857 13061 3903 13201
rect 4161 13061 4207 13201
rect 4305 13061 4351 13201
rect 4609 13061 4655 13201
rect 4753 13061 4799 13201
rect 5057 13061 5103 13201
rect 5537 13061 5583 13201
rect 5841 13061 5887 13201
rect 5985 13061 6031 13201
rect 6289 13061 6335 13201
rect 6433 13061 6479 13201
rect 6737 13061 6783 13201
rect 6881 13061 6927 13201
rect 7185 13061 7231 13201
rect 7329 13061 7375 13201
rect 7633 13061 7679 13201
rect 7777 13061 7823 13201
rect 8081 13061 8127 13201
rect 8225 13061 8271 13201
rect 8529 13061 8575 13201
rect 8673 13061 8719 13201
rect 8977 13061 9023 13201
rect 9121 13061 9167 13201
rect 9425 13061 9471 13201
rect 9569 13061 9615 13201
rect 9873 13061 9919 13201
rect 10017 13061 10063 13201
rect 10321 13061 10367 13201
rect 10465 13061 10511 13201
rect 10769 13061 10815 13201
rect 10913 13061 10959 13201
rect 11217 13061 11263 13201
rect 11361 13061 11407 13201
rect 11665 13061 11711 13201
rect 11809 13061 11855 13201
rect 12113 13061 12159 13201
rect 12257 13061 12303 13201
rect 12561 13061 12607 13201
rect 12705 13061 12751 13201
rect 13009 13061 13055 13201
rect 13489 13061 13535 13201
rect 13793 13061 13839 13201
rect 13937 13061 13983 13201
rect 14241 13061 14287 13201
rect 14741 13069 14787 13209
rect 14945 13069 14991 13209
rect 15413 13069 15459 13209
rect 15617 13069 15663 13209
rect 16085 13069 16131 13209
rect 16289 13069 16335 13209
rect 16757 13069 16803 13209
rect 16961 13069 17007 13209
rect 17429 13069 17475 13209
rect 17633 13069 17679 13209
rect 18101 13069 18147 13209
rect 18305 13069 18351 13209
rect 18773 13069 18819 13209
rect 18977 13069 19023 13209
rect 19445 13069 19491 13209
rect 19649 13069 19695 13209
rect 19873 13061 19919 13201
rect 20177 13061 20223 13201
rect 20321 13061 20367 13201
rect 20625 13061 20671 13201
rect 20769 13061 20815 13201
rect 21073 13061 21119 13201
rect 21441 13061 21487 13201
rect 21745 13061 21791 13201
rect 21889 13061 21935 13201
rect 22193 13061 22239 13201
rect 1617 11887 1663 12027
rect 1921 11887 1967 12027
rect 2065 11887 2111 12027
rect 2369 11887 2415 12027
rect 2513 11887 2559 12027
rect 2817 11887 2863 12027
rect 2961 11887 3007 12027
rect 3265 11887 3311 12027
rect 3409 11887 3455 12027
rect 3713 11887 3759 12027
rect 3857 11887 3903 12027
rect 4161 11887 4207 12027
rect 4305 11887 4351 12027
rect 4609 11887 4655 12027
rect 4753 11887 4799 12027
rect 5057 11887 5103 12027
rect 5201 11887 5247 12027
rect 5505 11887 5551 12027
rect 5649 11887 5695 12027
rect 5953 11887 5999 12027
rect 6097 11887 6143 12027
rect 6401 11887 6447 12027
rect 6545 11887 6591 12027
rect 6849 11887 6895 12027
rect 6993 11887 7039 12027
rect 7297 11887 7343 12027
rect 7441 11887 7487 12027
rect 7745 11887 7791 12027
rect 7889 11887 7935 12027
rect 8193 11887 8239 12027
rect 8337 11887 8383 12027
rect 8641 11887 8687 12027
rect 8785 11887 8831 12027
rect 9089 11887 9135 12027
rect 9569 11887 9615 12027
rect 9873 11887 9919 12027
rect 10017 11887 10063 12027
rect 10321 11887 10367 12027
rect 10465 11887 10511 12027
rect 10769 11887 10815 12027
rect 10913 11887 10959 12027
rect 11217 11887 11263 12027
rect 11361 11887 11407 12027
rect 11665 11887 11711 12027
rect 11809 11887 11855 12027
rect 12113 11887 12159 12027
rect 12257 11887 12303 12027
rect 12561 11887 12607 12027
rect 12705 11887 12751 12027
rect 13009 11887 13055 12027
rect 13153 11887 13199 12027
rect 13457 11887 13503 12027
rect 13601 11887 13647 12027
rect 13905 11887 13951 12027
rect 14069 11879 14115 12019
rect 14273 11879 14319 12019
rect 14741 11879 14787 12019
rect 14945 11879 14991 12019
rect 15413 11879 15459 12019
rect 15617 11879 15663 12019
rect 16085 11879 16131 12019
rect 16289 11879 16335 12019
rect 16757 11879 16803 12019
rect 16961 11879 17007 12019
rect 17653 11879 17699 12019
rect 17857 11879 17903 12019
rect 18325 11879 18371 12019
rect 18529 11879 18575 12019
rect 18997 11879 19043 12019
rect 19201 11879 19247 12019
rect 19669 11879 19715 12019
rect 19873 11879 19919 12019
rect 20341 11879 20387 12019
rect 20545 11879 20591 12019
rect 20769 11887 20815 12027
rect 21073 11887 21119 12027
rect 21217 11887 21263 12027
rect 21521 11887 21567 12027
rect 21665 11887 21711 12027
rect 21969 11887 22015 12027
rect 1617 11493 1663 11633
rect 1921 11493 1967 11633
rect 2065 11493 2111 11633
rect 2369 11493 2415 11633
rect 2513 11493 2559 11633
rect 2817 11493 2863 11633
rect 2961 11493 3007 11633
rect 3265 11493 3311 11633
rect 3409 11493 3455 11633
rect 3713 11493 3759 11633
rect 3857 11493 3903 11633
rect 4161 11493 4207 11633
rect 4305 11493 4351 11633
rect 4609 11493 4655 11633
rect 4753 11493 4799 11633
rect 5057 11493 5103 11633
rect 5537 11493 5583 11633
rect 5841 11493 5887 11633
rect 6065 11501 6111 11641
rect 6269 11501 6315 11641
rect 6849 11501 6895 11641
rect 7053 11501 7099 11641
rect 7521 11501 7567 11641
rect 7725 11501 7771 11641
rect 8193 11501 8239 11641
rect 8397 11501 8443 11641
rect 8561 11493 8607 11633
rect 8865 11493 8911 11633
rect 9141 11501 9187 11641
rect 9345 11501 9391 11641
rect 9813 11501 9859 11641
rect 10017 11501 10063 11641
rect 10485 11501 10531 11641
rect 10689 11501 10735 11641
rect 10913 11493 10959 11633
rect 11217 11493 11263 11633
rect 11361 11493 11407 11633
rect 11665 11493 11711 11633
rect 12053 11501 12099 11641
rect 12257 11501 12303 11641
rect 12725 11501 12771 11641
rect 12929 11501 12975 11641
rect 13621 11501 13667 11641
rect 13825 11501 13871 11641
rect 14049 11493 14095 11633
rect 14353 11493 14399 11633
rect 14741 11501 14787 11641
rect 14945 11501 14991 11641
rect 15413 11501 15459 11641
rect 15617 11501 15663 11641
rect 16085 11501 16131 11641
rect 16289 11501 16335 11641
rect 16757 11501 16803 11641
rect 16961 11501 17007 11641
rect 17429 11501 17475 11641
rect 17633 11501 17679 11641
rect 18101 11501 18147 11641
rect 18305 11501 18351 11641
rect 18773 11501 18819 11641
rect 18977 11501 19023 11641
rect 19445 11501 19491 11641
rect 19649 11501 19695 11641
rect 20117 11501 20163 11641
rect 20321 11501 20367 11641
rect 20545 11493 20591 11633
rect 20849 11493 20895 11633
rect 21441 11493 21487 11633
rect 21745 11493 21791 11633
rect 21889 11493 21935 11633
rect 22193 11493 22239 11633
rect 1617 10319 1663 10459
rect 1921 10319 1967 10459
rect 2065 10319 2111 10459
rect 2369 10319 2415 10459
rect 2513 10319 2559 10459
rect 2817 10319 2863 10459
rect 2961 10319 3007 10459
rect 3265 10319 3311 10459
rect 3409 10319 3455 10459
rect 3713 10319 3759 10459
rect 3857 10319 3903 10459
rect 4161 10319 4207 10459
rect 4305 10319 4351 10459
rect 4609 10319 4655 10459
rect 4753 10319 4799 10459
rect 5057 10319 5103 10459
rect 5333 10311 5379 10451
rect 5537 10311 5583 10451
rect 6005 10311 6051 10451
rect 6209 10311 6255 10451
rect 6677 10311 6723 10451
rect 6881 10311 6927 10451
rect 7349 10311 7395 10451
rect 7553 10311 7599 10451
rect 8021 10311 8067 10451
rect 8225 10311 8271 10451
rect 8805 10311 8851 10451
rect 9009 10311 9055 10451
rect 9813 10311 9859 10451
rect 10017 10311 10063 10451
rect 10485 10311 10531 10451
rect 10689 10311 10735 10451
rect 11157 10311 11203 10451
rect 11361 10311 11407 10451
rect 11941 10311 11987 10451
rect 12145 10311 12191 10451
rect 12613 10311 12659 10451
rect 12817 10311 12863 10451
rect 13285 10311 13331 10451
rect 13489 10311 13535 10451
rect 13957 10311 14003 10451
rect 14161 10311 14207 10451
rect 14629 10311 14675 10451
rect 14833 10311 14879 10451
rect 15301 10311 15347 10451
rect 15505 10311 15551 10451
rect 15973 10311 16019 10451
rect 16177 10311 16223 10451
rect 16645 10311 16691 10451
rect 16849 10311 16895 10451
rect 17653 10311 17699 10451
rect 17857 10311 17903 10451
rect 18325 10311 18371 10451
rect 18529 10311 18575 10451
rect 18997 10311 19043 10451
rect 19201 10311 19247 10451
rect 19669 10311 19715 10451
rect 19873 10311 19919 10451
rect 20341 10311 20387 10451
rect 20545 10311 20591 10451
rect 21013 10311 21059 10451
rect 21217 10311 21263 10451
rect 21685 10311 21731 10451
rect 21889 10311 21935 10451
rect 1617 9925 1663 10065
rect 1921 9925 1967 10065
rect 2065 9925 2111 10065
rect 2369 9925 2415 10065
rect 2513 9925 2559 10065
rect 2817 9925 2863 10065
rect 2961 9925 3007 10065
rect 3265 9925 3311 10065
rect 3409 9925 3455 10065
rect 3713 9925 3759 10065
rect 4101 9933 4147 10073
rect 4305 9933 4351 10073
rect 4773 9933 4819 10073
rect 4977 9933 5023 10073
rect 5781 9933 5827 10073
rect 5985 9933 6031 10073
rect 6453 9933 6499 10073
rect 6657 9933 6703 10073
rect 7125 9933 7171 10073
rect 7329 9933 7375 10073
rect 7797 9933 7843 10073
rect 8001 9933 8047 10073
rect 8469 9933 8515 10073
rect 8673 9933 8719 10073
rect 9141 9933 9187 10073
rect 9345 9933 9391 10073
rect 9813 9933 9859 10073
rect 10017 9933 10063 10073
rect 10485 9933 10531 10073
rect 10689 9933 10735 10073
rect 10913 9925 10959 10065
rect 11217 9925 11263 10065
rect 11381 9933 11427 10073
rect 11585 9933 11631 10073
rect 12053 9933 12099 10073
rect 12257 9933 12303 10073
rect 12725 9933 12771 10073
rect 12929 9933 12975 10073
rect 13621 9933 13667 10073
rect 13825 9933 13871 10073
rect 14293 9933 14339 10073
rect 14497 9933 14543 10073
rect 14965 9933 15011 10073
rect 15169 9933 15215 10073
rect 15637 9933 15683 10073
rect 15841 9933 15887 10073
rect 16309 9933 16355 10073
rect 16513 9933 16559 10073
rect 16981 9933 17027 10073
rect 17185 9933 17231 10073
rect 17713 9933 17759 10073
rect 17917 9933 17963 10073
rect 18325 9933 18371 10073
rect 18529 9933 18575 10073
rect 18997 9933 19043 10073
rect 19201 9933 19247 10073
rect 19669 9933 19715 10073
rect 19873 9933 19919 10073
rect 20341 9933 20387 10073
rect 20545 9933 20591 10073
rect 20769 9925 20815 10065
rect 21073 9925 21119 10065
rect 21573 9933 21619 10073
rect 21777 9933 21823 10073
rect 22001 9925 22047 10065
rect 22305 9925 22351 10065
rect 1617 8751 1663 8891
rect 1921 8751 1967 8891
rect 2065 8751 2111 8891
rect 2369 8751 2415 8891
rect 2513 8751 2559 8891
rect 2817 8751 2863 8891
rect 3317 8743 3363 8883
rect 3521 8743 3567 8883
rect 3989 8743 4035 8883
rect 4193 8743 4239 8883
rect 4661 8743 4707 8883
rect 4865 8743 4911 8883
rect 5333 8743 5379 8883
rect 5537 8743 5583 8883
rect 6005 8743 6051 8883
rect 6209 8743 6255 8883
rect 6677 8743 6723 8883
rect 6881 8743 6927 8883
rect 7349 8743 7395 8883
rect 7553 8743 7599 8883
rect 8133 8743 8179 8883
rect 8337 8743 8383 8883
rect 8805 8743 8851 8883
rect 9009 8743 9055 8883
rect 9569 8751 9615 8891
rect 9873 8751 9919 8891
rect 10261 8743 10307 8883
rect 10465 8743 10511 8883
rect 10933 8743 10979 8883
rect 11137 8743 11183 8883
rect 11605 8743 11651 8883
rect 11809 8743 11855 8883
rect 12277 8743 12323 8883
rect 12481 8743 12527 8883
rect 12949 8743 12995 8883
rect 13153 8743 13199 8883
rect 13621 8743 13667 8883
rect 13825 8743 13871 8883
rect 14293 8743 14339 8883
rect 14497 8743 14543 8883
rect 14965 8743 15011 8883
rect 15169 8743 15215 8883
rect 15637 8743 15683 8883
rect 15841 8743 15887 8883
rect 16309 8743 16355 8883
rect 16513 8743 16559 8883
rect 16737 8751 16783 8891
rect 17041 8751 17087 8891
rect 17653 8743 17699 8883
rect 17857 8743 17903 8883
rect 18325 8743 18371 8883
rect 18529 8743 18575 8883
rect 18997 8743 19043 8883
rect 19201 8743 19247 8883
rect 19669 8743 19715 8883
rect 19873 8743 19919 8883
rect 20341 8743 20387 8883
rect 20545 8743 20591 8883
rect 20769 8751 20815 8891
rect 21073 8751 21119 8891
rect 21217 8751 21263 8891
rect 21521 8751 21567 8891
rect 21665 8751 21711 8891
rect 21969 8751 22015 8891
rect 1617 8357 1663 8497
rect 1921 8357 1967 8497
rect 2065 8357 2111 8497
rect 2369 8357 2415 8497
rect 2817 8365 2863 8505
rect 3021 8365 3067 8505
rect 3429 8365 3475 8505
rect 3633 8365 3679 8505
rect 4101 8365 4147 8505
rect 4305 8365 4351 8505
rect 4773 8365 4819 8505
rect 4977 8365 5023 8505
rect 5781 8365 5827 8505
rect 5985 8365 6031 8505
rect 6453 8365 6499 8505
rect 6657 8365 6703 8505
rect 7125 8365 7171 8505
rect 7329 8365 7375 8505
rect 7797 8365 7843 8505
rect 8001 8365 8047 8505
rect 8469 8365 8515 8505
rect 8673 8365 8719 8505
rect 9141 8365 9187 8505
rect 9345 8365 9391 8505
rect 9813 8365 9859 8505
rect 10017 8365 10063 8505
rect 10485 8365 10531 8505
rect 10689 8365 10735 8505
rect 11217 8365 11263 8505
rect 11421 8365 11467 8505
rect 11585 8357 11631 8497
rect 11889 8357 11935 8497
rect 12053 8365 12099 8505
rect 12257 8365 12303 8505
rect 12725 8365 12771 8505
rect 12929 8365 12975 8505
rect 13621 8365 13667 8505
rect 13825 8365 13871 8505
rect 14293 8365 14339 8505
rect 14497 8365 14543 8505
rect 14965 8365 15011 8505
rect 15169 8365 15215 8505
rect 15637 8365 15683 8505
rect 15841 8365 15887 8505
rect 16309 8365 16355 8505
rect 16513 8365 16559 8505
rect 16981 8365 17027 8505
rect 17185 8365 17231 8505
rect 17653 8365 17699 8505
rect 17857 8365 17903 8505
rect 18325 8365 18371 8505
rect 18529 8365 18575 8505
rect 18997 8365 19043 8505
rect 19201 8365 19247 8505
rect 19669 8365 19715 8505
rect 19873 8365 19919 8505
rect 20401 8365 20447 8505
rect 20605 8365 20651 8505
rect 20769 8357 20815 8497
rect 21073 8357 21119 8497
rect 21441 8357 21487 8497
rect 21745 8357 21791 8497
rect 21889 8357 21935 8497
rect 22193 8357 22239 8497
rect 2033 7175 2079 7315
rect 2237 7175 2283 7315
rect 2645 7175 2691 7315
rect 2849 7175 2895 7315
rect 3317 7175 3363 7315
rect 3521 7175 3567 7315
rect 3989 7175 4035 7315
rect 4193 7175 4239 7315
rect 4661 7175 4707 7315
rect 4865 7175 4911 7315
rect 5333 7175 5379 7315
rect 5537 7175 5583 7315
rect 6005 7175 6051 7315
rect 6209 7175 6255 7315
rect 6677 7175 6723 7315
rect 6881 7175 6927 7315
rect 7349 7175 7395 7315
rect 7553 7175 7599 7315
rect 8133 7175 8179 7315
rect 8337 7175 8383 7315
rect 8805 7175 8851 7315
rect 9009 7175 9055 7315
rect 9813 7175 9859 7315
rect 10017 7175 10063 7315
rect 10485 7175 10531 7315
rect 10689 7175 10735 7315
rect 11217 7175 11263 7315
rect 11421 7175 11467 7315
rect 11829 7175 11875 7315
rect 12033 7175 12079 7315
rect 12501 7175 12547 7315
rect 12705 7175 12751 7315
rect 13173 7175 13219 7315
rect 13377 7175 13423 7315
rect 13845 7175 13891 7315
rect 14049 7175 14095 7315
rect 14517 7175 14563 7315
rect 14721 7175 14767 7315
rect 15189 7175 15235 7315
rect 15393 7175 15439 7315
rect 15861 7175 15907 7315
rect 16065 7175 16111 7315
rect 16533 7175 16579 7315
rect 16737 7175 16783 7315
rect 17653 7175 17699 7315
rect 17857 7175 17903 7315
rect 18325 7175 18371 7315
rect 18529 7175 18575 7315
rect 18997 7175 19043 7315
rect 19201 7175 19247 7315
rect 19669 7175 19715 7315
rect 19873 7175 19919 7315
rect 20341 7175 20387 7315
rect 20545 7175 20591 7315
rect 21013 7175 21059 7315
rect 21217 7175 21263 7315
rect 21441 7183 21487 7323
rect 21745 7183 21791 7323
rect 21889 7183 21935 7323
rect 22193 7183 22239 7323
rect 1617 6789 1663 6929
rect 1921 6789 1967 6929
rect 2085 6797 2131 6937
rect 2289 6797 2335 6937
rect 2757 6797 2803 6937
rect 2961 6797 3007 6937
rect 3429 6797 3475 6937
rect 3633 6797 3679 6937
rect 4101 6797 4147 6937
rect 4305 6797 4351 6937
rect 4773 6797 4819 6937
rect 4977 6797 5023 6937
rect 5669 6797 5715 6937
rect 5873 6797 5919 6937
rect 6341 6797 6387 6937
rect 6545 6797 6591 6937
rect 7013 6797 7059 6937
rect 7217 6797 7263 6937
rect 7685 6797 7731 6937
rect 7889 6797 7935 6937
rect 8357 6797 8403 6937
rect 8561 6797 8607 6937
rect 9029 6797 9075 6937
rect 9233 6797 9279 6937
rect 9701 6797 9747 6937
rect 9905 6797 9951 6937
rect 10373 6797 10419 6937
rect 10577 6797 10623 6937
rect 11045 6797 11091 6937
rect 11249 6797 11295 6937
rect 11717 6797 11763 6937
rect 11921 6797 11967 6937
rect 12389 6797 12435 6937
rect 12593 6797 12639 6937
rect 12817 6789 12863 6929
rect 13121 6789 13167 6929
rect 13489 6789 13535 6929
rect 13793 6789 13839 6929
rect 14069 6797 14115 6937
rect 14273 6797 14319 6937
rect 14741 6797 14787 6937
rect 14945 6797 14991 6937
rect 15413 6797 15459 6937
rect 15617 6797 15663 6937
rect 16085 6797 16131 6937
rect 16289 6797 16335 6937
rect 16757 6797 16803 6937
rect 16961 6797 17007 6937
rect 17429 6797 17475 6937
rect 17633 6797 17679 6937
rect 18101 6797 18147 6937
rect 18305 6797 18351 6937
rect 18773 6797 18819 6937
rect 18977 6797 19023 6937
rect 19445 6797 19491 6937
rect 19649 6797 19695 6937
rect 20177 6797 20223 6937
rect 20381 6797 20427 6937
rect 20545 6789 20591 6929
rect 20849 6789 20895 6929
rect 21573 6797 21619 6937
rect 21777 6797 21823 6937
rect 22001 6789 22047 6929
rect 22305 6789 22351 6929
rect 1973 5607 2019 5747
rect 2177 5607 2223 5747
rect 2645 5607 2691 5747
rect 2849 5607 2895 5747
rect 3317 5607 3363 5747
rect 3521 5607 3567 5747
rect 3989 5607 4035 5747
rect 4193 5607 4239 5747
rect 4661 5607 4707 5747
rect 4865 5607 4911 5747
rect 5333 5607 5379 5747
rect 5537 5607 5583 5747
rect 6005 5607 6051 5747
rect 6209 5607 6255 5747
rect 6677 5607 6723 5747
rect 6881 5607 6927 5747
rect 7349 5607 7395 5747
rect 7553 5607 7599 5747
rect 8021 5607 8067 5747
rect 8225 5607 8271 5747
rect 8693 5607 8739 5747
rect 8897 5607 8943 5747
rect 9701 5607 9747 5747
rect 9905 5607 9951 5747
rect 10373 5607 10419 5747
rect 10577 5607 10623 5747
rect 11045 5607 11091 5747
rect 11249 5607 11295 5747
rect 11717 5607 11763 5747
rect 11921 5607 11967 5747
rect 12501 5607 12547 5747
rect 12705 5607 12751 5747
rect 13173 5607 13219 5747
rect 13377 5607 13423 5747
rect 13845 5607 13891 5747
rect 14049 5607 14095 5747
rect 14517 5607 14563 5747
rect 14721 5607 14767 5747
rect 15189 5607 15235 5747
rect 15393 5607 15439 5747
rect 15861 5607 15907 5747
rect 16065 5607 16111 5747
rect 16533 5607 16579 5747
rect 16737 5607 16783 5747
rect 17653 5607 17699 5747
rect 17857 5607 17903 5747
rect 18325 5607 18371 5747
rect 18529 5607 18575 5747
rect 18997 5607 19043 5747
rect 19201 5607 19247 5747
rect 19669 5607 19715 5747
rect 19873 5607 19919 5747
rect 20341 5607 20387 5747
rect 20545 5607 20591 5747
rect 21013 5607 21059 5747
rect 21217 5607 21263 5747
rect 21745 5607 21791 5747
rect 21949 5607 21995 5747
rect 1617 5221 1663 5361
rect 1921 5221 1967 5361
rect 2085 5229 2131 5369
rect 2289 5229 2335 5369
rect 2757 5229 2803 5369
rect 2961 5229 3007 5369
rect 3429 5229 3475 5369
rect 3633 5229 3679 5369
rect 4101 5229 4147 5369
rect 4305 5229 4351 5369
rect 4773 5229 4819 5369
rect 4977 5229 5023 5369
rect 5669 5229 5715 5369
rect 5873 5229 5919 5369
rect 6341 5229 6387 5369
rect 6545 5229 6591 5369
rect 7013 5229 7059 5369
rect 7217 5229 7263 5369
rect 7685 5229 7731 5369
rect 7889 5229 7935 5369
rect 8357 5229 8403 5369
rect 8561 5229 8607 5369
rect 9029 5229 9075 5369
rect 9233 5229 9279 5369
rect 9701 5229 9747 5369
rect 9905 5229 9951 5369
rect 10373 5229 10419 5369
rect 10577 5229 10623 5369
rect 10801 5221 10847 5361
rect 11105 5221 11151 5361
rect 11381 5229 11427 5369
rect 11585 5229 11631 5369
rect 12053 5229 12099 5369
rect 12257 5229 12303 5369
rect 12725 5229 12771 5369
rect 12929 5229 12975 5369
rect 13489 5221 13535 5361
rect 13793 5221 13839 5361
rect 13957 5229 14003 5369
rect 14161 5229 14207 5369
rect 14629 5229 14675 5369
rect 14833 5229 14879 5369
rect 15301 5229 15347 5369
rect 15505 5229 15551 5369
rect 15973 5229 16019 5369
rect 16177 5229 16223 5369
rect 16645 5229 16691 5369
rect 16849 5229 16895 5369
rect 17317 5229 17363 5369
rect 17521 5229 17567 5369
rect 17989 5229 18035 5369
rect 18193 5229 18239 5369
rect 18661 5229 18707 5369
rect 18865 5229 18911 5369
rect 19333 5229 19379 5369
rect 19537 5229 19583 5369
rect 20005 5229 20051 5369
rect 20209 5229 20255 5369
rect 20677 5229 20723 5369
rect 20881 5229 20927 5369
rect 21573 5229 21619 5369
rect 21777 5229 21823 5369
rect 22001 5221 22047 5361
rect 22305 5221 22351 5361
rect 1617 4047 1663 4187
rect 1921 4047 1967 4187
rect 2309 4039 2355 4179
rect 2513 4039 2559 4179
rect 2981 4039 3027 4179
rect 3185 4039 3231 4179
rect 3653 4039 3699 4179
rect 3857 4039 3903 4179
rect 4325 4039 4371 4179
rect 4529 4039 4575 4179
rect 4997 4039 5043 4179
rect 5201 4039 5247 4179
rect 5669 4039 5715 4179
rect 5873 4039 5919 4179
rect 6341 4039 6387 4179
rect 6545 4039 6591 4179
rect 7013 4039 7059 4179
rect 7217 4039 7263 4179
rect 7685 4039 7731 4179
rect 7889 4039 7935 4179
rect 8357 4039 8403 4179
rect 8561 4039 8607 4179
rect 8785 4047 8831 4187
rect 9089 4047 9135 4187
rect 9701 4039 9747 4179
rect 9905 4039 9951 4179
rect 10373 4039 10419 4179
rect 10577 4039 10623 4179
rect 11045 4039 11091 4179
rect 11249 4039 11295 4179
rect 11473 4047 11519 4187
rect 11777 4047 11823 4187
rect 12277 4039 12323 4179
rect 12481 4039 12527 4179
rect 12949 4039 12995 4179
rect 13153 4039 13199 4179
rect 13621 4039 13667 4179
rect 13825 4039 13871 4179
rect 14293 4039 14339 4179
rect 14497 4039 14543 4179
rect 14965 4039 15011 4179
rect 15169 4039 15215 4179
rect 15637 4039 15683 4179
rect 15841 4039 15887 4179
rect 16309 4039 16355 4179
rect 16513 4039 16559 4179
rect 16737 4047 16783 4187
rect 17041 4047 17087 4187
rect 17653 4039 17699 4179
rect 17857 4039 17903 4179
rect 18325 4039 18371 4179
rect 18529 4039 18575 4179
rect 18997 4039 19043 4179
rect 19201 4039 19247 4179
rect 19669 4039 19715 4179
rect 19873 4039 19919 4179
rect 20341 4039 20387 4179
rect 20545 4039 20591 4179
rect 21013 4039 21059 4179
rect 21217 4039 21263 4179
rect 21745 4039 21791 4179
rect 21949 4039 21995 4179
rect 1617 3653 1663 3793
rect 1921 3653 1967 3793
rect 2065 3653 2111 3793
rect 2369 3653 2415 3793
rect 2757 3661 2803 3801
rect 2961 3661 3007 3801
rect 3429 3661 3475 3801
rect 3633 3661 3679 3801
rect 4101 3661 4147 3801
rect 4305 3661 4351 3801
rect 4773 3661 4819 3801
rect 4977 3661 5023 3801
rect 5729 3661 5775 3801
rect 5933 3661 5979 3801
rect 6401 3661 6447 3801
rect 6605 3661 6651 3801
rect 7073 3661 7119 3801
rect 7277 3661 7323 3801
rect 7685 3661 7731 3801
rect 7889 3661 7935 3801
rect 8417 3661 8463 3801
rect 8621 3661 8667 3801
rect 8785 3653 8831 3793
rect 9089 3653 9135 3793
rect 9649 3661 9695 3801
rect 9853 3661 9899 3801
rect 10261 3661 10307 3801
rect 10465 3661 10511 3801
rect 10933 3661 10979 3801
rect 11137 3661 11183 3801
rect 11665 3661 11711 3801
rect 11869 3661 11915 3801
rect 12033 3653 12079 3793
rect 12337 3653 12383 3793
rect 12481 3653 12527 3793
rect 12785 3653 12831 3793
rect 13377 3653 13423 3793
rect 13681 3653 13727 3793
rect 13845 3661 13891 3801
rect 14049 3661 14095 3801
rect 14517 3661 14563 3801
rect 14721 3661 14767 3801
rect 15189 3661 15235 3801
rect 15393 3661 15439 3801
rect 15861 3661 15907 3801
rect 16065 3661 16111 3801
rect 16533 3661 16579 3801
rect 16737 3661 16783 3801
rect 17429 3661 17475 3801
rect 17633 3661 17679 3801
rect 18101 3661 18147 3801
rect 18305 3661 18351 3801
rect 18773 3661 18819 3801
rect 18977 3661 19023 3801
rect 19445 3661 19491 3801
rect 19649 3661 19695 3801
rect 20117 3661 20163 3801
rect 20321 3661 20367 3801
rect 20545 3653 20591 3793
rect 20849 3653 20895 3793
rect 21217 3653 21263 3793
rect 21521 3653 21567 3793
rect 21665 3653 21711 3793
rect 21969 3653 22015 3793
<< mvpsubdiff >>
rect 1400 15906 1504 15936
rect 1400 15759 1429 15906
rect 1475 15759 1504 15906
rect 1400 15736 1504 15759
rect 5320 15906 5432 15936
rect 5320 15759 5353 15906
rect 5399 15759 5432 15906
rect 5320 15736 5432 15759
rect 9240 15906 9352 15936
rect 9240 15759 9273 15906
rect 9319 15759 9352 15906
rect 9240 15736 9352 15759
rect 13160 15906 13272 15936
rect 13160 15759 13193 15906
rect 13239 15759 13272 15906
rect 13160 15736 13272 15759
rect 17080 15906 17192 15936
rect 17080 15759 17113 15906
rect 17159 15759 17192 15906
rect 17080 15736 17192 15759
rect 21000 15906 21112 15936
rect 21000 15759 21033 15906
rect 21079 15759 21112 15906
rect 21000 15736 21112 15759
rect 22464 15906 22568 15936
rect 22464 15759 22493 15906
rect 22539 15759 22568 15906
rect 22464 15736 22568 15759
rect 1400 15601 1504 15624
rect 1400 15454 1429 15601
rect 1475 15454 1504 15601
rect 1400 15424 1504 15454
rect 9352 15601 9464 15624
rect 9352 15454 9385 15601
rect 9431 15454 9464 15601
rect 9352 15424 9464 15454
rect 17304 15601 17416 15624
rect 17304 15454 17337 15601
rect 17383 15454 17416 15601
rect 17304 15424 17416 15454
rect 22464 15601 22568 15624
rect 22464 15454 22493 15601
rect 22539 15454 22568 15601
rect 22464 15424 22568 15454
rect 1400 14338 1504 14368
rect 1400 14191 1429 14338
rect 1475 14191 1504 14338
rect 1400 14168 1504 14191
rect 5320 14338 5432 14368
rect 5320 14191 5353 14338
rect 5399 14191 5432 14338
rect 5320 14168 5432 14191
rect 13272 14338 13384 14368
rect 13272 14191 13305 14338
rect 13351 14191 13384 14338
rect 13272 14168 13384 14191
rect 21224 14338 21336 14368
rect 21224 14191 21257 14338
rect 21303 14191 21336 14338
rect 21224 14168 21336 14191
rect 22464 14338 22568 14368
rect 22464 14191 22493 14338
rect 22539 14191 22568 14338
rect 22464 14168 22568 14191
rect 1400 14033 1504 14056
rect 1400 13886 1429 14033
rect 1475 13886 1504 14033
rect 1400 13856 1504 13886
rect 9352 14033 9464 14056
rect 9352 13886 9385 14033
rect 9431 13886 9464 14033
rect 9352 13856 9464 13886
rect 17304 14033 17416 14056
rect 17304 13886 17337 14033
rect 17383 13886 17416 14033
rect 17304 13856 17416 13886
rect 22464 14033 22568 14056
rect 22464 13886 22493 14033
rect 22539 13886 22568 14033
rect 22464 13856 22568 13886
rect 1400 12770 1504 12800
rect 1400 12623 1429 12770
rect 1475 12623 1504 12770
rect 1400 12600 1504 12623
rect 5320 12770 5432 12800
rect 5320 12623 5353 12770
rect 5399 12623 5432 12770
rect 5320 12600 5432 12623
rect 13272 12770 13384 12800
rect 13272 12623 13305 12770
rect 13351 12623 13384 12770
rect 13272 12600 13384 12623
rect 21224 12770 21336 12800
rect 21224 12623 21257 12770
rect 21303 12623 21336 12770
rect 21224 12600 21336 12623
rect 22464 12770 22568 12800
rect 22464 12623 22493 12770
rect 22539 12623 22568 12770
rect 22464 12600 22568 12623
rect 1400 12465 1504 12488
rect 1400 12318 1429 12465
rect 1475 12318 1504 12465
rect 1400 12288 1504 12318
rect 9352 12465 9464 12488
rect 9352 12318 9385 12465
rect 9431 12318 9464 12465
rect 9352 12288 9464 12318
rect 17304 12465 17416 12488
rect 17304 12318 17337 12465
rect 17383 12318 17416 12465
rect 17304 12288 17416 12318
rect 22464 12465 22568 12488
rect 22464 12318 22493 12465
rect 22539 12318 22568 12465
rect 22464 12288 22568 12318
rect 1400 11202 1504 11232
rect 1400 11055 1429 11202
rect 1475 11055 1504 11202
rect 1400 11032 1504 11055
rect 5320 11202 5432 11232
rect 5320 11055 5353 11202
rect 5399 11055 5432 11202
rect 5320 11032 5432 11055
rect 13272 11202 13384 11232
rect 13272 11055 13305 11202
rect 13351 11055 13384 11202
rect 13272 11032 13384 11055
rect 21224 11202 21336 11232
rect 21224 11055 21257 11202
rect 21303 11055 21336 11202
rect 21224 11032 21336 11055
rect 22464 11202 22568 11232
rect 22464 11055 22493 11202
rect 22539 11055 22568 11202
rect 22464 11032 22568 11055
rect 1400 10897 1504 10920
rect 1400 10750 1429 10897
rect 1475 10750 1504 10897
rect 1400 10720 1504 10750
rect 9352 10897 9464 10920
rect 9352 10750 9385 10897
rect 9431 10750 9464 10897
rect 9352 10720 9464 10750
rect 17304 10897 17416 10920
rect 17304 10750 17337 10897
rect 17383 10750 17416 10897
rect 17304 10720 17416 10750
rect 22464 10897 22568 10920
rect 22464 10750 22493 10897
rect 22539 10750 22568 10897
rect 22464 10720 22568 10750
rect 1400 9634 1504 9664
rect 1400 9487 1429 9634
rect 1475 9487 1504 9634
rect 1400 9464 1504 9487
rect 5320 9634 5432 9664
rect 5320 9487 5353 9634
rect 5399 9487 5432 9634
rect 5320 9464 5432 9487
rect 13272 9634 13384 9664
rect 13272 9487 13305 9634
rect 13351 9487 13384 9634
rect 13272 9464 13384 9487
rect 21224 9634 21336 9664
rect 21224 9487 21257 9634
rect 21303 9487 21336 9634
rect 21224 9464 21336 9487
rect 22464 9634 22568 9664
rect 22464 9487 22493 9634
rect 22539 9487 22568 9634
rect 22464 9464 22568 9487
rect 1400 9329 1504 9352
rect 1400 9182 1429 9329
rect 1475 9182 1504 9329
rect 1400 9152 1504 9182
rect 9352 9329 9464 9352
rect 9352 9182 9385 9329
rect 9431 9182 9464 9329
rect 9352 9152 9464 9182
rect 17304 9329 17416 9352
rect 17304 9182 17337 9329
rect 17383 9182 17416 9329
rect 17304 9152 17416 9182
rect 22464 9329 22568 9352
rect 22464 9182 22493 9329
rect 22539 9182 22568 9329
rect 22464 9152 22568 9182
rect 1400 8066 1504 8096
rect 1400 7919 1429 8066
rect 1475 7919 1504 8066
rect 1400 7896 1504 7919
rect 5320 8066 5432 8096
rect 5320 7919 5353 8066
rect 5399 7919 5432 8066
rect 5320 7896 5432 7919
rect 13272 8066 13384 8096
rect 13272 7919 13305 8066
rect 13351 7919 13384 8066
rect 13272 7896 13384 7919
rect 21224 8066 21336 8096
rect 21224 7919 21257 8066
rect 21303 7919 21336 8066
rect 21224 7896 21336 7919
rect 22464 8066 22568 8096
rect 22464 7919 22493 8066
rect 22539 7919 22568 8066
rect 22464 7896 22568 7919
rect 1400 7761 1504 7784
rect 1400 7614 1429 7761
rect 1475 7614 1504 7761
rect 1400 7584 1504 7614
rect 9352 7761 9464 7784
rect 9352 7614 9385 7761
rect 9431 7614 9464 7761
rect 9352 7584 9464 7614
rect 17304 7761 17416 7784
rect 17304 7614 17337 7761
rect 17383 7614 17416 7761
rect 17304 7584 17416 7614
rect 22464 7761 22568 7784
rect 22464 7614 22493 7761
rect 22539 7614 22568 7761
rect 22464 7584 22568 7614
rect 1400 6498 1504 6528
rect 1400 6351 1429 6498
rect 1475 6351 1504 6498
rect 1400 6328 1504 6351
rect 5320 6498 5432 6528
rect 5320 6351 5353 6498
rect 5399 6351 5432 6498
rect 5320 6328 5432 6351
rect 13272 6498 13384 6528
rect 13272 6351 13305 6498
rect 13351 6351 13384 6498
rect 13272 6328 13384 6351
rect 21224 6498 21336 6528
rect 21224 6351 21257 6498
rect 21303 6351 21336 6498
rect 21224 6328 21336 6351
rect 22464 6498 22568 6528
rect 22464 6351 22493 6498
rect 22539 6351 22568 6498
rect 22464 6328 22568 6351
rect 1400 6193 1504 6216
rect 1400 6046 1429 6193
rect 1475 6046 1504 6193
rect 1400 6016 1504 6046
rect 9352 6193 9464 6216
rect 9352 6046 9385 6193
rect 9431 6046 9464 6193
rect 9352 6016 9464 6046
rect 17304 6193 17416 6216
rect 17304 6046 17337 6193
rect 17383 6046 17416 6193
rect 17304 6016 17416 6046
rect 22464 6193 22568 6216
rect 22464 6046 22493 6193
rect 22539 6046 22568 6193
rect 22464 6016 22568 6046
rect 1400 4930 1504 4960
rect 1400 4783 1429 4930
rect 1475 4783 1504 4930
rect 1400 4760 1504 4783
rect 5320 4930 5432 4960
rect 5320 4783 5353 4930
rect 5399 4783 5432 4930
rect 5320 4760 5432 4783
rect 13272 4930 13384 4960
rect 13272 4783 13305 4930
rect 13351 4783 13384 4930
rect 13272 4760 13384 4783
rect 21224 4930 21336 4960
rect 21224 4783 21257 4930
rect 21303 4783 21336 4930
rect 21224 4760 21336 4783
rect 22464 4930 22568 4960
rect 22464 4783 22493 4930
rect 22539 4783 22568 4930
rect 22464 4760 22568 4783
rect 1400 4625 1504 4648
rect 1400 4478 1429 4625
rect 1475 4478 1504 4625
rect 1400 4448 1504 4478
rect 9352 4625 9464 4648
rect 9352 4478 9385 4625
rect 9431 4478 9464 4625
rect 9352 4448 9464 4478
rect 17304 4625 17416 4648
rect 17304 4478 17337 4625
rect 17383 4478 17416 4625
rect 17304 4448 17416 4478
rect 22464 4625 22568 4648
rect 22464 4478 22493 4625
rect 22539 4478 22568 4625
rect 22464 4448 22568 4478
rect 1400 3362 1504 3392
rect 1400 3215 1429 3362
rect 1475 3215 1504 3362
rect 1400 3192 1504 3215
rect 5320 3362 5432 3392
rect 5320 3215 5353 3362
rect 5399 3215 5432 3362
rect 5320 3192 5432 3215
rect 9240 3362 9352 3392
rect 9240 3215 9273 3362
rect 9319 3215 9352 3362
rect 9240 3192 9352 3215
rect 13160 3362 13272 3392
rect 13160 3215 13193 3362
rect 13239 3215 13272 3362
rect 13160 3192 13272 3215
rect 17080 3362 17192 3392
rect 17080 3215 17113 3362
rect 17159 3215 17192 3362
rect 17080 3192 17192 3215
rect 21000 3362 21112 3392
rect 21000 3215 21033 3362
rect 21079 3215 21112 3362
rect 21000 3192 21112 3215
rect 22464 3362 22568 3392
rect 22464 3215 22493 3362
rect 22539 3215 22568 3362
rect 22464 3192 22568 3215
<< mvnsubdiff >>
rect 1416 16379 1488 16392
rect 1416 16333 1429 16379
rect 1475 16333 1488 16379
rect 1416 16251 1488 16333
rect 1416 16205 1429 16251
rect 1475 16205 1488 16251
rect 1416 16123 1488 16205
rect 5336 16379 5416 16392
rect 5336 16333 5353 16379
rect 5399 16333 5416 16379
rect 5336 16251 5416 16333
rect 5336 16205 5353 16251
rect 5399 16205 5416 16251
rect 1416 16077 1429 16123
rect 1475 16077 1488 16123
rect 1416 16064 1488 16077
rect 5336 16123 5416 16205
rect 9256 16379 9336 16392
rect 9256 16333 9273 16379
rect 9319 16333 9336 16379
rect 9256 16251 9336 16333
rect 9256 16205 9273 16251
rect 9319 16205 9336 16251
rect 5336 16077 5353 16123
rect 5399 16077 5416 16123
rect 5336 16064 5416 16077
rect 9256 16123 9336 16205
rect 13176 16379 13256 16392
rect 13176 16333 13193 16379
rect 13239 16333 13256 16379
rect 13176 16251 13256 16333
rect 13176 16205 13193 16251
rect 13239 16205 13256 16251
rect 9256 16077 9273 16123
rect 9319 16077 9336 16123
rect 9256 16064 9336 16077
rect 13176 16123 13256 16205
rect 17096 16379 17176 16392
rect 17096 16333 17113 16379
rect 17159 16333 17176 16379
rect 17096 16251 17176 16333
rect 17096 16205 17113 16251
rect 17159 16205 17176 16251
rect 13176 16077 13193 16123
rect 13239 16077 13256 16123
rect 13176 16064 13256 16077
rect 17096 16123 17176 16205
rect 21016 16379 21096 16392
rect 21016 16333 21033 16379
rect 21079 16333 21096 16379
rect 21016 16251 21096 16333
rect 21016 16205 21033 16251
rect 21079 16205 21096 16251
rect 17096 16077 17113 16123
rect 17159 16077 17176 16123
rect 17096 16064 17176 16077
rect 21016 16123 21096 16205
rect 22480 16379 22552 16392
rect 22480 16333 22493 16379
rect 22539 16333 22552 16379
rect 22480 16251 22552 16333
rect 22480 16205 22493 16251
rect 22539 16205 22552 16251
rect 21016 16077 21033 16123
rect 21079 16077 21096 16123
rect 21016 16064 21096 16077
rect 22480 16123 22552 16205
rect 22480 16077 22493 16123
rect 22539 16077 22552 16123
rect 22480 16064 22552 16077
rect 1416 15283 1488 15296
rect 1416 15237 1429 15283
rect 1475 15237 1488 15283
rect 1416 15155 1488 15237
rect 9368 15283 9448 15296
rect 9368 15237 9385 15283
rect 9431 15237 9448 15283
rect 1416 15109 1429 15155
rect 1475 15109 1488 15155
rect 1416 15027 1488 15109
rect 1416 14981 1429 15027
rect 1475 14981 1488 15027
rect 1416 14968 1488 14981
rect 9368 15155 9448 15237
rect 17320 15283 17400 15296
rect 17320 15237 17337 15283
rect 17383 15237 17400 15283
rect 9368 15109 9385 15155
rect 9431 15109 9448 15155
rect 9368 15027 9448 15109
rect 9368 14981 9385 15027
rect 9431 14981 9448 15027
rect 9368 14968 9448 14981
rect 17320 15155 17400 15237
rect 22480 15283 22552 15296
rect 22480 15237 22493 15283
rect 22539 15237 22552 15283
rect 17320 15109 17337 15155
rect 17383 15109 17400 15155
rect 17320 15027 17400 15109
rect 17320 14981 17337 15027
rect 17383 14981 17400 15027
rect 17320 14968 17400 14981
rect 22480 15155 22552 15237
rect 22480 15109 22493 15155
rect 22539 15109 22552 15155
rect 22480 15027 22552 15109
rect 22480 14981 22493 15027
rect 22539 14981 22552 15027
rect 22480 14968 22552 14981
rect 1416 14811 1488 14824
rect 1416 14765 1429 14811
rect 1475 14765 1488 14811
rect 1416 14683 1488 14765
rect 1416 14637 1429 14683
rect 1475 14637 1488 14683
rect 1416 14555 1488 14637
rect 5336 14811 5416 14824
rect 5336 14765 5353 14811
rect 5399 14765 5416 14811
rect 5336 14683 5416 14765
rect 5336 14637 5353 14683
rect 5399 14637 5416 14683
rect 1416 14509 1429 14555
rect 1475 14509 1488 14555
rect 1416 14496 1488 14509
rect 5336 14555 5416 14637
rect 13288 14811 13368 14824
rect 13288 14765 13305 14811
rect 13351 14765 13368 14811
rect 13288 14683 13368 14765
rect 13288 14637 13305 14683
rect 13351 14637 13368 14683
rect 5336 14509 5353 14555
rect 5399 14509 5416 14555
rect 5336 14496 5416 14509
rect 13288 14555 13368 14637
rect 21240 14811 21320 14824
rect 21240 14765 21257 14811
rect 21303 14765 21320 14811
rect 21240 14683 21320 14765
rect 21240 14637 21257 14683
rect 21303 14637 21320 14683
rect 13288 14509 13305 14555
rect 13351 14509 13368 14555
rect 13288 14496 13368 14509
rect 21240 14555 21320 14637
rect 22480 14811 22552 14824
rect 22480 14765 22493 14811
rect 22539 14765 22552 14811
rect 22480 14683 22552 14765
rect 22480 14637 22493 14683
rect 22539 14637 22552 14683
rect 21240 14509 21257 14555
rect 21303 14509 21320 14555
rect 21240 14496 21320 14509
rect 22480 14555 22552 14637
rect 22480 14509 22493 14555
rect 22539 14509 22552 14555
rect 22480 14496 22552 14509
rect 1416 13715 1488 13728
rect 1416 13669 1429 13715
rect 1475 13669 1488 13715
rect 1416 13587 1488 13669
rect 9368 13715 9448 13728
rect 9368 13669 9385 13715
rect 9431 13669 9448 13715
rect 1416 13541 1429 13587
rect 1475 13541 1488 13587
rect 1416 13459 1488 13541
rect 1416 13413 1429 13459
rect 1475 13413 1488 13459
rect 1416 13400 1488 13413
rect 9368 13587 9448 13669
rect 17320 13715 17400 13728
rect 17320 13669 17337 13715
rect 17383 13669 17400 13715
rect 9368 13541 9385 13587
rect 9431 13541 9448 13587
rect 9368 13459 9448 13541
rect 9368 13413 9385 13459
rect 9431 13413 9448 13459
rect 9368 13400 9448 13413
rect 17320 13587 17400 13669
rect 22480 13715 22552 13728
rect 22480 13669 22493 13715
rect 22539 13669 22552 13715
rect 17320 13541 17337 13587
rect 17383 13541 17400 13587
rect 17320 13459 17400 13541
rect 17320 13413 17337 13459
rect 17383 13413 17400 13459
rect 17320 13400 17400 13413
rect 22480 13587 22552 13669
rect 22480 13541 22493 13587
rect 22539 13541 22552 13587
rect 22480 13459 22552 13541
rect 22480 13413 22493 13459
rect 22539 13413 22552 13459
rect 22480 13400 22552 13413
rect 1416 13243 1488 13256
rect 1416 13197 1429 13243
rect 1475 13197 1488 13243
rect 1416 13115 1488 13197
rect 1416 13069 1429 13115
rect 1475 13069 1488 13115
rect 1416 12987 1488 13069
rect 5336 13243 5416 13256
rect 5336 13197 5353 13243
rect 5399 13197 5416 13243
rect 5336 13115 5416 13197
rect 5336 13069 5353 13115
rect 5399 13069 5416 13115
rect 1416 12941 1429 12987
rect 1475 12941 1488 12987
rect 1416 12928 1488 12941
rect 5336 12987 5416 13069
rect 13288 13243 13368 13256
rect 13288 13197 13305 13243
rect 13351 13197 13368 13243
rect 13288 13115 13368 13197
rect 13288 13069 13305 13115
rect 13351 13069 13368 13115
rect 5336 12941 5353 12987
rect 5399 12941 5416 12987
rect 5336 12928 5416 12941
rect 13288 12987 13368 13069
rect 21240 13243 21320 13256
rect 21240 13197 21257 13243
rect 21303 13197 21320 13243
rect 21240 13115 21320 13197
rect 21240 13069 21257 13115
rect 21303 13069 21320 13115
rect 13288 12941 13305 12987
rect 13351 12941 13368 12987
rect 13288 12928 13368 12941
rect 21240 12987 21320 13069
rect 22480 13243 22552 13256
rect 22480 13197 22493 13243
rect 22539 13197 22552 13243
rect 22480 13115 22552 13197
rect 22480 13069 22493 13115
rect 22539 13069 22552 13115
rect 21240 12941 21257 12987
rect 21303 12941 21320 12987
rect 21240 12928 21320 12941
rect 22480 12987 22552 13069
rect 22480 12941 22493 12987
rect 22539 12941 22552 12987
rect 22480 12928 22552 12941
rect 1416 12147 1488 12160
rect 1416 12101 1429 12147
rect 1475 12101 1488 12147
rect 1416 12019 1488 12101
rect 9368 12147 9448 12160
rect 9368 12101 9385 12147
rect 9431 12101 9448 12147
rect 1416 11973 1429 12019
rect 1475 11973 1488 12019
rect 1416 11891 1488 11973
rect 1416 11845 1429 11891
rect 1475 11845 1488 11891
rect 1416 11832 1488 11845
rect 9368 12019 9448 12101
rect 17320 12147 17400 12160
rect 17320 12101 17337 12147
rect 17383 12101 17400 12147
rect 9368 11973 9385 12019
rect 9431 11973 9448 12019
rect 9368 11891 9448 11973
rect 9368 11845 9385 11891
rect 9431 11845 9448 11891
rect 9368 11832 9448 11845
rect 17320 12019 17400 12101
rect 22480 12147 22552 12160
rect 22480 12101 22493 12147
rect 22539 12101 22552 12147
rect 17320 11973 17337 12019
rect 17383 11973 17400 12019
rect 17320 11891 17400 11973
rect 17320 11845 17337 11891
rect 17383 11845 17400 11891
rect 17320 11832 17400 11845
rect 22480 12019 22552 12101
rect 22480 11973 22493 12019
rect 22539 11973 22552 12019
rect 22480 11891 22552 11973
rect 22480 11845 22493 11891
rect 22539 11845 22552 11891
rect 22480 11832 22552 11845
rect 1416 11675 1488 11688
rect 1416 11629 1429 11675
rect 1475 11629 1488 11675
rect 1416 11547 1488 11629
rect 1416 11501 1429 11547
rect 1475 11501 1488 11547
rect 1416 11419 1488 11501
rect 5336 11675 5416 11688
rect 5336 11629 5353 11675
rect 5399 11629 5416 11675
rect 5336 11547 5416 11629
rect 5336 11501 5353 11547
rect 5399 11501 5416 11547
rect 1416 11373 1429 11419
rect 1475 11373 1488 11419
rect 1416 11360 1488 11373
rect 5336 11419 5416 11501
rect 13288 11675 13368 11688
rect 13288 11629 13305 11675
rect 13351 11629 13368 11675
rect 13288 11547 13368 11629
rect 13288 11501 13305 11547
rect 13351 11501 13368 11547
rect 5336 11373 5353 11419
rect 5399 11373 5416 11419
rect 5336 11360 5416 11373
rect 13288 11419 13368 11501
rect 21240 11675 21320 11688
rect 21240 11629 21257 11675
rect 21303 11629 21320 11675
rect 21240 11547 21320 11629
rect 21240 11501 21257 11547
rect 21303 11501 21320 11547
rect 13288 11373 13305 11419
rect 13351 11373 13368 11419
rect 13288 11360 13368 11373
rect 21240 11419 21320 11501
rect 22480 11675 22552 11688
rect 22480 11629 22493 11675
rect 22539 11629 22552 11675
rect 22480 11547 22552 11629
rect 22480 11501 22493 11547
rect 22539 11501 22552 11547
rect 21240 11373 21257 11419
rect 21303 11373 21320 11419
rect 21240 11360 21320 11373
rect 22480 11419 22552 11501
rect 22480 11373 22493 11419
rect 22539 11373 22552 11419
rect 22480 11360 22552 11373
rect 1416 10579 1488 10592
rect 1416 10533 1429 10579
rect 1475 10533 1488 10579
rect 1416 10451 1488 10533
rect 9368 10579 9448 10592
rect 9368 10533 9385 10579
rect 9431 10533 9448 10579
rect 1416 10405 1429 10451
rect 1475 10405 1488 10451
rect 1416 10323 1488 10405
rect 1416 10277 1429 10323
rect 1475 10277 1488 10323
rect 1416 10264 1488 10277
rect 9368 10451 9448 10533
rect 17320 10579 17400 10592
rect 17320 10533 17337 10579
rect 17383 10533 17400 10579
rect 9368 10405 9385 10451
rect 9431 10405 9448 10451
rect 9368 10323 9448 10405
rect 9368 10277 9385 10323
rect 9431 10277 9448 10323
rect 9368 10264 9448 10277
rect 17320 10451 17400 10533
rect 22480 10579 22552 10592
rect 22480 10533 22493 10579
rect 22539 10533 22552 10579
rect 17320 10405 17337 10451
rect 17383 10405 17400 10451
rect 17320 10323 17400 10405
rect 17320 10277 17337 10323
rect 17383 10277 17400 10323
rect 17320 10264 17400 10277
rect 22480 10451 22552 10533
rect 22480 10405 22493 10451
rect 22539 10405 22552 10451
rect 22480 10323 22552 10405
rect 22480 10277 22493 10323
rect 22539 10277 22552 10323
rect 22480 10264 22552 10277
rect 1416 10107 1488 10120
rect 1416 10061 1429 10107
rect 1475 10061 1488 10107
rect 1416 9979 1488 10061
rect 1416 9933 1429 9979
rect 1475 9933 1488 9979
rect 1416 9851 1488 9933
rect 5336 10107 5416 10120
rect 5336 10061 5353 10107
rect 5399 10061 5416 10107
rect 5336 9979 5416 10061
rect 5336 9933 5353 9979
rect 5399 9933 5416 9979
rect 1416 9805 1429 9851
rect 1475 9805 1488 9851
rect 1416 9792 1488 9805
rect 5336 9851 5416 9933
rect 13288 10107 13368 10120
rect 13288 10061 13305 10107
rect 13351 10061 13368 10107
rect 13288 9979 13368 10061
rect 13288 9933 13305 9979
rect 13351 9933 13368 9979
rect 5336 9805 5353 9851
rect 5399 9805 5416 9851
rect 5336 9792 5416 9805
rect 13288 9851 13368 9933
rect 21240 10107 21320 10120
rect 21240 10061 21257 10107
rect 21303 10061 21320 10107
rect 21240 9979 21320 10061
rect 21240 9933 21257 9979
rect 21303 9933 21320 9979
rect 13288 9805 13305 9851
rect 13351 9805 13368 9851
rect 13288 9792 13368 9805
rect 21240 9851 21320 9933
rect 22480 10107 22552 10120
rect 22480 10061 22493 10107
rect 22539 10061 22552 10107
rect 22480 9979 22552 10061
rect 22480 9933 22493 9979
rect 22539 9933 22552 9979
rect 21240 9805 21257 9851
rect 21303 9805 21320 9851
rect 21240 9792 21320 9805
rect 22480 9851 22552 9933
rect 22480 9805 22493 9851
rect 22539 9805 22552 9851
rect 22480 9792 22552 9805
rect 1416 9011 1488 9024
rect 1416 8965 1429 9011
rect 1475 8965 1488 9011
rect 1416 8883 1488 8965
rect 9368 9011 9448 9024
rect 9368 8965 9385 9011
rect 9431 8965 9448 9011
rect 1416 8837 1429 8883
rect 1475 8837 1488 8883
rect 1416 8755 1488 8837
rect 1416 8709 1429 8755
rect 1475 8709 1488 8755
rect 1416 8696 1488 8709
rect 9368 8883 9448 8965
rect 17320 9011 17400 9024
rect 17320 8965 17337 9011
rect 17383 8965 17400 9011
rect 9368 8837 9385 8883
rect 9431 8837 9448 8883
rect 9368 8755 9448 8837
rect 9368 8709 9385 8755
rect 9431 8709 9448 8755
rect 9368 8696 9448 8709
rect 17320 8883 17400 8965
rect 22480 9011 22552 9024
rect 22480 8965 22493 9011
rect 22539 8965 22552 9011
rect 17320 8837 17337 8883
rect 17383 8837 17400 8883
rect 17320 8755 17400 8837
rect 17320 8709 17337 8755
rect 17383 8709 17400 8755
rect 17320 8696 17400 8709
rect 22480 8883 22552 8965
rect 22480 8837 22493 8883
rect 22539 8837 22552 8883
rect 22480 8755 22552 8837
rect 22480 8709 22493 8755
rect 22539 8709 22552 8755
rect 22480 8696 22552 8709
rect 1416 8539 1488 8552
rect 1416 8493 1429 8539
rect 1475 8493 1488 8539
rect 1416 8411 1488 8493
rect 1416 8365 1429 8411
rect 1475 8365 1488 8411
rect 1416 8283 1488 8365
rect 5336 8539 5416 8552
rect 5336 8493 5353 8539
rect 5399 8493 5416 8539
rect 5336 8411 5416 8493
rect 5336 8365 5353 8411
rect 5399 8365 5416 8411
rect 1416 8237 1429 8283
rect 1475 8237 1488 8283
rect 1416 8224 1488 8237
rect 5336 8283 5416 8365
rect 13288 8539 13368 8552
rect 13288 8493 13305 8539
rect 13351 8493 13368 8539
rect 13288 8411 13368 8493
rect 13288 8365 13305 8411
rect 13351 8365 13368 8411
rect 5336 8237 5353 8283
rect 5399 8237 5416 8283
rect 5336 8224 5416 8237
rect 13288 8283 13368 8365
rect 21240 8539 21320 8552
rect 21240 8493 21257 8539
rect 21303 8493 21320 8539
rect 21240 8411 21320 8493
rect 21240 8365 21257 8411
rect 21303 8365 21320 8411
rect 13288 8237 13305 8283
rect 13351 8237 13368 8283
rect 13288 8224 13368 8237
rect 21240 8283 21320 8365
rect 22480 8539 22552 8552
rect 22480 8493 22493 8539
rect 22539 8493 22552 8539
rect 22480 8411 22552 8493
rect 22480 8365 22493 8411
rect 22539 8365 22552 8411
rect 21240 8237 21257 8283
rect 21303 8237 21320 8283
rect 21240 8224 21320 8237
rect 22480 8283 22552 8365
rect 22480 8237 22493 8283
rect 22539 8237 22552 8283
rect 22480 8224 22552 8237
rect 1416 7443 1488 7456
rect 1416 7397 1429 7443
rect 1475 7397 1488 7443
rect 1416 7315 1488 7397
rect 9368 7443 9448 7456
rect 9368 7397 9385 7443
rect 9431 7397 9448 7443
rect 1416 7269 1429 7315
rect 1475 7269 1488 7315
rect 1416 7187 1488 7269
rect 1416 7141 1429 7187
rect 1475 7141 1488 7187
rect 1416 7128 1488 7141
rect 9368 7315 9448 7397
rect 17320 7443 17400 7456
rect 17320 7397 17337 7443
rect 17383 7397 17400 7443
rect 9368 7269 9385 7315
rect 9431 7269 9448 7315
rect 9368 7187 9448 7269
rect 9368 7141 9385 7187
rect 9431 7141 9448 7187
rect 9368 7128 9448 7141
rect 17320 7315 17400 7397
rect 22480 7443 22552 7456
rect 22480 7397 22493 7443
rect 22539 7397 22552 7443
rect 17320 7269 17337 7315
rect 17383 7269 17400 7315
rect 17320 7187 17400 7269
rect 17320 7141 17337 7187
rect 17383 7141 17400 7187
rect 17320 7128 17400 7141
rect 22480 7315 22552 7397
rect 22480 7269 22493 7315
rect 22539 7269 22552 7315
rect 22480 7187 22552 7269
rect 22480 7141 22493 7187
rect 22539 7141 22552 7187
rect 22480 7128 22552 7141
rect 1416 6971 1488 6984
rect 1416 6925 1429 6971
rect 1475 6925 1488 6971
rect 1416 6843 1488 6925
rect 1416 6797 1429 6843
rect 1475 6797 1488 6843
rect 1416 6715 1488 6797
rect 5336 6971 5416 6984
rect 5336 6925 5353 6971
rect 5399 6925 5416 6971
rect 5336 6843 5416 6925
rect 5336 6797 5353 6843
rect 5399 6797 5416 6843
rect 1416 6669 1429 6715
rect 1475 6669 1488 6715
rect 1416 6656 1488 6669
rect 5336 6715 5416 6797
rect 13288 6971 13368 6984
rect 13288 6925 13305 6971
rect 13351 6925 13368 6971
rect 13288 6843 13368 6925
rect 13288 6797 13305 6843
rect 13351 6797 13368 6843
rect 5336 6669 5353 6715
rect 5399 6669 5416 6715
rect 5336 6656 5416 6669
rect 13288 6715 13368 6797
rect 21240 6971 21320 6984
rect 21240 6925 21257 6971
rect 21303 6925 21320 6971
rect 21240 6843 21320 6925
rect 21240 6797 21257 6843
rect 21303 6797 21320 6843
rect 13288 6669 13305 6715
rect 13351 6669 13368 6715
rect 13288 6656 13368 6669
rect 21240 6715 21320 6797
rect 22480 6971 22552 6984
rect 22480 6925 22493 6971
rect 22539 6925 22552 6971
rect 22480 6843 22552 6925
rect 22480 6797 22493 6843
rect 22539 6797 22552 6843
rect 21240 6669 21257 6715
rect 21303 6669 21320 6715
rect 21240 6656 21320 6669
rect 22480 6715 22552 6797
rect 22480 6669 22493 6715
rect 22539 6669 22552 6715
rect 22480 6656 22552 6669
rect 1416 5875 1488 5888
rect 1416 5829 1429 5875
rect 1475 5829 1488 5875
rect 1416 5747 1488 5829
rect 9368 5875 9448 5888
rect 9368 5829 9385 5875
rect 9431 5829 9448 5875
rect 1416 5701 1429 5747
rect 1475 5701 1488 5747
rect 1416 5619 1488 5701
rect 1416 5573 1429 5619
rect 1475 5573 1488 5619
rect 1416 5560 1488 5573
rect 9368 5747 9448 5829
rect 17320 5875 17400 5888
rect 17320 5829 17337 5875
rect 17383 5829 17400 5875
rect 9368 5701 9385 5747
rect 9431 5701 9448 5747
rect 9368 5619 9448 5701
rect 9368 5573 9385 5619
rect 9431 5573 9448 5619
rect 9368 5560 9448 5573
rect 17320 5747 17400 5829
rect 22480 5875 22552 5888
rect 22480 5829 22493 5875
rect 22539 5829 22552 5875
rect 17320 5701 17337 5747
rect 17383 5701 17400 5747
rect 17320 5619 17400 5701
rect 17320 5573 17337 5619
rect 17383 5573 17400 5619
rect 17320 5560 17400 5573
rect 22480 5747 22552 5829
rect 22480 5701 22493 5747
rect 22539 5701 22552 5747
rect 22480 5619 22552 5701
rect 22480 5573 22493 5619
rect 22539 5573 22552 5619
rect 22480 5560 22552 5573
rect 1416 5403 1488 5416
rect 1416 5357 1429 5403
rect 1475 5357 1488 5403
rect 1416 5275 1488 5357
rect 1416 5229 1429 5275
rect 1475 5229 1488 5275
rect 1416 5147 1488 5229
rect 5336 5403 5416 5416
rect 5336 5357 5353 5403
rect 5399 5357 5416 5403
rect 5336 5275 5416 5357
rect 5336 5229 5353 5275
rect 5399 5229 5416 5275
rect 1416 5101 1429 5147
rect 1475 5101 1488 5147
rect 1416 5088 1488 5101
rect 5336 5147 5416 5229
rect 13288 5403 13368 5416
rect 13288 5357 13305 5403
rect 13351 5357 13368 5403
rect 13288 5275 13368 5357
rect 13288 5229 13305 5275
rect 13351 5229 13368 5275
rect 5336 5101 5353 5147
rect 5399 5101 5416 5147
rect 5336 5088 5416 5101
rect 13288 5147 13368 5229
rect 21240 5403 21320 5416
rect 21240 5357 21257 5403
rect 21303 5357 21320 5403
rect 21240 5275 21320 5357
rect 21240 5229 21257 5275
rect 21303 5229 21320 5275
rect 13288 5101 13305 5147
rect 13351 5101 13368 5147
rect 13288 5088 13368 5101
rect 21240 5147 21320 5229
rect 22480 5403 22552 5416
rect 22480 5357 22493 5403
rect 22539 5357 22552 5403
rect 22480 5275 22552 5357
rect 22480 5229 22493 5275
rect 22539 5229 22552 5275
rect 21240 5101 21257 5147
rect 21303 5101 21320 5147
rect 21240 5088 21320 5101
rect 22480 5147 22552 5229
rect 22480 5101 22493 5147
rect 22539 5101 22552 5147
rect 22480 5088 22552 5101
rect 1416 4307 1488 4320
rect 1416 4261 1429 4307
rect 1475 4261 1488 4307
rect 1416 4179 1488 4261
rect 9368 4307 9448 4320
rect 9368 4261 9385 4307
rect 9431 4261 9448 4307
rect 1416 4133 1429 4179
rect 1475 4133 1488 4179
rect 1416 4051 1488 4133
rect 1416 4005 1429 4051
rect 1475 4005 1488 4051
rect 1416 3992 1488 4005
rect 9368 4179 9448 4261
rect 17320 4307 17400 4320
rect 17320 4261 17337 4307
rect 17383 4261 17400 4307
rect 9368 4133 9385 4179
rect 9431 4133 9448 4179
rect 9368 4051 9448 4133
rect 9368 4005 9385 4051
rect 9431 4005 9448 4051
rect 9368 3992 9448 4005
rect 17320 4179 17400 4261
rect 22480 4307 22552 4320
rect 22480 4261 22493 4307
rect 22539 4261 22552 4307
rect 17320 4133 17337 4179
rect 17383 4133 17400 4179
rect 17320 4051 17400 4133
rect 17320 4005 17337 4051
rect 17383 4005 17400 4051
rect 17320 3992 17400 4005
rect 22480 4179 22552 4261
rect 22480 4133 22493 4179
rect 22539 4133 22552 4179
rect 22480 4051 22552 4133
rect 22480 4005 22493 4051
rect 22539 4005 22552 4051
rect 22480 3992 22552 4005
rect 1416 3835 1488 3848
rect 1416 3789 1429 3835
rect 1475 3789 1488 3835
rect 1416 3707 1488 3789
rect 1416 3661 1429 3707
rect 1475 3661 1488 3707
rect 1416 3579 1488 3661
rect 5336 3835 5416 3848
rect 5336 3789 5353 3835
rect 5399 3789 5416 3835
rect 5336 3707 5416 3789
rect 5336 3661 5353 3707
rect 5399 3661 5416 3707
rect 1416 3533 1429 3579
rect 1475 3533 1488 3579
rect 1416 3520 1488 3533
rect 5336 3579 5416 3661
rect 9256 3835 9336 3848
rect 9256 3789 9273 3835
rect 9319 3789 9336 3835
rect 9256 3707 9336 3789
rect 9256 3661 9273 3707
rect 9319 3661 9336 3707
rect 5336 3533 5353 3579
rect 5399 3533 5416 3579
rect 5336 3520 5416 3533
rect 9256 3579 9336 3661
rect 13176 3835 13256 3848
rect 13176 3789 13193 3835
rect 13239 3789 13256 3835
rect 13176 3707 13256 3789
rect 13176 3661 13193 3707
rect 13239 3661 13256 3707
rect 9256 3533 9273 3579
rect 9319 3533 9336 3579
rect 9256 3520 9336 3533
rect 13176 3579 13256 3661
rect 17096 3835 17176 3848
rect 17096 3789 17113 3835
rect 17159 3789 17176 3835
rect 17096 3707 17176 3789
rect 17096 3661 17113 3707
rect 17159 3661 17176 3707
rect 13176 3533 13193 3579
rect 13239 3533 13256 3579
rect 13176 3520 13256 3533
rect 17096 3579 17176 3661
rect 21016 3835 21096 3848
rect 21016 3789 21033 3835
rect 21079 3789 21096 3835
rect 21016 3707 21096 3789
rect 21016 3661 21033 3707
rect 21079 3661 21096 3707
rect 17096 3533 17113 3579
rect 17159 3533 17176 3579
rect 17096 3520 17176 3533
rect 21016 3579 21096 3661
rect 22480 3835 22552 3848
rect 22480 3789 22493 3835
rect 22539 3789 22552 3835
rect 22480 3707 22552 3789
rect 22480 3661 22493 3707
rect 22539 3661 22552 3707
rect 21016 3533 21033 3579
rect 21079 3533 21096 3579
rect 21016 3520 21096 3533
rect 22480 3579 22552 3661
rect 22480 3533 22493 3579
rect 22539 3533 22552 3579
rect 22480 3520 22552 3533
<< mvpsubdiffcont >>
rect 1429 15759 1475 15906
rect 5353 15759 5399 15906
rect 9273 15759 9319 15906
rect 13193 15759 13239 15906
rect 17113 15759 17159 15906
rect 21033 15759 21079 15906
rect 22493 15759 22539 15906
rect 1429 15454 1475 15601
rect 9385 15454 9431 15601
rect 17337 15454 17383 15601
rect 22493 15454 22539 15601
rect 1429 14191 1475 14338
rect 5353 14191 5399 14338
rect 13305 14191 13351 14338
rect 21257 14191 21303 14338
rect 22493 14191 22539 14338
rect 1429 13886 1475 14033
rect 9385 13886 9431 14033
rect 17337 13886 17383 14033
rect 22493 13886 22539 14033
rect 1429 12623 1475 12770
rect 5353 12623 5399 12770
rect 13305 12623 13351 12770
rect 21257 12623 21303 12770
rect 22493 12623 22539 12770
rect 1429 12318 1475 12465
rect 9385 12318 9431 12465
rect 17337 12318 17383 12465
rect 22493 12318 22539 12465
rect 1429 11055 1475 11202
rect 5353 11055 5399 11202
rect 13305 11055 13351 11202
rect 21257 11055 21303 11202
rect 22493 11055 22539 11202
rect 1429 10750 1475 10897
rect 9385 10750 9431 10897
rect 17337 10750 17383 10897
rect 22493 10750 22539 10897
rect 1429 9487 1475 9634
rect 5353 9487 5399 9634
rect 13305 9487 13351 9634
rect 21257 9487 21303 9634
rect 22493 9487 22539 9634
rect 1429 9182 1475 9329
rect 9385 9182 9431 9329
rect 17337 9182 17383 9329
rect 22493 9182 22539 9329
rect 1429 7919 1475 8066
rect 5353 7919 5399 8066
rect 13305 7919 13351 8066
rect 21257 7919 21303 8066
rect 22493 7919 22539 8066
rect 1429 7614 1475 7761
rect 9385 7614 9431 7761
rect 17337 7614 17383 7761
rect 22493 7614 22539 7761
rect 1429 6351 1475 6498
rect 5353 6351 5399 6498
rect 13305 6351 13351 6498
rect 21257 6351 21303 6498
rect 22493 6351 22539 6498
rect 1429 6046 1475 6193
rect 9385 6046 9431 6193
rect 17337 6046 17383 6193
rect 22493 6046 22539 6193
rect 1429 4783 1475 4930
rect 5353 4783 5399 4930
rect 13305 4783 13351 4930
rect 21257 4783 21303 4930
rect 22493 4783 22539 4930
rect 1429 4478 1475 4625
rect 9385 4478 9431 4625
rect 17337 4478 17383 4625
rect 22493 4478 22539 4625
rect 1429 3215 1475 3362
rect 5353 3215 5399 3362
rect 9273 3215 9319 3362
rect 13193 3215 13239 3362
rect 17113 3215 17159 3362
rect 21033 3215 21079 3362
rect 22493 3215 22539 3362
<< mvnsubdiffcont >>
rect 1429 16333 1475 16379
rect 1429 16205 1475 16251
rect 5353 16333 5399 16379
rect 5353 16205 5399 16251
rect 1429 16077 1475 16123
rect 9273 16333 9319 16379
rect 9273 16205 9319 16251
rect 5353 16077 5399 16123
rect 13193 16333 13239 16379
rect 13193 16205 13239 16251
rect 9273 16077 9319 16123
rect 17113 16333 17159 16379
rect 17113 16205 17159 16251
rect 13193 16077 13239 16123
rect 21033 16333 21079 16379
rect 21033 16205 21079 16251
rect 17113 16077 17159 16123
rect 22493 16333 22539 16379
rect 22493 16205 22539 16251
rect 21033 16077 21079 16123
rect 22493 16077 22539 16123
rect 1429 15237 1475 15283
rect 9385 15237 9431 15283
rect 1429 15109 1475 15155
rect 1429 14981 1475 15027
rect 17337 15237 17383 15283
rect 9385 15109 9431 15155
rect 9385 14981 9431 15027
rect 22493 15237 22539 15283
rect 17337 15109 17383 15155
rect 17337 14981 17383 15027
rect 22493 15109 22539 15155
rect 22493 14981 22539 15027
rect 1429 14765 1475 14811
rect 1429 14637 1475 14683
rect 5353 14765 5399 14811
rect 5353 14637 5399 14683
rect 1429 14509 1475 14555
rect 13305 14765 13351 14811
rect 13305 14637 13351 14683
rect 5353 14509 5399 14555
rect 21257 14765 21303 14811
rect 21257 14637 21303 14683
rect 13305 14509 13351 14555
rect 22493 14765 22539 14811
rect 22493 14637 22539 14683
rect 21257 14509 21303 14555
rect 22493 14509 22539 14555
rect 1429 13669 1475 13715
rect 9385 13669 9431 13715
rect 1429 13541 1475 13587
rect 1429 13413 1475 13459
rect 17337 13669 17383 13715
rect 9385 13541 9431 13587
rect 9385 13413 9431 13459
rect 22493 13669 22539 13715
rect 17337 13541 17383 13587
rect 17337 13413 17383 13459
rect 22493 13541 22539 13587
rect 22493 13413 22539 13459
rect 1429 13197 1475 13243
rect 1429 13069 1475 13115
rect 5353 13197 5399 13243
rect 5353 13069 5399 13115
rect 1429 12941 1475 12987
rect 13305 13197 13351 13243
rect 13305 13069 13351 13115
rect 5353 12941 5399 12987
rect 21257 13197 21303 13243
rect 21257 13069 21303 13115
rect 13305 12941 13351 12987
rect 22493 13197 22539 13243
rect 22493 13069 22539 13115
rect 21257 12941 21303 12987
rect 22493 12941 22539 12987
rect 1429 12101 1475 12147
rect 9385 12101 9431 12147
rect 1429 11973 1475 12019
rect 1429 11845 1475 11891
rect 17337 12101 17383 12147
rect 9385 11973 9431 12019
rect 9385 11845 9431 11891
rect 22493 12101 22539 12147
rect 17337 11973 17383 12019
rect 17337 11845 17383 11891
rect 22493 11973 22539 12019
rect 22493 11845 22539 11891
rect 1429 11629 1475 11675
rect 1429 11501 1475 11547
rect 5353 11629 5399 11675
rect 5353 11501 5399 11547
rect 1429 11373 1475 11419
rect 13305 11629 13351 11675
rect 13305 11501 13351 11547
rect 5353 11373 5399 11419
rect 21257 11629 21303 11675
rect 21257 11501 21303 11547
rect 13305 11373 13351 11419
rect 22493 11629 22539 11675
rect 22493 11501 22539 11547
rect 21257 11373 21303 11419
rect 22493 11373 22539 11419
rect 1429 10533 1475 10579
rect 9385 10533 9431 10579
rect 1429 10405 1475 10451
rect 1429 10277 1475 10323
rect 17337 10533 17383 10579
rect 9385 10405 9431 10451
rect 9385 10277 9431 10323
rect 22493 10533 22539 10579
rect 17337 10405 17383 10451
rect 17337 10277 17383 10323
rect 22493 10405 22539 10451
rect 22493 10277 22539 10323
rect 1429 10061 1475 10107
rect 1429 9933 1475 9979
rect 5353 10061 5399 10107
rect 5353 9933 5399 9979
rect 1429 9805 1475 9851
rect 13305 10061 13351 10107
rect 13305 9933 13351 9979
rect 5353 9805 5399 9851
rect 21257 10061 21303 10107
rect 21257 9933 21303 9979
rect 13305 9805 13351 9851
rect 22493 10061 22539 10107
rect 22493 9933 22539 9979
rect 21257 9805 21303 9851
rect 22493 9805 22539 9851
rect 1429 8965 1475 9011
rect 9385 8965 9431 9011
rect 1429 8837 1475 8883
rect 1429 8709 1475 8755
rect 17337 8965 17383 9011
rect 9385 8837 9431 8883
rect 9385 8709 9431 8755
rect 22493 8965 22539 9011
rect 17337 8837 17383 8883
rect 17337 8709 17383 8755
rect 22493 8837 22539 8883
rect 22493 8709 22539 8755
rect 1429 8493 1475 8539
rect 1429 8365 1475 8411
rect 5353 8493 5399 8539
rect 5353 8365 5399 8411
rect 1429 8237 1475 8283
rect 13305 8493 13351 8539
rect 13305 8365 13351 8411
rect 5353 8237 5399 8283
rect 21257 8493 21303 8539
rect 21257 8365 21303 8411
rect 13305 8237 13351 8283
rect 22493 8493 22539 8539
rect 22493 8365 22539 8411
rect 21257 8237 21303 8283
rect 22493 8237 22539 8283
rect 1429 7397 1475 7443
rect 9385 7397 9431 7443
rect 1429 7269 1475 7315
rect 1429 7141 1475 7187
rect 17337 7397 17383 7443
rect 9385 7269 9431 7315
rect 9385 7141 9431 7187
rect 22493 7397 22539 7443
rect 17337 7269 17383 7315
rect 17337 7141 17383 7187
rect 22493 7269 22539 7315
rect 22493 7141 22539 7187
rect 1429 6925 1475 6971
rect 1429 6797 1475 6843
rect 5353 6925 5399 6971
rect 5353 6797 5399 6843
rect 1429 6669 1475 6715
rect 13305 6925 13351 6971
rect 13305 6797 13351 6843
rect 5353 6669 5399 6715
rect 21257 6925 21303 6971
rect 21257 6797 21303 6843
rect 13305 6669 13351 6715
rect 22493 6925 22539 6971
rect 22493 6797 22539 6843
rect 21257 6669 21303 6715
rect 22493 6669 22539 6715
rect 1429 5829 1475 5875
rect 9385 5829 9431 5875
rect 1429 5701 1475 5747
rect 1429 5573 1475 5619
rect 17337 5829 17383 5875
rect 9385 5701 9431 5747
rect 9385 5573 9431 5619
rect 22493 5829 22539 5875
rect 17337 5701 17383 5747
rect 17337 5573 17383 5619
rect 22493 5701 22539 5747
rect 22493 5573 22539 5619
rect 1429 5357 1475 5403
rect 1429 5229 1475 5275
rect 5353 5357 5399 5403
rect 5353 5229 5399 5275
rect 1429 5101 1475 5147
rect 13305 5357 13351 5403
rect 13305 5229 13351 5275
rect 5353 5101 5399 5147
rect 21257 5357 21303 5403
rect 21257 5229 21303 5275
rect 13305 5101 13351 5147
rect 22493 5357 22539 5403
rect 22493 5229 22539 5275
rect 21257 5101 21303 5147
rect 22493 5101 22539 5147
rect 1429 4261 1475 4307
rect 9385 4261 9431 4307
rect 1429 4133 1475 4179
rect 1429 4005 1475 4051
rect 17337 4261 17383 4307
rect 9385 4133 9431 4179
rect 9385 4005 9431 4051
rect 22493 4261 22539 4307
rect 17337 4133 17383 4179
rect 17337 4005 17383 4051
rect 22493 4133 22539 4179
rect 22493 4005 22539 4051
rect 1429 3789 1475 3835
rect 1429 3661 1475 3707
rect 5353 3789 5399 3835
rect 5353 3661 5399 3707
rect 1429 3533 1475 3579
rect 9273 3789 9319 3835
rect 9273 3661 9319 3707
rect 5353 3533 5399 3579
rect 13193 3789 13239 3835
rect 13193 3661 13239 3707
rect 9273 3533 9319 3579
rect 17113 3789 17159 3835
rect 17113 3661 17159 3707
rect 13193 3533 13239 3579
rect 21033 3789 21079 3835
rect 21033 3661 21079 3707
rect 17113 3533 17159 3579
rect 22493 3789 22539 3835
rect 22493 3661 22539 3707
rect 21033 3533 21079 3579
rect 22493 3533 22539 3579
<< polysilicon >>
rect 1692 16396 1892 16440
rect 2140 16396 2340 16440
rect 2588 16396 2788 16440
rect 3036 16396 3236 16440
rect 3484 16396 3684 16440
rect 3932 16396 4132 16440
rect 4380 16396 4580 16440
rect 4828 16396 5028 16440
rect 5612 16396 5812 16440
rect 6060 16396 6260 16440
rect 6508 16396 6708 16440
rect 6956 16396 7156 16440
rect 7404 16396 7604 16440
rect 7852 16396 8052 16440
rect 8300 16396 8500 16440
rect 8748 16396 8948 16440
rect 9532 16396 9732 16440
rect 9980 16396 10180 16440
rect 10428 16396 10628 16440
rect 10876 16396 11076 16440
rect 11324 16396 11524 16440
rect 11772 16396 11972 16440
rect 12220 16396 12420 16440
rect 12668 16396 12868 16440
rect 13452 16396 13652 16440
rect 13900 16396 14100 16440
rect 14348 16396 14548 16440
rect 14796 16396 14996 16440
rect 15244 16396 15444 16440
rect 15692 16396 15892 16440
rect 16140 16396 16340 16440
rect 16588 16396 16788 16440
rect 17372 16396 17572 16440
rect 17820 16396 18020 16440
rect 18268 16396 18468 16440
rect 18716 16396 18916 16440
rect 19164 16396 19364 16440
rect 19612 16396 19812 16440
rect 20060 16396 20260 16440
rect 20508 16396 20708 16440
rect 21292 16396 21492 16440
rect 21740 16396 21940 16440
rect 1692 16118 1892 16152
rect 1692 16072 1728 16118
rect 1868 16072 1892 16118
rect 1692 16055 1892 16072
rect 2140 16118 2340 16152
rect 2140 16072 2176 16118
rect 2316 16072 2340 16118
rect 2140 16055 2340 16072
rect 2588 16118 2788 16152
rect 2588 16072 2624 16118
rect 2764 16072 2788 16118
rect 2588 16055 2788 16072
rect 3036 16118 3236 16152
rect 3036 16072 3072 16118
rect 3212 16072 3236 16118
rect 3036 16055 3236 16072
rect 3484 16118 3684 16152
rect 3484 16072 3520 16118
rect 3660 16072 3684 16118
rect 3484 16055 3684 16072
rect 3932 16118 4132 16152
rect 3932 16072 3968 16118
rect 4108 16072 4132 16118
rect 3932 16055 4132 16072
rect 4380 16118 4580 16152
rect 4380 16072 4416 16118
rect 4556 16072 4580 16118
rect 4380 16055 4580 16072
rect 4828 16118 5028 16152
rect 4828 16072 4864 16118
rect 5004 16072 5028 16118
rect 4828 16055 5028 16072
rect 5612 16118 5812 16152
rect 5612 16072 5648 16118
rect 5788 16072 5812 16118
rect 5612 16055 5812 16072
rect 6060 16118 6260 16152
rect 6060 16072 6096 16118
rect 6236 16072 6260 16118
rect 6060 16055 6260 16072
rect 6508 16118 6708 16152
rect 6508 16072 6544 16118
rect 6684 16072 6708 16118
rect 6508 16055 6708 16072
rect 6956 16118 7156 16152
rect 6956 16072 6992 16118
rect 7132 16072 7156 16118
rect 6956 16055 7156 16072
rect 7404 16118 7604 16152
rect 7404 16072 7440 16118
rect 7580 16072 7604 16118
rect 7404 16055 7604 16072
rect 7852 16118 8052 16152
rect 7852 16072 7888 16118
rect 8028 16072 8052 16118
rect 7852 16055 8052 16072
rect 8300 16118 8500 16152
rect 8300 16072 8336 16118
rect 8476 16072 8500 16118
rect 8300 16055 8500 16072
rect 8748 16118 8948 16152
rect 8748 16072 8784 16118
rect 8924 16072 8948 16118
rect 8748 16055 8948 16072
rect 9532 16118 9732 16152
rect 9532 16072 9568 16118
rect 9708 16072 9732 16118
rect 9532 16055 9732 16072
rect 9980 16118 10180 16152
rect 9980 16072 10016 16118
rect 10156 16072 10180 16118
rect 9980 16055 10180 16072
rect 10428 16118 10628 16152
rect 10428 16072 10464 16118
rect 10604 16072 10628 16118
rect 10428 16055 10628 16072
rect 10876 16118 11076 16152
rect 10876 16072 10912 16118
rect 11052 16072 11076 16118
rect 10876 16055 11076 16072
rect 11324 16118 11524 16152
rect 11324 16072 11360 16118
rect 11500 16072 11524 16118
rect 11324 16055 11524 16072
rect 11772 16118 11972 16152
rect 11772 16072 11808 16118
rect 11948 16072 11972 16118
rect 11772 16055 11972 16072
rect 12220 16118 12420 16152
rect 12220 16072 12256 16118
rect 12396 16072 12420 16118
rect 12220 16055 12420 16072
rect 12668 16118 12868 16152
rect 12668 16072 12704 16118
rect 12844 16072 12868 16118
rect 12668 16055 12868 16072
rect 13452 16118 13652 16152
rect 13452 16072 13488 16118
rect 13628 16072 13652 16118
rect 13452 16055 13652 16072
rect 13900 16118 14100 16152
rect 13900 16072 13936 16118
rect 14076 16072 14100 16118
rect 13900 16055 14100 16072
rect 14348 16118 14548 16152
rect 14348 16072 14384 16118
rect 14524 16072 14548 16118
rect 14348 16055 14548 16072
rect 14796 16118 14996 16152
rect 14796 16072 14832 16118
rect 14972 16072 14996 16118
rect 14796 16055 14996 16072
rect 15244 16118 15444 16152
rect 15244 16072 15280 16118
rect 15420 16072 15444 16118
rect 15244 16055 15444 16072
rect 15692 16118 15892 16152
rect 15692 16072 15728 16118
rect 15868 16072 15892 16118
rect 15692 16055 15892 16072
rect 16140 16118 16340 16152
rect 16140 16072 16176 16118
rect 16316 16072 16340 16118
rect 16140 16055 16340 16072
rect 16588 16118 16788 16152
rect 16588 16072 16624 16118
rect 16764 16072 16788 16118
rect 16588 16055 16788 16072
rect 17372 16118 17572 16152
rect 17372 16072 17408 16118
rect 17548 16072 17572 16118
rect 17372 16055 17572 16072
rect 17820 16118 18020 16152
rect 17820 16072 17856 16118
rect 17996 16072 18020 16118
rect 17820 16055 18020 16072
rect 18268 16118 18468 16152
rect 18268 16072 18304 16118
rect 18444 16072 18468 16118
rect 18268 16055 18468 16072
rect 18716 16118 18916 16152
rect 18716 16072 18752 16118
rect 18892 16072 18916 16118
rect 18716 16055 18916 16072
rect 19164 16118 19364 16152
rect 19164 16072 19200 16118
rect 19340 16072 19364 16118
rect 19164 16055 19364 16072
rect 19612 16118 19812 16152
rect 19612 16072 19648 16118
rect 19788 16072 19812 16118
rect 19612 16055 19812 16072
rect 20060 16118 20260 16152
rect 20060 16072 20096 16118
rect 20236 16072 20260 16118
rect 20060 16055 20260 16072
rect 20508 16118 20708 16152
rect 20508 16072 20544 16118
rect 20684 16072 20708 16118
rect 20508 16055 20708 16072
rect 21292 16118 21492 16152
rect 21292 16072 21328 16118
rect 21468 16072 21492 16118
rect 21292 16055 21492 16072
rect 21740 16118 21940 16152
rect 21740 16072 21776 16118
rect 21916 16072 21940 16118
rect 21740 16055 21940 16072
rect 1692 15991 1892 16004
rect 1692 15945 1720 15991
rect 1860 15945 1892 15991
rect 1692 15912 1892 15945
rect 2140 15991 2340 16004
rect 2140 15945 2168 15991
rect 2308 15945 2340 15991
rect 2140 15912 2340 15945
rect 2588 15991 2788 16004
rect 2588 15945 2616 15991
rect 2756 15945 2788 15991
rect 2588 15912 2788 15945
rect 3036 15991 3236 16004
rect 3036 15945 3064 15991
rect 3204 15945 3236 15991
rect 3036 15912 3236 15945
rect 3484 15991 3684 16004
rect 3484 15945 3512 15991
rect 3652 15945 3684 15991
rect 3484 15912 3684 15945
rect 3932 15991 4132 16004
rect 3932 15945 3960 15991
rect 4100 15945 4132 15991
rect 3932 15912 4132 15945
rect 4380 15991 4580 16004
rect 4380 15945 4408 15991
rect 4548 15945 4580 15991
rect 4380 15912 4580 15945
rect 4828 15991 5028 16004
rect 4828 15945 4856 15991
rect 4996 15945 5028 15991
rect 4828 15912 5028 15945
rect 5612 15991 5812 16004
rect 5612 15945 5640 15991
rect 5780 15945 5812 15991
rect 5612 15912 5812 15945
rect 6060 15991 6260 16004
rect 6060 15945 6088 15991
rect 6228 15945 6260 15991
rect 6060 15912 6260 15945
rect 6508 15991 6708 16004
rect 6508 15945 6536 15991
rect 6676 15945 6708 15991
rect 6508 15912 6708 15945
rect 6956 15991 7156 16004
rect 6956 15945 6984 15991
rect 7124 15945 7156 15991
rect 6956 15912 7156 15945
rect 7404 15991 7604 16004
rect 7404 15945 7432 15991
rect 7572 15945 7604 15991
rect 7404 15912 7604 15945
rect 7852 15991 8052 16004
rect 7852 15945 7880 15991
rect 8020 15945 8052 15991
rect 7852 15912 8052 15945
rect 8300 15991 8500 16004
rect 8300 15945 8328 15991
rect 8468 15945 8500 15991
rect 8300 15912 8500 15945
rect 8748 15991 8948 16004
rect 8748 15945 8776 15991
rect 8916 15945 8948 15991
rect 8748 15912 8948 15945
rect 9532 15991 9732 16004
rect 9532 15945 9560 15991
rect 9700 15945 9732 15991
rect 1692 15704 1892 15748
rect 2140 15704 2340 15748
rect 2588 15704 2788 15748
rect 3036 15704 3236 15748
rect 3484 15704 3684 15748
rect 3932 15704 4132 15748
rect 4380 15704 4580 15748
rect 4828 15704 5028 15748
rect 9532 15912 9732 15945
rect 9980 15991 10180 16004
rect 9980 15945 10008 15991
rect 10148 15945 10180 15991
rect 9980 15912 10180 15945
rect 10428 15991 10628 16004
rect 10428 15945 10456 15991
rect 10596 15945 10628 15991
rect 10428 15912 10628 15945
rect 10876 15991 11076 16004
rect 10876 15945 10904 15991
rect 11044 15945 11076 15991
rect 10876 15912 11076 15945
rect 11324 15991 11524 16004
rect 11324 15945 11352 15991
rect 11492 15945 11524 15991
rect 11324 15912 11524 15945
rect 11772 15991 11972 16004
rect 11772 15945 11800 15991
rect 11940 15945 11972 15991
rect 11772 15912 11972 15945
rect 12220 15991 12420 16004
rect 12220 15945 12248 15991
rect 12388 15945 12420 15991
rect 12220 15912 12420 15945
rect 12668 15991 12868 16004
rect 12668 15945 12696 15991
rect 12836 15945 12868 15991
rect 12668 15912 12868 15945
rect 13452 15991 13652 16004
rect 13452 15945 13480 15991
rect 13620 15945 13652 15991
rect 5612 15704 5812 15748
rect 6060 15704 6260 15748
rect 6508 15704 6708 15748
rect 6956 15704 7156 15748
rect 7404 15704 7604 15748
rect 7852 15704 8052 15748
rect 8300 15704 8500 15748
rect 8748 15704 8948 15748
rect 13452 15912 13652 15945
rect 13900 15991 14100 16004
rect 13900 15945 13928 15991
rect 14068 15945 14100 15991
rect 13900 15912 14100 15945
rect 14348 15991 14548 16004
rect 14348 15945 14376 15991
rect 14516 15945 14548 15991
rect 14348 15912 14548 15945
rect 14796 15991 14996 16004
rect 14796 15945 14824 15991
rect 14964 15945 14996 15991
rect 14796 15912 14996 15945
rect 15244 15991 15444 16004
rect 15244 15945 15272 15991
rect 15412 15945 15444 15991
rect 15244 15912 15444 15945
rect 15692 15991 15892 16004
rect 15692 15945 15720 15991
rect 15860 15945 15892 15991
rect 15692 15912 15892 15945
rect 16140 15991 16340 16004
rect 16140 15945 16168 15991
rect 16308 15945 16340 15991
rect 16140 15912 16340 15945
rect 16588 15991 16788 16004
rect 16588 15945 16616 15991
rect 16756 15945 16788 15991
rect 16588 15912 16788 15945
rect 17372 15991 17572 16004
rect 17372 15945 17400 15991
rect 17540 15945 17572 15991
rect 9532 15704 9732 15748
rect 9980 15704 10180 15748
rect 10428 15704 10628 15748
rect 10876 15704 11076 15748
rect 11324 15704 11524 15748
rect 11772 15704 11972 15748
rect 12220 15704 12420 15748
rect 12668 15704 12868 15748
rect 17372 15912 17572 15945
rect 17820 15991 18020 16004
rect 17820 15945 17848 15991
rect 17988 15945 18020 15991
rect 17820 15912 18020 15945
rect 18268 15991 18468 16004
rect 18268 15945 18296 15991
rect 18436 15945 18468 15991
rect 18268 15912 18468 15945
rect 18716 15991 18916 16004
rect 18716 15945 18744 15991
rect 18884 15945 18916 15991
rect 18716 15912 18916 15945
rect 19164 15991 19364 16004
rect 19164 15945 19192 15991
rect 19332 15945 19364 15991
rect 19164 15912 19364 15945
rect 19612 15991 19812 16004
rect 19612 15945 19640 15991
rect 19780 15945 19812 15991
rect 19612 15912 19812 15945
rect 20060 15991 20260 16004
rect 20060 15945 20088 15991
rect 20228 15945 20260 15991
rect 20060 15912 20260 15945
rect 20508 15991 20708 16004
rect 20508 15945 20536 15991
rect 20676 15945 20708 15991
rect 20508 15912 20708 15945
rect 21292 15991 21492 16004
rect 21292 15945 21320 15991
rect 21460 15945 21492 15991
rect 13452 15704 13652 15748
rect 13900 15704 14100 15748
rect 14348 15704 14548 15748
rect 14796 15704 14996 15748
rect 15244 15704 15444 15748
rect 15692 15704 15892 15748
rect 16140 15704 16340 15748
rect 16588 15704 16788 15748
rect 21292 15912 21492 15945
rect 21740 15991 21940 16004
rect 21740 15945 21768 15991
rect 21908 15945 21940 15991
rect 21740 15912 21940 15945
rect 17372 15704 17572 15748
rect 17820 15704 18020 15748
rect 18268 15704 18468 15748
rect 18716 15704 18916 15748
rect 19164 15704 19364 15748
rect 19612 15704 19812 15748
rect 20060 15704 20260 15748
rect 20508 15704 20708 15748
rect 21292 15704 21492 15748
rect 21740 15704 21940 15748
rect 1692 15612 1892 15656
rect 2140 15612 2340 15656
rect 2588 15612 2788 15656
rect 3036 15612 3236 15656
rect 3484 15612 3684 15656
rect 3932 15612 4132 15656
rect 4380 15612 4580 15656
rect 4828 15612 5028 15656
rect 5276 15612 5476 15656
rect 5724 15612 5924 15656
rect 6172 15612 6372 15656
rect 6620 15612 6820 15656
rect 7068 15612 7268 15656
rect 7516 15612 7716 15656
rect 7964 15612 8164 15656
rect 8412 15612 8612 15656
rect 8860 15612 9060 15656
rect 9644 15612 9844 15656
rect 10092 15612 10292 15656
rect 10540 15612 10740 15656
rect 10988 15612 11188 15656
rect 11436 15612 11636 15656
rect 11884 15612 12084 15656
rect 12332 15612 12532 15656
rect 12780 15612 12980 15656
rect 13228 15612 13428 15656
rect 13676 15612 13876 15656
rect 14124 15612 14324 15656
rect 14572 15612 14772 15656
rect 15020 15612 15220 15656
rect 15468 15612 15668 15656
rect 15916 15612 16116 15656
rect 16364 15612 16564 15656
rect 16812 15612 17012 15656
rect 1692 15415 1892 15448
rect 1692 15369 1720 15415
rect 1860 15369 1892 15415
rect 1692 15356 1892 15369
rect 2140 15415 2340 15448
rect 2140 15369 2168 15415
rect 2308 15369 2340 15415
rect 2140 15356 2340 15369
rect 2588 15415 2788 15448
rect 2588 15369 2616 15415
rect 2756 15369 2788 15415
rect 2588 15356 2788 15369
rect 3036 15415 3236 15448
rect 3036 15369 3064 15415
rect 3204 15369 3236 15415
rect 3036 15356 3236 15369
rect 3484 15415 3684 15448
rect 3484 15369 3512 15415
rect 3652 15369 3684 15415
rect 3484 15356 3684 15369
rect 3932 15415 4132 15448
rect 3932 15369 3960 15415
rect 4100 15369 4132 15415
rect 3932 15356 4132 15369
rect 4380 15415 4580 15448
rect 4380 15369 4408 15415
rect 4548 15369 4580 15415
rect 4380 15356 4580 15369
rect 4828 15415 5028 15448
rect 4828 15369 4856 15415
rect 4996 15369 5028 15415
rect 4828 15356 5028 15369
rect 5276 15415 5476 15448
rect 5276 15369 5304 15415
rect 5444 15369 5476 15415
rect 5276 15356 5476 15369
rect 5724 15415 5924 15448
rect 5724 15369 5752 15415
rect 5892 15369 5924 15415
rect 5724 15356 5924 15369
rect 6172 15415 6372 15448
rect 6172 15369 6200 15415
rect 6340 15369 6372 15415
rect 6172 15356 6372 15369
rect 6620 15415 6820 15448
rect 6620 15369 6648 15415
rect 6788 15369 6820 15415
rect 6620 15356 6820 15369
rect 7068 15415 7268 15448
rect 7068 15369 7096 15415
rect 7236 15369 7268 15415
rect 7068 15356 7268 15369
rect 7516 15415 7716 15448
rect 7516 15369 7544 15415
rect 7684 15369 7716 15415
rect 7516 15356 7716 15369
rect 7964 15415 8164 15448
rect 7964 15369 7992 15415
rect 8132 15369 8164 15415
rect 7964 15356 8164 15369
rect 8412 15415 8612 15448
rect 8412 15369 8440 15415
rect 8580 15369 8612 15415
rect 8412 15356 8612 15369
rect 8860 15415 9060 15448
rect 17596 15612 17796 15656
rect 18044 15612 18244 15656
rect 18492 15612 18692 15656
rect 18940 15612 19140 15656
rect 19388 15612 19588 15656
rect 19836 15612 20036 15656
rect 20284 15612 20484 15656
rect 20732 15612 20932 15656
rect 21180 15612 21380 15656
rect 21628 15612 21828 15656
rect 22076 15612 22276 15656
rect 8860 15369 8888 15415
rect 9028 15369 9060 15415
rect 8860 15356 9060 15369
rect 9644 15415 9844 15448
rect 9644 15369 9672 15415
rect 9812 15369 9844 15415
rect 9644 15356 9844 15369
rect 10092 15415 10292 15448
rect 10092 15369 10120 15415
rect 10260 15369 10292 15415
rect 10092 15356 10292 15369
rect 10540 15415 10740 15448
rect 10540 15369 10568 15415
rect 10708 15369 10740 15415
rect 10540 15356 10740 15369
rect 10988 15415 11188 15448
rect 10988 15369 11016 15415
rect 11156 15369 11188 15415
rect 10988 15356 11188 15369
rect 11436 15415 11636 15448
rect 11436 15369 11464 15415
rect 11604 15369 11636 15415
rect 11436 15356 11636 15369
rect 11884 15415 12084 15448
rect 11884 15369 11912 15415
rect 12052 15369 12084 15415
rect 11884 15356 12084 15369
rect 12332 15415 12532 15448
rect 12332 15369 12360 15415
rect 12500 15369 12532 15415
rect 12332 15356 12532 15369
rect 12780 15415 12980 15448
rect 12780 15369 12808 15415
rect 12948 15369 12980 15415
rect 12780 15356 12980 15369
rect 13228 15415 13428 15448
rect 13228 15369 13256 15415
rect 13396 15369 13428 15415
rect 13228 15356 13428 15369
rect 13676 15415 13876 15448
rect 13676 15369 13704 15415
rect 13844 15369 13876 15415
rect 13676 15356 13876 15369
rect 14124 15415 14324 15448
rect 14124 15369 14152 15415
rect 14292 15369 14324 15415
rect 14124 15356 14324 15369
rect 14572 15415 14772 15448
rect 14572 15369 14600 15415
rect 14740 15369 14772 15415
rect 14572 15356 14772 15369
rect 15020 15415 15220 15448
rect 15020 15369 15048 15415
rect 15188 15369 15220 15415
rect 15020 15356 15220 15369
rect 15468 15415 15668 15448
rect 15468 15369 15496 15415
rect 15636 15369 15668 15415
rect 15468 15356 15668 15369
rect 15916 15415 16116 15448
rect 15916 15369 15944 15415
rect 16084 15369 16116 15415
rect 15916 15356 16116 15369
rect 16364 15415 16564 15448
rect 16364 15369 16392 15415
rect 16532 15369 16564 15415
rect 16364 15356 16564 15369
rect 16812 15415 17012 15448
rect 16812 15369 16840 15415
rect 16980 15369 17012 15415
rect 16812 15356 17012 15369
rect 17596 15415 17796 15448
rect 17596 15369 17624 15415
rect 17764 15369 17796 15415
rect 17596 15356 17796 15369
rect 18044 15415 18244 15448
rect 18044 15369 18072 15415
rect 18212 15369 18244 15415
rect 18044 15356 18244 15369
rect 18492 15415 18692 15448
rect 18492 15369 18520 15415
rect 18660 15369 18692 15415
rect 18492 15356 18692 15369
rect 18940 15415 19140 15448
rect 18940 15369 18968 15415
rect 19108 15369 19140 15415
rect 18940 15356 19140 15369
rect 19388 15415 19588 15448
rect 19388 15369 19416 15415
rect 19556 15369 19588 15415
rect 19388 15356 19588 15369
rect 19836 15415 20036 15448
rect 19836 15369 19864 15415
rect 20004 15369 20036 15415
rect 19836 15356 20036 15369
rect 20284 15415 20484 15448
rect 20284 15369 20312 15415
rect 20452 15369 20484 15415
rect 20284 15356 20484 15369
rect 20732 15415 20932 15448
rect 20732 15369 20760 15415
rect 20900 15369 20932 15415
rect 20732 15356 20932 15369
rect 21180 15415 21380 15448
rect 21180 15369 21208 15415
rect 21348 15369 21380 15415
rect 21180 15356 21380 15369
rect 21628 15415 21828 15448
rect 21628 15369 21656 15415
rect 21796 15369 21828 15415
rect 21628 15356 21828 15369
rect 22076 15415 22276 15448
rect 22076 15369 22104 15415
rect 22244 15369 22276 15415
rect 22076 15356 22276 15369
rect 1692 15288 1892 15305
rect 1692 15242 1728 15288
rect 1868 15242 1892 15288
rect 1692 15208 1892 15242
rect 2140 15288 2340 15305
rect 2140 15242 2176 15288
rect 2316 15242 2340 15288
rect 2140 15208 2340 15242
rect 2588 15288 2788 15305
rect 2588 15242 2624 15288
rect 2764 15242 2788 15288
rect 2588 15208 2788 15242
rect 3036 15288 3236 15305
rect 3036 15242 3072 15288
rect 3212 15242 3236 15288
rect 3036 15208 3236 15242
rect 3484 15288 3684 15305
rect 3484 15242 3520 15288
rect 3660 15242 3684 15288
rect 3484 15208 3684 15242
rect 3932 15288 4132 15305
rect 3932 15242 3968 15288
rect 4108 15242 4132 15288
rect 3932 15208 4132 15242
rect 4380 15288 4580 15305
rect 4380 15242 4416 15288
rect 4556 15242 4580 15288
rect 4380 15208 4580 15242
rect 4828 15288 5028 15305
rect 4828 15242 4864 15288
rect 5004 15242 5028 15288
rect 4828 15208 5028 15242
rect 5276 15288 5476 15305
rect 5276 15242 5312 15288
rect 5452 15242 5476 15288
rect 5276 15208 5476 15242
rect 5724 15288 5924 15305
rect 5724 15242 5760 15288
rect 5900 15242 5924 15288
rect 5724 15208 5924 15242
rect 6172 15288 6372 15305
rect 6172 15242 6208 15288
rect 6348 15242 6372 15288
rect 6172 15208 6372 15242
rect 6620 15288 6820 15305
rect 6620 15242 6656 15288
rect 6796 15242 6820 15288
rect 6620 15208 6820 15242
rect 7068 15288 7268 15305
rect 7068 15242 7104 15288
rect 7244 15242 7268 15288
rect 7068 15208 7268 15242
rect 7516 15288 7716 15305
rect 7516 15242 7552 15288
rect 7692 15242 7716 15288
rect 7516 15208 7716 15242
rect 7964 15288 8164 15305
rect 7964 15242 8000 15288
rect 8140 15242 8164 15288
rect 7964 15208 8164 15242
rect 8412 15288 8612 15305
rect 8412 15242 8448 15288
rect 8588 15242 8612 15288
rect 8412 15208 8612 15242
rect 8860 15288 9060 15305
rect 8860 15242 8896 15288
rect 9036 15242 9060 15288
rect 8860 15208 9060 15242
rect 9644 15288 9844 15305
rect 9644 15242 9680 15288
rect 9820 15242 9844 15288
rect 9644 15208 9844 15242
rect 10092 15288 10292 15305
rect 10092 15242 10128 15288
rect 10268 15242 10292 15288
rect 10092 15208 10292 15242
rect 10540 15288 10740 15305
rect 10540 15242 10576 15288
rect 10716 15242 10740 15288
rect 10540 15208 10740 15242
rect 10988 15288 11188 15305
rect 10988 15242 11024 15288
rect 11164 15242 11188 15288
rect 10988 15208 11188 15242
rect 11436 15288 11636 15305
rect 11436 15242 11472 15288
rect 11612 15242 11636 15288
rect 11436 15208 11636 15242
rect 11884 15288 12084 15305
rect 11884 15242 11920 15288
rect 12060 15242 12084 15288
rect 11884 15208 12084 15242
rect 12332 15288 12532 15305
rect 12332 15242 12368 15288
rect 12508 15242 12532 15288
rect 12332 15208 12532 15242
rect 12780 15288 12980 15305
rect 12780 15242 12816 15288
rect 12956 15242 12980 15288
rect 12780 15208 12980 15242
rect 13228 15288 13428 15305
rect 13228 15242 13264 15288
rect 13404 15242 13428 15288
rect 13228 15208 13428 15242
rect 13676 15288 13876 15305
rect 13676 15242 13712 15288
rect 13852 15242 13876 15288
rect 13676 15208 13876 15242
rect 14124 15288 14324 15305
rect 14124 15242 14160 15288
rect 14300 15242 14324 15288
rect 14124 15208 14324 15242
rect 14572 15288 14772 15305
rect 14572 15242 14608 15288
rect 14748 15242 14772 15288
rect 14572 15208 14772 15242
rect 15020 15288 15220 15305
rect 15020 15242 15056 15288
rect 15196 15242 15220 15288
rect 15020 15208 15220 15242
rect 15468 15288 15668 15305
rect 15468 15242 15504 15288
rect 15644 15242 15668 15288
rect 15468 15208 15668 15242
rect 15916 15288 16116 15305
rect 15916 15242 15952 15288
rect 16092 15242 16116 15288
rect 15916 15208 16116 15242
rect 16364 15288 16564 15305
rect 16364 15242 16400 15288
rect 16540 15242 16564 15288
rect 16364 15208 16564 15242
rect 16812 15288 17012 15305
rect 16812 15242 16848 15288
rect 16988 15242 17012 15288
rect 16812 15208 17012 15242
rect 17596 15288 17796 15305
rect 17596 15242 17632 15288
rect 17772 15242 17796 15288
rect 17596 15208 17796 15242
rect 18044 15288 18244 15305
rect 18044 15242 18080 15288
rect 18220 15242 18244 15288
rect 18044 15208 18244 15242
rect 18492 15288 18692 15305
rect 18492 15242 18528 15288
rect 18668 15242 18692 15288
rect 18492 15208 18692 15242
rect 18940 15288 19140 15305
rect 18940 15242 18976 15288
rect 19116 15242 19140 15288
rect 18940 15208 19140 15242
rect 19388 15288 19588 15305
rect 19388 15242 19424 15288
rect 19564 15242 19588 15288
rect 19388 15208 19588 15242
rect 19836 15288 20036 15305
rect 19836 15242 19872 15288
rect 20012 15242 20036 15288
rect 19836 15208 20036 15242
rect 20284 15288 20484 15305
rect 20284 15242 20320 15288
rect 20460 15242 20484 15288
rect 20284 15208 20484 15242
rect 20732 15288 20932 15305
rect 20732 15242 20768 15288
rect 20908 15242 20932 15288
rect 20732 15208 20932 15242
rect 21180 15288 21380 15305
rect 21180 15242 21216 15288
rect 21356 15242 21380 15288
rect 21180 15208 21380 15242
rect 21628 15288 21828 15305
rect 21628 15242 21664 15288
rect 21804 15242 21828 15288
rect 21628 15208 21828 15242
rect 22076 15288 22276 15305
rect 22076 15242 22112 15288
rect 22252 15242 22276 15288
rect 22076 15208 22276 15242
rect 1692 14920 1892 14964
rect 2140 14920 2340 14964
rect 2588 14920 2788 14964
rect 3036 14920 3236 14964
rect 3484 14920 3684 14964
rect 3932 14920 4132 14964
rect 4380 14920 4580 14964
rect 4828 14920 5028 14964
rect 5276 14920 5476 14964
rect 5724 14920 5924 14964
rect 6172 14920 6372 14964
rect 6620 14920 6820 14964
rect 7068 14920 7268 14964
rect 7516 14920 7716 14964
rect 7964 14920 8164 14964
rect 8412 14920 8612 14964
rect 8860 14920 9060 14964
rect 9644 14920 9844 14964
rect 10092 14920 10292 14964
rect 10540 14920 10740 14964
rect 10988 14920 11188 14964
rect 11436 14920 11636 14964
rect 11884 14920 12084 14964
rect 12332 14920 12532 14964
rect 12780 14920 12980 14964
rect 13228 14920 13428 14964
rect 13676 14920 13876 14964
rect 14124 14920 14324 14964
rect 14572 14920 14772 14964
rect 15020 14920 15220 14964
rect 15468 14920 15668 14964
rect 15916 14920 16116 14964
rect 16364 14920 16564 14964
rect 16812 14920 17012 14964
rect 17596 14920 17796 14964
rect 18044 14920 18244 14964
rect 18492 14920 18692 14964
rect 18940 14920 19140 14964
rect 19388 14920 19588 14964
rect 19836 14920 20036 14964
rect 20284 14920 20484 14964
rect 20732 14920 20932 14964
rect 21180 14920 21380 14964
rect 21628 14920 21828 14964
rect 22076 14920 22276 14964
rect 1692 14828 1892 14872
rect 2140 14828 2340 14872
rect 2588 14828 2788 14872
rect 3036 14828 3236 14872
rect 3484 14828 3684 14872
rect 3932 14828 4132 14872
rect 4380 14828 4580 14872
rect 4828 14828 5028 14872
rect 5612 14828 5812 14872
rect 6060 14828 6260 14872
rect 6508 14828 6708 14872
rect 6956 14828 7156 14872
rect 7404 14828 7604 14872
rect 7852 14828 8052 14872
rect 8300 14828 8500 14872
rect 8748 14828 8948 14872
rect 9196 14828 9396 14872
rect 9644 14828 9844 14872
rect 10092 14828 10292 14872
rect 10540 14828 10740 14872
rect 10988 14828 11188 14872
rect 11436 14828 11636 14872
rect 11884 14828 12084 14872
rect 12332 14828 12532 14872
rect 12780 14828 12980 14872
rect 13564 14828 13764 14872
rect 14012 14828 14212 14872
rect 14460 14828 14660 14872
rect 14908 14828 15108 14872
rect 15356 14828 15556 14872
rect 15804 14828 16004 14872
rect 16252 14828 16452 14872
rect 16892 14828 16992 14872
rect 17564 14828 17664 14872
rect 17932 14828 18132 14872
rect 18380 14828 18580 14872
rect 18828 14828 19028 14872
rect 19276 14828 19476 14872
rect 19724 14828 19924 14872
rect 20172 14828 20372 14872
rect 20620 14828 20820 14872
rect 21516 14828 21716 14872
rect 21964 14828 22164 14872
rect 1692 14550 1892 14584
rect 1692 14504 1728 14550
rect 1868 14504 1892 14550
rect 1692 14487 1892 14504
rect 2140 14550 2340 14584
rect 2140 14504 2176 14550
rect 2316 14504 2340 14550
rect 2140 14487 2340 14504
rect 2588 14550 2788 14584
rect 2588 14504 2624 14550
rect 2764 14504 2788 14550
rect 2588 14487 2788 14504
rect 3036 14550 3236 14584
rect 3036 14504 3072 14550
rect 3212 14504 3236 14550
rect 3036 14487 3236 14504
rect 3484 14550 3684 14584
rect 3484 14504 3520 14550
rect 3660 14504 3684 14550
rect 3484 14487 3684 14504
rect 3932 14550 4132 14584
rect 3932 14504 3968 14550
rect 4108 14504 4132 14550
rect 3932 14487 4132 14504
rect 4380 14550 4580 14584
rect 4380 14504 4416 14550
rect 4556 14504 4580 14550
rect 4380 14487 4580 14504
rect 4828 14550 5028 14584
rect 4828 14504 4864 14550
rect 5004 14504 5028 14550
rect 4828 14487 5028 14504
rect 5612 14550 5812 14584
rect 5612 14504 5648 14550
rect 5788 14504 5812 14550
rect 5612 14487 5812 14504
rect 6060 14550 6260 14584
rect 6060 14504 6096 14550
rect 6236 14504 6260 14550
rect 6060 14487 6260 14504
rect 6508 14550 6708 14584
rect 6508 14504 6544 14550
rect 6684 14504 6708 14550
rect 6508 14487 6708 14504
rect 6956 14550 7156 14584
rect 6956 14504 6992 14550
rect 7132 14504 7156 14550
rect 6956 14487 7156 14504
rect 7404 14550 7604 14584
rect 7404 14504 7440 14550
rect 7580 14504 7604 14550
rect 7404 14487 7604 14504
rect 7852 14550 8052 14584
rect 7852 14504 7888 14550
rect 8028 14504 8052 14550
rect 7852 14487 8052 14504
rect 8300 14550 8500 14584
rect 8300 14504 8336 14550
rect 8476 14504 8500 14550
rect 8300 14487 8500 14504
rect 8748 14550 8948 14584
rect 8748 14504 8784 14550
rect 8924 14504 8948 14550
rect 8748 14487 8948 14504
rect 9196 14550 9396 14584
rect 9196 14504 9232 14550
rect 9372 14504 9396 14550
rect 9196 14487 9396 14504
rect 9644 14550 9844 14584
rect 9644 14504 9680 14550
rect 9820 14504 9844 14550
rect 9644 14487 9844 14504
rect 10092 14550 10292 14584
rect 10092 14504 10128 14550
rect 10268 14504 10292 14550
rect 10092 14487 10292 14504
rect 10540 14550 10740 14584
rect 10540 14504 10576 14550
rect 10716 14504 10740 14550
rect 10540 14487 10740 14504
rect 10988 14550 11188 14584
rect 10988 14504 11024 14550
rect 11164 14504 11188 14550
rect 10988 14487 11188 14504
rect 11436 14550 11636 14584
rect 11436 14504 11472 14550
rect 11612 14504 11636 14550
rect 11436 14487 11636 14504
rect 11884 14550 12084 14584
rect 11884 14504 11920 14550
rect 12060 14504 12084 14550
rect 11884 14487 12084 14504
rect 12332 14550 12532 14584
rect 12332 14504 12368 14550
rect 12508 14504 12532 14550
rect 12332 14487 12532 14504
rect 12780 14550 12980 14584
rect 12780 14504 12816 14550
rect 12956 14504 12980 14550
rect 12780 14487 12980 14504
rect 13564 14550 13764 14584
rect 13564 14504 13600 14550
rect 13740 14504 13764 14550
rect 13564 14487 13764 14504
rect 14012 14550 14212 14584
rect 14012 14504 14048 14550
rect 14188 14504 14212 14550
rect 14012 14487 14212 14504
rect 14460 14550 14660 14584
rect 14460 14504 14496 14550
rect 14636 14504 14660 14550
rect 14460 14487 14660 14504
rect 14908 14550 15108 14584
rect 14908 14504 14944 14550
rect 15084 14504 15108 14550
rect 14908 14487 15108 14504
rect 15356 14550 15556 14584
rect 15356 14504 15392 14550
rect 15532 14504 15556 14550
rect 15356 14487 15556 14504
rect 15804 14550 16004 14584
rect 15804 14504 15840 14550
rect 15980 14504 16004 14550
rect 15804 14487 16004 14504
rect 16252 14550 16452 14584
rect 16252 14504 16288 14550
rect 16428 14504 16452 14550
rect 16252 14487 16452 14504
rect 16892 14535 16992 14584
rect 1692 14423 1892 14436
rect 1692 14377 1720 14423
rect 1860 14377 1892 14423
rect 1692 14344 1892 14377
rect 2140 14423 2340 14436
rect 2140 14377 2168 14423
rect 2308 14377 2340 14423
rect 2140 14344 2340 14377
rect 2588 14423 2788 14436
rect 2588 14377 2616 14423
rect 2756 14377 2788 14423
rect 2588 14344 2788 14377
rect 3036 14423 3236 14436
rect 3036 14377 3064 14423
rect 3204 14377 3236 14423
rect 3036 14344 3236 14377
rect 3484 14423 3684 14436
rect 3484 14377 3512 14423
rect 3652 14377 3684 14423
rect 3484 14344 3684 14377
rect 3932 14423 4132 14436
rect 3932 14377 3960 14423
rect 4100 14377 4132 14423
rect 3932 14344 4132 14377
rect 4380 14423 4580 14436
rect 4380 14377 4408 14423
rect 4548 14377 4580 14423
rect 4380 14344 4580 14377
rect 4828 14423 5028 14436
rect 4828 14377 4856 14423
rect 4996 14377 5028 14423
rect 4828 14344 5028 14377
rect 5612 14423 5812 14436
rect 5612 14377 5640 14423
rect 5780 14377 5812 14423
rect 5612 14344 5812 14377
rect 6060 14423 6260 14436
rect 6060 14377 6088 14423
rect 6228 14377 6260 14423
rect 6060 14344 6260 14377
rect 6508 14423 6708 14436
rect 6508 14377 6536 14423
rect 6676 14377 6708 14423
rect 6508 14344 6708 14377
rect 6956 14423 7156 14436
rect 6956 14377 6984 14423
rect 7124 14377 7156 14423
rect 6956 14344 7156 14377
rect 7404 14423 7604 14436
rect 7404 14377 7432 14423
rect 7572 14377 7604 14423
rect 7404 14344 7604 14377
rect 7852 14423 8052 14436
rect 7852 14377 7880 14423
rect 8020 14377 8052 14423
rect 7852 14344 8052 14377
rect 8300 14423 8500 14436
rect 8300 14377 8328 14423
rect 8468 14377 8500 14423
rect 8300 14344 8500 14377
rect 8748 14423 8948 14436
rect 8748 14377 8776 14423
rect 8916 14377 8948 14423
rect 8748 14344 8948 14377
rect 9196 14423 9396 14436
rect 9196 14377 9224 14423
rect 9364 14377 9396 14423
rect 9196 14344 9396 14377
rect 9644 14423 9844 14436
rect 9644 14377 9672 14423
rect 9812 14377 9844 14423
rect 9644 14344 9844 14377
rect 10092 14423 10292 14436
rect 10092 14377 10120 14423
rect 10260 14377 10292 14423
rect 10092 14344 10292 14377
rect 10540 14423 10740 14436
rect 10540 14377 10568 14423
rect 10708 14377 10740 14423
rect 10540 14344 10740 14377
rect 10988 14423 11188 14436
rect 10988 14377 11016 14423
rect 11156 14377 11188 14423
rect 10988 14344 11188 14377
rect 11436 14423 11636 14436
rect 11436 14377 11464 14423
rect 11604 14377 11636 14423
rect 11436 14344 11636 14377
rect 11884 14423 12084 14436
rect 11884 14377 11912 14423
rect 12052 14377 12084 14423
rect 11884 14344 12084 14377
rect 12332 14423 12532 14436
rect 12332 14377 12360 14423
rect 12500 14377 12532 14423
rect 12332 14344 12532 14377
rect 12780 14423 12980 14436
rect 12780 14377 12808 14423
rect 12948 14377 12980 14423
rect 12780 14344 12980 14377
rect 13564 14423 13764 14436
rect 13564 14377 13592 14423
rect 13732 14377 13764 14423
rect 1692 14136 1892 14180
rect 2140 14136 2340 14180
rect 2588 14136 2788 14180
rect 3036 14136 3236 14180
rect 3484 14136 3684 14180
rect 3932 14136 4132 14180
rect 4380 14136 4580 14180
rect 4828 14136 5028 14180
rect 13564 14344 13764 14377
rect 14012 14423 14212 14436
rect 14012 14377 14040 14423
rect 14180 14377 14212 14423
rect 14012 14344 14212 14377
rect 14460 14423 14660 14436
rect 14460 14377 14488 14423
rect 14628 14377 14660 14423
rect 14460 14344 14660 14377
rect 14908 14423 15108 14436
rect 14908 14377 14936 14423
rect 15076 14377 15108 14423
rect 14908 14344 15108 14377
rect 15356 14423 15556 14436
rect 15356 14377 15384 14423
rect 15524 14377 15556 14423
rect 15356 14344 15556 14377
rect 15804 14423 16004 14436
rect 15804 14377 15832 14423
rect 15972 14377 16004 14423
rect 15804 14344 16004 14377
rect 16252 14423 16452 14436
rect 16252 14377 16280 14423
rect 16420 14377 16452 14423
rect 16252 14344 16452 14377
rect 16892 14395 16933 14535
rect 16979 14498 16992 14535
rect 17564 14535 17664 14584
rect 16979 14395 17012 14498
rect 16892 14344 17012 14395
rect 17564 14395 17605 14535
rect 17651 14498 17664 14535
rect 17932 14550 18132 14584
rect 17932 14504 17968 14550
rect 18108 14504 18132 14550
rect 17651 14395 17684 14498
rect 17932 14487 18132 14504
rect 18380 14550 18580 14584
rect 18380 14504 18416 14550
rect 18556 14504 18580 14550
rect 18380 14487 18580 14504
rect 18828 14550 19028 14584
rect 18828 14504 18864 14550
rect 19004 14504 19028 14550
rect 18828 14487 19028 14504
rect 19276 14550 19476 14584
rect 19276 14504 19312 14550
rect 19452 14504 19476 14550
rect 19276 14487 19476 14504
rect 19724 14550 19924 14584
rect 19724 14504 19760 14550
rect 19900 14504 19924 14550
rect 19724 14487 19924 14504
rect 20172 14550 20372 14584
rect 20172 14504 20208 14550
rect 20348 14504 20372 14550
rect 20172 14487 20372 14504
rect 20620 14550 20820 14584
rect 20620 14504 20656 14550
rect 20796 14504 20820 14550
rect 20620 14487 20820 14504
rect 21516 14550 21716 14584
rect 21516 14504 21552 14550
rect 21692 14504 21716 14550
rect 21516 14487 21716 14504
rect 21964 14550 22164 14584
rect 21964 14504 22000 14550
rect 22140 14504 22164 14550
rect 21964 14487 22164 14504
rect 17564 14344 17684 14395
rect 17932 14423 18132 14436
rect 17932 14377 17960 14423
rect 18100 14377 18132 14423
rect 17932 14344 18132 14377
rect 18380 14423 18580 14436
rect 18380 14377 18408 14423
rect 18548 14377 18580 14423
rect 18380 14344 18580 14377
rect 18828 14423 19028 14436
rect 18828 14377 18856 14423
rect 18996 14377 19028 14423
rect 18828 14344 19028 14377
rect 19276 14423 19476 14436
rect 19276 14377 19304 14423
rect 19444 14377 19476 14423
rect 19276 14344 19476 14377
rect 19724 14423 19924 14436
rect 19724 14377 19752 14423
rect 19892 14377 19924 14423
rect 19724 14344 19924 14377
rect 20172 14423 20372 14436
rect 20172 14377 20200 14423
rect 20340 14377 20372 14423
rect 20172 14344 20372 14377
rect 20620 14423 20820 14436
rect 20620 14377 20648 14423
rect 20788 14377 20820 14423
rect 20620 14344 20820 14377
rect 21516 14423 21716 14436
rect 21516 14377 21544 14423
rect 21684 14377 21716 14423
rect 5612 14136 5812 14180
rect 6060 14136 6260 14180
rect 6508 14136 6708 14180
rect 6956 14136 7156 14180
rect 7404 14136 7604 14180
rect 7852 14136 8052 14180
rect 8300 14136 8500 14180
rect 8748 14136 8948 14180
rect 9196 14136 9396 14180
rect 9644 14136 9844 14180
rect 10092 14136 10292 14180
rect 10540 14136 10740 14180
rect 10988 14136 11188 14180
rect 11436 14136 11636 14180
rect 11884 14136 12084 14180
rect 12332 14136 12532 14180
rect 12780 14136 12980 14180
rect 21516 14344 21716 14377
rect 21964 14423 22164 14436
rect 21964 14377 21992 14423
rect 22132 14377 22164 14423
rect 21964 14344 22164 14377
rect 13564 14136 13764 14180
rect 14012 14136 14212 14180
rect 14460 14136 14660 14180
rect 14908 14136 15108 14180
rect 15356 14136 15556 14180
rect 15804 14136 16004 14180
rect 16252 14136 16452 14180
rect 16892 14136 17012 14180
rect 17564 14136 17684 14180
rect 17932 14136 18132 14180
rect 18380 14136 18580 14180
rect 18828 14136 19028 14180
rect 19276 14136 19476 14180
rect 19724 14136 19924 14180
rect 20172 14136 20372 14180
rect 20620 14136 20820 14180
rect 21516 14136 21716 14180
rect 21964 14136 22164 14180
rect 1692 14044 1892 14088
rect 2140 14044 2340 14088
rect 2588 14044 2788 14088
rect 3036 14044 3236 14088
rect 3484 14044 3684 14088
rect 3932 14044 4132 14088
rect 4380 14044 4580 14088
rect 4828 14044 5028 14088
rect 5276 14044 5476 14088
rect 5724 14044 5924 14088
rect 6172 14044 6372 14088
rect 6620 14044 6820 14088
rect 7068 14044 7268 14088
rect 7516 14044 7716 14088
rect 7964 14044 8164 14088
rect 8412 14044 8612 14088
rect 8860 14044 9060 14088
rect 9644 14044 9844 14088
rect 10092 14044 10292 14088
rect 10540 14044 10740 14088
rect 10988 14044 11188 14088
rect 11436 14044 11636 14088
rect 11884 14044 12084 14088
rect 12332 14044 12532 14088
rect 12780 14044 12980 14088
rect 13228 14044 13428 14088
rect 13676 14044 13876 14088
rect 14124 14044 14324 14088
rect 14572 14044 14772 14088
rect 15020 14044 15220 14088
rect 15468 14044 15668 14088
rect 16140 14044 16260 14088
rect 16812 14044 16932 14088
rect 1692 13847 1892 13880
rect 1692 13801 1720 13847
rect 1860 13801 1892 13847
rect 1692 13788 1892 13801
rect 2140 13847 2340 13880
rect 2140 13801 2168 13847
rect 2308 13801 2340 13847
rect 2140 13788 2340 13801
rect 2588 13847 2788 13880
rect 2588 13801 2616 13847
rect 2756 13801 2788 13847
rect 2588 13788 2788 13801
rect 3036 13847 3236 13880
rect 3036 13801 3064 13847
rect 3204 13801 3236 13847
rect 3036 13788 3236 13801
rect 3484 13847 3684 13880
rect 3484 13801 3512 13847
rect 3652 13801 3684 13847
rect 3484 13788 3684 13801
rect 3932 13847 4132 13880
rect 3932 13801 3960 13847
rect 4100 13801 4132 13847
rect 3932 13788 4132 13801
rect 4380 13847 4580 13880
rect 4380 13801 4408 13847
rect 4548 13801 4580 13847
rect 4380 13788 4580 13801
rect 4828 13847 5028 13880
rect 4828 13801 4856 13847
rect 4996 13801 5028 13847
rect 4828 13788 5028 13801
rect 5276 13847 5476 13880
rect 5276 13801 5304 13847
rect 5444 13801 5476 13847
rect 5276 13788 5476 13801
rect 5724 13847 5924 13880
rect 5724 13801 5752 13847
rect 5892 13801 5924 13847
rect 5724 13788 5924 13801
rect 6172 13847 6372 13880
rect 6172 13801 6200 13847
rect 6340 13801 6372 13847
rect 6172 13788 6372 13801
rect 6620 13847 6820 13880
rect 6620 13801 6648 13847
rect 6788 13801 6820 13847
rect 6620 13788 6820 13801
rect 7068 13847 7268 13880
rect 7068 13801 7096 13847
rect 7236 13801 7268 13847
rect 7068 13788 7268 13801
rect 7516 13847 7716 13880
rect 7516 13801 7544 13847
rect 7684 13801 7716 13847
rect 7516 13788 7716 13801
rect 7964 13847 8164 13880
rect 7964 13801 7992 13847
rect 8132 13801 8164 13847
rect 7964 13788 8164 13801
rect 8412 13847 8612 13880
rect 8412 13801 8440 13847
rect 8580 13801 8612 13847
rect 8412 13788 8612 13801
rect 8860 13847 9060 13880
rect 17708 14044 17828 14088
rect 18380 14044 18500 14088
rect 18828 14044 19028 14088
rect 19276 14044 19476 14088
rect 19724 14044 19924 14088
rect 20172 14044 20372 14088
rect 20620 14044 20820 14088
rect 21068 14044 21268 14088
rect 21516 14044 21716 14088
rect 21964 14044 22164 14088
rect 8860 13801 8888 13847
rect 9028 13801 9060 13847
rect 8860 13788 9060 13801
rect 9644 13847 9844 13880
rect 9644 13801 9672 13847
rect 9812 13801 9844 13847
rect 9644 13788 9844 13801
rect 10092 13847 10292 13880
rect 10092 13801 10120 13847
rect 10260 13801 10292 13847
rect 10092 13788 10292 13801
rect 10540 13847 10740 13880
rect 10540 13801 10568 13847
rect 10708 13801 10740 13847
rect 10540 13788 10740 13801
rect 10988 13847 11188 13880
rect 10988 13801 11016 13847
rect 11156 13801 11188 13847
rect 10988 13788 11188 13801
rect 11436 13847 11636 13880
rect 11436 13801 11464 13847
rect 11604 13801 11636 13847
rect 11436 13788 11636 13801
rect 11884 13847 12084 13880
rect 11884 13801 11912 13847
rect 12052 13801 12084 13847
rect 11884 13788 12084 13801
rect 12332 13847 12532 13880
rect 12332 13801 12360 13847
rect 12500 13801 12532 13847
rect 12332 13788 12532 13801
rect 12780 13847 12980 13880
rect 12780 13801 12808 13847
rect 12948 13801 12980 13847
rect 12780 13788 12980 13801
rect 13228 13847 13428 13880
rect 13228 13801 13256 13847
rect 13396 13801 13428 13847
rect 13228 13788 13428 13801
rect 13676 13847 13876 13880
rect 13676 13801 13704 13847
rect 13844 13801 13876 13847
rect 13676 13788 13876 13801
rect 14124 13847 14324 13880
rect 14124 13801 14152 13847
rect 14292 13801 14324 13847
rect 14124 13788 14324 13801
rect 14572 13847 14772 13880
rect 14572 13801 14600 13847
rect 14740 13801 14772 13847
rect 14572 13788 14772 13801
rect 15020 13847 15220 13880
rect 15020 13801 15048 13847
rect 15188 13801 15220 13847
rect 15020 13788 15220 13801
rect 15468 13847 15668 13880
rect 15468 13801 15496 13847
rect 15636 13801 15668 13847
rect 15468 13788 15668 13801
rect 16140 13829 16260 13880
rect 1692 13720 1892 13737
rect 1692 13674 1728 13720
rect 1868 13674 1892 13720
rect 1692 13640 1892 13674
rect 2140 13720 2340 13737
rect 2140 13674 2176 13720
rect 2316 13674 2340 13720
rect 2140 13640 2340 13674
rect 2588 13720 2788 13737
rect 2588 13674 2624 13720
rect 2764 13674 2788 13720
rect 2588 13640 2788 13674
rect 3036 13720 3236 13737
rect 3036 13674 3072 13720
rect 3212 13674 3236 13720
rect 3036 13640 3236 13674
rect 3484 13720 3684 13737
rect 3484 13674 3520 13720
rect 3660 13674 3684 13720
rect 3484 13640 3684 13674
rect 3932 13720 4132 13737
rect 3932 13674 3968 13720
rect 4108 13674 4132 13720
rect 3932 13640 4132 13674
rect 4380 13720 4580 13737
rect 4380 13674 4416 13720
rect 4556 13674 4580 13720
rect 4380 13640 4580 13674
rect 4828 13720 5028 13737
rect 4828 13674 4864 13720
rect 5004 13674 5028 13720
rect 4828 13640 5028 13674
rect 5276 13720 5476 13737
rect 5276 13674 5312 13720
rect 5452 13674 5476 13720
rect 5276 13640 5476 13674
rect 5724 13720 5924 13737
rect 5724 13674 5760 13720
rect 5900 13674 5924 13720
rect 5724 13640 5924 13674
rect 6172 13720 6372 13737
rect 6172 13674 6208 13720
rect 6348 13674 6372 13720
rect 6172 13640 6372 13674
rect 6620 13720 6820 13737
rect 6620 13674 6656 13720
rect 6796 13674 6820 13720
rect 6620 13640 6820 13674
rect 7068 13720 7268 13737
rect 7068 13674 7104 13720
rect 7244 13674 7268 13720
rect 7068 13640 7268 13674
rect 7516 13720 7716 13737
rect 7516 13674 7552 13720
rect 7692 13674 7716 13720
rect 7516 13640 7716 13674
rect 7964 13720 8164 13737
rect 7964 13674 8000 13720
rect 8140 13674 8164 13720
rect 7964 13640 8164 13674
rect 8412 13720 8612 13737
rect 8412 13674 8448 13720
rect 8588 13674 8612 13720
rect 8412 13640 8612 13674
rect 8860 13720 9060 13737
rect 8860 13674 8896 13720
rect 9036 13674 9060 13720
rect 8860 13640 9060 13674
rect 9644 13720 9844 13737
rect 9644 13674 9680 13720
rect 9820 13674 9844 13720
rect 9644 13640 9844 13674
rect 10092 13720 10292 13737
rect 10092 13674 10128 13720
rect 10268 13674 10292 13720
rect 10092 13640 10292 13674
rect 10540 13720 10740 13737
rect 10540 13674 10576 13720
rect 10716 13674 10740 13720
rect 10540 13640 10740 13674
rect 10988 13720 11188 13737
rect 10988 13674 11024 13720
rect 11164 13674 11188 13720
rect 10988 13640 11188 13674
rect 11436 13720 11636 13737
rect 11436 13674 11472 13720
rect 11612 13674 11636 13720
rect 11436 13640 11636 13674
rect 11884 13720 12084 13737
rect 11884 13674 11920 13720
rect 12060 13674 12084 13720
rect 11884 13640 12084 13674
rect 12332 13720 12532 13737
rect 12332 13674 12368 13720
rect 12508 13674 12532 13720
rect 12332 13640 12532 13674
rect 12780 13720 12980 13737
rect 12780 13674 12816 13720
rect 12956 13674 12980 13720
rect 12780 13640 12980 13674
rect 13228 13720 13428 13737
rect 13228 13674 13264 13720
rect 13404 13674 13428 13720
rect 13228 13640 13428 13674
rect 13676 13720 13876 13737
rect 13676 13674 13712 13720
rect 13852 13674 13876 13720
rect 13676 13640 13876 13674
rect 14124 13720 14324 13737
rect 14124 13674 14160 13720
rect 14300 13674 14324 13720
rect 14124 13640 14324 13674
rect 14572 13720 14772 13737
rect 14572 13674 14608 13720
rect 14748 13674 14772 13720
rect 14572 13640 14772 13674
rect 15020 13720 15220 13737
rect 15020 13674 15056 13720
rect 15196 13674 15220 13720
rect 15020 13640 15220 13674
rect 15468 13720 15668 13737
rect 16140 13726 16173 13829
rect 15468 13674 15504 13720
rect 15644 13674 15668 13720
rect 15468 13640 15668 13674
rect 16160 13689 16173 13726
rect 16219 13689 16260 13829
rect 16812 13829 16932 13880
rect 16812 13726 16845 13829
rect 16160 13640 16260 13689
rect 16832 13689 16845 13726
rect 16891 13689 16932 13829
rect 17708 13829 17828 13880
rect 16832 13640 16932 13689
rect 17708 13726 17741 13829
rect 17728 13689 17741 13726
rect 17787 13689 17828 13829
rect 18380 13829 18500 13880
rect 18380 13726 18413 13829
rect 17728 13640 17828 13689
rect 18400 13689 18413 13726
rect 18459 13689 18500 13829
rect 18828 13847 19028 13880
rect 18828 13801 18856 13847
rect 18996 13801 19028 13847
rect 18828 13788 19028 13801
rect 19276 13847 19476 13880
rect 19276 13801 19304 13847
rect 19444 13801 19476 13847
rect 19276 13788 19476 13801
rect 19724 13847 19924 13880
rect 19724 13801 19752 13847
rect 19892 13801 19924 13847
rect 19724 13788 19924 13801
rect 20172 13847 20372 13880
rect 20172 13801 20200 13847
rect 20340 13801 20372 13847
rect 20172 13788 20372 13801
rect 20620 13847 20820 13880
rect 20620 13801 20648 13847
rect 20788 13801 20820 13847
rect 20620 13788 20820 13801
rect 21068 13847 21268 13880
rect 21068 13801 21096 13847
rect 21236 13801 21268 13847
rect 21068 13788 21268 13801
rect 21516 13847 21716 13880
rect 21516 13801 21544 13847
rect 21684 13801 21716 13847
rect 21516 13788 21716 13801
rect 21964 13847 22164 13880
rect 21964 13801 21992 13847
rect 22132 13801 22164 13847
rect 21964 13788 22164 13801
rect 18400 13640 18500 13689
rect 18828 13720 19028 13737
rect 18828 13674 18864 13720
rect 19004 13674 19028 13720
rect 18828 13640 19028 13674
rect 19276 13720 19476 13737
rect 19276 13674 19312 13720
rect 19452 13674 19476 13720
rect 19276 13640 19476 13674
rect 19724 13720 19924 13737
rect 19724 13674 19760 13720
rect 19900 13674 19924 13720
rect 19724 13640 19924 13674
rect 20172 13720 20372 13737
rect 20172 13674 20208 13720
rect 20348 13674 20372 13720
rect 20172 13640 20372 13674
rect 20620 13720 20820 13737
rect 20620 13674 20656 13720
rect 20796 13674 20820 13720
rect 20620 13640 20820 13674
rect 21068 13720 21268 13737
rect 21068 13674 21104 13720
rect 21244 13674 21268 13720
rect 21068 13640 21268 13674
rect 21516 13720 21716 13737
rect 21516 13674 21552 13720
rect 21692 13674 21716 13720
rect 21516 13640 21716 13674
rect 21964 13720 22164 13737
rect 21964 13674 22000 13720
rect 22140 13674 22164 13720
rect 21964 13640 22164 13674
rect 1692 13352 1892 13396
rect 2140 13352 2340 13396
rect 2588 13352 2788 13396
rect 3036 13352 3236 13396
rect 3484 13352 3684 13396
rect 3932 13352 4132 13396
rect 4380 13352 4580 13396
rect 4828 13352 5028 13396
rect 5276 13352 5476 13396
rect 5724 13352 5924 13396
rect 6172 13352 6372 13396
rect 6620 13352 6820 13396
rect 7068 13352 7268 13396
rect 7516 13352 7716 13396
rect 7964 13352 8164 13396
rect 8412 13352 8612 13396
rect 8860 13352 9060 13396
rect 9644 13352 9844 13396
rect 10092 13352 10292 13396
rect 10540 13352 10740 13396
rect 10988 13352 11188 13396
rect 11436 13352 11636 13396
rect 11884 13352 12084 13396
rect 12332 13352 12532 13396
rect 12780 13352 12980 13396
rect 13228 13352 13428 13396
rect 13676 13352 13876 13396
rect 14124 13352 14324 13396
rect 14572 13352 14772 13396
rect 15020 13352 15220 13396
rect 15468 13352 15668 13396
rect 16160 13352 16260 13396
rect 16832 13352 16932 13396
rect 17728 13352 17828 13396
rect 18400 13352 18500 13396
rect 18828 13352 19028 13396
rect 19276 13352 19476 13396
rect 19724 13352 19924 13396
rect 20172 13352 20372 13396
rect 20620 13352 20820 13396
rect 21068 13352 21268 13396
rect 21516 13352 21716 13396
rect 21964 13352 22164 13396
rect 1692 13260 1892 13304
rect 2140 13260 2340 13304
rect 2588 13260 2788 13304
rect 3036 13260 3236 13304
rect 3484 13260 3684 13304
rect 3932 13260 4132 13304
rect 4380 13260 4580 13304
rect 4828 13260 5028 13304
rect 5612 13260 5812 13304
rect 6060 13260 6260 13304
rect 6508 13260 6708 13304
rect 6956 13260 7156 13304
rect 7404 13260 7604 13304
rect 7852 13260 8052 13304
rect 8300 13260 8500 13304
rect 8748 13260 8948 13304
rect 9196 13260 9396 13304
rect 9644 13260 9844 13304
rect 10092 13260 10292 13304
rect 10540 13260 10740 13304
rect 10988 13260 11188 13304
rect 11436 13260 11636 13304
rect 11884 13260 12084 13304
rect 12332 13260 12532 13304
rect 12780 13260 12980 13304
rect 13564 13260 13764 13304
rect 14012 13260 14212 13304
rect 14816 13260 14916 13304
rect 15488 13260 15588 13304
rect 16160 13260 16260 13304
rect 16832 13260 16932 13304
rect 17504 13260 17604 13304
rect 18176 13260 18276 13304
rect 18848 13260 18948 13304
rect 19520 13260 19620 13304
rect 19948 13260 20148 13304
rect 20396 13260 20596 13304
rect 20844 13260 21044 13304
rect 21516 13260 21716 13304
rect 21964 13260 22164 13304
rect 1692 12982 1892 13016
rect 1692 12936 1728 12982
rect 1868 12936 1892 12982
rect 1692 12919 1892 12936
rect 2140 12982 2340 13016
rect 2140 12936 2176 12982
rect 2316 12936 2340 12982
rect 2140 12919 2340 12936
rect 2588 12982 2788 13016
rect 2588 12936 2624 12982
rect 2764 12936 2788 12982
rect 2588 12919 2788 12936
rect 3036 12982 3236 13016
rect 3036 12936 3072 12982
rect 3212 12936 3236 12982
rect 3036 12919 3236 12936
rect 3484 12982 3684 13016
rect 3484 12936 3520 12982
rect 3660 12936 3684 12982
rect 3484 12919 3684 12936
rect 3932 12982 4132 13016
rect 3932 12936 3968 12982
rect 4108 12936 4132 12982
rect 3932 12919 4132 12936
rect 4380 12982 4580 13016
rect 4380 12936 4416 12982
rect 4556 12936 4580 12982
rect 4380 12919 4580 12936
rect 4828 12982 5028 13016
rect 4828 12936 4864 12982
rect 5004 12936 5028 12982
rect 4828 12919 5028 12936
rect 5612 12982 5812 13016
rect 5612 12936 5648 12982
rect 5788 12936 5812 12982
rect 5612 12919 5812 12936
rect 6060 12982 6260 13016
rect 6060 12936 6096 12982
rect 6236 12936 6260 12982
rect 6060 12919 6260 12936
rect 6508 12982 6708 13016
rect 6508 12936 6544 12982
rect 6684 12936 6708 12982
rect 6508 12919 6708 12936
rect 6956 12982 7156 13016
rect 6956 12936 6992 12982
rect 7132 12936 7156 12982
rect 6956 12919 7156 12936
rect 7404 12982 7604 13016
rect 7404 12936 7440 12982
rect 7580 12936 7604 12982
rect 7404 12919 7604 12936
rect 7852 12982 8052 13016
rect 7852 12936 7888 12982
rect 8028 12936 8052 12982
rect 7852 12919 8052 12936
rect 8300 12982 8500 13016
rect 8300 12936 8336 12982
rect 8476 12936 8500 12982
rect 8300 12919 8500 12936
rect 8748 12982 8948 13016
rect 8748 12936 8784 12982
rect 8924 12936 8948 12982
rect 8748 12919 8948 12936
rect 9196 12982 9396 13016
rect 9196 12936 9232 12982
rect 9372 12936 9396 12982
rect 9196 12919 9396 12936
rect 9644 12982 9844 13016
rect 9644 12936 9680 12982
rect 9820 12936 9844 12982
rect 9644 12919 9844 12936
rect 10092 12982 10292 13016
rect 10092 12936 10128 12982
rect 10268 12936 10292 12982
rect 10092 12919 10292 12936
rect 10540 12982 10740 13016
rect 10540 12936 10576 12982
rect 10716 12936 10740 12982
rect 10540 12919 10740 12936
rect 10988 12982 11188 13016
rect 10988 12936 11024 12982
rect 11164 12936 11188 12982
rect 10988 12919 11188 12936
rect 11436 12982 11636 13016
rect 11436 12936 11472 12982
rect 11612 12936 11636 12982
rect 11436 12919 11636 12936
rect 11884 12982 12084 13016
rect 11884 12936 11920 12982
rect 12060 12936 12084 12982
rect 11884 12919 12084 12936
rect 12332 12982 12532 13016
rect 12332 12936 12368 12982
rect 12508 12936 12532 12982
rect 12332 12919 12532 12936
rect 12780 12982 12980 13016
rect 12780 12936 12816 12982
rect 12956 12936 12980 12982
rect 12780 12919 12980 12936
rect 13564 12982 13764 13016
rect 13564 12936 13600 12982
rect 13740 12936 13764 12982
rect 13564 12919 13764 12936
rect 14012 12982 14212 13016
rect 14012 12936 14048 12982
rect 14188 12936 14212 12982
rect 14012 12919 14212 12936
rect 14816 12967 14916 13016
rect 14816 12930 14829 12967
rect 1692 12855 1892 12868
rect 1692 12809 1720 12855
rect 1860 12809 1892 12855
rect 1692 12776 1892 12809
rect 2140 12855 2340 12868
rect 2140 12809 2168 12855
rect 2308 12809 2340 12855
rect 2140 12776 2340 12809
rect 2588 12855 2788 12868
rect 2588 12809 2616 12855
rect 2756 12809 2788 12855
rect 2588 12776 2788 12809
rect 3036 12855 3236 12868
rect 3036 12809 3064 12855
rect 3204 12809 3236 12855
rect 3036 12776 3236 12809
rect 3484 12855 3684 12868
rect 3484 12809 3512 12855
rect 3652 12809 3684 12855
rect 3484 12776 3684 12809
rect 3932 12855 4132 12868
rect 3932 12809 3960 12855
rect 4100 12809 4132 12855
rect 3932 12776 4132 12809
rect 4380 12855 4580 12868
rect 4380 12809 4408 12855
rect 4548 12809 4580 12855
rect 4380 12776 4580 12809
rect 4828 12855 5028 12868
rect 4828 12809 4856 12855
rect 4996 12809 5028 12855
rect 4828 12776 5028 12809
rect 5612 12855 5812 12868
rect 5612 12809 5640 12855
rect 5780 12809 5812 12855
rect 5612 12776 5812 12809
rect 6060 12855 6260 12868
rect 6060 12809 6088 12855
rect 6228 12809 6260 12855
rect 6060 12776 6260 12809
rect 6508 12855 6708 12868
rect 6508 12809 6536 12855
rect 6676 12809 6708 12855
rect 6508 12776 6708 12809
rect 6956 12855 7156 12868
rect 6956 12809 6984 12855
rect 7124 12809 7156 12855
rect 6956 12776 7156 12809
rect 7404 12855 7604 12868
rect 7404 12809 7432 12855
rect 7572 12809 7604 12855
rect 7404 12776 7604 12809
rect 7852 12855 8052 12868
rect 7852 12809 7880 12855
rect 8020 12809 8052 12855
rect 7852 12776 8052 12809
rect 8300 12855 8500 12868
rect 8300 12809 8328 12855
rect 8468 12809 8500 12855
rect 8300 12776 8500 12809
rect 8748 12855 8948 12868
rect 8748 12809 8776 12855
rect 8916 12809 8948 12855
rect 8748 12776 8948 12809
rect 9196 12855 9396 12868
rect 9196 12809 9224 12855
rect 9364 12809 9396 12855
rect 9196 12776 9396 12809
rect 9644 12855 9844 12868
rect 9644 12809 9672 12855
rect 9812 12809 9844 12855
rect 9644 12776 9844 12809
rect 10092 12855 10292 12868
rect 10092 12809 10120 12855
rect 10260 12809 10292 12855
rect 10092 12776 10292 12809
rect 10540 12855 10740 12868
rect 10540 12809 10568 12855
rect 10708 12809 10740 12855
rect 10540 12776 10740 12809
rect 10988 12855 11188 12868
rect 10988 12809 11016 12855
rect 11156 12809 11188 12855
rect 10988 12776 11188 12809
rect 11436 12855 11636 12868
rect 11436 12809 11464 12855
rect 11604 12809 11636 12855
rect 11436 12776 11636 12809
rect 11884 12855 12084 12868
rect 11884 12809 11912 12855
rect 12052 12809 12084 12855
rect 11884 12776 12084 12809
rect 12332 12855 12532 12868
rect 12332 12809 12360 12855
rect 12500 12809 12532 12855
rect 12332 12776 12532 12809
rect 12780 12855 12980 12868
rect 12780 12809 12808 12855
rect 12948 12809 12980 12855
rect 12780 12776 12980 12809
rect 13564 12855 13764 12868
rect 13564 12809 13592 12855
rect 13732 12809 13764 12855
rect 1692 12568 1892 12612
rect 2140 12568 2340 12612
rect 2588 12568 2788 12612
rect 3036 12568 3236 12612
rect 3484 12568 3684 12612
rect 3932 12568 4132 12612
rect 4380 12568 4580 12612
rect 4828 12568 5028 12612
rect 13564 12776 13764 12809
rect 14012 12855 14212 12868
rect 14012 12809 14040 12855
rect 14180 12809 14212 12855
rect 14012 12776 14212 12809
rect 14796 12827 14829 12930
rect 14875 12827 14916 12967
rect 15488 12967 15588 13016
rect 15488 12930 15501 12967
rect 14796 12776 14916 12827
rect 15468 12827 15501 12930
rect 15547 12827 15588 12967
rect 16160 12967 16260 13016
rect 16160 12930 16173 12967
rect 15468 12776 15588 12827
rect 16140 12827 16173 12930
rect 16219 12827 16260 12967
rect 16832 12967 16932 13016
rect 16832 12930 16845 12967
rect 16140 12776 16260 12827
rect 16812 12827 16845 12930
rect 16891 12827 16932 12967
rect 17504 12967 17604 13016
rect 17504 12930 17517 12967
rect 16812 12776 16932 12827
rect 17484 12827 17517 12930
rect 17563 12827 17604 12967
rect 18176 12967 18276 13016
rect 18176 12930 18189 12967
rect 17484 12776 17604 12827
rect 18156 12827 18189 12930
rect 18235 12827 18276 12967
rect 18848 12967 18948 13016
rect 18848 12930 18861 12967
rect 18156 12776 18276 12827
rect 18828 12827 18861 12930
rect 18907 12827 18948 12967
rect 19520 12967 19620 13016
rect 19520 12930 19533 12967
rect 18828 12776 18948 12827
rect 19500 12827 19533 12930
rect 19579 12827 19620 12967
rect 19948 12982 20148 13016
rect 19948 12936 19984 12982
rect 20124 12936 20148 12982
rect 19948 12919 20148 12936
rect 20396 12982 20596 13016
rect 20396 12936 20432 12982
rect 20572 12936 20596 12982
rect 20396 12919 20596 12936
rect 20844 12982 21044 13016
rect 20844 12936 20880 12982
rect 21020 12936 21044 12982
rect 20844 12919 21044 12936
rect 21516 12982 21716 13016
rect 21516 12936 21552 12982
rect 21692 12936 21716 12982
rect 21516 12919 21716 12936
rect 21964 12982 22164 13016
rect 21964 12936 22000 12982
rect 22140 12936 22164 12982
rect 21964 12919 22164 12936
rect 19500 12776 19620 12827
rect 19948 12855 20148 12868
rect 19948 12809 19976 12855
rect 20116 12809 20148 12855
rect 19948 12776 20148 12809
rect 20396 12855 20596 12868
rect 20396 12809 20424 12855
rect 20564 12809 20596 12855
rect 20396 12776 20596 12809
rect 20844 12855 21044 12868
rect 20844 12809 20872 12855
rect 21012 12809 21044 12855
rect 20844 12776 21044 12809
rect 21516 12855 21716 12868
rect 21516 12809 21544 12855
rect 21684 12809 21716 12855
rect 5612 12568 5812 12612
rect 6060 12568 6260 12612
rect 6508 12568 6708 12612
rect 6956 12568 7156 12612
rect 7404 12568 7604 12612
rect 7852 12568 8052 12612
rect 8300 12568 8500 12612
rect 8748 12568 8948 12612
rect 9196 12568 9396 12612
rect 9644 12568 9844 12612
rect 10092 12568 10292 12612
rect 10540 12568 10740 12612
rect 10988 12568 11188 12612
rect 11436 12568 11636 12612
rect 11884 12568 12084 12612
rect 12332 12568 12532 12612
rect 12780 12568 12980 12612
rect 21516 12776 21716 12809
rect 21964 12855 22164 12868
rect 21964 12809 21992 12855
rect 22132 12809 22164 12855
rect 21964 12776 22164 12809
rect 13564 12568 13764 12612
rect 14012 12568 14212 12612
rect 14796 12568 14916 12612
rect 15468 12568 15588 12612
rect 16140 12568 16260 12612
rect 16812 12568 16932 12612
rect 17484 12568 17604 12612
rect 18156 12568 18276 12612
rect 18828 12568 18948 12612
rect 19500 12568 19620 12612
rect 19948 12568 20148 12612
rect 20396 12568 20596 12612
rect 20844 12568 21044 12612
rect 21516 12568 21716 12612
rect 21964 12568 22164 12612
rect 1692 12476 1892 12520
rect 2140 12476 2340 12520
rect 2588 12476 2788 12520
rect 3036 12476 3236 12520
rect 3484 12476 3684 12520
rect 3932 12476 4132 12520
rect 4380 12476 4580 12520
rect 4828 12476 5028 12520
rect 5276 12476 5476 12520
rect 5724 12476 5924 12520
rect 6172 12476 6372 12520
rect 6620 12476 6820 12520
rect 7068 12476 7268 12520
rect 7516 12476 7716 12520
rect 7964 12476 8164 12520
rect 8412 12476 8612 12520
rect 8860 12476 9060 12520
rect 9644 12476 9844 12520
rect 10092 12476 10292 12520
rect 10540 12476 10740 12520
rect 10988 12476 11188 12520
rect 11436 12476 11636 12520
rect 11884 12476 12084 12520
rect 12332 12476 12532 12520
rect 12780 12476 12980 12520
rect 13228 12476 13428 12520
rect 13676 12476 13876 12520
rect 14124 12476 14244 12520
rect 14796 12476 14916 12520
rect 15468 12476 15588 12520
rect 16140 12476 16260 12520
rect 16812 12476 16932 12520
rect 1692 12279 1892 12312
rect 1692 12233 1720 12279
rect 1860 12233 1892 12279
rect 1692 12220 1892 12233
rect 2140 12279 2340 12312
rect 2140 12233 2168 12279
rect 2308 12233 2340 12279
rect 2140 12220 2340 12233
rect 2588 12279 2788 12312
rect 2588 12233 2616 12279
rect 2756 12233 2788 12279
rect 2588 12220 2788 12233
rect 3036 12279 3236 12312
rect 3036 12233 3064 12279
rect 3204 12233 3236 12279
rect 3036 12220 3236 12233
rect 3484 12279 3684 12312
rect 3484 12233 3512 12279
rect 3652 12233 3684 12279
rect 3484 12220 3684 12233
rect 3932 12279 4132 12312
rect 3932 12233 3960 12279
rect 4100 12233 4132 12279
rect 3932 12220 4132 12233
rect 4380 12279 4580 12312
rect 4380 12233 4408 12279
rect 4548 12233 4580 12279
rect 4380 12220 4580 12233
rect 4828 12279 5028 12312
rect 4828 12233 4856 12279
rect 4996 12233 5028 12279
rect 4828 12220 5028 12233
rect 5276 12279 5476 12312
rect 5276 12233 5304 12279
rect 5444 12233 5476 12279
rect 5276 12220 5476 12233
rect 5724 12279 5924 12312
rect 5724 12233 5752 12279
rect 5892 12233 5924 12279
rect 5724 12220 5924 12233
rect 6172 12279 6372 12312
rect 6172 12233 6200 12279
rect 6340 12233 6372 12279
rect 6172 12220 6372 12233
rect 6620 12279 6820 12312
rect 6620 12233 6648 12279
rect 6788 12233 6820 12279
rect 6620 12220 6820 12233
rect 7068 12279 7268 12312
rect 7068 12233 7096 12279
rect 7236 12233 7268 12279
rect 7068 12220 7268 12233
rect 7516 12279 7716 12312
rect 7516 12233 7544 12279
rect 7684 12233 7716 12279
rect 7516 12220 7716 12233
rect 7964 12279 8164 12312
rect 7964 12233 7992 12279
rect 8132 12233 8164 12279
rect 7964 12220 8164 12233
rect 8412 12279 8612 12312
rect 8412 12233 8440 12279
rect 8580 12233 8612 12279
rect 8412 12220 8612 12233
rect 8860 12279 9060 12312
rect 17708 12476 17828 12520
rect 18380 12476 18500 12520
rect 19052 12476 19172 12520
rect 19724 12476 19844 12520
rect 20396 12476 20516 12520
rect 20844 12476 21044 12520
rect 21292 12476 21492 12520
rect 21740 12476 21940 12520
rect 8860 12233 8888 12279
rect 9028 12233 9060 12279
rect 8860 12220 9060 12233
rect 9644 12279 9844 12312
rect 9644 12233 9672 12279
rect 9812 12233 9844 12279
rect 9644 12220 9844 12233
rect 10092 12279 10292 12312
rect 10092 12233 10120 12279
rect 10260 12233 10292 12279
rect 10092 12220 10292 12233
rect 10540 12279 10740 12312
rect 10540 12233 10568 12279
rect 10708 12233 10740 12279
rect 10540 12220 10740 12233
rect 10988 12279 11188 12312
rect 10988 12233 11016 12279
rect 11156 12233 11188 12279
rect 10988 12220 11188 12233
rect 11436 12279 11636 12312
rect 11436 12233 11464 12279
rect 11604 12233 11636 12279
rect 11436 12220 11636 12233
rect 11884 12279 12084 12312
rect 11884 12233 11912 12279
rect 12052 12233 12084 12279
rect 11884 12220 12084 12233
rect 12332 12279 12532 12312
rect 12332 12233 12360 12279
rect 12500 12233 12532 12279
rect 12332 12220 12532 12233
rect 12780 12279 12980 12312
rect 12780 12233 12808 12279
rect 12948 12233 12980 12279
rect 12780 12220 12980 12233
rect 13228 12279 13428 12312
rect 13228 12233 13256 12279
rect 13396 12233 13428 12279
rect 13228 12220 13428 12233
rect 13676 12279 13876 12312
rect 13676 12233 13704 12279
rect 13844 12233 13876 12279
rect 13676 12220 13876 12233
rect 14124 12261 14244 12312
rect 1692 12152 1892 12169
rect 1692 12106 1728 12152
rect 1868 12106 1892 12152
rect 1692 12072 1892 12106
rect 2140 12152 2340 12169
rect 2140 12106 2176 12152
rect 2316 12106 2340 12152
rect 2140 12072 2340 12106
rect 2588 12152 2788 12169
rect 2588 12106 2624 12152
rect 2764 12106 2788 12152
rect 2588 12072 2788 12106
rect 3036 12152 3236 12169
rect 3036 12106 3072 12152
rect 3212 12106 3236 12152
rect 3036 12072 3236 12106
rect 3484 12152 3684 12169
rect 3484 12106 3520 12152
rect 3660 12106 3684 12152
rect 3484 12072 3684 12106
rect 3932 12152 4132 12169
rect 3932 12106 3968 12152
rect 4108 12106 4132 12152
rect 3932 12072 4132 12106
rect 4380 12152 4580 12169
rect 4380 12106 4416 12152
rect 4556 12106 4580 12152
rect 4380 12072 4580 12106
rect 4828 12152 5028 12169
rect 4828 12106 4864 12152
rect 5004 12106 5028 12152
rect 4828 12072 5028 12106
rect 5276 12152 5476 12169
rect 5276 12106 5312 12152
rect 5452 12106 5476 12152
rect 5276 12072 5476 12106
rect 5724 12152 5924 12169
rect 5724 12106 5760 12152
rect 5900 12106 5924 12152
rect 5724 12072 5924 12106
rect 6172 12152 6372 12169
rect 6172 12106 6208 12152
rect 6348 12106 6372 12152
rect 6172 12072 6372 12106
rect 6620 12152 6820 12169
rect 6620 12106 6656 12152
rect 6796 12106 6820 12152
rect 6620 12072 6820 12106
rect 7068 12152 7268 12169
rect 7068 12106 7104 12152
rect 7244 12106 7268 12152
rect 7068 12072 7268 12106
rect 7516 12152 7716 12169
rect 7516 12106 7552 12152
rect 7692 12106 7716 12152
rect 7516 12072 7716 12106
rect 7964 12152 8164 12169
rect 7964 12106 8000 12152
rect 8140 12106 8164 12152
rect 7964 12072 8164 12106
rect 8412 12152 8612 12169
rect 8412 12106 8448 12152
rect 8588 12106 8612 12152
rect 8412 12072 8612 12106
rect 8860 12152 9060 12169
rect 8860 12106 8896 12152
rect 9036 12106 9060 12152
rect 8860 12072 9060 12106
rect 9644 12152 9844 12169
rect 9644 12106 9680 12152
rect 9820 12106 9844 12152
rect 9644 12072 9844 12106
rect 10092 12152 10292 12169
rect 10092 12106 10128 12152
rect 10268 12106 10292 12152
rect 10092 12072 10292 12106
rect 10540 12152 10740 12169
rect 10540 12106 10576 12152
rect 10716 12106 10740 12152
rect 10540 12072 10740 12106
rect 10988 12152 11188 12169
rect 10988 12106 11024 12152
rect 11164 12106 11188 12152
rect 10988 12072 11188 12106
rect 11436 12152 11636 12169
rect 11436 12106 11472 12152
rect 11612 12106 11636 12152
rect 11436 12072 11636 12106
rect 11884 12152 12084 12169
rect 11884 12106 11920 12152
rect 12060 12106 12084 12152
rect 11884 12072 12084 12106
rect 12332 12152 12532 12169
rect 12332 12106 12368 12152
rect 12508 12106 12532 12152
rect 12332 12072 12532 12106
rect 12780 12152 12980 12169
rect 12780 12106 12816 12152
rect 12956 12106 12980 12152
rect 12780 12072 12980 12106
rect 13228 12152 13428 12169
rect 13228 12106 13264 12152
rect 13404 12106 13428 12152
rect 13228 12072 13428 12106
rect 13676 12152 13876 12169
rect 14124 12158 14157 12261
rect 13676 12106 13712 12152
rect 13852 12106 13876 12152
rect 13676 12072 13876 12106
rect 14144 12121 14157 12158
rect 14203 12121 14244 12261
rect 14796 12261 14916 12312
rect 14796 12158 14829 12261
rect 14144 12072 14244 12121
rect 14816 12121 14829 12158
rect 14875 12121 14916 12261
rect 15468 12261 15588 12312
rect 15468 12158 15501 12261
rect 14816 12072 14916 12121
rect 15488 12121 15501 12158
rect 15547 12121 15588 12261
rect 16140 12261 16260 12312
rect 16140 12158 16173 12261
rect 15488 12072 15588 12121
rect 16160 12121 16173 12158
rect 16219 12121 16260 12261
rect 16812 12261 16932 12312
rect 16812 12158 16845 12261
rect 16160 12072 16260 12121
rect 16832 12121 16845 12158
rect 16891 12121 16932 12261
rect 17708 12261 17828 12312
rect 16832 12072 16932 12121
rect 17708 12158 17741 12261
rect 17728 12121 17741 12158
rect 17787 12121 17828 12261
rect 18380 12261 18500 12312
rect 18380 12158 18413 12261
rect 17728 12072 17828 12121
rect 18400 12121 18413 12158
rect 18459 12121 18500 12261
rect 19052 12261 19172 12312
rect 19052 12158 19085 12261
rect 18400 12072 18500 12121
rect 19072 12121 19085 12158
rect 19131 12121 19172 12261
rect 19724 12261 19844 12312
rect 19724 12158 19757 12261
rect 19072 12072 19172 12121
rect 19744 12121 19757 12158
rect 19803 12121 19844 12261
rect 20396 12261 20516 12312
rect 20396 12158 20429 12261
rect 19744 12072 19844 12121
rect 20416 12121 20429 12158
rect 20475 12121 20516 12261
rect 20844 12279 21044 12312
rect 20844 12233 20872 12279
rect 21012 12233 21044 12279
rect 20844 12220 21044 12233
rect 21292 12279 21492 12312
rect 21292 12233 21320 12279
rect 21460 12233 21492 12279
rect 21292 12220 21492 12233
rect 21740 12279 21940 12312
rect 21740 12233 21768 12279
rect 21908 12233 21940 12279
rect 21740 12220 21940 12233
rect 20416 12072 20516 12121
rect 20844 12152 21044 12169
rect 20844 12106 20880 12152
rect 21020 12106 21044 12152
rect 20844 12072 21044 12106
rect 21292 12152 21492 12169
rect 21292 12106 21328 12152
rect 21468 12106 21492 12152
rect 21292 12072 21492 12106
rect 21740 12152 21940 12169
rect 21740 12106 21776 12152
rect 21916 12106 21940 12152
rect 21740 12072 21940 12106
rect 1692 11784 1892 11828
rect 2140 11784 2340 11828
rect 2588 11784 2788 11828
rect 3036 11784 3236 11828
rect 3484 11784 3684 11828
rect 3932 11784 4132 11828
rect 4380 11784 4580 11828
rect 4828 11784 5028 11828
rect 5276 11784 5476 11828
rect 5724 11784 5924 11828
rect 6172 11784 6372 11828
rect 6620 11784 6820 11828
rect 7068 11784 7268 11828
rect 7516 11784 7716 11828
rect 7964 11784 8164 11828
rect 8412 11784 8612 11828
rect 8860 11784 9060 11828
rect 9644 11784 9844 11828
rect 10092 11784 10292 11828
rect 10540 11784 10740 11828
rect 10988 11784 11188 11828
rect 11436 11784 11636 11828
rect 11884 11784 12084 11828
rect 12332 11784 12532 11828
rect 12780 11784 12980 11828
rect 13228 11784 13428 11828
rect 13676 11784 13876 11828
rect 14144 11784 14244 11828
rect 14816 11784 14916 11828
rect 15488 11784 15588 11828
rect 16160 11784 16260 11828
rect 16832 11784 16932 11828
rect 17728 11784 17828 11828
rect 18400 11784 18500 11828
rect 19072 11784 19172 11828
rect 19744 11784 19844 11828
rect 20416 11784 20516 11828
rect 20844 11784 21044 11828
rect 21292 11784 21492 11828
rect 21740 11784 21940 11828
rect 1692 11692 1892 11736
rect 2140 11692 2340 11736
rect 2588 11692 2788 11736
rect 3036 11692 3236 11736
rect 3484 11692 3684 11736
rect 3932 11692 4132 11736
rect 4380 11692 4580 11736
rect 4828 11692 5028 11736
rect 5612 11692 5812 11736
rect 6140 11692 6240 11736
rect 6924 11692 7024 11736
rect 7596 11692 7696 11736
rect 8268 11692 8368 11736
rect 8636 11692 8836 11736
rect 9216 11692 9316 11736
rect 9888 11692 9988 11736
rect 10560 11692 10660 11736
rect 10988 11692 11188 11736
rect 11436 11692 11636 11736
rect 12128 11692 12228 11736
rect 12800 11692 12900 11736
rect 13696 11692 13796 11736
rect 14124 11692 14324 11736
rect 14816 11692 14916 11736
rect 15488 11692 15588 11736
rect 16160 11692 16260 11736
rect 16832 11692 16932 11736
rect 17504 11692 17604 11736
rect 18176 11692 18276 11736
rect 18848 11692 18948 11736
rect 19520 11692 19620 11736
rect 20192 11692 20292 11736
rect 20620 11692 20820 11736
rect 21516 11692 21716 11736
rect 21964 11692 22164 11736
rect 1692 11414 1892 11448
rect 1692 11368 1728 11414
rect 1868 11368 1892 11414
rect 1692 11351 1892 11368
rect 2140 11414 2340 11448
rect 2140 11368 2176 11414
rect 2316 11368 2340 11414
rect 2140 11351 2340 11368
rect 2588 11414 2788 11448
rect 2588 11368 2624 11414
rect 2764 11368 2788 11414
rect 2588 11351 2788 11368
rect 3036 11414 3236 11448
rect 3036 11368 3072 11414
rect 3212 11368 3236 11414
rect 3036 11351 3236 11368
rect 3484 11414 3684 11448
rect 3484 11368 3520 11414
rect 3660 11368 3684 11414
rect 3484 11351 3684 11368
rect 3932 11414 4132 11448
rect 3932 11368 3968 11414
rect 4108 11368 4132 11414
rect 3932 11351 4132 11368
rect 4380 11414 4580 11448
rect 4380 11368 4416 11414
rect 4556 11368 4580 11414
rect 4380 11351 4580 11368
rect 4828 11414 5028 11448
rect 4828 11368 4864 11414
rect 5004 11368 5028 11414
rect 4828 11351 5028 11368
rect 5612 11414 5812 11448
rect 5612 11368 5648 11414
rect 5788 11368 5812 11414
rect 5612 11351 5812 11368
rect 6140 11399 6240 11448
rect 1692 11287 1892 11300
rect 1692 11241 1720 11287
rect 1860 11241 1892 11287
rect 1692 11208 1892 11241
rect 2140 11287 2340 11300
rect 2140 11241 2168 11287
rect 2308 11241 2340 11287
rect 2140 11208 2340 11241
rect 2588 11287 2788 11300
rect 2588 11241 2616 11287
rect 2756 11241 2788 11287
rect 2588 11208 2788 11241
rect 3036 11287 3236 11300
rect 3036 11241 3064 11287
rect 3204 11241 3236 11287
rect 3036 11208 3236 11241
rect 3484 11287 3684 11300
rect 3484 11241 3512 11287
rect 3652 11241 3684 11287
rect 3484 11208 3684 11241
rect 3932 11287 4132 11300
rect 3932 11241 3960 11287
rect 4100 11241 4132 11287
rect 3932 11208 4132 11241
rect 4380 11287 4580 11300
rect 4380 11241 4408 11287
rect 4548 11241 4580 11287
rect 4380 11208 4580 11241
rect 4828 11287 5028 11300
rect 4828 11241 4856 11287
rect 4996 11241 5028 11287
rect 4828 11208 5028 11241
rect 5612 11287 5812 11300
rect 5612 11241 5640 11287
rect 5780 11241 5812 11287
rect 5612 11208 5812 11241
rect 6140 11259 6181 11399
rect 6227 11362 6240 11399
rect 6924 11399 7024 11448
rect 6227 11259 6260 11362
rect 6140 11208 6260 11259
rect 6924 11259 6965 11399
rect 7011 11362 7024 11399
rect 7596 11399 7696 11448
rect 7011 11259 7044 11362
rect 6924 11208 7044 11259
rect 7596 11259 7637 11399
rect 7683 11362 7696 11399
rect 8268 11399 8368 11448
rect 7683 11259 7716 11362
rect 7596 11208 7716 11259
rect 8268 11259 8309 11399
rect 8355 11362 8368 11399
rect 8636 11414 8836 11448
rect 8636 11368 8672 11414
rect 8812 11368 8836 11414
rect 8355 11259 8388 11362
rect 8636 11351 8836 11368
rect 9216 11399 9316 11448
rect 9216 11362 9229 11399
rect 8268 11208 8388 11259
rect 8636 11287 8836 11300
rect 8636 11241 8664 11287
rect 8804 11241 8836 11287
rect 8636 11208 8836 11241
rect 9196 11259 9229 11362
rect 9275 11259 9316 11399
rect 9888 11399 9988 11448
rect 9888 11362 9901 11399
rect 9196 11208 9316 11259
rect 9868 11259 9901 11362
rect 9947 11259 9988 11399
rect 10560 11399 10660 11448
rect 10560 11362 10573 11399
rect 9868 11208 9988 11259
rect 10540 11259 10573 11362
rect 10619 11259 10660 11399
rect 10988 11414 11188 11448
rect 10988 11368 11024 11414
rect 11164 11368 11188 11414
rect 10988 11351 11188 11368
rect 11436 11414 11636 11448
rect 11436 11368 11472 11414
rect 11612 11368 11636 11414
rect 11436 11351 11636 11368
rect 12128 11399 12228 11448
rect 12128 11362 12141 11399
rect 10540 11208 10660 11259
rect 10988 11287 11188 11300
rect 10988 11241 11016 11287
rect 11156 11241 11188 11287
rect 10988 11208 11188 11241
rect 11436 11287 11636 11300
rect 11436 11241 11464 11287
rect 11604 11241 11636 11287
rect 11436 11208 11636 11241
rect 12108 11259 12141 11362
rect 12187 11259 12228 11399
rect 12800 11399 12900 11448
rect 12800 11362 12813 11399
rect 12108 11208 12228 11259
rect 12780 11259 12813 11362
rect 12859 11259 12900 11399
rect 13696 11399 13796 11448
rect 13696 11362 13709 11399
rect 12780 11208 12900 11259
rect 13676 11259 13709 11362
rect 13755 11259 13796 11399
rect 14124 11414 14324 11448
rect 14124 11368 14160 11414
rect 14300 11368 14324 11414
rect 14124 11351 14324 11368
rect 14816 11399 14916 11448
rect 14816 11362 14829 11399
rect 1692 11000 1892 11044
rect 2140 11000 2340 11044
rect 2588 11000 2788 11044
rect 3036 11000 3236 11044
rect 3484 11000 3684 11044
rect 3932 11000 4132 11044
rect 4380 11000 4580 11044
rect 4828 11000 5028 11044
rect 13676 11208 13796 11259
rect 14124 11287 14324 11300
rect 14124 11241 14152 11287
rect 14292 11241 14324 11287
rect 14124 11208 14324 11241
rect 14796 11259 14829 11362
rect 14875 11259 14916 11399
rect 15488 11399 15588 11448
rect 15488 11362 15501 11399
rect 14796 11208 14916 11259
rect 15468 11259 15501 11362
rect 15547 11259 15588 11399
rect 16160 11399 16260 11448
rect 16160 11362 16173 11399
rect 15468 11208 15588 11259
rect 16140 11259 16173 11362
rect 16219 11259 16260 11399
rect 16832 11399 16932 11448
rect 16832 11362 16845 11399
rect 16140 11208 16260 11259
rect 16812 11259 16845 11362
rect 16891 11259 16932 11399
rect 17504 11399 17604 11448
rect 17504 11362 17517 11399
rect 16812 11208 16932 11259
rect 17484 11259 17517 11362
rect 17563 11259 17604 11399
rect 18176 11399 18276 11448
rect 18176 11362 18189 11399
rect 17484 11208 17604 11259
rect 18156 11259 18189 11362
rect 18235 11259 18276 11399
rect 18848 11399 18948 11448
rect 18848 11362 18861 11399
rect 18156 11208 18276 11259
rect 18828 11259 18861 11362
rect 18907 11259 18948 11399
rect 19520 11399 19620 11448
rect 19520 11362 19533 11399
rect 18828 11208 18948 11259
rect 19500 11259 19533 11362
rect 19579 11259 19620 11399
rect 20192 11399 20292 11448
rect 20192 11362 20205 11399
rect 19500 11208 19620 11259
rect 20172 11259 20205 11362
rect 20251 11259 20292 11399
rect 20620 11414 20820 11448
rect 20620 11368 20656 11414
rect 20796 11368 20820 11414
rect 20620 11351 20820 11368
rect 21516 11414 21716 11448
rect 21516 11368 21552 11414
rect 21692 11368 21716 11414
rect 21516 11351 21716 11368
rect 21964 11414 22164 11448
rect 21964 11368 22000 11414
rect 22140 11368 22164 11414
rect 21964 11351 22164 11368
rect 20172 11208 20292 11259
rect 20620 11287 20820 11300
rect 20620 11241 20648 11287
rect 20788 11241 20820 11287
rect 20620 11208 20820 11241
rect 21516 11287 21716 11300
rect 21516 11241 21544 11287
rect 21684 11241 21716 11287
rect 5612 11000 5812 11044
rect 6140 11000 6260 11044
rect 6924 11000 7044 11044
rect 7596 11000 7716 11044
rect 8268 11000 8388 11044
rect 8636 11000 8836 11044
rect 9196 11000 9316 11044
rect 9868 11000 9988 11044
rect 10540 11000 10660 11044
rect 10988 11000 11188 11044
rect 11436 11000 11636 11044
rect 12108 11000 12228 11044
rect 12780 11000 12900 11044
rect 21516 11208 21716 11241
rect 21964 11287 22164 11300
rect 21964 11241 21992 11287
rect 22132 11241 22164 11287
rect 21964 11208 22164 11241
rect 13676 11000 13796 11044
rect 14124 11000 14324 11044
rect 14796 11000 14916 11044
rect 15468 11000 15588 11044
rect 16140 11000 16260 11044
rect 16812 11000 16932 11044
rect 17484 11000 17604 11044
rect 18156 11000 18276 11044
rect 18828 11000 18948 11044
rect 19500 11000 19620 11044
rect 20172 11000 20292 11044
rect 20620 11000 20820 11044
rect 21516 11000 21716 11044
rect 21964 11000 22164 11044
rect 1692 10908 1892 10952
rect 2140 10908 2340 10952
rect 2588 10908 2788 10952
rect 3036 10908 3236 10952
rect 3484 10908 3684 10952
rect 3932 10908 4132 10952
rect 4380 10908 4580 10952
rect 4828 10908 5028 10952
rect 5388 10908 5508 10952
rect 6060 10908 6180 10952
rect 6732 10908 6852 10952
rect 7404 10908 7524 10952
rect 8076 10908 8196 10952
rect 8860 10908 8980 10952
rect 9868 10908 9988 10952
rect 10540 10908 10660 10952
rect 11212 10908 11332 10952
rect 11996 10908 12116 10952
rect 12668 10908 12788 10952
rect 13340 10908 13460 10952
rect 14012 10908 14132 10952
rect 14684 10908 14804 10952
rect 15356 10908 15476 10952
rect 16028 10908 16148 10952
rect 16700 10908 16820 10952
rect 1692 10711 1892 10744
rect 1692 10665 1720 10711
rect 1860 10665 1892 10711
rect 1692 10652 1892 10665
rect 2140 10711 2340 10744
rect 2140 10665 2168 10711
rect 2308 10665 2340 10711
rect 2140 10652 2340 10665
rect 2588 10711 2788 10744
rect 2588 10665 2616 10711
rect 2756 10665 2788 10711
rect 2588 10652 2788 10665
rect 3036 10711 3236 10744
rect 3036 10665 3064 10711
rect 3204 10665 3236 10711
rect 3036 10652 3236 10665
rect 3484 10711 3684 10744
rect 3484 10665 3512 10711
rect 3652 10665 3684 10711
rect 3484 10652 3684 10665
rect 3932 10711 4132 10744
rect 3932 10665 3960 10711
rect 4100 10665 4132 10711
rect 3932 10652 4132 10665
rect 4380 10711 4580 10744
rect 4380 10665 4408 10711
rect 4548 10665 4580 10711
rect 4380 10652 4580 10665
rect 4828 10711 5028 10744
rect 4828 10665 4856 10711
rect 4996 10665 5028 10711
rect 4828 10652 5028 10665
rect 5388 10693 5508 10744
rect 1692 10584 1892 10601
rect 1692 10538 1728 10584
rect 1868 10538 1892 10584
rect 1692 10504 1892 10538
rect 2140 10584 2340 10601
rect 2140 10538 2176 10584
rect 2316 10538 2340 10584
rect 2140 10504 2340 10538
rect 2588 10584 2788 10601
rect 2588 10538 2624 10584
rect 2764 10538 2788 10584
rect 2588 10504 2788 10538
rect 3036 10584 3236 10601
rect 3036 10538 3072 10584
rect 3212 10538 3236 10584
rect 3036 10504 3236 10538
rect 3484 10584 3684 10601
rect 3484 10538 3520 10584
rect 3660 10538 3684 10584
rect 3484 10504 3684 10538
rect 3932 10584 4132 10601
rect 3932 10538 3968 10584
rect 4108 10538 4132 10584
rect 3932 10504 4132 10538
rect 4380 10584 4580 10601
rect 4380 10538 4416 10584
rect 4556 10538 4580 10584
rect 4380 10504 4580 10538
rect 4828 10584 5028 10601
rect 5388 10590 5421 10693
rect 4828 10538 4864 10584
rect 5004 10538 5028 10584
rect 4828 10504 5028 10538
rect 5408 10553 5421 10590
rect 5467 10553 5508 10693
rect 6060 10693 6180 10744
rect 6060 10590 6093 10693
rect 5408 10504 5508 10553
rect 6080 10553 6093 10590
rect 6139 10553 6180 10693
rect 6732 10693 6852 10744
rect 6732 10590 6765 10693
rect 6080 10504 6180 10553
rect 6752 10553 6765 10590
rect 6811 10553 6852 10693
rect 7404 10693 7524 10744
rect 7404 10590 7437 10693
rect 6752 10504 6852 10553
rect 7424 10553 7437 10590
rect 7483 10553 7524 10693
rect 8076 10693 8196 10744
rect 8076 10590 8109 10693
rect 7424 10504 7524 10553
rect 8096 10553 8109 10590
rect 8155 10553 8196 10693
rect 8860 10693 8980 10744
rect 17708 10908 17828 10952
rect 18380 10908 18500 10952
rect 19052 10908 19172 10952
rect 19724 10908 19844 10952
rect 20396 10908 20516 10952
rect 21068 10908 21188 10952
rect 21740 10908 21860 10952
rect 8860 10590 8893 10693
rect 8096 10504 8196 10553
rect 8880 10553 8893 10590
rect 8939 10553 8980 10693
rect 9868 10693 9988 10744
rect 8880 10504 8980 10553
rect 9868 10590 9901 10693
rect 9888 10553 9901 10590
rect 9947 10553 9988 10693
rect 10540 10693 10660 10744
rect 10540 10590 10573 10693
rect 9888 10504 9988 10553
rect 10560 10553 10573 10590
rect 10619 10553 10660 10693
rect 11212 10693 11332 10744
rect 11212 10590 11245 10693
rect 10560 10504 10660 10553
rect 11232 10553 11245 10590
rect 11291 10553 11332 10693
rect 11996 10693 12116 10744
rect 11996 10590 12029 10693
rect 11232 10504 11332 10553
rect 12016 10553 12029 10590
rect 12075 10553 12116 10693
rect 12668 10693 12788 10744
rect 12668 10590 12701 10693
rect 12016 10504 12116 10553
rect 12688 10553 12701 10590
rect 12747 10553 12788 10693
rect 13340 10693 13460 10744
rect 13340 10590 13373 10693
rect 12688 10504 12788 10553
rect 13360 10553 13373 10590
rect 13419 10553 13460 10693
rect 14012 10693 14132 10744
rect 14012 10590 14045 10693
rect 13360 10504 13460 10553
rect 14032 10553 14045 10590
rect 14091 10553 14132 10693
rect 14684 10693 14804 10744
rect 14684 10590 14717 10693
rect 14032 10504 14132 10553
rect 14704 10553 14717 10590
rect 14763 10553 14804 10693
rect 15356 10693 15476 10744
rect 15356 10590 15389 10693
rect 14704 10504 14804 10553
rect 15376 10553 15389 10590
rect 15435 10553 15476 10693
rect 16028 10693 16148 10744
rect 16028 10590 16061 10693
rect 15376 10504 15476 10553
rect 16048 10553 16061 10590
rect 16107 10553 16148 10693
rect 16700 10693 16820 10744
rect 16700 10590 16733 10693
rect 16048 10504 16148 10553
rect 16720 10553 16733 10590
rect 16779 10553 16820 10693
rect 17708 10693 17828 10744
rect 16720 10504 16820 10553
rect 17708 10590 17741 10693
rect 17728 10553 17741 10590
rect 17787 10553 17828 10693
rect 18380 10693 18500 10744
rect 18380 10590 18413 10693
rect 17728 10504 17828 10553
rect 18400 10553 18413 10590
rect 18459 10553 18500 10693
rect 19052 10693 19172 10744
rect 19052 10590 19085 10693
rect 18400 10504 18500 10553
rect 19072 10553 19085 10590
rect 19131 10553 19172 10693
rect 19724 10693 19844 10744
rect 19724 10590 19757 10693
rect 19072 10504 19172 10553
rect 19744 10553 19757 10590
rect 19803 10553 19844 10693
rect 20396 10693 20516 10744
rect 20396 10590 20429 10693
rect 19744 10504 19844 10553
rect 20416 10553 20429 10590
rect 20475 10553 20516 10693
rect 21068 10693 21188 10744
rect 21068 10590 21101 10693
rect 20416 10504 20516 10553
rect 21088 10553 21101 10590
rect 21147 10553 21188 10693
rect 21740 10693 21860 10744
rect 21740 10590 21773 10693
rect 21088 10504 21188 10553
rect 21760 10553 21773 10590
rect 21819 10553 21860 10693
rect 21760 10504 21860 10553
rect 1692 10216 1892 10260
rect 2140 10216 2340 10260
rect 2588 10216 2788 10260
rect 3036 10216 3236 10260
rect 3484 10216 3684 10260
rect 3932 10216 4132 10260
rect 4380 10216 4580 10260
rect 4828 10216 5028 10260
rect 5408 10216 5508 10260
rect 6080 10216 6180 10260
rect 6752 10216 6852 10260
rect 7424 10216 7524 10260
rect 8096 10216 8196 10260
rect 8880 10216 8980 10260
rect 9888 10216 9988 10260
rect 10560 10216 10660 10260
rect 11232 10216 11332 10260
rect 12016 10216 12116 10260
rect 12688 10216 12788 10260
rect 13360 10216 13460 10260
rect 14032 10216 14132 10260
rect 14704 10216 14804 10260
rect 15376 10216 15476 10260
rect 16048 10216 16148 10260
rect 16720 10216 16820 10260
rect 17728 10216 17828 10260
rect 18400 10216 18500 10260
rect 19072 10216 19172 10260
rect 19744 10216 19844 10260
rect 20416 10216 20516 10260
rect 21088 10216 21188 10260
rect 21760 10216 21860 10260
rect 1692 10124 1892 10168
rect 2140 10124 2340 10168
rect 2588 10124 2788 10168
rect 3036 10124 3236 10168
rect 3484 10124 3684 10168
rect 4176 10124 4276 10168
rect 4848 10124 4948 10168
rect 5856 10124 5956 10168
rect 6528 10124 6628 10168
rect 7200 10124 7300 10168
rect 7872 10124 7972 10168
rect 8544 10124 8644 10168
rect 9216 10124 9316 10168
rect 9888 10124 9988 10168
rect 10560 10124 10660 10168
rect 10988 10124 11188 10168
rect 11456 10124 11556 10168
rect 12128 10124 12228 10168
rect 12800 10124 12900 10168
rect 13696 10124 13796 10168
rect 14368 10124 14468 10168
rect 15040 10124 15140 10168
rect 15712 10124 15812 10168
rect 16384 10124 16484 10168
rect 17056 10124 17156 10168
rect 17788 10124 17888 10168
rect 18400 10124 18500 10168
rect 19072 10124 19172 10168
rect 19744 10124 19844 10168
rect 20416 10124 20516 10168
rect 20844 10124 21044 10168
rect 21648 10124 21748 10168
rect 22076 10124 22276 10168
rect 1692 9846 1892 9880
rect 1692 9800 1728 9846
rect 1868 9800 1892 9846
rect 1692 9783 1892 9800
rect 2140 9846 2340 9880
rect 2140 9800 2176 9846
rect 2316 9800 2340 9846
rect 2140 9783 2340 9800
rect 2588 9846 2788 9880
rect 2588 9800 2624 9846
rect 2764 9800 2788 9846
rect 2588 9783 2788 9800
rect 3036 9846 3236 9880
rect 3036 9800 3072 9846
rect 3212 9800 3236 9846
rect 3036 9783 3236 9800
rect 3484 9846 3684 9880
rect 3484 9800 3520 9846
rect 3660 9800 3684 9846
rect 3484 9783 3684 9800
rect 4176 9831 4276 9880
rect 4176 9794 4189 9831
rect 1692 9719 1892 9732
rect 1692 9673 1720 9719
rect 1860 9673 1892 9719
rect 1692 9640 1892 9673
rect 2140 9719 2340 9732
rect 2140 9673 2168 9719
rect 2308 9673 2340 9719
rect 2140 9640 2340 9673
rect 2588 9719 2788 9732
rect 2588 9673 2616 9719
rect 2756 9673 2788 9719
rect 2588 9640 2788 9673
rect 3036 9719 3236 9732
rect 3036 9673 3064 9719
rect 3204 9673 3236 9719
rect 3036 9640 3236 9673
rect 3484 9719 3684 9732
rect 3484 9673 3512 9719
rect 3652 9673 3684 9719
rect 3484 9640 3684 9673
rect 4156 9691 4189 9794
rect 4235 9691 4276 9831
rect 4848 9831 4948 9880
rect 4848 9794 4861 9831
rect 4156 9640 4276 9691
rect 4828 9691 4861 9794
rect 4907 9691 4948 9831
rect 5856 9831 5956 9880
rect 5856 9794 5869 9831
rect 4828 9640 4948 9691
rect 5836 9691 5869 9794
rect 5915 9691 5956 9831
rect 6528 9831 6628 9880
rect 6528 9794 6541 9831
rect 5836 9640 5956 9691
rect 6508 9691 6541 9794
rect 6587 9691 6628 9831
rect 7200 9831 7300 9880
rect 7200 9794 7213 9831
rect 6508 9640 6628 9691
rect 7180 9691 7213 9794
rect 7259 9691 7300 9831
rect 7872 9831 7972 9880
rect 7872 9794 7885 9831
rect 7180 9640 7300 9691
rect 7852 9691 7885 9794
rect 7931 9691 7972 9831
rect 8544 9831 8644 9880
rect 8544 9794 8557 9831
rect 7852 9640 7972 9691
rect 8524 9691 8557 9794
rect 8603 9691 8644 9831
rect 9216 9831 9316 9880
rect 9216 9794 9229 9831
rect 8524 9640 8644 9691
rect 9196 9691 9229 9794
rect 9275 9691 9316 9831
rect 9888 9831 9988 9880
rect 9888 9794 9901 9831
rect 9196 9640 9316 9691
rect 9868 9691 9901 9794
rect 9947 9691 9988 9831
rect 10560 9831 10660 9880
rect 10560 9794 10573 9831
rect 9868 9640 9988 9691
rect 10540 9691 10573 9794
rect 10619 9691 10660 9831
rect 10988 9846 11188 9880
rect 10988 9800 11024 9846
rect 11164 9800 11188 9846
rect 10988 9783 11188 9800
rect 11456 9831 11556 9880
rect 11456 9794 11469 9831
rect 10540 9640 10660 9691
rect 10988 9719 11188 9732
rect 10988 9673 11016 9719
rect 11156 9673 11188 9719
rect 10988 9640 11188 9673
rect 11436 9691 11469 9794
rect 11515 9691 11556 9831
rect 12128 9831 12228 9880
rect 12128 9794 12141 9831
rect 11436 9640 11556 9691
rect 12108 9691 12141 9794
rect 12187 9691 12228 9831
rect 12800 9831 12900 9880
rect 12800 9794 12813 9831
rect 12108 9640 12228 9691
rect 12780 9691 12813 9794
rect 12859 9691 12900 9831
rect 13696 9831 13796 9880
rect 13696 9794 13709 9831
rect 12780 9640 12900 9691
rect 13676 9691 13709 9794
rect 13755 9691 13796 9831
rect 14368 9831 14468 9880
rect 14368 9794 14381 9831
rect 1692 9432 1892 9476
rect 2140 9432 2340 9476
rect 2588 9432 2788 9476
rect 3036 9432 3236 9476
rect 3484 9432 3684 9476
rect 4156 9432 4276 9476
rect 4828 9432 4948 9476
rect 13676 9640 13796 9691
rect 14348 9691 14381 9794
rect 14427 9691 14468 9831
rect 15040 9831 15140 9880
rect 15040 9794 15053 9831
rect 14348 9640 14468 9691
rect 15020 9691 15053 9794
rect 15099 9691 15140 9831
rect 15712 9831 15812 9880
rect 15712 9794 15725 9831
rect 15020 9640 15140 9691
rect 15692 9691 15725 9794
rect 15771 9691 15812 9831
rect 16384 9831 16484 9880
rect 16384 9794 16397 9831
rect 15692 9640 15812 9691
rect 16364 9691 16397 9794
rect 16443 9691 16484 9831
rect 17056 9831 17156 9880
rect 17056 9794 17069 9831
rect 16364 9640 16484 9691
rect 17036 9691 17069 9794
rect 17115 9691 17156 9831
rect 17036 9640 17156 9691
rect 17788 9831 17888 9880
rect 17788 9691 17829 9831
rect 17875 9794 17888 9831
rect 18400 9831 18500 9880
rect 18400 9794 18413 9831
rect 17875 9691 17908 9794
rect 17788 9640 17908 9691
rect 18380 9691 18413 9794
rect 18459 9691 18500 9831
rect 19072 9831 19172 9880
rect 19072 9794 19085 9831
rect 18380 9640 18500 9691
rect 19052 9691 19085 9794
rect 19131 9691 19172 9831
rect 19744 9831 19844 9880
rect 19744 9794 19757 9831
rect 19052 9640 19172 9691
rect 19724 9691 19757 9794
rect 19803 9691 19844 9831
rect 20416 9831 20516 9880
rect 20416 9794 20429 9831
rect 19724 9640 19844 9691
rect 20396 9691 20429 9794
rect 20475 9691 20516 9831
rect 20844 9846 21044 9880
rect 20844 9800 20880 9846
rect 21020 9800 21044 9846
rect 20844 9783 21044 9800
rect 21648 9831 21748 9880
rect 21648 9794 21661 9831
rect 20396 9640 20516 9691
rect 20844 9719 21044 9732
rect 20844 9673 20872 9719
rect 21012 9673 21044 9719
rect 20844 9640 21044 9673
rect 21628 9691 21661 9794
rect 21707 9691 21748 9831
rect 22076 9846 22276 9880
rect 22076 9800 22112 9846
rect 22252 9800 22276 9846
rect 22076 9783 22276 9800
rect 5836 9432 5956 9476
rect 6508 9432 6628 9476
rect 7180 9432 7300 9476
rect 7852 9432 7972 9476
rect 8524 9432 8644 9476
rect 9196 9432 9316 9476
rect 9868 9432 9988 9476
rect 10540 9432 10660 9476
rect 10988 9432 11188 9476
rect 11436 9432 11556 9476
rect 12108 9432 12228 9476
rect 12780 9432 12900 9476
rect 21628 9640 21748 9691
rect 22076 9719 22276 9732
rect 22076 9673 22104 9719
rect 22244 9673 22276 9719
rect 22076 9640 22276 9673
rect 13676 9432 13796 9476
rect 14348 9432 14468 9476
rect 15020 9432 15140 9476
rect 15692 9432 15812 9476
rect 16364 9432 16484 9476
rect 17036 9432 17156 9476
rect 17788 9432 17908 9476
rect 18380 9432 18500 9476
rect 19052 9432 19172 9476
rect 19724 9432 19844 9476
rect 20396 9432 20516 9476
rect 20844 9432 21044 9476
rect 21628 9432 21748 9476
rect 22076 9432 22276 9476
rect 1692 9340 1892 9384
rect 2140 9340 2340 9384
rect 2588 9340 2788 9384
rect 3372 9340 3492 9384
rect 4044 9340 4164 9384
rect 4716 9340 4836 9384
rect 5388 9340 5508 9384
rect 6060 9340 6180 9384
rect 6732 9340 6852 9384
rect 7404 9340 7524 9384
rect 8188 9340 8308 9384
rect 8860 9340 8980 9384
rect 9644 9340 9844 9384
rect 10316 9340 10436 9384
rect 10988 9340 11108 9384
rect 11660 9340 11780 9384
rect 12332 9340 12452 9384
rect 13004 9340 13124 9384
rect 13676 9340 13796 9384
rect 14348 9340 14468 9384
rect 15020 9340 15140 9384
rect 15692 9340 15812 9384
rect 16364 9340 16484 9384
rect 16812 9340 17012 9384
rect 1692 9143 1892 9176
rect 1692 9097 1720 9143
rect 1860 9097 1892 9143
rect 1692 9084 1892 9097
rect 2140 9143 2340 9176
rect 2140 9097 2168 9143
rect 2308 9097 2340 9143
rect 2140 9084 2340 9097
rect 2588 9143 2788 9176
rect 2588 9097 2616 9143
rect 2756 9097 2788 9143
rect 2588 9084 2788 9097
rect 3372 9125 3492 9176
rect 1692 9016 1892 9033
rect 1692 8970 1728 9016
rect 1868 8970 1892 9016
rect 1692 8936 1892 8970
rect 2140 9016 2340 9033
rect 2140 8970 2176 9016
rect 2316 8970 2340 9016
rect 2140 8936 2340 8970
rect 2588 9016 2788 9033
rect 3372 9022 3405 9125
rect 2588 8970 2624 9016
rect 2764 8970 2788 9016
rect 2588 8936 2788 8970
rect 3392 8985 3405 9022
rect 3451 8985 3492 9125
rect 4044 9125 4164 9176
rect 4044 9022 4077 9125
rect 3392 8936 3492 8985
rect 4064 8985 4077 9022
rect 4123 8985 4164 9125
rect 4716 9125 4836 9176
rect 4716 9022 4749 9125
rect 4064 8936 4164 8985
rect 4736 8985 4749 9022
rect 4795 8985 4836 9125
rect 5388 9125 5508 9176
rect 5388 9022 5421 9125
rect 4736 8936 4836 8985
rect 5408 8985 5421 9022
rect 5467 8985 5508 9125
rect 6060 9125 6180 9176
rect 6060 9022 6093 9125
rect 5408 8936 5508 8985
rect 6080 8985 6093 9022
rect 6139 8985 6180 9125
rect 6732 9125 6852 9176
rect 6732 9022 6765 9125
rect 6080 8936 6180 8985
rect 6752 8985 6765 9022
rect 6811 8985 6852 9125
rect 7404 9125 7524 9176
rect 7404 9022 7437 9125
rect 6752 8936 6852 8985
rect 7424 8985 7437 9022
rect 7483 8985 7524 9125
rect 8188 9125 8308 9176
rect 8188 9022 8221 9125
rect 7424 8936 7524 8985
rect 8208 8985 8221 9022
rect 8267 8985 8308 9125
rect 8860 9125 8980 9176
rect 17708 9340 17828 9384
rect 18380 9340 18500 9384
rect 19052 9340 19172 9384
rect 19724 9340 19844 9384
rect 20396 9340 20516 9384
rect 20844 9340 21044 9384
rect 21292 9340 21492 9384
rect 21740 9340 21940 9384
rect 8860 9022 8893 9125
rect 8208 8936 8308 8985
rect 8880 8985 8893 9022
rect 8939 8985 8980 9125
rect 9644 9143 9844 9176
rect 9644 9097 9672 9143
rect 9812 9097 9844 9143
rect 9644 9084 9844 9097
rect 10316 9125 10436 9176
rect 8880 8936 8980 8985
rect 9644 9016 9844 9033
rect 10316 9022 10349 9125
rect 9644 8970 9680 9016
rect 9820 8970 9844 9016
rect 9644 8936 9844 8970
rect 10336 8985 10349 9022
rect 10395 8985 10436 9125
rect 10988 9125 11108 9176
rect 10988 9022 11021 9125
rect 10336 8936 10436 8985
rect 11008 8985 11021 9022
rect 11067 8985 11108 9125
rect 11660 9125 11780 9176
rect 11660 9022 11693 9125
rect 11008 8936 11108 8985
rect 11680 8985 11693 9022
rect 11739 8985 11780 9125
rect 12332 9125 12452 9176
rect 12332 9022 12365 9125
rect 11680 8936 11780 8985
rect 12352 8985 12365 9022
rect 12411 8985 12452 9125
rect 13004 9125 13124 9176
rect 13004 9022 13037 9125
rect 12352 8936 12452 8985
rect 13024 8985 13037 9022
rect 13083 8985 13124 9125
rect 13676 9125 13796 9176
rect 13676 9022 13709 9125
rect 13024 8936 13124 8985
rect 13696 8985 13709 9022
rect 13755 8985 13796 9125
rect 14348 9125 14468 9176
rect 14348 9022 14381 9125
rect 13696 8936 13796 8985
rect 14368 8985 14381 9022
rect 14427 8985 14468 9125
rect 15020 9125 15140 9176
rect 15020 9022 15053 9125
rect 14368 8936 14468 8985
rect 15040 8985 15053 9022
rect 15099 8985 15140 9125
rect 15692 9125 15812 9176
rect 15692 9022 15725 9125
rect 15040 8936 15140 8985
rect 15712 8985 15725 9022
rect 15771 8985 15812 9125
rect 16364 9125 16484 9176
rect 16364 9022 16397 9125
rect 15712 8936 15812 8985
rect 16384 8985 16397 9022
rect 16443 8985 16484 9125
rect 16812 9143 17012 9176
rect 16812 9097 16840 9143
rect 16980 9097 17012 9143
rect 16812 9084 17012 9097
rect 17708 9125 17828 9176
rect 16384 8936 16484 8985
rect 16812 9016 17012 9033
rect 16812 8970 16848 9016
rect 16988 8970 17012 9016
rect 16812 8936 17012 8970
rect 17708 9022 17741 9125
rect 17728 8985 17741 9022
rect 17787 8985 17828 9125
rect 18380 9125 18500 9176
rect 18380 9022 18413 9125
rect 17728 8936 17828 8985
rect 18400 8985 18413 9022
rect 18459 8985 18500 9125
rect 19052 9125 19172 9176
rect 19052 9022 19085 9125
rect 18400 8936 18500 8985
rect 19072 8985 19085 9022
rect 19131 8985 19172 9125
rect 19724 9125 19844 9176
rect 19724 9022 19757 9125
rect 19072 8936 19172 8985
rect 19744 8985 19757 9022
rect 19803 8985 19844 9125
rect 20396 9125 20516 9176
rect 20396 9022 20429 9125
rect 19744 8936 19844 8985
rect 20416 8985 20429 9022
rect 20475 8985 20516 9125
rect 20844 9143 21044 9176
rect 20844 9097 20872 9143
rect 21012 9097 21044 9143
rect 20844 9084 21044 9097
rect 21292 9143 21492 9176
rect 21292 9097 21320 9143
rect 21460 9097 21492 9143
rect 21292 9084 21492 9097
rect 21740 9143 21940 9176
rect 21740 9097 21768 9143
rect 21908 9097 21940 9143
rect 21740 9084 21940 9097
rect 20416 8936 20516 8985
rect 20844 9016 21044 9033
rect 20844 8970 20880 9016
rect 21020 8970 21044 9016
rect 20844 8936 21044 8970
rect 21292 9016 21492 9033
rect 21292 8970 21328 9016
rect 21468 8970 21492 9016
rect 21292 8936 21492 8970
rect 21740 9016 21940 9033
rect 21740 8970 21776 9016
rect 21916 8970 21940 9016
rect 21740 8936 21940 8970
rect 1692 8648 1892 8692
rect 2140 8648 2340 8692
rect 2588 8648 2788 8692
rect 3392 8648 3492 8692
rect 4064 8648 4164 8692
rect 4736 8648 4836 8692
rect 5408 8648 5508 8692
rect 6080 8648 6180 8692
rect 6752 8648 6852 8692
rect 7424 8648 7524 8692
rect 8208 8648 8308 8692
rect 8880 8648 8980 8692
rect 9644 8648 9844 8692
rect 10336 8648 10436 8692
rect 11008 8648 11108 8692
rect 11680 8648 11780 8692
rect 12352 8648 12452 8692
rect 13024 8648 13124 8692
rect 13696 8648 13796 8692
rect 14368 8648 14468 8692
rect 15040 8648 15140 8692
rect 15712 8648 15812 8692
rect 16384 8648 16484 8692
rect 16812 8648 17012 8692
rect 17728 8648 17828 8692
rect 18400 8648 18500 8692
rect 19072 8648 19172 8692
rect 19744 8648 19844 8692
rect 20416 8648 20516 8692
rect 20844 8648 21044 8692
rect 21292 8648 21492 8692
rect 21740 8648 21940 8692
rect 1692 8556 1892 8600
rect 2140 8556 2340 8600
rect 2892 8556 2992 8600
rect 3504 8556 3604 8600
rect 4176 8556 4276 8600
rect 4848 8556 4948 8600
rect 5856 8556 5956 8600
rect 6528 8556 6628 8600
rect 7200 8556 7300 8600
rect 7872 8556 7972 8600
rect 8544 8556 8644 8600
rect 9216 8556 9316 8600
rect 9888 8556 9988 8600
rect 10560 8556 10660 8600
rect 11292 8556 11392 8600
rect 11660 8556 11860 8600
rect 12128 8556 12228 8600
rect 12800 8556 12900 8600
rect 13696 8556 13796 8600
rect 14368 8556 14468 8600
rect 15040 8556 15140 8600
rect 15712 8556 15812 8600
rect 16384 8556 16484 8600
rect 17056 8556 17156 8600
rect 17728 8556 17828 8600
rect 18400 8556 18500 8600
rect 19072 8556 19172 8600
rect 19744 8556 19844 8600
rect 20476 8556 20576 8600
rect 20844 8556 21044 8600
rect 21516 8556 21716 8600
rect 21964 8556 22164 8600
rect 1692 8278 1892 8312
rect 1692 8232 1728 8278
rect 1868 8232 1892 8278
rect 1692 8215 1892 8232
rect 2140 8278 2340 8312
rect 2140 8232 2176 8278
rect 2316 8232 2340 8278
rect 2140 8215 2340 8232
rect 2892 8263 2992 8312
rect 1692 8151 1892 8164
rect 1692 8105 1720 8151
rect 1860 8105 1892 8151
rect 1692 8072 1892 8105
rect 2140 8151 2340 8164
rect 2140 8105 2168 8151
rect 2308 8105 2340 8151
rect 2140 8072 2340 8105
rect 2892 8123 2933 8263
rect 2979 8226 2992 8263
rect 3504 8263 3604 8312
rect 3504 8226 3517 8263
rect 2979 8123 3012 8226
rect 2892 8072 3012 8123
rect 3484 8123 3517 8226
rect 3563 8123 3604 8263
rect 4176 8263 4276 8312
rect 4176 8226 4189 8263
rect 3484 8072 3604 8123
rect 4156 8123 4189 8226
rect 4235 8123 4276 8263
rect 4848 8263 4948 8312
rect 4848 8226 4861 8263
rect 4156 8072 4276 8123
rect 4828 8123 4861 8226
rect 4907 8123 4948 8263
rect 5856 8263 5956 8312
rect 5856 8226 5869 8263
rect 4828 8072 4948 8123
rect 5836 8123 5869 8226
rect 5915 8123 5956 8263
rect 6528 8263 6628 8312
rect 6528 8226 6541 8263
rect 5836 8072 5956 8123
rect 6508 8123 6541 8226
rect 6587 8123 6628 8263
rect 7200 8263 7300 8312
rect 7200 8226 7213 8263
rect 6508 8072 6628 8123
rect 7180 8123 7213 8226
rect 7259 8123 7300 8263
rect 7872 8263 7972 8312
rect 7872 8226 7885 8263
rect 7180 8072 7300 8123
rect 7852 8123 7885 8226
rect 7931 8123 7972 8263
rect 8544 8263 8644 8312
rect 8544 8226 8557 8263
rect 7852 8072 7972 8123
rect 8524 8123 8557 8226
rect 8603 8123 8644 8263
rect 9216 8263 9316 8312
rect 9216 8226 9229 8263
rect 8524 8072 8644 8123
rect 9196 8123 9229 8226
rect 9275 8123 9316 8263
rect 9888 8263 9988 8312
rect 9888 8226 9901 8263
rect 9196 8072 9316 8123
rect 9868 8123 9901 8226
rect 9947 8123 9988 8263
rect 10560 8263 10660 8312
rect 10560 8226 10573 8263
rect 9868 8072 9988 8123
rect 10540 8123 10573 8226
rect 10619 8123 10660 8263
rect 10540 8072 10660 8123
rect 11292 8263 11392 8312
rect 11292 8123 11333 8263
rect 11379 8226 11392 8263
rect 11660 8278 11860 8312
rect 11660 8232 11696 8278
rect 11836 8232 11860 8278
rect 11379 8123 11412 8226
rect 11660 8215 11860 8232
rect 12128 8263 12228 8312
rect 12128 8226 12141 8263
rect 11292 8072 11412 8123
rect 11660 8151 11860 8164
rect 11660 8105 11688 8151
rect 11828 8105 11860 8151
rect 11660 8072 11860 8105
rect 12108 8123 12141 8226
rect 12187 8123 12228 8263
rect 12800 8263 12900 8312
rect 12800 8226 12813 8263
rect 12108 8072 12228 8123
rect 12780 8123 12813 8226
rect 12859 8123 12900 8263
rect 13696 8263 13796 8312
rect 13696 8226 13709 8263
rect 12780 8072 12900 8123
rect 13676 8123 13709 8226
rect 13755 8123 13796 8263
rect 14368 8263 14468 8312
rect 14368 8226 14381 8263
rect 1692 7864 1892 7908
rect 2140 7864 2340 7908
rect 2892 7864 3012 7908
rect 3484 7864 3604 7908
rect 4156 7864 4276 7908
rect 4828 7864 4948 7908
rect 13676 8072 13796 8123
rect 14348 8123 14381 8226
rect 14427 8123 14468 8263
rect 15040 8263 15140 8312
rect 15040 8226 15053 8263
rect 14348 8072 14468 8123
rect 15020 8123 15053 8226
rect 15099 8123 15140 8263
rect 15712 8263 15812 8312
rect 15712 8226 15725 8263
rect 15020 8072 15140 8123
rect 15692 8123 15725 8226
rect 15771 8123 15812 8263
rect 16384 8263 16484 8312
rect 16384 8226 16397 8263
rect 15692 8072 15812 8123
rect 16364 8123 16397 8226
rect 16443 8123 16484 8263
rect 17056 8263 17156 8312
rect 17056 8226 17069 8263
rect 16364 8072 16484 8123
rect 17036 8123 17069 8226
rect 17115 8123 17156 8263
rect 17728 8263 17828 8312
rect 17728 8226 17741 8263
rect 17036 8072 17156 8123
rect 17708 8123 17741 8226
rect 17787 8123 17828 8263
rect 18400 8263 18500 8312
rect 18400 8226 18413 8263
rect 17708 8072 17828 8123
rect 18380 8123 18413 8226
rect 18459 8123 18500 8263
rect 19072 8263 19172 8312
rect 19072 8226 19085 8263
rect 18380 8072 18500 8123
rect 19052 8123 19085 8226
rect 19131 8123 19172 8263
rect 19744 8263 19844 8312
rect 19744 8226 19757 8263
rect 19052 8072 19172 8123
rect 19724 8123 19757 8226
rect 19803 8123 19844 8263
rect 19724 8072 19844 8123
rect 20476 8263 20576 8312
rect 20476 8123 20517 8263
rect 20563 8226 20576 8263
rect 20844 8278 21044 8312
rect 20844 8232 20880 8278
rect 21020 8232 21044 8278
rect 20563 8123 20596 8226
rect 20844 8215 21044 8232
rect 21516 8278 21716 8312
rect 21516 8232 21552 8278
rect 21692 8232 21716 8278
rect 21516 8215 21716 8232
rect 21964 8278 22164 8312
rect 21964 8232 22000 8278
rect 22140 8232 22164 8278
rect 21964 8215 22164 8232
rect 20476 8072 20596 8123
rect 20844 8151 21044 8164
rect 20844 8105 20872 8151
rect 21012 8105 21044 8151
rect 20844 8072 21044 8105
rect 21516 8151 21716 8164
rect 21516 8105 21544 8151
rect 21684 8105 21716 8151
rect 5836 7864 5956 7908
rect 6508 7864 6628 7908
rect 7180 7864 7300 7908
rect 7852 7864 7972 7908
rect 8524 7864 8644 7908
rect 9196 7864 9316 7908
rect 9868 7864 9988 7908
rect 10540 7864 10660 7908
rect 11292 7864 11412 7908
rect 11660 7864 11860 7908
rect 12108 7864 12228 7908
rect 12780 7864 12900 7908
rect 21516 8072 21716 8105
rect 21964 8151 22164 8164
rect 21964 8105 21992 8151
rect 22132 8105 22164 8151
rect 21964 8072 22164 8105
rect 13676 7864 13796 7908
rect 14348 7864 14468 7908
rect 15020 7864 15140 7908
rect 15692 7864 15812 7908
rect 16364 7864 16484 7908
rect 17036 7864 17156 7908
rect 17708 7864 17828 7908
rect 18380 7864 18500 7908
rect 19052 7864 19172 7908
rect 19724 7864 19844 7908
rect 20476 7864 20596 7908
rect 20844 7864 21044 7908
rect 21516 7864 21716 7908
rect 21964 7864 22164 7908
rect 2108 7772 2228 7816
rect 2700 7772 2820 7816
rect 3372 7772 3492 7816
rect 4044 7772 4164 7816
rect 4716 7772 4836 7816
rect 5388 7772 5508 7816
rect 6060 7772 6180 7816
rect 6732 7772 6852 7816
rect 7404 7772 7524 7816
rect 8188 7772 8308 7816
rect 8860 7772 8980 7816
rect 9868 7772 9988 7816
rect 10540 7772 10660 7816
rect 11292 7772 11412 7816
rect 11884 7772 12004 7816
rect 12556 7772 12676 7816
rect 13228 7772 13348 7816
rect 13900 7772 14020 7816
rect 14572 7772 14692 7816
rect 15244 7772 15364 7816
rect 15916 7772 16036 7816
rect 16588 7772 16708 7816
rect 2108 7557 2228 7608
rect 2108 7417 2149 7557
rect 2195 7454 2228 7557
rect 2700 7557 2820 7608
rect 2700 7454 2733 7557
rect 2195 7417 2208 7454
rect 2108 7368 2208 7417
rect 2720 7417 2733 7454
rect 2779 7417 2820 7557
rect 3372 7557 3492 7608
rect 3372 7454 3405 7557
rect 2720 7368 2820 7417
rect 3392 7417 3405 7454
rect 3451 7417 3492 7557
rect 4044 7557 4164 7608
rect 4044 7454 4077 7557
rect 3392 7368 3492 7417
rect 4064 7417 4077 7454
rect 4123 7417 4164 7557
rect 4716 7557 4836 7608
rect 4716 7454 4749 7557
rect 4064 7368 4164 7417
rect 4736 7417 4749 7454
rect 4795 7417 4836 7557
rect 5388 7557 5508 7608
rect 5388 7454 5421 7557
rect 4736 7368 4836 7417
rect 5408 7417 5421 7454
rect 5467 7417 5508 7557
rect 6060 7557 6180 7608
rect 6060 7454 6093 7557
rect 5408 7368 5508 7417
rect 6080 7417 6093 7454
rect 6139 7417 6180 7557
rect 6732 7557 6852 7608
rect 6732 7454 6765 7557
rect 6080 7368 6180 7417
rect 6752 7417 6765 7454
rect 6811 7417 6852 7557
rect 7404 7557 7524 7608
rect 7404 7454 7437 7557
rect 6752 7368 6852 7417
rect 7424 7417 7437 7454
rect 7483 7417 7524 7557
rect 8188 7557 8308 7608
rect 8188 7454 8221 7557
rect 7424 7368 7524 7417
rect 8208 7417 8221 7454
rect 8267 7417 8308 7557
rect 8860 7557 8980 7608
rect 17708 7772 17828 7816
rect 18380 7772 18500 7816
rect 19052 7772 19172 7816
rect 19724 7772 19844 7816
rect 20396 7772 20516 7816
rect 21068 7772 21188 7816
rect 21516 7772 21716 7816
rect 21964 7772 22164 7816
rect 8860 7454 8893 7557
rect 8208 7368 8308 7417
rect 8880 7417 8893 7454
rect 8939 7417 8980 7557
rect 9868 7557 9988 7608
rect 8880 7368 8980 7417
rect 9868 7454 9901 7557
rect 9888 7417 9901 7454
rect 9947 7417 9988 7557
rect 10540 7557 10660 7608
rect 10540 7454 10573 7557
rect 9888 7368 9988 7417
rect 10560 7417 10573 7454
rect 10619 7417 10660 7557
rect 10560 7368 10660 7417
rect 11292 7557 11412 7608
rect 11292 7417 11333 7557
rect 11379 7454 11412 7557
rect 11884 7557 12004 7608
rect 11884 7454 11917 7557
rect 11379 7417 11392 7454
rect 11292 7368 11392 7417
rect 11904 7417 11917 7454
rect 11963 7417 12004 7557
rect 12556 7557 12676 7608
rect 12556 7454 12589 7557
rect 11904 7368 12004 7417
rect 12576 7417 12589 7454
rect 12635 7417 12676 7557
rect 13228 7557 13348 7608
rect 13228 7454 13261 7557
rect 12576 7368 12676 7417
rect 13248 7417 13261 7454
rect 13307 7417 13348 7557
rect 13900 7557 14020 7608
rect 13900 7454 13933 7557
rect 13248 7368 13348 7417
rect 13920 7417 13933 7454
rect 13979 7417 14020 7557
rect 14572 7557 14692 7608
rect 14572 7454 14605 7557
rect 13920 7368 14020 7417
rect 14592 7417 14605 7454
rect 14651 7417 14692 7557
rect 15244 7557 15364 7608
rect 15244 7454 15277 7557
rect 14592 7368 14692 7417
rect 15264 7417 15277 7454
rect 15323 7417 15364 7557
rect 15916 7557 16036 7608
rect 15916 7454 15949 7557
rect 15264 7368 15364 7417
rect 15936 7417 15949 7454
rect 15995 7417 16036 7557
rect 16588 7557 16708 7608
rect 16588 7454 16621 7557
rect 15936 7368 16036 7417
rect 16608 7417 16621 7454
rect 16667 7417 16708 7557
rect 17708 7557 17828 7608
rect 16608 7368 16708 7417
rect 17708 7454 17741 7557
rect 17728 7417 17741 7454
rect 17787 7417 17828 7557
rect 18380 7557 18500 7608
rect 18380 7454 18413 7557
rect 17728 7368 17828 7417
rect 18400 7417 18413 7454
rect 18459 7417 18500 7557
rect 19052 7557 19172 7608
rect 19052 7454 19085 7557
rect 18400 7368 18500 7417
rect 19072 7417 19085 7454
rect 19131 7417 19172 7557
rect 19724 7557 19844 7608
rect 19724 7454 19757 7557
rect 19072 7368 19172 7417
rect 19744 7417 19757 7454
rect 19803 7417 19844 7557
rect 20396 7557 20516 7608
rect 20396 7454 20429 7557
rect 19744 7368 19844 7417
rect 20416 7417 20429 7454
rect 20475 7417 20516 7557
rect 21068 7557 21188 7608
rect 21068 7454 21101 7557
rect 20416 7368 20516 7417
rect 21088 7417 21101 7454
rect 21147 7417 21188 7557
rect 21516 7575 21716 7608
rect 21516 7529 21544 7575
rect 21684 7529 21716 7575
rect 21516 7516 21716 7529
rect 21964 7575 22164 7608
rect 21964 7529 21992 7575
rect 22132 7529 22164 7575
rect 21964 7516 22164 7529
rect 21088 7368 21188 7417
rect 21516 7448 21716 7465
rect 21516 7402 21552 7448
rect 21692 7402 21716 7448
rect 21516 7368 21716 7402
rect 21964 7448 22164 7465
rect 21964 7402 22000 7448
rect 22140 7402 22164 7448
rect 21964 7368 22164 7402
rect 2108 7080 2208 7124
rect 2720 7080 2820 7124
rect 3392 7080 3492 7124
rect 4064 7080 4164 7124
rect 4736 7080 4836 7124
rect 5408 7080 5508 7124
rect 6080 7080 6180 7124
rect 6752 7080 6852 7124
rect 7424 7080 7524 7124
rect 8208 7080 8308 7124
rect 8880 7080 8980 7124
rect 9888 7080 9988 7124
rect 10560 7080 10660 7124
rect 11292 7080 11392 7124
rect 11904 7080 12004 7124
rect 12576 7080 12676 7124
rect 13248 7080 13348 7124
rect 13920 7080 14020 7124
rect 14592 7080 14692 7124
rect 15264 7080 15364 7124
rect 15936 7080 16036 7124
rect 16608 7080 16708 7124
rect 17728 7080 17828 7124
rect 18400 7080 18500 7124
rect 19072 7080 19172 7124
rect 19744 7080 19844 7124
rect 20416 7080 20516 7124
rect 21088 7080 21188 7124
rect 21516 7080 21716 7124
rect 21964 7080 22164 7124
rect 1692 6988 1892 7032
rect 2160 6988 2260 7032
rect 2832 6988 2932 7032
rect 3504 6988 3604 7032
rect 4176 6988 4276 7032
rect 4848 6988 4948 7032
rect 5744 6988 5844 7032
rect 6416 6988 6516 7032
rect 7088 6988 7188 7032
rect 7760 6988 7860 7032
rect 8432 6988 8532 7032
rect 9104 6988 9204 7032
rect 9776 6988 9876 7032
rect 10448 6988 10548 7032
rect 11120 6988 11220 7032
rect 11792 6988 11892 7032
rect 12464 6988 12564 7032
rect 12892 6988 13092 7032
rect 13564 6988 13764 7032
rect 14144 6988 14244 7032
rect 14816 6988 14916 7032
rect 15488 6988 15588 7032
rect 16160 6988 16260 7032
rect 16832 6988 16932 7032
rect 17504 6988 17604 7032
rect 18176 6988 18276 7032
rect 18848 6988 18948 7032
rect 19520 6988 19620 7032
rect 20252 6988 20352 7032
rect 20620 6988 20820 7032
rect 21648 6988 21748 7032
rect 22076 6988 22276 7032
rect 1692 6710 1892 6744
rect 1692 6664 1728 6710
rect 1868 6664 1892 6710
rect 1692 6647 1892 6664
rect 2160 6695 2260 6744
rect 2160 6658 2173 6695
rect 1692 6583 1892 6596
rect 1692 6537 1720 6583
rect 1860 6537 1892 6583
rect 1692 6504 1892 6537
rect 2140 6555 2173 6658
rect 2219 6555 2260 6695
rect 2832 6695 2932 6744
rect 2832 6658 2845 6695
rect 2140 6504 2260 6555
rect 2812 6555 2845 6658
rect 2891 6555 2932 6695
rect 3504 6695 3604 6744
rect 3504 6658 3517 6695
rect 2812 6504 2932 6555
rect 3484 6555 3517 6658
rect 3563 6555 3604 6695
rect 4176 6695 4276 6744
rect 4176 6658 4189 6695
rect 3484 6504 3604 6555
rect 4156 6555 4189 6658
rect 4235 6555 4276 6695
rect 4848 6695 4948 6744
rect 4848 6658 4861 6695
rect 4156 6504 4276 6555
rect 4828 6555 4861 6658
rect 4907 6555 4948 6695
rect 5744 6695 5844 6744
rect 5744 6658 5757 6695
rect 4828 6504 4948 6555
rect 5724 6555 5757 6658
rect 5803 6555 5844 6695
rect 6416 6695 6516 6744
rect 6416 6658 6429 6695
rect 5724 6504 5844 6555
rect 6396 6555 6429 6658
rect 6475 6555 6516 6695
rect 7088 6695 7188 6744
rect 7088 6658 7101 6695
rect 6396 6504 6516 6555
rect 7068 6555 7101 6658
rect 7147 6555 7188 6695
rect 7760 6695 7860 6744
rect 7760 6658 7773 6695
rect 7068 6504 7188 6555
rect 7740 6555 7773 6658
rect 7819 6555 7860 6695
rect 8432 6695 8532 6744
rect 8432 6658 8445 6695
rect 7740 6504 7860 6555
rect 8412 6555 8445 6658
rect 8491 6555 8532 6695
rect 9104 6695 9204 6744
rect 9104 6658 9117 6695
rect 8412 6504 8532 6555
rect 9084 6555 9117 6658
rect 9163 6555 9204 6695
rect 9776 6695 9876 6744
rect 9776 6658 9789 6695
rect 9084 6504 9204 6555
rect 9756 6555 9789 6658
rect 9835 6555 9876 6695
rect 10448 6695 10548 6744
rect 10448 6658 10461 6695
rect 9756 6504 9876 6555
rect 10428 6555 10461 6658
rect 10507 6555 10548 6695
rect 11120 6695 11220 6744
rect 11120 6658 11133 6695
rect 10428 6504 10548 6555
rect 11100 6555 11133 6658
rect 11179 6555 11220 6695
rect 11792 6695 11892 6744
rect 11792 6658 11805 6695
rect 11100 6504 11220 6555
rect 11772 6555 11805 6658
rect 11851 6555 11892 6695
rect 12464 6695 12564 6744
rect 12464 6658 12477 6695
rect 11772 6504 11892 6555
rect 12444 6555 12477 6658
rect 12523 6555 12564 6695
rect 12892 6710 13092 6744
rect 12892 6664 12928 6710
rect 13068 6664 13092 6710
rect 12892 6647 13092 6664
rect 13564 6710 13764 6744
rect 13564 6664 13600 6710
rect 13740 6664 13764 6710
rect 13564 6647 13764 6664
rect 14144 6695 14244 6744
rect 14144 6658 14157 6695
rect 12444 6504 12564 6555
rect 12892 6583 13092 6596
rect 12892 6537 12920 6583
rect 13060 6537 13092 6583
rect 12892 6504 13092 6537
rect 13564 6583 13764 6596
rect 13564 6537 13592 6583
rect 13732 6537 13764 6583
rect 1692 6296 1892 6340
rect 2140 6296 2260 6340
rect 2812 6296 2932 6340
rect 3484 6296 3604 6340
rect 4156 6296 4276 6340
rect 4828 6296 4948 6340
rect 13564 6504 13764 6537
rect 14124 6555 14157 6658
rect 14203 6555 14244 6695
rect 14816 6695 14916 6744
rect 14816 6658 14829 6695
rect 14124 6504 14244 6555
rect 14796 6555 14829 6658
rect 14875 6555 14916 6695
rect 15488 6695 15588 6744
rect 15488 6658 15501 6695
rect 14796 6504 14916 6555
rect 15468 6555 15501 6658
rect 15547 6555 15588 6695
rect 16160 6695 16260 6744
rect 16160 6658 16173 6695
rect 15468 6504 15588 6555
rect 16140 6555 16173 6658
rect 16219 6555 16260 6695
rect 16832 6695 16932 6744
rect 16832 6658 16845 6695
rect 16140 6504 16260 6555
rect 16812 6555 16845 6658
rect 16891 6555 16932 6695
rect 17504 6695 17604 6744
rect 17504 6658 17517 6695
rect 16812 6504 16932 6555
rect 17484 6555 17517 6658
rect 17563 6555 17604 6695
rect 18176 6695 18276 6744
rect 18176 6658 18189 6695
rect 17484 6504 17604 6555
rect 18156 6555 18189 6658
rect 18235 6555 18276 6695
rect 18848 6695 18948 6744
rect 18848 6658 18861 6695
rect 18156 6504 18276 6555
rect 18828 6555 18861 6658
rect 18907 6555 18948 6695
rect 19520 6695 19620 6744
rect 19520 6658 19533 6695
rect 18828 6504 18948 6555
rect 19500 6555 19533 6658
rect 19579 6555 19620 6695
rect 19500 6504 19620 6555
rect 20252 6695 20352 6744
rect 20252 6555 20293 6695
rect 20339 6658 20352 6695
rect 20620 6710 20820 6744
rect 20620 6664 20656 6710
rect 20796 6664 20820 6710
rect 20339 6555 20372 6658
rect 20620 6647 20820 6664
rect 21648 6695 21748 6744
rect 21648 6658 21661 6695
rect 20252 6504 20372 6555
rect 20620 6583 20820 6596
rect 20620 6537 20648 6583
rect 20788 6537 20820 6583
rect 20620 6504 20820 6537
rect 21628 6555 21661 6658
rect 21707 6555 21748 6695
rect 22076 6710 22276 6744
rect 22076 6664 22112 6710
rect 22252 6664 22276 6710
rect 22076 6647 22276 6664
rect 5724 6296 5844 6340
rect 6396 6296 6516 6340
rect 7068 6296 7188 6340
rect 7740 6296 7860 6340
rect 8412 6296 8532 6340
rect 9084 6296 9204 6340
rect 9756 6296 9876 6340
rect 10428 6296 10548 6340
rect 11100 6296 11220 6340
rect 11772 6296 11892 6340
rect 12444 6296 12564 6340
rect 12892 6296 13092 6340
rect 21628 6504 21748 6555
rect 22076 6583 22276 6596
rect 22076 6537 22104 6583
rect 22244 6537 22276 6583
rect 22076 6504 22276 6537
rect 13564 6296 13764 6340
rect 14124 6296 14244 6340
rect 14796 6296 14916 6340
rect 15468 6296 15588 6340
rect 16140 6296 16260 6340
rect 16812 6296 16932 6340
rect 17484 6296 17604 6340
rect 18156 6296 18276 6340
rect 18828 6296 18948 6340
rect 19500 6296 19620 6340
rect 20252 6296 20372 6340
rect 20620 6296 20820 6340
rect 21628 6296 21748 6340
rect 22076 6296 22276 6340
rect 2028 6204 2148 6248
rect 2700 6204 2820 6248
rect 3372 6204 3492 6248
rect 4044 6204 4164 6248
rect 4716 6204 4836 6248
rect 5388 6204 5508 6248
rect 6060 6204 6180 6248
rect 6732 6204 6852 6248
rect 7404 6204 7524 6248
rect 8076 6204 8196 6248
rect 8748 6204 8868 6248
rect 9756 6204 9876 6248
rect 10428 6204 10548 6248
rect 11100 6204 11220 6248
rect 11772 6204 11892 6248
rect 12556 6204 12676 6248
rect 13228 6204 13348 6248
rect 13900 6204 14020 6248
rect 14572 6204 14692 6248
rect 15244 6204 15364 6248
rect 15916 6204 16036 6248
rect 16588 6204 16708 6248
rect 2028 5989 2148 6040
rect 2028 5886 2061 5989
rect 2048 5849 2061 5886
rect 2107 5849 2148 5989
rect 2700 5989 2820 6040
rect 2700 5886 2733 5989
rect 2048 5800 2148 5849
rect 2720 5849 2733 5886
rect 2779 5849 2820 5989
rect 3372 5989 3492 6040
rect 3372 5886 3405 5989
rect 2720 5800 2820 5849
rect 3392 5849 3405 5886
rect 3451 5849 3492 5989
rect 4044 5989 4164 6040
rect 4044 5886 4077 5989
rect 3392 5800 3492 5849
rect 4064 5849 4077 5886
rect 4123 5849 4164 5989
rect 4716 5989 4836 6040
rect 4716 5886 4749 5989
rect 4064 5800 4164 5849
rect 4736 5849 4749 5886
rect 4795 5849 4836 5989
rect 5388 5989 5508 6040
rect 5388 5886 5421 5989
rect 4736 5800 4836 5849
rect 5408 5849 5421 5886
rect 5467 5849 5508 5989
rect 6060 5989 6180 6040
rect 6060 5886 6093 5989
rect 5408 5800 5508 5849
rect 6080 5849 6093 5886
rect 6139 5849 6180 5989
rect 6732 5989 6852 6040
rect 6732 5886 6765 5989
rect 6080 5800 6180 5849
rect 6752 5849 6765 5886
rect 6811 5849 6852 5989
rect 7404 5989 7524 6040
rect 7404 5886 7437 5989
rect 6752 5800 6852 5849
rect 7424 5849 7437 5886
rect 7483 5849 7524 5989
rect 8076 5989 8196 6040
rect 8076 5886 8109 5989
rect 7424 5800 7524 5849
rect 8096 5849 8109 5886
rect 8155 5849 8196 5989
rect 8748 5989 8868 6040
rect 17708 6204 17828 6248
rect 18380 6204 18500 6248
rect 19052 6204 19172 6248
rect 19724 6204 19844 6248
rect 20396 6204 20516 6248
rect 21068 6204 21188 6248
rect 21820 6204 21940 6248
rect 8748 5886 8781 5989
rect 8096 5800 8196 5849
rect 8768 5849 8781 5886
rect 8827 5849 8868 5989
rect 9756 5989 9876 6040
rect 8768 5800 8868 5849
rect 9756 5886 9789 5989
rect 9776 5849 9789 5886
rect 9835 5849 9876 5989
rect 10428 5989 10548 6040
rect 10428 5886 10461 5989
rect 9776 5800 9876 5849
rect 10448 5849 10461 5886
rect 10507 5849 10548 5989
rect 11100 5989 11220 6040
rect 11100 5886 11133 5989
rect 10448 5800 10548 5849
rect 11120 5849 11133 5886
rect 11179 5849 11220 5989
rect 11772 5989 11892 6040
rect 11772 5886 11805 5989
rect 11120 5800 11220 5849
rect 11792 5849 11805 5886
rect 11851 5849 11892 5989
rect 12556 5989 12676 6040
rect 12556 5886 12589 5989
rect 11792 5800 11892 5849
rect 12576 5849 12589 5886
rect 12635 5849 12676 5989
rect 13228 5989 13348 6040
rect 13228 5886 13261 5989
rect 12576 5800 12676 5849
rect 13248 5849 13261 5886
rect 13307 5849 13348 5989
rect 13900 5989 14020 6040
rect 13900 5886 13933 5989
rect 13248 5800 13348 5849
rect 13920 5849 13933 5886
rect 13979 5849 14020 5989
rect 14572 5989 14692 6040
rect 14572 5886 14605 5989
rect 13920 5800 14020 5849
rect 14592 5849 14605 5886
rect 14651 5849 14692 5989
rect 15244 5989 15364 6040
rect 15244 5886 15277 5989
rect 14592 5800 14692 5849
rect 15264 5849 15277 5886
rect 15323 5849 15364 5989
rect 15916 5989 16036 6040
rect 15916 5886 15949 5989
rect 15264 5800 15364 5849
rect 15936 5849 15949 5886
rect 15995 5849 16036 5989
rect 16588 5989 16708 6040
rect 16588 5886 16621 5989
rect 15936 5800 16036 5849
rect 16608 5849 16621 5886
rect 16667 5849 16708 5989
rect 17708 5989 17828 6040
rect 16608 5800 16708 5849
rect 17708 5886 17741 5989
rect 17728 5849 17741 5886
rect 17787 5849 17828 5989
rect 18380 5989 18500 6040
rect 18380 5886 18413 5989
rect 17728 5800 17828 5849
rect 18400 5849 18413 5886
rect 18459 5849 18500 5989
rect 19052 5989 19172 6040
rect 19052 5886 19085 5989
rect 18400 5800 18500 5849
rect 19072 5849 19085 5886
rect 19131 5849 19172 5989
rect 19724 5989 19844 6040
rect 19724 5886 19757 5989
rect 19072 5800 19172 5849
rect 19744 5849 19757 5886
rect 19803 5849 19844 5989
rect 20396 5989 20516 6040
rect 20396 5886 20429 5989
rect 19744 5800 19844 5849
rect 20416 5849 20429 5886
rect 20475 5849 20516 5989
rect 21068 5989 21188 6040
rect 21068 5886 21101 5989
rect 20416 5800 20516 5849
rect 21088 5849 21101 5886
rect 21147 5849 21188 5989
rect 21088 5800 21188 5849
rect 21820 5989 21940 6040
rect 21820 5849 21861 5989
rect 21907 5886 21940 5989
rect 21907 5849 21920 5886
rect 21820 5800 21920 5849
rect 2048 5512 2148 5556
rect 2720 5512 2820 5556
rect 3392 5512 3492 5556
rect 4064 5512 4164 5556
rect 4736 5512 4836 5556
rect 5408 5512 5508 5556
rect 6080 5512 6180 5556
rect 6752 5512 6852 5556
rect 7424 5512 7524 5556
rect 8096 5512 8196 5556
rect 8768 5512 8868 5556
rect 9776 5512 9876 5556
rect 10448 5512 10548 5556
rect 11120 5512 11220 5556
rect 11792 5512 11892 5556
rect 12576 5512 12676 5556
rect 13248 5512 13348 5556
rect 13920 5512 14020 5556
rect 14592 5512 14692 5556
rect 15264 5512 15364 5556
rect 15936 5512 16036 5556
rect 16608 5512 16708 5556
rect 17728 5512 17828 5556
rect 18400 5512 18500 5556
rect 19072 5512 19172 5556
rect 19744 5512 19844 5556
rect 20416 5512 20516 5556
rect 21088 5512 21188 5556
rect 21820 5512 21920 5556
rect 1692 5420 1892 5464
rect 2160 5420 2260 5464
rect 2832 5420 2932 5464
rect 3504 5420 3604 5464
rect 4176 5420 4276 5464
rect 4848 5420 4948 5464
rect 5744 5420 5844 5464
rect 6416 5420 6516 5464
rect 7088 5420 7188 5464
rect 7760 5420 7860 5464
rect 8432 5420 8532 5464
rect 9104 5420 9204 5464
rect 9776 5420 9876 5464
rect 10448 5420 10548 5464
rect 10876 5420 11076 5464
rect 11456 5420 11556 5464
rect 12128 5420 12228 5464
rect 12800 5420 12900 5464
rect 13564 5420 13764 5464
rect 14032 5420 14132 5464
rect 14704 5420 14804 5464
rect 15376 5420 15476 5464
rect 16048 5420 16148 5464
rect 16720 5420 16820 5464
rect 17392 5420 17492 5464
rect 18064 5420 18164 5464
rect 18736 5420 18836 5464
rect 19408 5420 19508 5464
rect 20080 5420 20180 5464
rect 20752 5420 20852 5464
rect 21648 5420 21748 5464
rect 22076 5420 22276 5464
rect 1692 5142 1892 5176
rect 1692 5096 1728 5142
rect 1868 5096 1892 5142
rect 1692 5079 1892 5096
rect 2160 5127 2260 5176
rect 2160 5090 2173 5127
rect 1692 5015 1892 5028
rect 1692 4969 1720 5015
rect 1860 4969 1892 5015
rect 1692 4936 1892 4969
rect 2140 4987 2173 5090
rect 2219 4987 2260 5127
rect 2832 5127 2932 5176
rect 2832 5090 2845 5127
rect 2140 4936 2260 4987
rect 2812 4987 2845 5090
rect 2891 4987 2932 5127
rect 3504 5127 3604 5176
rect 3504 5090 3517 5127
rect 2812 4936 2932 4987
rect 3484 4987 3517 5090
rect 3563 4987 3604 5127
rect 4176 5127 4276 5176
rect 4176 5090 4189 5127
rect 3484 4936 3604 4987
rect 4156 4987 4189 5090
rect 4235 4987 4276 5127
rect 4848 5127 4948 5176
rect 4848 5090 4861 5127
rect 4156 4936 4276 4987
rect 4828 4987 4861 5090
rect 4907 4987 4948 5127
rect 5744 5127 5844 5176
rect 5744 5090 5757 5127
rect 4828 4936 4948 4987
rect 5724 4987 5757 5090
rect 5803 4987 5844 5127
rect 6416 5127 6516 5176
rect 6416 5090 6429 5127
rect 5724 4936 5844 4987
rect 6396 4987 6429 5090
rect 6475 4987 6516 5127
rect 7088 5127 7188 5176
rect 7088 5090 7101 5127
rect 6396 4936 6516 4987
rect 7068 4987 7101 5090
rect 7147 4987 7188 5127
rect 7760 5127 7860 5176
rect 7760 5090 7773 5127
rect 7068 4936 7188 4987
rect 7740 4987 7773 5090
rect 7819 4987 7860 5127
rect 8432 5127 8532 5176
rect 8432 5090 8445 5127
rect 7740 4936 7860 4987
rect 8412 4987 8445 5090
rect 8491 4987 8532 5127
rect 9104 5127 9204 5176
rect 9104 5090 9117 5127
rect 8412 4936 8532 4987
rect 9084 4987 9117 5090
rect 9163 4987 9204 5127
rect 9776 5127 9876 5176
rect 9776 5090 9789 5127
rect 9084 4936 9204 4987
rect 9756 4987 9789 5090
rect 9835 4987 9876 5127
rect 10448 5127 10548 5176
rect 10448 5090 10461 5127
rect 9756 4936 9876 4987
rect 10428 4987 10461 5090
rect 10507 4987 10548 5127
rect 10876 5142 11076 5176
rect 10876 5096 10912 5142
rect 11052 5096 11076 5142
rect 10876 5079 11076 5096
rect 11456 5127 11556 5176
rect 11456 5090 11469 5127
rect 10428 4936 10548 4987
rect 10876 5015 11076 5028
rect 10876 4969 10904 5015
rect 11044 4969 11076 5015
rect 10876 4936 11076 4969
rect 11436 4987 11469 5090
rect 11515 4987 11556 5127
rect 12128 5127 12228 5176
rect 12128 5090 12141 5127
rect 11436 4936 11556 4987
rect 12108 4987 12141 5090
rect 12187 4987 12228 5127
rect 12800 5127 12900 5176
rect 12800 5090 12813 5127
rect 12108 4936 12228 4987
rect 12780 4987 12813 5090
rect 12859 4987 12900 5127
rect 13564 5142 13764 5176
rect 13564 5096 13600 5142
rect 13740 5096 13764 5142
rect 13564 5079 13764 5096
rect 14032 5127 14132 5176
rect 14032 5090 14045 5127
rect 12780 4936 12900 4987
rect 13564 5015 13764 5028
rect 13564 4969 13592 5015
rect 13732 4969 13764 5015
rect 1692 4728 1892 4772
rect 2140 4728 2260 4772
rect 2812 4728 2932 4772
rect 3484 4728 3604 4772
rect 4156 4728 4276 4772
rect 4828 4728 4948 4772
rect 13564 4936 13764 4969
rect 14012 4987 14045 5090
rect 14091 4987 14132 5127
rect 14704 5127 14804 5176
rect 14704 5090 14717 5127
rect 14012 4936 14132 4987
rect 14684 4987 14717 5090
rect 14763 4987 14804 5127
rect 15376 5127 15476 5176
rect 15376 5090 15389 5127
rect 14684 4936 14804 4987
rect 15356 4987 15389 5090
rect 15435 4987 15476 5127
rect 16048 5127 16148 5176
rect 16048 5090 16061 5127
rect 15356 4936 15476 4987
rect 16028 4987 16061 5090
rect 16107 4987 16148 5127
rect 16720 5127 16820 5176
rect 16720 5090 16733 5127
rect 16028 4936 16148 4987
rect 16700 4987 16733 5090
rect 16779 4987 16820 5127
rect 17392 5127 17492 5176
rect 17392 5090 17405 5127
rect 16700 4936 16820 4987
rect 17372 4987 17405 5090
rect 17451 4987 17492 5127
rect 18064 5127 18164 5176
rect 18064 5090 18077 5127
rect 17372 4936 17492 4987
rect 18044 4987 18077 5090
rect 18123 4987 18164 5127
rect 18736 5127 18836 5176
rect 18736 5090 18749 5127
rect 18044 4936 18164 4987
rect 18716 4987 18749 5090
rect 18795 4987 18836 5127
rect 19408 5127 19508 5176
rect 19408 5090 19421 5127
rect 18716 4936 18836 4987
rect 19388 4987 19421 5090
rect 19467 4987 19508 5127
rect 20080 5127 20180 5176
rect 20080 5090 20093 5127
rect 19388 4936 19508 4987
rect 20060 4987 20093 5090
rect 20139 4987 20180 5127
rect 20752 5127 20852 5176
rect 20752 5090 20765 5127
rect 20060 4936 20180 4987
rect 20732 4987 20765 5090
rect 20811 4987 20852 5127
rect 21648 5127 21748 5176
rect 21648 5090 21661 5127
rect 20732 4936 20852 4987
rect 21628 4987 21661 5090
rect 21707 4987 21748 5127
rect 22076 5142 22276 5176
rect 22076 5096 22112 5142
rect 22252 5096 22276 5142
rect 22076 5079 22276 5096
rect 5724 4728 5844 4772
rect 6396 4728 6516 4772
rect 7068 4728 7188 4772
rect 7740 4728 7860 4772
rect 8412 4728 8532 4772
rect 9084 4728 9204 4772
rect 9756 4728 9876 4772
rect 10428 4728 10548 4772
rect 10876 4728 11076 4772
rect 11436 4728 11556 4772
rect 12108 4728 12228 4772
rect 12780 4728 12900 4772
rect 21628 4936 21748 4987
rect 22076 5015 22276 5028
rect 22076 4969 22104 5015
rect 22244 4969 22276 5015
rect 22076 4936 22276 4969
rect 13564 4728 13764 4772
rect 14012 4728 14132 4772
rect 14684 4728 14804 4772
rect 15356 4728 15476 4772
rect 16028 4728 16148 4772
rect 16700 4728 16820 4772
rect 17372 4728 17492 4772
rect 18044 4728 18164 4772
rect 18716 4728 18836 4772
rect 19388 4728 19508 4772
rect 20060 4728 20180 4772
rect 20732 4728 20852 4772
rect 21628 4728 21748 4772
rect 22076 4728 22276 4772
rect 1692 4636 1892 4680
rect 2364 4636 2484 4680
rect 3036 4636 3156 4680
rect 3708 4636 3828 4680
rect 4380 4636 4500 4680
rect 5052 4636 5172 4680
rect 5724 4636 5844 4680
rect 6396 4636 6516 4680
rect 7068 4636 7188 4680
rect 7740 4636 7860 4680
rect 8412 4636 8532 4680
rect 8860 4636 9060 4680
rect 9756 4636 9876 4680
rect 10428 4636 10548 4680
rect 11100 4636 11220 4680
rect 11548 4636 11748 4680
rect 12332 4636 12452 4680
rect 13004 4636 13124 4680
rect 13676 4636 13796 4680
rect 14348 4636 14468 4680
rect 15020 4636 15140 4680
rect 15692 4636 15812 4680
rect 16364 4636 16484 4680
rect 16812 4636 17012 4680
rect 1692 4439 1892 4472
rect 1692 4393 1720 4439
rect 1860 4393 1892 4439
rect 1692 4380 1892 4393
rect 2364 4421 2484 4472
rect 1692 4312 1892 4329
rect 2364 4318 2397 4421
rect 1692 4266 1728 4312
rect 1868 4266 1892 4312
rect 1692 4232 1892 4266
rect 2384 4281 2397 4318
rect 2443 4281 2484 4421
rect 3036 4421 3156 4472
rect 3036 4318 3069 4421
rect 2384 4232 2484 4281
rect 3056 4281 3069 4318
rect 3115 4281 3156 4421
rect 3708 4421 3828 4472
rect 3708 4318 3741 4421
rect 3056 4232 3156 4281
rect 3728 4281 3741 4318
rect 3787 4281 3828 4421
rect 4380 4421 4500 4472
rect 4380 4318 4413 4421
rect 3728 4232 3828 4281
rect 4400 4281 4413 4318
rect 4459 4281 4500 4421
rect 5052 4421 5172 4472
rect 5052 4318 5085 4421
rect 4400 4232 4500 4281
rect 5072 4281 5085 4318
rect 5131 4281 5172 4421
rect 5724 4421 5844 4472
rect 5724 4318 5757 4421
rect 5072 4232 5172 4281
rect 5744 4281 5757 4318
rect 5803 4281 5844 4421
rect 6396 4421 6516 4472
rect 6396 4318 6429 4421
rect 5744 4232 5844 4281
rect 6416 4281 6429 4318
rect 6475 4281 6516 4421
rect 7068 4421 7188 4472
rect 7068 4318 7101 4421
rect 6416 4232 6516 4281
rect 7088 4281 7101 4318
rect 7147 4281 7188 4421
rect 7740 4421 7860 4472
rect 7740 4318 7773 4421
rect 7088 4232 7188 4281
rect 7760 4281 7773 4318
rect 7819 4281 7860 4421
rect 8412 4421 8532 4472
rect 8412 4318 8445 4421
rect 7760 4232 7860 4281
rect 8432 4281 8445 4318
rect 8491 4281 8532 4421
rect 8860 4439 9060 4472
rect 17708 4636 17828 4680
rect 18380 4636 18500 4680
rect 19052 4636 19172 4680
rect 19724 4636 19844 4680
rect 20396 4636 20516 4680
rect 21068 4636 21188 4680
rect 21820 4636 21940 4680
rect 8860 4393 8888 4439
rect 9028 4393 9060 4439
rect 8860 4380 9060 4393
rect 9756 4421 9876 4472
rect 8432 4232 8532 4281
rect 8860 4312 9060 4329
rect 8860 4266 8896 4312
rect 9036 4266 9060 4312
rect 8860 4232 9060 4266
rect 9756 4318 9789 4421
rect 9776 4281 9789 4318
rect 9835 4281 9876 4421
rect 10428 4421 10548 4472
rect 10428 4318 10461 4421
rect 9776 4232 9876 4281
rect 10448 4281 10461 4318
rect 10507 4281 10548 4421
rect 11100 4421 11220 4472
rect 11100 4318 11133 4421
rect 10448 4232 10548 4281
rect 11120 4281 11133 4318
rect 11179 4281 11220 4421
rect 11548 4439 11748 4472
rect 11548 4393 11576 4439
rect 11716 4393 11748 4439
rect 11548 4380 11748 4393
rect 12332 4421 12452 4472
rect 11120 4232 11220 4281
rect 11548 4312 11748 4329
rect 12332 4318 12365 4421
rect 11548 4266 11584 4312
rect 11724 4266 11748 4312
rect 11548 4232 11748 4266
rect 12352 4281 12365 4318
rect 12411 4281 12452 4421
rect 13004 4421 13124 4472
rect 13004 4318 13037 4421
rect 12352 4232 12452 4281
rect 13024 4281 13037 4318
rect 13083 4281 13124 4421
rect 13676 4421 13796 4472
rect 13676 4318 13709 4421
rect 13024 4232 13124 4281
rect 13696 4281 13709 4318
rect 13755 4281 13796 4421
rect 14348 4421 14468 4472
rect 14348 4318 14381 4421
rect 13696 4232 13796 4281
rect 14368 4281 14381 4318
rect 14427 4281 14468 4421
rect 15020 4421 15140 4472
rect 15020 4318 15053 4421
rect 14368 4232 14468 4281
rect 15040 4281 15053 4318
rect 15099 4281 15140 4421
rect 15692 4421 15812 4472
rect 15692 4318 15725 4421
rect 15040 4232 15140 4281
rect 15712 4281 15725 4318
rect 15771 4281 15812 4421
rect 16364 4421 16484 4472
rect 16364 4318 16397 4421
rect 15712 4232 15812 4281
rect 16384 4281 16397 4318
rect 16443 4281 16484 4421
rect 16812 4439 17012 4472
rect 16812 4393 16840 4439
rect 16980 4393 17012 4439
rect 16812 4380 17012 4393
rect 17708 4421 17828 4472
rect 16384 4232 16484 4281
rect 16812 4312 17012 4329
rect 16812 4266 16848 4312
rect 16988 4266 17012 4312
rect 16812 4232 17012 4266
rect 17708 4318 17741 4421
rect 17728 4281 17741 4318
rect 17787 4281 17828 4421
rect 18380 4421 18500 4472
rect 18380 4318 18413 4421
rect 17728 4232 17828 4281
rect 18400 4281 18413 4318
rect 18459 4281 18500 4421
rect 19052 4421 19172 4472
rect 19052 4318 19085 4421
rect 18400 4232 18500 4281
rect 19072 4281 19085 4318
rect 19131 4281 19172 4421
rect 19724 4421 19844 4472
rect 19724 4318 19757 4421
rect 19072 4232 19172 4281
rect 19744 4281 19757 4318
rect 19803 4281 19844 4421
rect 20396 4421 20516 4472
rect 20396 4318 20429 4421
rect 19744 4232 19844 4281
rect 20416 4281 20429 4318
rect 20475 4281 20516 4421
rect 21068 4421 21188 4472
rect 21068 4318 21101 4421
rect 20416 4232 20516 4281
rect 21088 4281 21101 4318
rect 21147 4281 21188 4421
rect 21088 4232 21188 4281
rect 21820 4421 21940 4472
rect 21820 4281 21861 4421
rect 21907 4318 21940 4421
rect 21907 4281 21920 4318
rect 21820 4232 21920 4281
rect 1692 3944 1892 3988
rect 2384 3944 2484 3988
rect 3056 3944 3156 3988
rect 3728 3944 3828 3988
rect 4400 3944 4500 3988
rect 5072 3944 5172 3988
rect 5744 3944 5844 3988
rect 6416 3944 6516 3988
rect 7088 3944 7188 3988
rect 7760 3944 7860 3988
rect 8432 3944 8532 3988
rect 8860 3944 9060 3988
rect 9776 3944 9876 3988
rect 10448 3944 10548 3988
rect 11120 3944 11220 3988
rect 11548 3944 11748 3988
rect 12352 3944 12452 3988
rect 13024 3944 13124 3988
rect 13696 3944 13796 3988
rect 14368 3944 14468 3988
rect 15040 3944 15140 3988
rect 15712 3944 15812 3988
rect 16384 3944 16484 3988
rect 16812 3944 17012 3988
rect 17728 3944 17828 3988
rect 18400 3944 18500 3988
rect 19072 3944 19172 3988
rect 19744 3944 19844 3988
rect 20416 3944 20516 3988
rect 21088 3944 21188 3988
rect 21820 3944 21920 3988
rect 1692 3852 1892 3896
rect 2140 3852 2340 3896
rect 2832 3852 2932 3896
rect 3504 3852 3604 3896
rect 4176 3852 4276 3896
rect 4848 3852 4948 3896
rect 5804 3852 5904 3896
rect 6476 3852 6576 3896
rect 7148 3852 7248 3896
rect 7760 3852 7860 3896
rect 8492 3852 8592 3896
rect 8860 3852 9060 3896
rect 9724 3852 9824 3896
rect 10336 3852 10436 3896
rect 11008 3852 11108 3896
rect 11740 3852 11840 3896
rect 12108 3852 12308 3896
rect 12556 3852 12756 3896
rect 13452 3852 13652 3896
rect 13920 3852 14020 3896
rect 14592 3852 14692 3896
rect 15264 3852 15364 3896
rect 15936 3852 16036 3896
rect 16608 3852 16708 3896
rect 17504 3852 17604 3896
rect 18176 3852 18276 3896
rect 18848 3852 18948 3896
rect 19520 3852 19620 3896
rect 20192 3852 20292 3896
rect 20620 3852 20820 3896
rect 21292 3852 21492 3896
rect 21740 3852 21940 3896
rect 1692 3574 1892 3608
rect 1692 3528 1728 3574
rect 1868 3528 1892 3574
rect 1692 3511 1892 3528
rect 2140 3574 2340 3608
rect 2140 3528 2176 3574
rect 2316 3528 2340 3574
rect 2140 3511 2340 3528
rect 2832 3559 2932 3608
rect 2832 3522 2845 3559
rect 1692 3447 1892 3460
rect 1692 3401 1720 3447
rect 1860 3401 1892 3447
rect 1692 3368 1892 3401
rect 2140 3447 2340 3460
rect 2140 3401 2168 3447
rect 2308 3401 2340 3447
rect 2140 3368 2340 3401
rect 2812 3419 2845 3522
rect 2891 3419 2932 3559
rect 3504 3559 3604 3608
rect 3504 3522 3517 3559
rect 2812 3368 2932 3419
rect 3484 3419 3517 3522
rect 3563 3419 3604 3559
rect 4176 3559 4276 3608
rect 4176 3522 4189 3559
rect 3484 3368 3604 3419
rect 4156 3419 4189 3522
rect 4235 3419 4276 3559
rect 4848 3559 4948 3608
rect 4848 3522 4861 3559
rect 4156 3368 4276 3419
rect 4828 3419 4861 3522
rect 4907 3419 4948 3559
rect 5804 3559 5904 3608
rect 4828 3368 4948 3419
rect 5804 3419 5845 3559
rect 5891 3522 5904 3559
rect 6476 3559 6576 3608
rect 5891 3419 5924 3522
rect 5804 3368 5924 3419
rect 6476 3419 6517 3559
rect 6563 3522 6576 3559
rect 7148 3559 7248 3608
rect 6563 3419 6596 3522
rect 6476 3368 6596 3419
rect 7148 3419 7189 3559
rect 7235 3522 7248 3559
rect 7760 3559 7860 3608
rect 7760 3522 7773 3559
rect 7235 3419 7268 3522
rect 7148 3368 7268 3419
rect 7740 3419 7773 3522
rect 7819 3419 7860 3559
rect 7740 3368 7860 3419
rect 8492 3559 8592 3608
rect 8492 3419 8533 3559
rect 8579 3522 8592 3559
rect 8860 3574 9060 3608
rect 8860 3528 8896 3574
rect 9036 3528 9060 3574
rect 8579 3419 8612 3522
rect 8860 3511 9060 3528
rect 9724 3559 9824 3608
rect 8492 3368 8612 3419
rect 8860 3447 9060 3460
rect 8860 3401 8888 3447
rect 9028 3401 9060 3447
rect 8860 3368 9060 3401
rect 9724 3419 9765 3559
rect 9811 3522 9824 3559
rect 10336 3559 10436 3608
rect 10336 3522 10349 3559
rect 9811 3419 9844 3522
rect 1692 3160 1892 3204
rect 2140 3160 2340 3204
rect 2812 3160 2932 3204
rect 3484 3160 3604 3204
rect 4156 3160 4276 3204
rect 4828 3160 4948 3204
rect 9724 3368 9844 3419
rect 10316 3419 10349 3522
rect 10395 3419 10436 3559
rect 11008 3559 11108 3608
rect 11008 3522 11021 3559
rect 10316 3368 10436 3419
rect 10988 3419 11021 3522
rect 11067 3419 11108 3559
rect 10988 3368 11108 3419
rect 11740 3559 11840 3608
rect 11740 3419 11781 3559
rect 11827 3522 11840 3559
rect 12108 3574 12308 3608
rect 12108 3528 12144 3574
rect 12284 3528 12308 3574
rect 11827 3419 11860 3522
rect 12108 3511 12308 3528
rect 12556 3574 12756 3608
rect 12556 3528 12592 3574
rect 12732 3528 12756 3574
rect 12556 3511 12756 3528
rect 13452 3574 13652 3608
rect 13452 3528 13488 3574
rect 13628 3528 13652 3574
rect 13452 3511 13652 3528
rect 13920 3559 14020 3608
rect 13920 3522 13933 3559
rect 11740 3368 11860 3419
rect 12108 3447 12308 3460
rect 12108 3401 12136 3447
rect 12276 3401 12308 3447
rect 12108 3368 12308 3401
rect 12556 3447 12756 3460
rect 12556 3401 12584 3447
rect 12724 3401 12756 3447
rect 12556 3368 12756 3401
rect 13452 3447 13652 3460
rect 13452 3401 13480 3447
rect 13620 3401 13652 3447
rect 5804 3160 5924 3204
rect 6476 3160 6596 3204
rect 7148 3160 7268 3204
rect 7740 3160 7860 3204
rect 8492 3160 8612 3204
rect 8860 3160 9060 3204
rect 13452 3368 13652 3401
rect 13900 3419 13933 3522
rect 13979 3419 14020 3559
rect 14592 3559 14692 3608
rect 14592 3522 14605 3559
rect 13900 3368 14020 3419
rect 14572 3419 14605 3522
rect 14651 3419 14692 3559
rect 15264 3559 15364 3608
rect 15264 3522 15277 3559
rect 14572 3368 14692 3419
rect 15244 3419 15277 3522
rect 15323 3419 15364 3559
rect 15936 3559 16036 3608
rect 15936 3522 15949 3559
rect 15244 3368 15364 3419
rect 15916 3419 15949 3522
rect 15995 3419 16036 3559
rect 16608 3559 16708 3608
rect 16608 3522 16621 3559
rect 15916 3368 16036 3419
rect 16588 3419 16621 3522
rect 16667 3419 16708 3559
rect 17504 3559 17604 3608
rect 17504 3522 17517 3559
rect 16588 3368 16708 3419
rect 17484 3419 17517 3522
rect 17563 3419 17604 3559
rect 18176 3559 18276 3608
rect 18176 3522 18189 3559
rect 9724 3160 9844 3204
rect 10316 3160 10436 3204
rect 10988 3160 11108 3204
rect 11740 3160 11860 3204
rect 12108 3160 12308 3204
rect 12556 3160 12756 3204
rect 17484 3368 17604 3419
rect 18156 3419 18189 3522
rect 18235 3419 18276 3559
rect 18848 3559 18948 3608
rect 18848 3522 18861 3559
rect 18156 3368 18276 3419
rect 18828 3419 18861 3522
rect 18907 3419 18948 3559
rect 19520 3559 19620 3608
rect 19520 3522 19533 3559
rect 18828 3368 18948 3419
rect 19500 3419 19533 3522
rect 19579 3419 19620 3559
rect 20192 3559 20292 3608
rect 20192 3522 20205 3559
rect 19500 3368 19620 3419
rect 20172 3419 20205 3522
rect 20251 3419 20292 3559
rect 20620 3574 20820 3608
rect 20620 3528 20656 3574
rect 20796 3528 20820 3574
rect 20620 3511 20820 3528
rect 21292 3574 21492 3608
rect 21292 3528 21328 3574
rect 21468 3528 21492 3574
rect 21292 3511 21492 3528
rect 21740 3574 21940 3608
rect 21740 3528 21776 3574
rect 21916 3528 21940 3574
rect 21740 3511 21940 3528
rect 20172 3368 20292 3419
rect 20620 3447 20820 3460
rect 20620 3401 20648 3447
rect 20788 3401 20820 3447
rect 20620 3368 20820 3401
rect 21292 3447 21492 3460
rect 21292 3401 21320 3447
rect 21460 3401 21492 3447
rect 13452 3160 13652 3204
rect 13900 3160 14020 3204
rect 14572 3160 14692 3204
rect 15244 3160 15364 3204
rect 15916 3160 16036 3204
rect 16588 3160 16708 3204
rect 21292 3368 21492 3401
rect 21740 3447 21940 3460
rect 21740 3401 21768 3447
rect 21908 3401 21940 3447
rect 21740 3368 21940 3401
rect 17484 3160 17604 3204
rect 18156 3160 18276 3204
rect 18828 3160 18948 3204
rect 19500 3160 19620 3204
rect 20172 3160 20292 3204
rect 20620 3160 20820 3204
rect 21292 3160 21492 3204
rect 21740 3160 21940 3204
<< polycontact >>
rect 1728 16072 1868 16118
rect 2176 16072 2316 16118
rect 2624 16072 2764 16118
rect 3072 16072 3212 16118
rect 3520 16072 3660 16118
rect 3968 16072 4108 16118
rect 4416 16072 4556 16118
rect 4864 16072 5004 16118
rect 5648 16072 5788 16118
rect 6096 16072 6236 16118
rect 6544 16072 6684 16118
rect 6992 16072 7132 16118
rect 7440 16072 7580 16118
rect 7888 16072 8028 16118
rect 8336 16072 8476 16118
rect 8784 16072 8924 16118
rect 9568 16072 9708 16118
rect 10016 16072 10156 16118
rect 10464 16072 10604 16118
rect 10912 16072 11052 16118
rect 11360 16072 11500 16118
rect 11808 16072 11948 16118
rect 12256 16072 12396 16118
rect 12704 16072 12844 16118
rect 13488 16072 13628 16118
rect 13936 16072 14076 16118
rect 14384 16072 14524 16118
rect 14832 16072 14972 16118
rect 15280 16072 15420 16118
rect 15728 16072 15868 16118
rect 16176 16072 16316 16118
rect 16624 16072 16764 16118
rect 17408 16072 17548 16118
rect 17856 16072 17996 16118
rect 18304 16072 18444 16118
rect 18752 16072 18892 16118
rect 19200 16072 19340 16118
rect 19648 16072 19788 16118
rect 20096 16072 20236 16118
rect 20544 16072 20684 16118
rect 21328 16072 21468 16118
rect 21776 16072 21916 16118
rect 1720 15945 1860 15991
rect 2168 15945 2308 15991
rect 2616 15945 2756 15991
rect 3064 15945 3204 15991
rect 3512 15945 3652 15991
rect 3960 15945 4100 15991
rect 4408 15945 4548 15991
rect 4856 15945 4996 15991
rect 5640 15945 5780 15991
rect 6088 15945 6228 15991
rect 6536 15945 6676 15991
rect 6984 15945 7124 15991
rect 7432 15945 7572 15991
rect 7880 15945 8020 15991
rect 8328 15945 8468 15991
rect 8776 15945 8916 15991
rect 9560 15945 9700 15991
rect 10008 15945 10148 15991
rect 10456 15945 10596 15991
rect 10904 15945 11044 15991
rect 11352 15945 11492 15991
rect 11800 15945 11940 15991
rect 12248 15945 12388 15991
rect 12696 15945 12836 15991
rect 13480 15945 13620 15991
rect 13928 15945 14068 15991
rect 14376 15945 14516 15991
rect 14824 15945 14964 15991
rect 15272 15945 15412 15991
rect 15720 15945 15860 15991
rect 16168 15945 16308 15991
rect 16616 15945 16756 15991
rect 17400 15945 17540 15991
rect 17848 15945 17988 15991
rect 18296 15945 18436 15991
rect 18744 15945 18884 15991
rect 19192 15945 19332 15991
rect 19640 15945 19780 15991
rect 20088 15945 20228 15991
rect 20536 15945 20676 15991
rect 21320 15945 21460 15991
rect 21768 15945 21908 15991
rect 1720 15369 1860 15415
rect 2168 15369 2308 15415
rect 2616 15369 2756 15415
rect 3064 15369 3204 15415
rect 3512 15369 3652 15415
rect 3960 15369 4100 15415
rect 4408 15369 4548 15415
rect 4856 15369 4996 15415
rect 5304 15369 5444 15415
rect 5752 15369 5892 15415
rect 6200 15369 6340 15415
rect 6648 15369 6788 15415
rect 7096 15369 7236 15415
rect 7544 15369 7684 15415
rect 7992 15369 8132 15415
rect 8440 15369 8580 15415
rect 8888 15369 9028 15415
rect 9672 15369 9812 15415
rect 10120 15369 10260 15415
rect 10568 15369 10708 15415
rect 11016 15369 11156 15415
rect 11464 15369 11604 15415
rect 11912 15369 12052 15415
rect 12360 15369 12500 15415
rect 12808 15369 12948 15415
rect 13256 15369 13396 15415
rect 13704 15369 13844 15415
rect 14152 15369 14292 15415
rect 14600 15369 14740 15415
rect 15048 15369 15188 15415
rect 15496 15369 15636 15415
rect 15944 15369 16084 15415
rect 16392 15369 16532 15415
rect 16840 15369 16980 15415
rect 17624 15369 17764 15415
rect 18072 15369 18212 15415
rect 18520 15369 18660 15415
rect 18968 15369 19108 15415
rect 19416 15369 19556 15415
rect 19864 15369 20004 15415
rect 20312 15369 20452 15415
rect 20760 15369 20900 15415
rect 21208 15369 21348 15415
rect 21656 15369 21796 15415
rect 22104 15369 22244 15415
rect 1728 15242 1868 15288
rect 2176 15242 2316 15288
rect 2624 15242 2764 15288
rect 3072 15242 3212 15288
rect 3520 15242 3660 15288
rect 3968 15242 4108 15288
rect 4416 15242 4556 15288
rect 4864 15242 5004 15288
rect 5312 15242 5452 15288
rect 5760 15242 5900 15288
rect 6208 15242 6348 15288
rect 6656 15242 6796 15288
rect 7104 15242 7244 15288
rect 7552 15242 7692 15288
rect 8000 15242 8140 15288
rect 8448 15242 8588 15288
rect 8896 15242 9036 15288
rect 9680 15242 9820 15288
rect 10128 15242 10268 15288
rect 10576 15242 10716 15288
rect 11024 15242 11164 15288
rect 11472 15242 11612 15288
rect 11920 15242 12060 15288
rect 12368 15242 12508 15288
rect 12816 15242 12956 15288
rect 13264 15242 13404 15288
rect 13712 15242 13852 15288
rect 14160 15242 14300 15288
rect 14608 15242 14748 15288
rect 15056 15242 15196 15288
rect 15504 15242 15644 15288
rect 15952 15242 16092 15288
rect 16400 15242 16540 15288
rect 16848 15242 16988 15288
rect 17632 15242 17772 15288
rect 18080 15242 18220 15288
rect 18528 15242 18668 15288
rect 18976 15242 19116 15288
rect 19424 15242 19564 15288
rect 19872 15242 20012 15288
rect 20320 15242 20460 15288
rect 20768 15242 20908 15288
rect 21216 15242 21356 15288
rect 21664 15242 21804 15288
rect 22112 15242 22252 15288
rect 1728 14504 1868 14550
rect 2176 14504 2316 14550
rect 2624 14504 2764 14550
rect 3072 14504 3212 14550
rect 3520 14504 3660 14550
rect 3968 14504 4108 14550
rect 4416 14504 4556 14550
rect 4864 14504 5004 14550
rect 5648 14504 5788 14550
rect 6096 14504 6236 14550
rect 6544 14504 6684 14550
rect 6992 14504 7132 14550
rect 7440 14504 7580 14550
rect 7888 14504 8028 14550
rect 8336 14504 8476 14550
rect 8784 14504 8924 14550
rect 9232 14504 9372 14550
rect 9680 14504 9820 14550
rect 10128 14504 10268 14550
rect 10576 14504 10716 14550
rect 11024 14504 11164 14550
rect 11472 14504 11612 14550
rect 11920 14504 12060 14550
rect 12368 14504 12508 14550
rect 12816 14504 12956 14550
rect 13600 14504 13740 14550
rect 14048 14504 14188 14550
rect 14496 14504 14636 14550
rect 14944 14504 15084 14550
rect 15392 14504 15532 14550
rect 15840 14504 15980 14550
rect 16288 14504 16428 14550
rect 1720 14377 1860 14423
rect 2168 14377 2308 14423
rect 2616 14377 2756 14423
rect 3064 14377 3204 14423
rect 3512 14377 3652 14423
rect 3960 14377 4100 14423
rect 4408 14377 4548 14423
rect 4856 14377 4996 14423
rect 5640 14377 5780 14423
rect 6088 14377 6228 14423
rect 6536 14377 6676 14423
rect 6984 14377 7124 14423
rect 7432 14377 7572 14423
rect 7880 14377 8020 14423
rect 8328 14377 8468 14423
rect 8776 14377 8916 14423
rect 9224 14377 9364 14423
rect 9672 14377 9812 14423
rect 10120 14377 10260 14423
rect 10568 14377 10708 14423
rect 11016 14377 11156 14423
rect 11464 14377 11604 14423
rect 11912 14377 12052 14423
rect 12360 14377 12500 14423
rect 12808 14377 12948 14423
rect 13592 14377 13732 14423
rect 14040 14377 14180 14423
rect 14488 14377 14628 14423
rect 14936 14377 15076 14423
rect 15384 14377 15524 14423
rect 15832 14377 15972 14423
rect 16280 14377 16420 14423
rect 16933 14395 16979 14535
rect 17605 14395 17651 14535
rect 17968 14504 18108 14550
rect 18416 14504 18556 14550
rect 18864 14504 19004 14550
rect 19312 14504 19452 14550
rect 19760 14504 19900 14550
rect 20208 14504 20348 14550
rect 20656 14504 20796 14550
rect 21552 14504 21692 14550
rect 22000 14504 22140 14550
rect 17960 14377 18100 14423
rect 18408 14377 18548 14423
rect 18856 14377 18996 14423
rect 19304 14377 19444 14423
rect 19752 14377 19892 14423
rect 20200 14377 20340 14423
rect 20648 14377 20788 14423
rect 21544 14377 21684 14423
rect 21992 14377 22132 14423
rect 1720 13801 1860 13847
rect 2168 13801 2308 13847
rect 2616 13801 2756 13847
rect 3064 13801 3204 13847
rect 3512 13801 3652 13847
rect 3960 13801 4100 13847
rect 4408 13801 4548 13847
rect 4856 13801 4996 13847
rect 5304 13801 5444 13847
rect 5752 13801 5892 13847
rect 6200 13801 6340 13847
rect 6648 13801 6788 13847
rect 7096 13801 7236 13847
rect 7544 13801 7684 13847
rect 7992 13801 8132 13847
rect 8440 13801 8580 13847
rect 8888 13801 9028 13847
rect 9672 13801 9812 13847
rect 10120 13801 10260 13847
rect 10568 13801 10708 13847
rect 11016 13801 11156 13847
rect 11464 13801 11604 13847
rect 11912 13801 12052 13847
rect 12360 13801 12500 13847
rect 12808 13801 12948 13847
rect 13256 13801 13396 13847
rect 13704 13801 13844 13847
rect 14152 13801 14292 13847
rect 14600 13801 14740 13847
rect 15048 13801 15188 13847
rect 15496 13801 15636 13847
rect 1728 13674 1868 13720
rect 2176 13674 2316 13720
rect 2624 13674 2764 13720
rect 3072 13674 3212 13720
rect 3520 13674 3660 13720
rect 3968 13674 4108 13720
rect 4416 13674 4556 13720
rect 4864 13674 5004 13720
rect 5312 13674 5452 13720
rect 5760 13674 5900 13720
rect 6208 13674 6348 13720
rect 6656 13674 6796 13720
rect 7104 13674 7244 13720
rect 7552 13674 7692 13720
rect 8000 13674 8140 13720
rect 8448 13674 8588 13720
rect 8896 13674 9036 13720
rect 9680 13674 9820 13720
rect 10128 13674 10268 13720
rect 10576 13674 10716 13720
rect 11024 13674 11164 13720
rect 11472 13674 11612 13720
rect 11920 13674 12060 13720
rect 12368 13674 12508 13720
rect 12816 13674 12956 13720
rect 13264 13674 13404 13720
rect 13712 13674 13852 13720
rect 14160 13674 14300 13720
rect 14608 13674 14748 13720
rect 15056 13674 15196 13720
rect 15504 13674 15644 13720
rect 16173 13689 16219 13829
rect 16845 13689 16891 13829
rect 17741 13689 17787 13829
rect 18413 13689 18459 13829
rect 18856 13801 18996 13847
rect 19304 13801 19444 13847
rect 19752 13801 19892 13847
rect 20200 13801 20340 13847
rect 20648 13801 20788 13847
rect 21096 13801 21236 13847
rect 21544 13801 21684 13847
rect 21992 13801 22132 13847
rect 18864 13674 19004 13720
rect 19312 13674 19452 13720
rect 19760 13674 19900 13720
rect 20208 13674 20348 13720
rect 20656 13674 20796 13720
rect 21104 13674 21244 13720
rect 21552 13674 21692 13720
rect 22000 13674 22140 13720
rect 1728 12936 1868 12982
rect 2176 12936 2316 12982
rect 2624 12936 2764 12982
rect 3072 12936 3212 12982
rect 3520 12936 3660 12982
rect 3968 12936 4108 12982
rect 4416 12936 4556 12982
rect 4864 12936 5004 12982
rect 5648 12936 5788 12982
rect 6096 12936 6236 12982
rect 6544 12936 6684 12982
rect 6992 12936 7132 12982
rect 7440 12936 7580 12982
rect 7888 12936 8028 12982
rect 8336 12936 8476 12982
rect 8784 12936 8924 12982
rect 9232 12936 9372 12982
rect 9680 12936 9820 12982
rect 10128 12936 10268 12982
rect 10576 12936 10716 12982
rect 11024 12936 11164 12982
rect 11472 12936 11612 12982
rect 11920 12936 12060 12982
rect 12368 12936 12508 12982
rect 12816 12936 12956 12982
rect 13600 12936 13740 12982
rect 14048 12936 14188 12982
rect 1720 12809 1860 12855
rect 2168 12809 2308 12855
rect 2616 12809 2756 12855
rect 3064 12809 3204 12855
rect 3512 12809 3652 12855
rect 3960 12809 4100 12855
rect 4408 12809 4548 12855
rect 4856 12809 4996 12855
rect 5640 12809 5780 12855
rect 6088 12809 6228 12855
rect 6536 12809 6676 12855
rect 6984 12809 7124 12855
rect 7432 12809 7572 12855
rect 7880 12809 8020 12855
rect 8328 12809 8468 12855
rect 8776 12809 8916 12855
rect 9224 12809 9364 12855
rect 9672 12809 9812 12855
rect 10120 12809 10260 12855
rect 10568 12809 10708 12855
rect 11016 12809 11156 12855
rect 11464 12809 11604 12855
rect 11912 12809 12052 12855
rect 12360 12809 12500 12855
rect 12808 12809 12948 12855
rect 13592 12809 13732 12855
rect 14040 12809 14180 12855
rect 14829 12827 14875 12967
rect 15501 12827 15547 12967
rect 16173 12827 16219 12967
rect 16845 12827 16891 12967
rect 17517 12827 17563 12967
rect 18189 12827 18235 12967
rect 18861 12827 18907 12967
rect 19533 12827 19579 12967
rect 19984 12936 20124 12982
rect 20432 12936 20572 12982
rect 20880 12936 21020 12982
rect 21552 12936 21692 12982
rect 22000 12936 22140 12982
rect 19976 12809 20116 12855
rect 20424 12809 20564 12855
rect 20872 12809 21012 12855
rect 21544 12809 21684 12855
rect 21992 12809 22132 12855
rect 1720 12233 1860 12279
rect 2168 12233 2308 12279
rect 2616 12233 2756 12279
rect 3064 12233 3204 12279
rect 3512 12233 3652 12279
rect 3960 12233 4100 12279
rect 4408 12233 4548 12279
rect 4856 12233 4996 12279
rect 5304 12233 5444 12279
rect 5752 12233 5892 12279
rect 6200 12233 6340 12279
rect 6648 12233 6788 12279
rect 7096 12233 7236 12279
rect 7544 12233 7684 12279
rect 7992 12233 8132 12279
rect 8440 12233 8580 12279
rect 8888 12233 9028 12279
rect 9672 12233 9812 12279
rect 10120 12233 10260 12279
rect 10568 12233 10708 12279
rect 11016 12233 11156 12279
rect 11464 12233 11604 12279
rect 11912 12233 12052 12279
rect 12360 12233 12500 12279
rect 12808 12233 12948 12279
rect 13256 12233 13396 12279
rect 13704 12233 13844 12279
rect 1728 12106 1868 12152
rect 2176 12106 2316 12152
rect 2624 12106 2764 12152
rect 3072 12106 3212 12152
rect 3520 12106 3660 12152
rect 3968 12106 4108 12152
rect 4416 12106 4556 12152
rect 4864 12106 5004 12152
rect 5312 12106 5452 12152
rect 5760 12106 5900 12152
rect 6208 12106 6348 12152
rect 6656 12106 6796 12152
rect 7104 12106 7244 12152
rect 7552 12106 7692 12152
rect 8000 12106 8140 12152
rect 8448 12106 8588 12152
rect 8896 12106 9036 12152
rect 9680 12106 9820 12152
rect 10128 12106 10268 12152
rect 10576 12106 10716 12152
rect 11024 12106 11164 12152
rect 11472 12106 11612 12152
rect 11920 12106 12060 12152
rect 12368 12106 12508 12152
rect 12816 12106 12956 12152
rect 13264 12106 13404 12152
rect 13712 12106 13852 12152
rect 14157 12121 14203 12261
rect 14829 12121 14875 12261
rect 15501 12121 15547 12261
rect 16173 12121 16219 12261
rect 16845 12121 16891 12261
rect 17741 12121 17787 12261
rect 18413 12121 18459 12261
rect 19085 12121 19131 12261
rect 19757 12121 19803 12261
rect 20429 12121 20475 12261
rect 20872 12233 21012 12279
rect 21320 12233 21460 12279
rect 21768 12233 21908 12279
rect 20880 12106 21020 12152
rect 21328 12106 21468 12152
rect 21776 12106 21916 12152
rect 1728 11368 1868 11414
rect 2176 11368 2316 11414
rect 2624 11368 2764 11414
rect 3072 11368 3212 11414
rect 3520 11368 3660 11414
rect 3968 11368 4108 11414
rect 4416 11368 4556 11414
rect 4864 11368 5004 11414
rect 5648 11368 5788 11414
rect 1720 11241 1860 11287
rect 2168 11241 2308 11287
rect 2616 11241 2756 11287
rect 3064 11241 3204 11287
rect 3512 11241 3652 11287
rect 3960 11241 4100 11287
rect 4408 11241 4548 11287
rect 4856 11241 4996 11287
rect 5640 11241 5780 11287
rect 6181 11259 6227 11399
rect 6965 11259 7011 11399
rect 7637 11259 7683 11399
rect 8309 11259 8355 11399
rect 8672 11368 8812 11414
rect 8664 11241 8804 11287
rect 9229 11259 9275 11399
rect 9901 11259 9947 11399
rect 10573 11259 10619 11399
rect 11024 11368 11164 11414
rect 11472 11368 11612 11414
rect 11016 11241 11156 11287
rect 11464 11241 11604 11287
rect 12141 11259 12187 11399
rect 12813 11259 12859 11399
rect 13709 11259 13755 11399
rect 14160 11368 14300 11414
rect 14152 11241 14292 11287
rect 14829 11259 14875 11399
rect 15501 11259 15547 11399
rect 16173 11259 16219 11399
rect 16845 11259 16891 11399
rect 17517 11259 17563 11399
rect 18189 11259 18235 11399
rect 18861 11259 18907 11399
rect 19533 11259 19579 11399
rect 20205 11259 20251 11399
rect 20656 11368 20796 11414
rect 21552 11368 21692 11414
rect 22000 11368 22140 11414
rect 20648 11241 20788 11287
rect 21544 11241 21684 11287
rect 21992 11241 22132 11287
rect 1720 10665 1860 10711
rect 2168 10665 2308 10711
rect 2616 10665 2756 10711
rect 3064 10665 3204 10711
rect 3512 10665 3652 10711
rect 3960 10665 4100 10711
rect 4408 10665 4548 10711
rect 4856 10665 4996 10711
rect 1728 10538 1868 10584
rect 2176 10538 2316 10584
rect 2624 10538 2764 10584
rect 3072 10538 3212 10584
rect 3520 10538 3660 10584
rect 3968 10538 4108 10584
rect 4416 10538 4556 10584
rect 4864 10538 5004 10584
rect 5421 10553 5467 10693
rect 6093 10553 6139 10693
rect 6765 10553 6811 10693
rect 7437 10553 7483 10693
rect 8109 10553 8155 10693
rect 8893 10553 8939 10693
rect 9901 10553 9947 10693
rect 10573 10553 10619 10693
rect 11245 10553 11291 10693
rect 12029 10553 12075 10693
rect 12701 10553 12747 10693
rect 13373 10553 13419 10693
rect 14045 10553 14091 10693
rect 14717 10553 14763 10693
rect 15389 10553 15435 10693
rect 16061 10553 16107 10693
rect 16733 10553 16779 10693
rect 17741 10553 17787 10693
rect 18413 10553 18459 10693
rect 19085 10553 19131 10693
rect 19757 10553 19803 10693
rect 20429 10553 20475 10693
rect 21101 10553 21147 10693
rect 21773 10553 21819 10693
rect 1728 9800 1868 9846
rect 2176 9800 2316 9846
rect 2624 9800 2764 9846
rect 3072 9800 3212 9846
rect 3520 9800 3660 9846
rect 1720 9673 1860 9719
rect 2168 9673 2308 9719
rect 2616 9673 2756 9719
rect 3064 9673 3204 9719
rect 3512 9673 3652 9719
rect 4189 9691 4235 9831
rect 4861 9691 4907 9831
rect 5869 9691 5915 9831
rect 6541 9691 6587 9831
rect 7213 9691 7259 9831
rect 7885 9691 7931 9831
rect 8557 9691 8603 9831
rect 9229 9691 9275 9831
rect 9901 9691 9947 9831
rect 10573 9691 10619 9831
rect 11024 9800 11164 9846
rect 11016 9673 11156 9719
rect 11469 9691 11515 9831
rect 12141 9691 12187 9831
rect 12813 9691 12859 9831
rect 13709 9691 13755 9831
rect 14381 9691 14427 9831
rect 15053 9691 15099 9831
rect 15725 9691 15771 9831
rect 16397 9691 16443 9831
rect 17069 9691 17115 9831
rect 17829 9691 17875 9831
rect 18413 9691 18459 9831
rect 19085 9691 19131 9831
rect 19757 9691 19803 9831
rect 20429 9691 20475 9831
rect 20880 9800 21020 9846
rect 20872 9673 21012 9719
rect 21661 9691 21707 9831
rect 22112 9800 22252 9846
rect 22104 9673 22244 9719
rect 1720 9097 1860 9143
rect 2168 9097 2308 9143
rect 2616 9097 2756 9143
rect 1728 8970 1868 9016
rect 2176 8970 2316 9016
rect 2624 8970 2764 9016
rect 3405 8985 3451 9125
rect 4077 8985 4123 9125
rect 4749 8985 4795 9125
rect 5421 8985 5467 9125
rect 6093 8985 6139 9125
rect 6765 8985 6811 9125
rect 7437 8985 7483 9125
rect 8221 8985 8267 9125
rect 8893 8985 8939 9125
rect 9672 9097 9812 9143
rect 9680 8970 9820 9016
rect 10349 8985 10395 9125
rect 11021 8985 11067 9125
rect 11693 8985 11739 9125
rect 12365 8985 12411 9125
rect 13037 8985 13083 9125
rect 13709 8985 13755 9125
rect 14381 8985 14427 9125
rect 15053 8985 15099 9125
rect 15725 8985 15771 9125
rect 16397 8985 16443 9125
rect 16840 9097 16980 9143
rect 16848 8970 16988 9016
rect 17741 8985 17787 9125
rect 18413 8985 18459 9125
rect 19085 8985 19131 9125
rect 19757 8985 19803 9125
rect 20429 8985 20475 9125
rect 20872 9097 21012 9143
rect 21320 9097 21460 9143
rect 21768 9097 21908 9143
rect 20880 8970 21020 9016
rect 21328 8970 21468 9016
rect 21776 8970 21916 9016
rect 1728 8232 1868 8278
rect 2176 8232 2316 8278
rect 1720 8105 1860 8151
rect 2168 8105 2308 8151
rect 2933 8123 2979 8263
rect 3517 8123 3563 8263
rect 4189 8123 4235 8263
rect 4861 8123 4907 8263
rect 5869 8123 5915 8263
rect 6541 8123 6587 8263
rect 7213 8123 7259 8263
rect 7885 8123 7931 8263
rect 8557 8123 8603 8263
rect 9229 8123 9275 8263
rect 9901 8123 9947 8263
rect 10573 8123 10619 8263
rect 11333 8123 11379 8263
rect 11696 8232 11836 8278
rect 11688 8105 11828 8151
rect 12141 8123 12187 8263
rect 12813 8123 12859 8263
rect 13709 8123 13755 8263
rect 14381 8123 14427 8263
rect 15053 8123 15099 8263
rect 15725 8123 15771 8263
rect 16397 8123 16443 8263
rect 17069 8123 17115 8263
rect 17741 8123 17787 8263
rect 18413 8123 18459 8263
rect 19085 8123 19131 8263
rect 19757 8123 19803 8263
rect 20517 8123 20563 8263
rect 20880 8232 21020 8278
rect 21552 8232 21692 8278
rect 22000 8232 22140 8278
rect 20872 8105 21012 8151
rect 21544 8105 21684 8151
rect 21992 8105 22132 8151
rect 2149 7417 2195 7557
rect 2733 7417 2779 7557
rect 3405 7417 3451 7557
rect 4077 7417 4123 7557
rect 4749 7417 4795 7557
rect 5421 7417 5467 7557
rect 6093 7417 6139 7557
rect 6765 7417 6811 7557
rect 7437 7417 7483 7557
rect 8221 7417 8267 7557
rect 8893 7417 8939 7557
rect 9901 7417 9947 7557
rect 10573 7417 10619 7557
rect 11333 7417 11379 7557
rect 11917 7417 11963 7557
rect 12589 7417 12635 7557
rect 13261 7417 13307 7557
rect 13933 7417 13979 7557
rect 14605 7417 14651 7557
rect 15277 7417 15323 7557
rect 15949 7417 15995 7557
rect 16621 7417 16667 7557
rect 17741 7417 17787 7557
rect 18413 7417 18459 7557
rect 19085 7417 19131 7557
rect 19757 7417 19803 7557
rect 20429 7417 20475 7557
rect 21101 7417 21147 7557
rect 21544 7529 21684 7575
rect 21992 7529 22132 7575
rect 21552 7402 21692 7448
rect 22000 7402 22140 7448
rect 1728 6664 1868 6710
rect 1720 6537 1860 6583
rect 2173 6555 2219 6695
rect 2845 6555 2891 6695
rect 3517 6555 3563 6695
rect 4189 6555 4235 6695
rect 4861 6555 4907 6695
rect 5757 6555 5803 6695
rect 6429 6555 6475 6695
rect 7101 6555 7147 6695
rect 7773 6555 7819 6695
rect 8445 6555 8491 6695
rect 9117 6555 9163 6695
rect 9789 6555 9835 6695
rect 10461 6555 10507 6695
rect 11133 6555 11179 6695
rect 11805 6555 11851 6695
rect 12477 6555 12523 6695
rect 12928 6664 13068 6710
rect 13600 6664 13740 6710
rect 12920 6537 13060 6583
rect 13592 6537 13732 6583
rect 14157 6555 14203 6695
rect 14829 6555 14875 6695
rect 15501 6555 15547 6695
rect 16173 6555 16219 6695
rect 16845 6555 16891 6695
rect 17517 6555 17563 6695
rect 18189 6555 18235 6695
rect 18861 6555 18907 6695
rect 19533 6555 19579 6695
rect 20293 6555 20339 6695
rect 20656 6664 20796 6710
rect 20648 6537 20788 6583
rect 21661 6555 21707 6695
rect 22112 6664 22252 6710
rect 22104 6537 22244 6583
rect 2061 5849 2107 5989
rect 2733 5849 2779 5989
rect 3405 5849 3451 5989
rect 4077 5849 4123 5989
rect 4749 5849 4795 5989
rect 5421 5849 5467 5989
rect 6093 5849 6139 5989
rect 6765 5849 6811 5989
rect 7437 5849 7483 5989
rect 8109 5849 8155 5989
rect 8781 5849 8827 5989
rect 9789 5849 9835 5989
rect 10461 5849 10507 5989
rect 11133 5849 11179 5989
rect 11805 5849 11851 5989
rect 12589 5849 12635 5989
rect 13261 5849 13307 5989
rect 13933 5849 13979 5989
rect 14605 5849 14651 5989
rect 15277 5849 15323 5989
rect 15949 5849 15995 5989
rect 16621 5849 16667 5989
rect 17741 5849 17787 5989
rect 18413 5849 18459 5989
rect 19085 5849 19131 5989
rect 19757 5849 19803 5989
rect 20429 5849 20475 5989
rect 21101 5849 21147 5989
rect 21861 5849 21907 5989
rect 1728 5096 1868 5142
rect 1720 4969 1860 5015
rect 2173 4987 2219 5127
rect 2845 4987 2891 5127
rect 3517 4987 3563 5127
rect 4189 4987 4235 5127
rect 4861 4987 4907 5127
rect 5757 4987 5803 5127
rect 6429 4987 6475 5127
rect 7101 4987 7147 5127
rect 7773 4987 7819 5127
rect 8445 4987 8491 5127
rect 9117 4987 9163 5127
rect 9789 4987 9835 5127
rect 10461 4987 10507 5127
rect 10912 5096 11052 5142
rect 10904 4969 11044 5015
rect 11469 4987 11515 5127
rect 12141 4987 12187 5127
rect 12813 4987 12859 5127
rect 13600 5096 13740 5142
rect 13592 4969 13732 5015
rect 14045 4987 14091 5127
rect 14717 4987 14763 5127
rect 15389 4987 15435 5127
rect 16061 4987 16107 5127
rect 16733 4987 16779 5127
rect 17405 4987 17451 5127
rect 18077 4987 18123 5127
rect 18749 4987 18795 5127
rect 19421 4987 19467 5127
rect 20093 4987 20139 5127
rect 20765 4987 20811 5127
rect 21661 4987 21707 5127
rect 22112 5096 22252 5142
rect 22104 4969 22244 5015
rect 1720 4393 1860 4439
rect 1728 4266 1868 4312
rect 2397 4281 2443 4421
rect 3069 4281 3115 4421
rect 3741 4281 3787 4421
rect 4413 4281 4459 4421
rect 5085 4281 5131 4421
rect 5757 4281 5803 4421
rect 6429 4281 6475 4421
rect 7101 4281 7147 4421
rect 7773 4281 7819 4421
rect 8445 4281 8491 4421
rect 8888 4393 9028 4439
rect 8896 4266 9036 4312
rect 9789 4281 9835 4421
rect 10461 4281 10507 4421
rect 11133 4281 11179 4421
rect 11576 4393 11716 4439
rect 11584 4266 11724 4312
rect 12365 4281 12411 4421
rect 13037 4281 13083 4421
rect 13709 4281 13755 4421
rect 14381 4281 14427 4421
rect 15053 4281 15099 4421
rect 15725 4281 15771 4421
rect 16397 4281 16443 4421
rect 16840 4393 16980 4439
rect 16848 4266 16988 4312
rect 17741 4281 17787 4421
rect 18413 4281 18459 4421
rect 19085 4281 19131 4421
rect 19757 4281 19803 4421
rect 20429 4281 20475 4421
rect 21101 4281 21147 4421
rect 21861 4281 21907 4421
rect 1728 3528 1868 3574
rect 2176 3528 2316 3574
rect 1720 3401 1860 3447
rect 2168 3401 2308 3447
rect 2845 3419 2891 3559
rect 3517 3419 3563 3559
rect 4189 3419 4235 3559
rect 4861 3419 4907 3559
rect 5845 3419 5891 3559
rect 6517 3419 6563 3559
rect 7189 3419 7235 3559
rect 7773 3419 7819 3559
rect 8533 3419 8579 3559
rect 8896 3528 9036 3574
rect 8888 3401 9028 3447
rect 9765 3419 9811 3559
rect 10349 3419 10395 3559
rect 11021 3419 11067 3559
rect 11781 3419 11827 3559
rect 12144 3528 12284 3574
rect 12592 3528 12732 3574
rect 13488 3528 13628 3574
rect 12136 3401 12276 3447
rect 12584 3401 12724 3447
rect 13480 3401 13620 3447
rect 13933 3419 13979 3559
rect 14605 3419 14651 3559
rect 15277 3419 15323 3559
rect 15949 3419 15995 3559
rect 16621 3419 16667 3559
rect 17517 3419 17563 3559
rect 18189 3419 18235 3559
rect 18861 3419 18907 3559
rect 19533 3419 19579 3559
rect 20205 3419 20251 3559
rect 20656 3528 20796 3574
rect 21328 3528 21468 3574
rect 21776 3528 21916 3574
rect 20648 3401 20788 3447
rect 21320 3401 21460 3447
rect 21768 3401 21908 3447
<< metal1 >>
rect 1344 16490 22624 16524
rect 1344 16438 3874 16490
rect 4134 16438 9194 16490
rect 9454 16438 14514 16490
rect 14774 16438 19834 16490
rect 20094 16438 22624 16490
rect 1344 16404 22624 16438
rect 1418 16379 1486 16404
rect 1418 16333 1429 16379
rect 1475 16333 1486 16379
rect 1418 16251 1486 16333
rect 1418 16205 1429 16251
rect 1475 16205 1486 16251
rect 1418 16123 1486 16205
rect 1418 16077 1429 16123
rect 1475 16077 1486 16123
rect 1418 16064 1486 16077
rect 1617 16337 1663 16358
rect 1617 15991 1663 16197
rect 1921 16337 1967 16404
rect 1921 16178 1967 16197
rect 2065 16337 2111 16358
rect 1714 16072 1728 16118
rect 1868 16072 1967 16118
rect 1617 15945 1720 15991
rect 1860 15945 1872 15991
rect 1418 15906 1486 15918
rect 1418 15759 1429 15906
rect 1475 15759 1486 15906
rect 1418 15740 1486 15759
rect 1617 15872 1663 15889
rect 1617 15740 1663 15826
rect 1921 15872 1967 16072
rect 2065 15991 2111 16197
rect 2369 16337 2415 16404
rect 2369 16178 2415 16197
rect 2513 16337 2559 16358
rect 2162 16072 2176 16118
rect 2316 16072 2415 16118
rect 2065 15945 2168 15991
rect 2308 15945 2320 15991
rect 1921 15786 1967 15826
rect 2065 15872 2111 15889
rect 2065 15740 2111 15826
rect 2369 15872 2415 16072
rect 2513 15991 2559 16197
rect 2817 16337 2863 16404
rect 2817 16178 2863 16197
rect 2961 16337 3007 16358
rect 2610 16072 2624 16118
rect 2764 16072 2863 16118
rect 2513 15945 2616 15991
rect 2756 15945 2768 15991
rect 2369 15786 2415 15826
rect 2513 15872 2559 15889
rect 2513 15740 2559 15826
rect 2817 15872 2863 16072
rect 2961 15991 3007 16197
rect 3265 16337 3311 16404
rect 3265 16178 3311 16197
rect 3409 16337 3455 16358
rect 3058 16072 3072 16118
rect 3212 16072 3311 16118
rect 2961 15945 3064 15991
rect 3204 15945 3216 15991
rect 2817 15786 2863 15826
rect 2961 15872 3007 15889
rect 2961 15740 3007 15826
rect 3265 15872 3311 16072
rect 3409 15991 3455 16197
rect 3713 16337 3759 16404
rect 3713 16178 3759 16197
rect 3857 16337 3903 16358
rect 3506 16072 3520 16118
rect 3660 16072 3759 16118
rect 3409 15945 3512 15991
rect 3652 15945 3664 15991
rect 3265 15786 3311 15826
rect 3409 15872 3455 15889
rect 3409 15740 3455 15826
rect 3713 15872 3759 16072
rect 3857 15991 3903 16197
rect 4161 16337 4207 16404
rect 4161 16178 4207 16197
rect 4305 16337 4351 16358
rect 3954 16072 3968 16118
rect 4108 16072 4207 16118
rect 3857 15945 3960 15991
rect 4100 15945 4112 15991
rect 3713 15786 3759 15826
rect 3857 15872 3903 15889
rect 3857 15740 3903 15826
rect 4161 15872 4207 16072
rect 4305 15991 4351 16197
rect 4609 16337 4655 16404
rect 4609 16178 4655 16197
rect 4753 16337 4799 16358
rect 4402 16072 4416 16118
rect 4556 16072 4655 16118
rect 4305 15945 4408 15991
rect 4548 15945 4560 15991
rect 4161 15786 4207 15826
rect 4305 15872 4351 15889
rect 4305 15740 4351 15826
rect 4609 15872 4655 16072
rect 4753 15991 4799 16197
rect 5057 16337 5103 16404
rect 5057 16178 5103 16197
rect 5342 16379 5410 16404
rect 5342 16333 5353 16379
rect 5399 16333 5410 16379
rect 5342 16251 5410 16333
rect 5342 16205 5353 16251
rect 5399 16205 5410 16251
rect 5342 16123 5410 16205
rect 4850 16072 4864 16118
rect 5004 16072 5103 16118
rect 4753 15945 4856 15991
rect 4996 15945 5008 15991
rect 4609 15786 4655 15826
rect 4753 15872 4799 15889
rect 4753 15740 4799 15826
rect 5057 15872 5103 16072
rect 5342 16077 5353 16123
rect 5399 16077 5410 16123
rect 5342 16066 5410 16077
rect 5537 16337 5583 16358
rect 5537 15991 5583 16197
rect 5841 16337 5887 16404
rect 5841 16178 5887 16197
rect 5985 16337 6031 16358
rect 5634 16072 5648 16118
rect 5788 16072 5887 16118
rect 5537 15945 5640 15991
rect 5780 15945 5792 15991
rect 5057 15786 5103 15826
rect 5342 15906 5410 15917
rect 5342 15759 5353 15906
rect 5399 15759 5410 15906
rect 5342 15740 5410 15759
rect 5537 15872 5583 15889
rect 5537 15740 5583 15826
rect 5841 15872 5887 16072
rect 5985 15991 6031 16197
rect 6289 16337 6335 16404
rect 6289 16178 6335 16197
rect 6433 16337 6479 16358
rect 6082 16072 6096 16118
rect 6236 16072 6335 16118
rect 5985 15945 6088 15991
rect 6228 15945 6240 15991
rect 5841 15786 5887 15826
rect 5985 15872 6031 15889
rect 5985 15740 6031 15826
rect 6289 15872 6335 16072
rect 6433 15991 6479 16197
rect 6737 16337 6783 16404
rect 6737 16178 6783 16197
rect 6881 16337 6927 16358
rect 6530 16072 6544 16118
rect 6684 16072 6783 16118
rect 6433 15945 6536 15991
rect 6676 15945 6688 15991
rect 6289 15786 6335 15826
rect 6433 15872 6479 15889
rect 6433 15740 6479 15826
rect 6737 15872 6783 16072
rect 6881 15991 6927 16197
rect 7185 16337 7231 16404
rect 7185 16178 7231 16197
rect 7329 16337 7375 16358
rect 6978 16072 6992 16118
rect 7132 16072 7231 16118
rect 6881 15945 6984 15991
rect 7124 15945 7136 15991
rect 6737 15786 6783 15826
rect 6881 15872 6927 15889
rect 6881 15740 6927 15826
rect 7185 15872 7231 16072
rect 7329 15991 7375 16197
rect 7633 16337 7679 16404
rect 7633 16178 7679 16197
rect 7777 16337 7823 16358
rect 7426 16072 7440 16118
rect 7580 16072 7679 16118
rect 7329 15945 7432 15991
rect 7572 15945 7584 15991
rect 7185 15786 7231 15826
rect 7329 15872 7375 15889
rect 7329 15740 7375 15826
rect 7633 15872 7679 16072
rect 7777 15991 7823 16197
rect 8081 16337 8127 16404
rect 8081 16178 8127 16197
rect 8225 16337 8271 16358
rect 7874 16072 7888 16118
rect 8028 16072 8127 16118
rect 7777 15945 7880 15991
rect 8020 15945 8032 15991
rect 7633 15786 7679 15826
rect 7777 15872 7823 15889
rect 7777 15740 7823 15826
rect 8081 15872 8127 16072
rect 8225 15991 8271 16197
rect 8529 16337 8575 16404
rect 8529 16178 8575 16197
rect 8673 16337 8719 16358
rect 8322 16072 8336 16118
rect 8476 16072 8575 16118
rect 8225 15945 8328 15991
rect 8468 15945 8480 15991
rect 8081 15786 8127 15826
rect 8225 15872 8271 15889
rect 8225 15740 8271 15826
rect 8529 15872 8575 16072
rect 8673 15991 8719 16197
rect 8977 16337 9023 16404
rect 8977 16178 9023 16197
rect 9262 16379 9330 16404
rect 9262 16333 9273 16379
rect 9319 16333 9330 16379
rect 9262 16251 9330 16333
rect 9262 16205 9273 16251
rect 9319 16205 9330 16251
rect 9262 16123 9330 16205
rect 8770 16072 8784 16118
rect 8924 16072 9023 16118
rect 8673 15945 8776 15991
rect 8916 15945 8928 15991
rect 8529 15786 8575 15826
rect 8673 15872 8719 15889
rect 8673 15740 8719 15826
rect 8977 15872 9023 16072
rect 9262 16077 9273 16123
rect 9319 16077 9330 16123
rect 9262 16066 9330 16077
rect 9457 16337 9503 16358
rect 9457 15991 9503 16197
rect 9761 16337 9807 16404
rect 9761 16178 9807 16197
rect 9905 16337 9951 16358
rect 9554 16072 9568 16118
rect 9708 16072 9807 16118
rect 9457 15945 9560 15991
rect 9700 15945 9712 15991
rect 8977 15786 9023 15826
rect 9262 15906 9330 15917
rect 9262 15759 9273 15906
rect 9319 15759 9330 15906
rect 9262 15740 9330 15759
rect 9457 15872 9503 15889
rect 9457 15740 9503 15826
rect 9761 15872 9807 16072
rect 9905 15991 9951 16197
rect 10209 16337 10255 16404
rect 10209 16178 10255 16197
rect 10353 16337 10399 16358
rect 10002 16072 10016 16118
rect 10156 16072 10255 16118
rect 9905 15945 10008 15991
rect 10148 15945 10160 15991
rect 9761 15786 9807 15826
rect 9905 15872 9951 15889
rect 9905 15740 9951 15826
rect 10209 15872 10255 16072
rect 10353 15991 10399 16197
rect 10657 16337 10703 16404
rect 10657 16178 10703 16197
rect 10801 16337 10847 16358
rect 10450 16072 10464 16118
rect 10604 16072 10703 16118
rect 10353 15945 10456 15991
rect 10596 15945 10608 15991
rect 10209 15786 10255 15826
rect 10353 15872 10399 15889
rect 10353 15740 10399 15826
rect 10657 15872 10703 16072
rect 10801 15991 10847 16197
rect 11105 16337 11151 16404
rect 11105 16178 11151 16197
rect 11249 16337 11295 16358
rect 10898 16072 10912 16118
rect 11052 16072 11151 16118
rect 10801 15945 10904 15991
rect 11044 15945 11056 15991
rect 10657 15786 10703 15826
rect 10801 15872 10847 15889
rect 10801 15740 10847 15826
rect 11105 15872 11151 16072
rect 11249 15991 11295 16197
rect 11553 16337 11599 16404
rect 11553 16178 11599 16197
rect 11697 16337 11743 16358
rect 11346 16072 11360 16118
rect 11500 16072 11599 16118
rect 11249 15945 11352 15991
rect 11492 15945 11504 15991
rect 11105 15786 11151 15826
rect 11249 15872 11295 15889
rect 11249 15740 11295 15826
rect 11553 15872 11599 16072
rect 11697 15991 11743 16197
rect 12001 16337 12047 16404
rect 12001 16178 12047 16197
rect 12145 16337 12191 16358
rect 11794 16072 11808 16118
rect 11948 16072 12047 16118
rect 11697 15945 11800 15991
rect 11940 15945 11952 15991
rect 11553 15786 11599 15826
rect 11697 15872 11743 15889
rect 11697 15740 11743 15826
rect 12001 15872 12047 16072
rect 12145 15991 12191 16197
rect 12449 16337 12495 16404
rect 12449 16178 12495 16197
rect 12593 16337 12639 16358
rect 12242 16072 12256 16118
rect 12396 16072 12495 16118
rect 12145 15945 12248 15991
rect 12388 15945 12400 15991
rect 12001 15786 12047 15826
rect 12145 15872 12191 15889
rect 12145 15740 12191 15826
rect 12449 15872 12495 16072
rect 12593 15991 12639 16197
rect 12897 16337 12943 16404
rect 12897 16178 12943 16197
rect 13182 16379 13250 16404
rect 13182 16333 13193 16379
rect 13239 16333 13250 16379
rect 13182 16251 13250 16333
rect 13182 16205 13193 16251
rect 13239 16205 13250 16251
rect 13182 16123 13250 16205
rect 12690 16072 12704 16118
rect 12844 16072 12943 16118
rect 12593 15945 12696 15991
rect 12836 15945 12848 15991
rect 12449 15786 12495 15826
rect 12593 15872 12639 15889
rect 12593 15740 12639 15826
rect 12897 15872 12943 16072
rect 13182 16077 13193 16123
rect 13239 16077 13250 16123
rect 13182 16066 13250 16077
rect 13377 16337 13423 16358
rect 13377 15991 13423 16197
rect 13681 16337 13727 16404
rect 13681 16178 13727 16197
rect 13825 16337 13871 16358
rect 13474 16072 13488 16118
rect 13628 16072 13727 16118
rect 13377 15945 13480 15991
rect 13620 15945 13632 15991
rect 12897 15786 12943 15826
rect 13182 15906 13250 15917
rect 13182 15759 13193 15906
rect 13239 15759 13250 15906
rect 13182 15740 13250 15759
rect 13377 15872 13423 15889
rect 13377 15740 13423 15826
rect 13681 15872 13727 16072
rect 13825 15991 13871 16197
rect 14129 16337 14175 16404
rect 14129 16178 14175 16197
rect 14273 16337 14319 16358
rect 13922 16072 13936 16118
rect 14076 16072 14175 16118
rect 13825 15945 13928 15991
rect 14068 15945 14080 15991
rect 13681 15786 13727 15826
rect 13825 15872 13871 15889
rect 13825 15740 13871 15826
rect 14129 15872 14175 16072
rect 14273 15991 14319 16197
rect 14577 16337 14623 16404
rect 14577 16178 14623 16197
rect 14721 16337 14767 16358
rect 14370 16072 14384 16118
rect 14524 16072 14623 16118
rect 14273 15945 14376 15991
rect 14516 15945 14528 15991
rect 14129 15786 14175 15826
rect 14273 15872 14319 15889
rect 14273 15740 14319 15826
rect 14577 15872 14623 16072
rect 14721 15991 14767 16197
rect 15025 16337 15071 16404
rect 15025 16178 15071 16197
rect 15169 16337 15215 16358
rect 14818 16072 14832 16118
rect 14972 16072 15071 16118
rect 14721 15945 14824 15991
rect 14964 15945 14976 15991
rect 14577 15786 14623 15826
rect 14721 15872 14767 15889
rect 14721 15740 14767 15826
rect 15025 15872 15071 16072
rect 15169 15991 15215 16197
rect 15473 16337 15519 16404
rect 15473 16178 15519 16197
rect 15617 16337 15663 16358
rect 15266 16072 15280 16118
rect 15420 16072 15519 16118
rect 15169 15945 15272 15991
rect 15412 15945 15424 15991
rect 15025 15786 15071 15826
rect 15169 15872 15215 15889
rect 15169 15740 15215 15826
rect 15473 15872 15519 16072
rect 15617 15991 15663 16197
rect 15921 16337 15967 16404
rect 15921 16178 15967 16197
rect 16065 16337 16111 16358
rect 15714 16072 15728 16118
rect 15868 16072 15967 16118
rect 15617 15945 15720 15991
rect 15860 15945 15872 15991
rect 15473 15786 15519 15826
rect 15617 15872 15663 15889
rect 15617 15740 15663 15826
rect 15921 15872 15967 16072
rect 16065 15991 16111 16197
rect 16369 16337 16415 16404
rect 16369 16178 16415 16197
rect 16513 16337 16559 16358
rect 16162 16072 16176 16118
rect 16316 16072 16415 16118
rect 16065 15945 16168 15991
rect 16308 15945 16320 15991
rect 15921 15786 15967 15826
rect 16065 15872 16111 15889
rect 16065 15740 16111 15826
rect 16369 15872 16415 16072
rect 16513 15991 16559 16197
rect 16817 16337 16863 16404
rect 16817 16178 16863 16197
rect 17102 16379 17170 16404
rect 17102 16333 17113 16379
rect 17159 16333 17170 16379
rect 17102 16251 17170 16333
rect 17102 16205 17113 16251
rect 17159 16205 17170 16251
rect 17102 16123 17170 16205
rect 16610 16072 16624 16118
rect 16764 16072 16863 16118
rect 16513 15945 16616 15991
rect 16756 15945 16768 15991
rect 16369 15786 16415 15826
rect 16513 15872 16559 15889
rect 16513 15740 16559 15826
rect 16817 15872 16863 16072
rect 17102 16077 17113 16123
rect 17159 16077 17170 16123
rect 17102 16066 17170 16077
rect 17297 16337 17343 16358
rect 17297 15991 17343 16197
rect 17601 16337 17647 16404
rect 17601 16178 17647 16197
rect 17745 16337 17791 16358
rect 17394 16072 17408 16118
rect 17548 16072 17647 16118
rect 17297 15945 17400 15991
rect 17540 15945 17552 15991
rect 16817 15786 16863 15826
rect 17102 15906 17170 15917
rect 17102 15759 17113 15906
rect 17159 15759 17170 15906
rect 17102 15740 17170 15759
rect 17297 15872 17343 15889
rect 17297 15740 17343 15826
rect 17601 15872 17647 16072
rect 17745 15991 17791 16197
rect 18049 16337 18095 16404
rect 18049 16178 18095 16197
rect 18193 16337 18239 16358
rect 17842 16072 17856 16118
rect 17996 16072 18095 16118
rect 17745 15945 17848 15991
rect 17988 15945 18000 15991
rect 17601 15786 17647 15826
rect 17745 15872 17791 15889
rect 17745 15740 17791 15826
rect 18049 15872 18095 16072
rect 18193 15991 18239 16197
rect 18497 16337 18543 16404
rect 18497 16178 18543 16197
rect 18641 16337 18687 16358
rect 18290 16072 18304 16118
rect 18444 16072 18543 16118
rect 18193 15945 18296 15991
rect 18436 15945 18448 15991
rect 18049 15786 18095 15826
rect 18193 15872 18239 15889
rect 18193 15740 18239 15826
rect 18497 15872 18543 16072
rect 18641 15991 18687 16197
rect 18945 16337 18991 16404
rect 18945 16178 18991 16197
rect 19089 16337 19135 16358
rect 18738 16072 18752 16118
rect 18892 16072 18991 16118
rect 18641 15945 18744 15991
rect 18884 15945 18896 15991
rect 18497 15786 18543 15826
rect 18641 15872 18687 15889
rect 18641 15740 18687 15826
rect 18945 15872 18991 16072
rect 19089 15991 19135 16197
rect 19393 16337 19439 16404
rect 19393 16178 19439 16197
rect 19537 16337 19583 16358
rect 19186 16072 19200 16118
rect 19340 16072 19439 16118
rect 19089 15945 19192 15991
rect 19332 15945 19344 15991
rect 18945 15786 18991 15826
rect 19089 15872 19135 15889
rect 19089 15740 19135 15826
rect 19393 15872 19439 16072
rect 19537 15991 19583 16197
rect 19841 16337 19887 16404
rect 19841 16178 19887 16197
rect 19985 16337 20031 16358
rect 19634 16072 19648 16118
rect 19788 16072 19887 16118
rect 19537 15945 19640 15991
rect 19780 15945 19792 15991
rect 19393 15786 19439 15826
rect 19537 15872 19583 15889
rect 19537 15740 19583 15826
rect 19841 15872 19887 16072
rect 19985 15991 20031 16197
rect 20289 16337 20335 16404
rect 20289 16178 20335 16197
rect 20433 16337 20479 16358
rect 20082 16072 20096 16118
rect 20236 16072 20335 16118
rect 19985 15945 20088 15991
rect 20228 15945 20240 15991
rect 19841 15786 19887 15826
rect 19985 15872 20031 15889
rect 19985 15740 20031 15826
rect 20289 15872 20335 16072
rect 20433 15991 20479 16197
rect 20737 16337 20783 16404
rect 20737 16178 20783 16197
rect 21022 16379 21090 16404
rect 21022 16333 21033 16379
rect 21079 16333 21090 16379
rect 21022 16251 21090 16333
rect 21022 16205 21033 16251
rect 21079 16205 21090 16251
rect 21022 16123 21090 16205
rect 20530 16072 20544 16118
rect 20684 16072 20783 16118
rect 20433 15945 20536 15991
rect 20676 15945 20688 15991
rect 20289 15786 20335 15826
rect 20433 15872 20479 15889
rect 20433 15740 20479 15826
rect 20737 15872 20783 16072
rect 21022 16077 21033 16123
rect 21079 16077 21090 16123
rect 21022 16066 21090 16077
rect 21217 16337 21263 16358
rect 21217 15991 21263 16197
rect 21521 16337 21567 16404
rect 21521 16178 21567 16197
rect 21665 16337 21711 16358
rect 21314 16072 21328 16118
rect 21468 16072 21567 16118
rect 21217 15945 21320 15991
rect 21460 15945 21472 15991
rect 20737 15786 20783 15826
rect 21022 15906 21090 15917
rect 21022 15759 21033 15906
rect 21079 15759 21090 15906
rect 21022 15740 21090 15759
rect 21217 15872 21263 15897
rect 21217 15740 21263 15826
rect 21521 15872 21567 16072
rect 21665 15991 21711 16197
rect 21969 16337 22015 16404
rect 21969 16178 22015 16197
rect 22482 16379 22550 16404
rect 22482 16333 22493 16379
rect 22539 16333 22550 16379
rect 22482 16251 22550 16333
rect 22482 16205 22493 16251
rect 22539 16205 22550 16251
rect 22482 16123 22550 16205
rect 21762 16072 21776 16118
rect 21916 16072 22015 16118
rect 21665 15945 21768 15991
rect 21908 15945 21920 15991
rect 21521 15786 21567 15826
rect 21665 15872 21711 15897
rect 21665 15740 21711 15826
rect 21969 15872 22015 16072
rect 22482 16077 22493 16123
rect 22539 16077 22550 16123
rect 22482 16064 22550 16077
rect 21969 15786 22015 15826
rect 22482 15906 22550 15918
rect 22482 15759 22493 15906
rect 22539 15759 22550 15906
rect 22482 15740 22550 15759
rect 1344 15706 22784 15740
rect 1344 15654 6534 15706
rect 6794 15654 11854 15706
rect 12114 15654 17174 15706
rect 17434 15654 22494 15706
rect 22754 15654 22784 15706
rect 1344 15620 22784 15654
rect 1418 15601 1486 15620
rect 1418 15454 1429 15601
rect 1475 15454 1486 15601
rect 1617 15534 1663 15620
rect 1617 15469 1663 15488
rect 1921 15534 1967 15574
rect 1418 15442 1486 15454
rect 1617 15369 1720 15415
rect 1860 15369 1872 15415
rect 1418 15283 1486 15296
rect 1418 15237 1429 15283
rect 1475 15237 1486 15283
rect 1418 15155 1486 15237
rect 1418 15109 1429 15155
rect 1475 15109 1486 15155
rect 1418 15027 1486 15109
rect 1418 14981 1429 15027
rect 1475 14981 1486 15027
rect 1617 15163 1663 15369
rect 1921 15288 1967 15488
rect 2065 15534 2111 15620
rect 2065 15469 2111 15488
rect 2369 15534 2415 15574
rect 1714 15242 1728 15288
rect 1868 15242 1967 15288
rect 2065 15369 2168 15415
rect 2308 15369 2320 15415
rect 1617 15002 1663 15023
rect 1921 15163 1967 15182
rect 1418 14956 1486 14981
rect 1921 14956 1967 15023
rect 2065 15163 2111 15369
rect 2369 15288 2415 15488
rect 2513 15534 2559 15620
rect 2513 15469 2559 15488
rect 2817 15534 2863 15574
rect 2162 15242 2176 15288
rect 2316 15242 2415 15288
rect 2513 15369 2616 15415
rect 2756 15369 2768 15415
rect 2065 15002 2111 15023
rect 2369 15163 2415 15182
rect 2369 14956 2415 15023
rect 2513 15163 2559 15369
rect 2817 15288 2863 15488
rect 2961 15534 3007 15620
rect 2961 15469 3007 15488
rect 3265 15534 3311 15574
rect 2610 15242 2624 15288
rect 2764 15242 2863 15288
rect 2961 15369 3064 15415
rect 3204 15369 3216 15415
rect 2513 15002 2559 15023
rect 2817 15163 2863 15182
rect 2817 14956 2863 15023
rect 2961 15163 3007 15369
rect 3265 15288 3311 15488
rect 3409 15534 3455 15620
rect 3409 15469 3455 15488
rect 3713 15534 3759 15574
rect 3058 15242 3072 15288
rect 3212 15242 3311 15288
rect 3409 15369 3512 15415
rect 3652 15369 3664 15415
rect 2961 15002 3007 15023
rect 3265 15163 3311 15182
rect 3265 14956 3311 15023
rect 3409 15163 3455 15369
rect 3713 15288 3759 15488
rect 3857 15534 3903 15620
rect 3857 15469 3903 15488
rect 4161 15534 4207 15574
rect 3506 15242 3520 15288
rect 3660 15242 3759 15288
rect 3857 15369 3960 15415
rect 4100 15369 4112 15415
rect 3409 15002 3455 15023
rect 3713 15163 3759 15182
rect 3713 14956 3759 15023
rect 3857 15163 3903 15369
rect 4161 15288 4207 15488
rect 4305 15534 4351 15620
rect 4305 15469 4351 15488
rect 4609 15534 4655 15574
rect 3954 15242 3968 15288
rect 4108 15242 4207 15288
rect 4305 15369 4408 15415
rect 4548 15369 4560 15415
rect 3857 15002 3903 15023
rect 4161 15163 4207 15182
rect 4161 14956 4207 15023
rect 4305 15163 4351 15369
rect 4609 15288 4655 15488
rect 4753 15534 4799 15620
rect 4753 15469 4799 15488
rect 5057 15534 5103 15574
rect 4402 15242 4416 15288
rect 4556 15242 4655 15288
rect 4753 15369 4856 15415
rect 4996 15369 5008 15415
rect 4305 15002 4351 15023
rect 4609 15163 4655 15182
rect 4609 14956 4655 15023
rect 4753 15163 4799 15369
rect 5057 15288 5103 15488
rect 5201 15534 5247 15620
rect 5201 15469 5247 15488
rect 5505 15534 5551 15574
rect 4850 15242 4864 15288
rect 5004 15242 5103 15288
rect 5201 15369 5304 15415
rect 5444 15369 5456 15415
rect 4753 15002 4799 15023
rect 5057 15163 5103 15182
rect 5057 14956 5103 15023
rect 5201 15163 5247 15369
rect 5505 15288 5551 15488
rect 5649 15534 5695 15620
rect 5649 15469 5695 15488
rect 5953 15534 5999 15574
rect 5298 15242 5312 15288
rect 5452 15242 5551 15288
rect 5649 15369 5752 15415
rect 5892 15369 5904 15415
rect 5201 15002 5247 15023
rect 5505 15163 5551 15182
rect 5505 14956 5551 15023
rect 5649 15163 5695 15369
rect 5953 15288 5999 15488
rect 6097 15534 6143 15620
rect 6097 15469 6143 15488
rect 6401 15534 6447 15574
rect 5746 15242 5760 15288
rect 5900 15242 5999 15288
rect 6097 15369 6200 15415
rect 6340 15369 6352 15415
rect 5649 15002 5695 15023
rect 5953 15163 5999 15182
rect 5953 14956 5999 15023
rect 6097 15163 6143 15369
rect 6401 15288 6447 15488
rect 6545 15534 6591 15620
rect 6545 15469 6591 15488
rect 6849 15534 6895 15574
rect 6194 15242 6208 15288
rect 6348 15242 6447 15288
rect 6545 15369 6648 15415
rect 6788 15369 6800 15415
rect 6097 15002 6143 15023
rect 6401 15163 6447 15182
rect 6401 14956 6447 15023
rect 6545 15163 6591 15369
rect 6849 15288 6895 15488
rect 6993 15534 7039 15620
rect 6993 15469 7039 15488
rect 7297 15534 7343 15574
rect 6642 15242 6656 15288
rect 6796 15242 6895 15288
rect 6993 15369 7096 15415
rect 7236 15369 7248 15415
rect 6545 15002 6591 15023
rect 6849 15163 6895 15182
rect 6849 14956 6895 15023
rect 6993 15163 7039 15369
rect 7297 15288 7343 15488
rect 7441 15534 7487 15620
rect 7441 15469 7487 15488
rect 7745 15534 7791 15574
rect 7090 15242 7104 15288
rect 7244 15242 7343 15288
rect 7441 15369 7544 15415
rect 7684 15369 7696 15415
rect 6993 15002 7039 15023
rect 7297 15163 7343 15182
rect 7297 14956 7343 15023
rect 7441 15163 7487 15369
rect 7745 15288 7791 15488
rect 7889 15534 7935 15620
rect 7889 15469 7935 15488
rect 8193 15534 8239 15574
rect 7538 15242 7552 15288
rect 7692 15242 7791 15288
rect 7889 15369 7992 15415
rect 8132 15369 8144 15415
rect 7441 15002 7487 15023
rect 7745 15163 7791 15182
rect 7745 14956 7791 15023
rect 7889 15163 7935 15369
rect 8193 15288 8239 15488
rect 8337 15534 8383 15620
rect 8337 15469 8383 15488
rect 8641 15534 8687 15574
rect 7986 15242 8000 15288
rect 8140 15242 8239 15288
rect 8337 15369 8440 15415
rect 8580 15369 8592 15415
rect 7889 15002 7935 15023
rect 8193 15163 8239 15182
rect 8193 14956 8239 15023
rect 8337 15163 8383 15369
rect 8641 15288 8687 15488
rect 8785 15534 8831 15620
rect 9374 15601 9442 15620
rect 8785 15461 8831 15488
rect 9089 15534 9135 15574
rect 8434 15242 8448 15288
rect 8588 15242 8687 15288
rect 8785 15369 8888 15415
rect 9028 15369 9040 15415
rect 8337 15002 8383 15023
rect 8641 15163 8687 15182
rect 8641 14956 8687 15023
rect 8785 15163 8831 15369
rect 9089 15288 9135 15488
rect 9374 15454 9385 15601
rect 9431 15454 9442 15601
rect 9569 15534 9615 15620
rect 9569 15469 9615 15488
rect 9873 15534 9919 15574
rect 9374 15443 9442 15454
rect 9569 15369 9672 15415
rect 9812 15369 9824 15415
rect 8882 15242 8896 15288
rect 9036 15242 9135 15288
rect 9374 15283 9442 15294
rect 9374 15237 9385 15283
rect 9431 15237 9442 15283
rect 8785 15002 8831 15023
rect 9089 15163 9135 15182
rect 9089 14956 9135 15023
rect 9374 15155 9442 15237
rect 9374 15109 9385 15155
rect 9431 15109 9442 15155
rect 9374 15027 9442 15109
rect 9374 14981 9385 15027
rect 9431 14981 9442 15027
rect 9569 15163 9615 15369
rect 9873 15288 9919 15488
rect 10017 15534 10063 15620
rect 10017 15469 10063 15488
rect 10321 15534 10367 15574
rect 9666 15242 9680 15288
rect 9820 15242 9919 15288
rect 10017 15369 10120 15415
rect 10260 15369 10272 15415
rect 9569 15002 9615 15023
rect 9873 15163 9919 15182
rect 9374 14956 9442 14981
rect 9873 14956 9919 15023
rect 10017 15163 10063 15369
rect 10321 15288 10367 15488
rect 10465 15534 10511 15620
rect 10465 15469 10511 15488
rect 10769 15534 10815 15574
rect 10114 15242 10128 15288
rect 10268 15242 10367 15288
rect 10465 15369 10568 15415
rect 10708 15369 10720 15415
rect 10017 15002 10063 15023
rect 10321 15163 10367 15182
rect 10321 14956 10367 15023
rect 10465 15163 10511 15369
rect 10769 15288 10815 15488
rect 10913 15534 10959 15620
rect 10913 15469 10959 15488
rect 11217 15534 11263 15574
rect 10562 15242 10576 15288
rect 10716 15242 10815 15288
rect 10913 15369 11016 15415
rect 11156 15369 11168 15415
rect 10465 15002 10511 15023
rect 10769 15163 10815 15182
rect 10769 14956 10815 15023
rect 10913 15163 10959 15369
rect 11217 15288 11263 15488
rect 11361 15534 11407 15620
rect 11361 15469 11407 15488
rect 11665 15534 11711 15574
rect 11010 15242 11024 15288
rect 11164 15242 11263 15288
rect 11361 15369 11464 15415
rect 11604 15369 11616 15415
rect 10913 15002 10959 15023
rect 11217 15163 11263 15182
rect 11217 14956 11263 15023
rect 11361 15163 11407 15369
rect 11665 15288 11711 15488
rect 11809 15534 11855 15620
rect 11809 15469 11855 15488
rect 12113 15534 12159 15574
rect 11458 15242 11472 15288
rect 11612 15242 11711 15288
rect 11809 15369 11912 15415
rect 12052 15369 12064 15415
rect 11361 15002 11407 15023
rect 11665 15163 11711 15182
rect 11665 14956 11711 15023
rect 11809 15163 11855 15369
rect 12113 15288 12159 15488
rect 12257 15534 12303 15620
rect 12257 15469 12303 15488
rect 12561 15534 12607 15574
rect 11906 15242 11920 15288
rect 12060 15242 12159 15288
rect 12257 15369 12360 15415
rect 12500 15369 12512 15415
rect 11809 15002 11855 15023
rect 12113 15163 12159 15182
rect 12113 14956 12159 15023
rect 12257 15163 12303 15369
rect 12561 15288 12607 15488
rect 12705 15534 12751 15620
rect 12705 15469 12751 15488
rect 13009 15534 13055 15574
rect 12354 15242 12368 15288
rect 12508 15242 12607 15288
rect 12705 15369 12808 15415
rect 12948 15369 12960 15415
rect 12257 15002 12303 15023
rect 12561 15163 12607 15182
rect 12561 14956 12607 15023
rect 12705 15163 12751 15369
rect 13009 15288 13055 15488
rect 13153 15534 13199 15620
rect 13153 15469 13199 15488
rect 13457 15534 13503 15574
rect 12802 15242 12816 15288
rect 12956 15242 13055 15288
rect 13153 15369 13256 15415
rect 13396 15369 13408 15415
rect 12705 15002 12751 15023
rect 13009 15163 13055 15182
rect 13009 14956 13055 15023
rect 13153 15163 13199 15369
rect 13457 15288 13503 15488
rect 13601 15534 13647 15620
rect 13601 15469 13647 15488
rect 13905 15534 13951 15574
rect 13250 15242 13264 15288
rect 13404 15242 13503 15288
rect 13601 15369 13704 15415
rect 13844 15369 13856 15415
rect 13153 15002 13199 15023
rect 13457 15163 13503 15182
rect 13457 14956 13503 15023
rect 13601 15163 13647 15369
rect 13905 15288 13951 15488
rect 14049 15534 14095 15620
rect 14049 15469 14095 15488
rect 14353 15534 14399 15574
rect 13698 15242 13712 15288
rect 13852 15242 13951 15288
rect 14049 15369 14152 15415
rect 14292 15369 14304 15415
rect 13601 15002 13647 15023
rect 13905 15163 13951 15182
rect 13905 14956 13951 15023
rect 14049 15163 14095 15369
rect 14353 15288 14399 15488
rect 14497 15534 14543 15620
rect 14497 15469 14543 15488
rect 14801 15534 14847 15574
rect 14146 15242 14160 15288
rect 14300 15242 14399 15288
rect 14497 15369 14600 15415
rect 14740 15369 14752 15415
rect 14049 15002 14095 15023
rect 14353 15163 14399 15182
rect 14353 14956 14399 15023
rect 14497 15163 14543 15369
rect 14801 15288 14847 15488
rect 14945 15534 14991 15620
rect 14945 15469 14991 15488
rect 15249 15534 15295 15574
rect 14594 15242 14608 15288
rect 14748 15242 14847 15288
rect 14945 15369 15048 15415
rect 15188 15369 15200 15415
rect 14497 15002 14543 15023
rect 14801 15163 14847 15182
rect 14801 14956 14847 15023
rect 14945 15163 14991 15369
rect 15249 15288 15295 15488
rect 15393 15534 15439 15620
rect 15393 15469 15439 15488
rect 15697 15534 15743 15574
rect 15042 15242 15056 15288
rect 15196 15242 15295 15288
rect 15393 15369 15496 15415
rect 15636 15369 15648 15415
rect 14945 15002 14991 15023
rect 15249 15163 15295 15182
rect 15249 14956 15295 15023
rect 15393 15163 15439 15369
rect 15697 15288 15743 15488
rect 15841 15534 15887 15620
rect 15841 15469 15887 15488
rect 16145 15534 16191 15574
rect 15490 15242 15504 15288
rect 15644 15242 15743 15288
rect 15841 15369 15944 15415
rect 16084 15369 16096 15415
rect 15393 15002 15439 15023
rect 15697 15163 15743 15182
rect 15697 14956 15743 15023
rect 15841 15163 15887 15369
rect 16145 15288 16191 15488
rect 16289 15534 16335 15620
rect 16289 15469 16335 15488
rect 16593 15534 16639 15574
rect 15938 15242 15952 15288
rect 16092 15242 16191 15288
rect 16289 15369 16392 15415
rect 16532 15369 16544 15415
rect 15841 15002 15887 15023
rect 16145 15163 16191 15182
rect 16145 14956 16191 15023
rect 16289 15163 16335 15369
rect 16593 15288 16639 15488
rect 16737 15534 16783 15620
rect 17326 15601 17394 15620
rect 16737 15461 16783 15488
rect 17041 15534 17087 15574
rect 16386 15242 16400 15288
rect 16540 15242 16639 15288
rect 16737 15369 16840 15415
rect 16980 15369 16992 15415
rect 16289 15002 16335 15023
rect 16593 15163 16639 15182
rect 16593 14956 16639 15023
rect 16737 15163 16783 15369
rect 17041 15288 17087 15488
rect 17326 15454 17337 15601
rect 17383 15454 17394 15601
rect 17521 15534 17567 15620
rect 17521 15471 17567 15488
rect 17825 15534 17871 15574
rect 17326 15443 17394 15454
rect 17521 15369 17624 15415
rect 17764 15369 17776 15415
rect 16834 15242 16848 15288
rect 16988 15242 17087 15288
rect 17326 15283 17394 15294
rect 17326 15237 17337 15283
rect 17383 15237 17394 15283
rect 16737 15002 16783 15023
rect 17041 15163 17087 15182
rect 17041 14956 17087 15023
rect 17326 15155 17394 15237
rect 17326 15109 17337 15155
rect 17383 15109 17394 15155
rect 17326 15027 17394 15109
rect 17326 14981 17337 15027
rect 17383 14981 17394 15027
rect 17521 15163 17567 15369
rect 17825 15288 17871 15488
rect 17969 15534 18015 15620
rect 17969 15471 18015 15488
rect 18273 15534 18319 15574
rect 17618 15242 17632 15288
rect 17772 15242 17871 15288
rect 17969 15369 18072 15415
rect 18212 15369 18224 15415
rect 17521 15002 17567 15023
rect 17825 15163 17871 15182
rect 17326 14956 17394 14981
rect 17825 14956 17871 15023
rect 17969 15163 18015 15369
rect 18273 15288 18319 15488
rect 18417 15534 18463 15620
rect 18417 15471 18463 15488
rect 18721 15534 18767 15574
rect 18066 15242 18080 15288
rect 18220 15242 18319 15288
rect 18417 15369 18520 15415
rect 18660 15369 18672 15415
rect 17969 15002 18015 15023
rect 18273 15163 18319 15182
rect 18273 14956 18319 15023
rect 18417 15163 18463 15369
rect 18721 15288 18767 15488
rect 18865 15534 18911 15620
rect 18865 15471 18911 15488
rect 19169 15534 19215 15574
rect 18514 15242 18528 15288
rect 18668 15242 18767 15288
rect 18865 15369 18968 15415
rect 19108 15369 19120 15415
rect 18417 15002 18463 15023
rect 18721 15163 18767 15182
rect 18721 14956 18767 15023
rect 18865 15163 18911 15369
rect 19169 15288 19215 15488
rect 19313 15534 19359 15620
rect 19313 15471 19359 15488
rect 19617 15534 19663 15574
rect 18962 15242 18976 15288
rect 19116 15242 19215 15288
rect 19313 15369 19416 15415
rect 19556 15369 19568 15415
rect 18865 15002 18911 15023
rect 19169 15163 19215 15182
rect 19169 14956 19215 15023
rect 19313 15163 19359 15369
rect 19617 15288 19663 15488
rect 19761 15534 19807 15620
rect 19761 15471 19807 15488
rect 20065 15534 20111 15574
rect 19410 15242 19424 15288
rect 19564 15242 19663 15288
rect 19761 15369 19864 15415
rect 20004 15369 20016 15415
rect 19313 15002 19359 15023
rect 19617 15163 19663 15182
rect 19617 14956 19663 15023
rect 19761 15163 19807 15369
rect 20065 15288 20111 15488
rect 20209 15534 20255 15620
rect 20209 15471 20255 15488
rect 20513 15534 20559 15574
rect 19858 15242 19872 15288
rect 20012 15242 20111 15288
rect 20209 15369 20312 15415
rect 20452 15369 20464 15415
rect 19761 15002 19807 15023
rect 20065 15163 20111 15182
rect 20065 14956 20111 15023
rect 20209 15163 20255 15369
rect 20513 15288 20559 15488
rect 20657 15534 20703 15620
rect 20657 15471 20703 15488
rect 20961 15534 21007 15574
rect 20306 15242 20320 15288
rect 20460 15242 20559 15288
rect 20657 15369 20760 15415
rect 20900 15369 20912 15415
rect 20209 15002 20255 15023
rect 20513 15163 20559 15182
rect 20513 14956 20559 15023
rect 20657 15163 20703 15369
rect 20961 15288 21007 15488
rect 21105 15534 21151 15620
rect 21105 15463 21151 15488
rect 21409 15534 21455 15574
rect 20754 15242 20768 15288
rect 20908 15242 21007 15288
rect 21105 15369 21208 15415
rect 21348 15369 21360 15415
rect 20657 15002 20703 15023
rect 20961 15163 21007 15182
rect 20961 14956 21007 15023
rect 21105 15163 21151 15369
rect 21409 15288 21455 15488
rect 21553 15534 21599 15620
rect 21553 15463 21599 15488
rect 21857 15534 21903 15574
rect 21202 15242 21216 15288
rect 21356 15242 21455 15288
rect 21553 15369 21656 15415
rect 21796 15369 21808 15415
rect 21105 15002 21151 15023
rect 21409 15163 21455 15182
rect 21409 14956 21455 15023
rect 21553 15163 21599 15369
rect 21857 15288 21903 15488
rect 22001 15534 22047 15620
rect 22482 15601 22550 15620
rect 22001 15461 22047 15488
rect 22305 15534 22351 15574
rect 21650 15242 21664 15288
rect 21804 15242 21903 15288
rect 22001 15369 22104 15415
rect 22244 15369 22256 15415
rect 21553 15002 21599 15023
rect 21857 15163 21903 15182
rect 21857 14956 21903 15023
rect 22001 15163 22047 15369
rect 22305 15288 22351 15488
rect 22482 15454 22493 15601
rect 22539 15454 22550 15601
rect 22482 15442 22550 15454
rect 22098 15242 22112 15288
rect 22252 15242 22351 15288
rect 22482 15283 22550 15296
rect 22482 15237 22493 15283
rect 22539 15237 22550 15283
rect 22001 15002 22047 15023
rect 22305 15163 22351 15182
rect 22305 14956 22351 15023
rect 22482 15155 22550 15237
rect 22482 15109 22493 15155
rect 22539 15109 22550 15155
rect 22482 15027 22550 15109
rect 22482 14981 22493 15027
rect 22539 14981 22550 15027
rect 22482 14956 22550 14981
rect 1344 14922 22624 14956
rect 1344 14870 3874 14922
rect 4134 14870 9194 14922
rect 9454 14870 14514 14922
rect 14774 14870 19834 14922
rect 20094 14870 22624 14922
rect 1344 14836 22624 14870
rect 1418 14811 1486 14836
rect 1418 14765 1429 14811
rect 1475 14765 1486 14811
rect 1418 14683 1486 14765
rect 1418 14637 1429 14683
rect 1475 14637 1486 14683
rect 1418 14555 1486 14637
rect 1418 14509 1429 14555
rect 1475 14509 1486 14555
rect 1418 14496 1486 14509
rect 1617 14769 1663 14790
rect 1617 14423 1663 14629
rect 1921 14769 1967 14836
rect 1921 14610 1967 14629
rect 2065 14769 2111 14790
rect 1714 14504 1728 14550
rect 1868 14504 1967 14550
rect 1617 14377 1720 14423
rect 1860 14377 1872 14423
rect 1418 14338 1486 14350
rect 1418 14191 1429 14338
rect 1475 14191 1486 14338
rect 1418 14172 1486 14191
rect 1617 14304 1663 14321
rect 1617 14172 1663 14258
rect 1921 14304 1967 14504
rect 2065 14423 2111 14629
rect 2369 14769 2415 14836
rect 2369 14610 2415 14629
rect 2513 14769 2559 14790
rect 2162 14504 2176 14550
rect 2316 14504 2415 14550
rect 2065 14377 2168 14423
rect 2308 14377 2320 14423
rect 1921 14218 1967 14258
rect 2065 14304 2111 14321
rect 2065 14172 2111 14258
rect 2369 14304 2415 14504
rect 2513 14423 2559 14629
rect 2817 14769 2863 14836
rect 2817 14610 2863 14629
rect 2961 14769 3007 14790
rect 2610 14504 2624 14550
rect 2764 14504 2863 14550
rect 2513 14377 2616 14423
rect 2756 14377 2768 14423
rect 2369 14218 2415 14258
rect 2513 14304 2559 14321
rect 2513 14172 2559 14258
rect 2817 14304 2863 14504
rect 2961 14423 3007 14629
rect 3265 14769 3311 14836
rect 3265 14610 3311 14629
rect 3409 14769 3455 14790
rect 3058 14504 3072 14550
rect 3212 14504 3311 14550
rect 2961 14377 3064 14423
rect 3204 14377 3216 14423
rect 2817 14218 2863 14258
rect 2961 14304 3007 14321
rect 2961 14172 3007 14258
rect 3265 14304 3311 14504
rect 3409 14423 3455 14629
rect 3713 14769 3759 14836
rect 3713 14610 3759 14629
rect 3857 14769 3903 14790
rect 3506 14504 3520 14550
rect 3660 14504 3759 14550
rect 3409 14377 3512 14423
rect 3652 14377 3664 14423
rect 3265 14218 3311 14258
rect 3409 14304 3455 14321
rect 3409 14172 3455 14258
rect 3713 14304 3759 14504
rect 3857 14423 3903 14629
rect 4161 14769 4207 14836
rect 4161 14610 4207 14629
rect 4305 14769 4351 14790
rect 3954 14504 3968 14550
rect 4108 14504 4207 14550
rect 3857 14377 3960 14423
rect 4100 14377 4112 14423
rect 3713 14218 3759 14258
rect 3857 14304 3903 14321
rect 3857 14172 3903 14258
rect 4161 14304 4207 14504
rect 4305 14423 4351 14629
rect 4609 14769 4655 14836
rect 4609 14610 4655 14629
rect 4753 14769 4799 14790
rect 4402 14504 4416 14550
rect 4556 14504 4655 14550
rect 4305 14377 4408 14423
rect 4548 14377 4560 14423
rect 4161 14218 4207 14258
rect 4305 14304 4351 14321
rect 4305 14172 4351 14258
rect 4609 14304 4655 14504
rect 4753 14423 4799 14629
rect 5057 14769 5103 14836
rect 5057 14610 5103 14629
rect 5342 14811 5410 14836
rect 5342 14765 5353 14811
rect 5399 14765 5410 14811
rect 5342 14683 5410 14765
rect 5342 14637 5353 14683
rect 5399 14637 5410 14683
rect 5342 14555 5410 14637
rect 4850 14504 4864 14550
rect 5004 14504 5103 14550
rect 4753 14377 4856 14423
rect 4996 14377 5008 14423
rect 4609 14218 4655 14258
rect 4753 14304 4799 14321
rect 4753 14172 4799 14258
rect 5057 14304 5103 14504
rect 5342 14509 5353 14555
rect 5399 14509 5410 14555
rect 5342 14498 5410 14509
rect 5537 14769 5583 14790
rect 5537 14423 5583 14629
rect 5841 14769 5887 14836
rect 5841 14610 5887 14629
rect 5985 14769 6031 14790
rect 5634 14504 5648 14550
rect 5788 14504 5887 14550
rect 5537 14377 5640 14423
rect 5780 14377 5792 14423
rect 5057 14218 5103 14258
rect 5342 14338 5410 14349
rect 5342 14191 5353 14338
rect 5399 14191 5410 14338
rect 5342 14172 5410 14191
rect 5537 14304 5583 14323
rect 5537 14172 5583 14258
rect 5841 14304 5887 14504
rect 5985 14423 6031 14629
rect 6289 14769 6335 14836
rect 6289 14610 6335 14629
rect 6433 14769 6479 14790
rect 6082 14504 6096 14550
rect 6236 14504 6335 14550
rect 5985 14377 6088 14423
rect 6228 14377 6240 14423
rect 5841 14218 5887 14258
rect 5985 14304 6031 14323
rect 5985 14172 6031 14258
rect 6289 14304 6335 14504
rect 6433 14423 6479 14629
rect 6737 14769 6783 14836
rect 6737 14610 6783 14629
rect 6881 14769 6927 14790
rect 6530 14504 6544 14550
rect 6684 14504 6783 14550
rect 6433 14377 6536 14423
rect 6676 14377 6688 14423
rect 6289 14218 6335 14258
rect 6433 14304 6479 14323
rect 6433 14172 6479 14258
rect 6737 14304 6783 14504
rect 6881 14423 6927 14629
rect 7185 14769 7231 14836
rect 7185 14610 7231 14629
rect 7329 14769 7375 14790
rect 6978 14504 6992 14550
rect 7132 14504 7231 14550
rect 6881 14377 6984 14423
rect 7124 14377 7136 14423
rect 6737 14218 6783 14258
rect 6881 14304 6927 14323
rect 6881 14172 6927 14258
rect 7185 14304 7231 14504
rect 7329 14423 7375 14629
rect 7633 14769 7679 14836
rect 7633 14610 7679 14629
rect 7777 14769 7823 14790
rect 7426 14504 7440 14550
rect 7580 14504 7679 14550
rect 7329 14377 7432 14423
rect 7572 14377 7584 14423
rect 7185 14218 7231 14258
rect 7329 14304 7375 14323
rect 7329 14172 7375 14258
rect 7633 14304 7679 14504
rect 7777 14423 7823 14629
rect 8081 14769 8127 14836
rect 8081 14610 8127 14629
rect 8225 14769 8271 14790
rect 7874 14504 7888 14550
rect 8028 14504 8127 14550
rect 7777 14377 7880 14423
rect 8020 14377 8032 14423
rect 7633 14218 7679 14258
rect 7777 14304 7823 14323
rect 7777 14172 7823 14258
rect 8081 14304 8127 14504
rect 8225 14423 8271 14629
rect 8529 14769 8575 14836
rect 8529 14610 8575 14629
rect 8673 14769 8719 14790
rect 8322 14504 8336 14550
rect 8476 14504 8575 14550
rect 8225 14377 8328 14423
rect 8468 14377 8480 14423
rect 8081 14218 8127 14258
rect 8225 14304 8271 14323
rect 8225 14172 8271 14258
rect 8529 14304 8575 14504
rect 8673 14423 8719 14629
rect 8977 14769 9023 14836
rect 8977 14610 9023 14629
rect 9121 14769 9167 14790
rect 8770 14504 8784 14550
rect 8924 14504 9023 14550
rect 8673 14377 8776 14423
rect 8916 14377 8928 14423
rect 8529 14218 8575 14258
rect 8673 14304 8719 14323
rect 8673 14172 8719 14258
rect 8977 14304 9023 14504
rect 9121 14423 9167 14629
rect 9425 14769 9471 14836
rect 9425 14610 9471 14629
rect 9569 14769 9615 14790
rect 9218 14504 9232 14550
rect 9372 14504 9471 14550
rect 9121 14377 9224 14423
rect 9364 14377 9376 14423
rect 8977 14218 9023 14258
rect 9121 14304 9167 14323
rect 9121 14172 9167 14258
rect 9425 14304 9471 14504
rect 9569 14423 9615 14629
rect 9873 14769 9919 14836
rect 9873 14610 9919 14629
rect 10017 14769 10063 14790
rect 9666 14504 9680 14550
rect 9820 14504 9919 14550
rect 9569 14377 9672 14423
rect 9812 14377 9824 14423
rect 9425 14218 9471 14258
rect 9569 14304 9615 14323
rect 9569 14172 9615 14258
rect 9873 14304 9919 14504
rect 10017 14423 10063 14629
rect 10321 14769 10367 14836
rect 10321 14610 10367 14629
rect 10465 14769 10511 14790
rect 10114 14504 10128 14550
rect 10268 14504 10367 14550
rect 10017 14377 10120 14423
rect 10260 14377 10272 14423
rect 9873 14218 9919 14258
rect 10017 14304 10063 14323
rect 10017 14172 10063 14258
rect 10321 14304 10367 14504
rect 10465 14423 10511 14629
rect 10769 14769 10815 14836
rect 10769 14610 10815 14629
rect 10913 14769 10959 14790
rect 10562 14504 10576 14550
rect 10716 14504 10815 14550
rect 10465 14377 10568 14423
rect 10708 14377 10720 14423
rect 10321 14218 10367 14258
rect 10465 14304 10511 14323
rect 10465 14172 10511 14258
rect 10769 14304 10815 14504
rect 10913 14423 10959 14629
rect 11217 14769 11263 14836
rect 11217 14610 11263 14629
rect 11361 14769 11407 14790
rect 11010 14504 11024 14550
rect 11164 14504 11263 14550
rect 10913 14377 11016 14423
rect 11156 14377 11168 14423
rect 10769 14218 10815 14258
rect 10913 14304 10959 14323
rect 10913 14172 10959 14258
rect 11217 14304 11263 14504
rect 11361 14423 11407 14629
rect 11665 14769 11711 14836
rect 11665 14610 11711 14629
rect 11809 14769 11855 14790
rect 11458 14504 11472 14550
rect 11612 14504 11711 14550
rect 11361 14377 11464 14423
rect 11604 14377 11616 14423
rect 11217 14218 11263 14258
rect 11361 14304 11407 14323
rect 11361 14172 11407 14258
rect 11665 14304 11711 14504
rect 11809 14423 11855 14629
rect 12113 14769 12159 14836
rect 12113 14610 12159 14629
rect 12257 14769 12303 14790
rect 11906 14504 11920 14550
rect 12060 14504 12159 14550
rect 11809 14377 11912 14423
rect 12052 14377 12064 14423
rect 11665 14218 11711 14258
rect 11809 14304 11855 14323
rect 11809 14172 11855 14258
rect 12113 14304 12159 14504
rect 12257 14423 12303 14629
rect 12561 14769 12607 14836
rect 12561 14610 12607 14629
rect 12705 14769 12751 14790
rect 12354 14504 12368 14550
rect 12508 14504 12607 14550
rect 12257 14377 12360 14423
rect 12500 14377 12512 14423
rect 12113 14218 12159 14258
rect 12257 14304 12303 14323
rect 12257 14172 12303 14258
rect 12561 14304 12607 14504
rect 12705 14423 12751 14629
rect 13009 14769 13055 14836
rect 13009 14610 13055 14629
rect 13294 14811 13362 14836
rect 13294 14765 13305 14811
rect 13351 14765 13362 14811
rect 13294 14683 13362 14765
rect 13294 14637 13305 14683
rect 13351 14637 13362 14683
rect 13294 14555 13362 14637
rect 12802 14504 12816 14550
rect 12956 14504 13055 14550
rect 12705 14377 12808 14423
rect 12948 14377 12960 14423
rect 12561 14218 12607 14258
rect 12705 14304 12751 14331
rect 12705 14172 12751 14258
rect 13009 14304 13055 14504
rect 13294 14509 13305 14555
rect 13351 14509 13362 14555
rect 13294 14498 13362 14509
rect 13489 14769 13535 14790
rect 13489 14423 13535 14629
rect 13793 14769 13839 14836
rect 13793 14610 13839 14629
rect 13937 14769 13983 14790
rect 13586 14504 13600 14550
rect 13740 14504 13839 14550
rect 13489 14377 13592 14423
rect 13732 14377 13744 14423
rect 13009 14218 13055 14258
rect 13294 14338 13362 14349
rect 13294 14191 13305 14338
rect 13351 14191 13362 14338
rect 13294 14172 13362 14191
rect 13489 14304 13535 14326
rect 13489 14172 13535 14258
rect 13793 14304 13839 14504
rect 13937 14423 13983 14629
rect 14241 14769 14287 14836
rect 14241 14610 14287 14629
rect 14385 14769 14431 14790
rect 14034 14504 14048 14550
rect 14188 14504 14287 14550
rect 13937 14377 14040 14423
rect 14180 14377 14192 14423
rect 13793 14218 13839 14258
rect 13937 14304 13983 14326
rect 13937 14172 13983 14258
rect 14241 14304 14287 14504
rect 14385 14423 14431 14629
rect 14689 14769 14735 14836
rect 14689 14610 14735 14629
rect 14833 14769 14879 14790
rect 14482 14504 14496 14550
rect 14636 14504 14735 14550
rect 14385 14377 14488 14423
rect 14628 14377 14640 14423
rect 14241 14218 14287 14258
rect 14385 14304 14431 14326
rect 14385 14172 14431 14258
rect 14689 14304 14735 14504
rect 14833 14423 14879 14629
rect 15137 14769 15183 14836
rect 15137 14610 15183 14629
rect 15281 14769 15327 14790
rect 14930 14504 14944 14550
rect 15084 14504 15183 14550
rect 14833 14377 14936 14423
rect 15076 14377 15088 14423
rect 14689 14218 14735 14258
rect 14833 14304 14879 14326
rect 14833 14172 14879 14258
rect 15137 14304 15183 14504
rect 15281 14423 15327 14629
rect 15585 14769 15631 14836
rect 15585 14610 15631 14629
rect 15729 14769 15775 14790
rect 15378 14504 15392 14550
rect 15532 14504 15631 14550
rect 15281 14377 15384 14423
rect 15524 14377 15536 14423
rect 15137 14218 15183 14258
rect 15281 14304 15327 14329
rect 15281 14172 15327 14258
rect 15585 14304 15631 14504
rect 15729 14423 15775 14629
rect 16033 14769 16079 14836
rect 16033 14610 16079 14629
rect 16177 14769 16223 14790
rect 15826 14504 15840 14550
rect 15980 14504 16079 14550
rect 15729 14377 15832 14423
rect 15972 14377 15984 14423
rect 15585 14218 15631 14258
rect 15729 14304 15775 14329
rect 15729 14172 15775 14258
rect 16033 14304 16079 14504
rect 16177 14423 16223 14629
rect 16481 14769 16527 14836
rect 16481 14610 16527 14629
rect 16817 14777 16883 14790
rect 16863 14642 16883 14777
rect 16817 14590 16830 14637
rect 16882 14590 16883 14642
rect 17021 14777 17067 14836
rect 17021 14618 17067 14637
rect 17489 14777 17555 14790
rect 17535 14637 17555 14777
rect 16274 14504 16288 14550
rect 16428 14504 16527 14550
rect 16177 14377 16280 14423
rect 16420 14377 16432 14423
rect 16033 14218 16079 14258
rect 16177 14304 16223 14331
rect 16177 14172 16223 14258
rect 16481 14304 16527 14504
rect 16481 14218 16527 14258
rect 16817 14304 16883 14590
rect 16929 14535 16994 14552
rect 16929 14395 16933 14535
rect 16979 14418 16994 14535
rect 16929 14366 16942 14395
rect 16929 14352 16994 14366
rect 16863 14258 16883 14304
rect 16817 14218 16883 14258
rect 17041 14304 17087 14344
rect 17041 14172 17087 14258
rect 17489 14306 17555 14637
rect 17693 14777 17739 14836
rect 17693 14618 17739 14637
rect 17857 14769 17903 14790
rect 17601 14535 17666 14552
rect 17601 14395 17605 14535
rect 17651 14418 17666 14535
rect 17601 14366 17614 14395
rect 17857 14423 17903 14629
rect 18161 14769 18207 14836
rect 18161 14610 18207 14629
rect 18305 14769 18351 14790
rect 17954 14504 17968 14550
rect 18108 14504 18207 14550
rect 17857 14377 17960 14423
rect 18100 14377 18112 14423
rect 17601 14352 17666 14366
rect 17489 14304 17502 14306
rect 17489 14254 17502 14258
rect 17554 14254 17555 14306
rect 17489 14218 17555 14254
rect 17713 14304 17759 14344
rect 17713 14172 17759 14258
rect 17857 14304 17903 14326
rect 17857 14172 17903 14258
rect 18161 14304 18207 14504
rect 18305 14423 18351 14629
rect 18609 14769 18655 14836
rect 18609 14610 18655 14629
rect 18753 14769 18799 14790
rect 18402 14504 18416 14550
rect 18556 14504 18655 14550
rect 18305 14377 18408 14423
rect 18548 14377 18560 14423
rect 18161 14218 18207 14258
rect 18305 14304 18351 14326
rect 18305 14172 18351 14258
rect 18609 14304 18655 14504
rect 18753 14423 18799 14629
rect 19057 14769 19103 14836
rect 19057 14610 19103 14629
rect 19201 14769 19247 14790
rect 18850 14504 18864 14550
rect 19004 14504 19103 14550
rect 18753 14377 18856 14423
rect 18996 14377 19008 14423
rect 18609 14218 18655 14258
rect 18753 14304 18799 14326
rect 18753 14172 18799 14258
rect 19057 14304 19103 14504
rect 19201 14423 19247 14629
rect 19505 14769 19551 14836
rect 19505 14610 19551 14629
rect 19649 14769 19695 14790
rect 19298 14504 19312 14550
rect 19452 14504 19551 14550
rect 19201 14377 19304 14423
rect 19444 14377 19456 14423
rect 19057 14218 19103 14258
rect 19201 14304 19247 14326
rect 19201 14172 19247 14258
rect 19505 14304 19551 14504
rect 19649 14423 19695 14629
rect 19953 14769 19999 14836
rect 19953 14610 19999 14629
rect 20097 14769 20143 14790
rect 19746 14504 19760 14550
rect 19900 14504 19999 14550
rect 19649 14377 19752 14423
rect 19892 14377 19904 14423
rect 19505 14218 19551 14258
rect 19649 14304 19695 14329
rect 19649 14172 19695 14258
rect 19953 14304 19999 14504
rect 20097 14423 20143 14629
rect 20401 14769 20447 14836
rect 20401 14610 20447 14629
rect 20545 14769 20591 14790
rect 20194 14504 20208 14550
rect 20348 14504 20447 14550
rect 20097 14377 20200 14423
rect 20340 14377 20352 14423
rect 19953 14218 19999 14258
rect 20097 14304 20143 14329
rect 20097 14172 20143 14258
rect 20401 14304 20447 14504
rect 20545 14423 20591 14629
rect 20849 14769 20895 14836
rect 20849 14610 20895 14629
rect 21246 14811 21314 14836
rect 21246 14765 21257 14811
rect 21303 14765 21314 14811
rect 21246 14683 21314 14765
rect 21246 14637 21257 14683
rect 21303 14637 21314 14683
rect 21246 14555 21314 14637
rect 20642 14504 20656 14550
rect 20796 14504 20895 14550
rect 20545 14377 20648 14423
rect 20788 14377 20800 14423
rect 20401 14218 20447 14258
rect 20545 14304 20591 14331
rect 20545 14172 20591 14258
rect 20849 14304 20895 14504
rect 21246 14509 21257 14555
rect 21303 14509 21314 14555
rect 21246 14498 21314 14509
rect 21441 14769 21487 14790
rect 21441 14423 21487 14629
rect 21745 14769 21791 14836
rect 21745 14610 21791 14629
rect 21889 14769 21935 14790
rect 21538 14504 21552 14550
rect 21692 14504 21791 14550
rect 21441 14377 21544 14423
rect 21684 14377 21696 14423
rect 20849 14218 20895 14258
rect 21246 14338 21314 14349
rect 21246 14191 21257 14338
rect 21303 14191 21314 14338
rect 21246 14172 21314 14191
rect 21441 14304 21487 14329
rect 21441 14172 21487 14258
rect 21745 14304 21791 14504
rect 21889 14423 21935 14629
rect 22193 14769 22239 14836
rect 22193 14610 22239 14629
rect 22482 14811 22550 14836
rect 22482 14765 22493 14811
rect 22539 14765 22550 14811
rect 22482 14683 22550 14765
rect 22482 14637 22493 14683
rect 22539 14637 22550 14683
rect 22482 14555 22550 14637
rect 21986 14504 22000 14550
rect 22140 14504 22239 14550
rect 21889 14377 21992 14423
rect 22132 14377 22144 14423
rect 21745 14218 21791 14258
rect 21889 14304 21935 14329
rect 21889 14172 21935 14258
rect 22193 14304 22239 14504
rect 22482 14509 22493 14555
rect 22539 14509 22550 14555
rect 22482 14496 22550 14509
rect 22193 14218 22239 14258
rect 22482 14338 22550 14350
rect 22482 14191 22493 14338
rect 22539 14191 22550 14338
rect 22482 14172 22550 14191
rect 1344 14138 22784 14172
rect 1344 14086 6534 14138
rect 6794 14086 11854 14138
rect 12114 14086 17174 14138
rect 17434 14086 22494 14138
rect 22754 14086 22784 14138
rect 1344 14052 22784 14086
rect 1418 14033 1486 14052
rect 1418 13886 1429 14033
rect 1475 13886 1486 14033
rect 1617 13966 1663 14052
rect 1617 13901 1663 13920
rect 1921 13966 1967 14006
rect 1418 13874 1486 13886
rect 1617 13801 1720 13847
rect 1860 13801 1872 13847
rect 1418 13715 1486 13728
rect 1418 13669 1429 13715
rect 1475 13669 1486 13715
rect 1418 13587 1486 13669
rect 1418 13541 1429 13587
rect 1475 13541 1486 13587
rect 1418 13459 1486 13541
rect 1418 13413 1429 13459
rect 1475 13413 1486 13459
rect 1617 13595 1663 13801
rect 1921 13720 1967 13920
rect 2065 13966 2111 14052
rect 2065 13901 2111 13920
rect 2369 13966 2415 14006
rect 1714 13674 1728 13720
rect 1868 13674 1967 13720
rect 2065 13801 2168 13847
rect 2308 13801 2320 13847
rect 1617 13434 1663 13455
rect 1921 13595 1967 13614
rect 1418 13388 1486 13413
rect 1921 13388 1967 13455
rect 2065 13595 2111 13801
rect 2369 13720 2415 13920
rect 2513 13966 2559 14052
rect 2513 13901 2559 13920
rect 2817 13966 2863 14006
rect 2162 13674 2176 13720
rect 2316 13674 2415 13720
rect 2513 13801 2616 13847
rect 2756 13801 2768 13847
rect 2065 13434 2111 13455
rect 2369 13595 2415 13614
rect 2369 13388 2415 13455
rect 2513 13595 2559 13801
rect 2817 13720 2863 13920
rect 2961 13966 3007 14052
rect 2961 13901 3007 13920
rect 3265 13966 3311 14006
rect 2610 13674 2624 13720
rect 2764 13674 2863 13720
rect 2961 13801 3064 13847
rect 3204 13801 3216 13847
rect 2513 13434 2559 13455
rect 2817 13595 2863 13614
rect 2817 13388 2863 13455
rect 2961 13595 3007 13801
rect 3265 13720 3311 13920
rect 3409 13966 3455 14052
rect 3409 13901 3455 13920
rect 3713 13966 3759 14006
rect 3058 13674 3072 13720
rect 3212 13674 3311 13720
rect 3409 13801 3512 13847
rect 3652 13801 3664 13847
rect 2961 13434 3007 13455
rect 3265 13595 3311 13614
rect 3265 13388 3311 13455
rect 3409 13595 3455 13801
rect 3713 13720 3759 13920
rect 3857 13966 3903 14052
rect 3857 13901 3903 13920
rect 4161 13966 4207 14006
rect 3506 13674 3520 13720
rect 3660 13674 3759 13720
rect 3857 13801 3960 13847
rect 4100 13801 4112 13847
rect 3409 13434 3455 13455
rect 3713 13595 3759 13614
rect 3713 13388 3759 13455
rect 3857 13595 3903 13801
rect 4161 13720 4207 13920
rect 4305 13966 4351 14052
rect 4305 13901 4351 13920
rect 4609 13966 4655 14006
rect 3954 13674 3968 13720
rect 4108 13674 4207 13720
rect 4305 13801 4408 13847
rect 4548 13801 4560 13847
rect 3857 13434 3903 13455
rect 4161 13595 4207 13614
rect 4161 13388 4207 13455
rect 4305 13595 4351 13801
rect 4609 13720 4655 13920
rect 4753 13966 4799 14052
rect 4753 13901 4799 13920
rect 5057 13966 5103 14006
rect 4402 13674 4416 13720
rect 4556 13674 4655 13720
rect 4753 13801 4856 13847
rect 4996 13801 5008 13847
rect 4305 13434 4351 13455
rect 4609 13595 4655 13614
rect 4609 13388 4655 13455
rect 4753 13595 4799 13801
rect 5057 13720 5103 13920
rect 5201 13966 5247 14052
rect 5201 13901 5247 13920
rect 5505 13966 5551 14006
rect 4850 13674 4864 13720
rect 5004 13674 5103 13720
rect 5201 13801 5304 13847
rect 5444 13801 5456 13847
rect 4753 13434 4799 13455
rect 5057 13595 5103 13614
rect 5057 13388 5103 13455
rect 5201 13595 5247 13801
rect 5505 13720 5551 13920
rect 5649 13966 5695 14052
rect 5649 13901 5695 13920
rect 5953 13966 5999 14006
rect 5298 13674 5312 13720
rect 5452 13674 5551 13720
rect 5649 13801 5752 13847
rect 5892 13801 5904 13847
rect 5201 13434 5247 13455
rect 5505 13595 5551 13614
rect 5505 13388 5551 13455
rect 5649 13595 5695 13801
rect 5953 13720 5999 13920
rect 6097 13966 6143 14052
rect 6097 13901 6143 13920
rect 6401 13966 6447 14006
rect 5746 13674 5760 13720
rect 5900 13674 5999 13720
rect 6097 13801 6200 13847
rect 6340 13801 6352 13847
rect 5649 13434 5695 13455
rect 5953 13595 5999 13614
rect 5953 13388 5999 13455
rect 6097 13595 6143 13801
rect 6401 13720 6447 13920
rect 6545 13966 6591 14052
rect 6545 13901 6591 13920
rect 6849 13966 6895 14006
rect 6194 13674 6208 13720
rect 6348 13674 6447 13720
rect 6545 13801 6648 13847
rect 6788 13801 6800 13847
rect 6097 13434 6143 13455
rect 6401 13595 6447 13614
rect 6401 13388 6447 13455
rect 6545 13595 6591 13801
rect 6849 13720 6895 13920
rect 6993 13966 7039 14052
rect 6993 13901 7039 13920
rect 7297 13966 7343 14006
rect 6642 13674 6656 13720
rect 6796 13674 6895 13720
rect 6993 13801 7096 13847
rect 7236 13801 7248 13847
rect 6545 13434 6591 13455
rect 6849 13595 6895 13614
rect 6849 13388 6895 13455
rect 6993 13595 7039 13801
rect 7297 13720 7343 13920
rect 7441 13966 7487 14052
rect 7441 13901 7487 13920
rect 7745 13966 7791 14006
rect 7090 13674 7104 13720
rect 7244 13674 7343 13720
rect 7441 13801 7544 13847
rect 7684 13801 7696 13847
rect 6993 13434 7039 13455
rect 7297 13595 7343 13614
rect 7297 13388 7343 13455
rect 7441 13595 7487 13801
rect 7745 13720 7791 13920
rect 7889 13966 7935 14052
rect 7889 13901 7935 13920
rect 8193 13966 8239 14006
rect 7538 13674 7552 13720
rect 7692 13674 7791 13720
rect 7889 13801 7992 13847
rect 8132 13801 8144 13847
rect 7441 13434 7487 13455
rect 7745 13595 7791 13614
rect 7745 13388 7791 13455
rect 7889 13595 7935 13801
rect 8193 13720 8239 13920
rect 8337 13966 8383 14052
rect 8337 13901 8383 13920
rect 8641 13966 8687 14006
rect 7986 13674 8000 13720
rect 8140 13674 8239 13720
rect 8337 13801 8440 13847
rect 8580 13801 8592 13847
rect 7889 13434 7935 13455
rect 8193 13595 8239 13614
rect 8193 13388 8239 13455
rect 8337 13595 8383 13801
rect 8641 13720 8687 13920
rect 8785 13966 8831 14052
rect 9374 14033 9442 14052
rect 8785 13893 8831 13920
rect 9089 13966 9135 14006
rect 8434 13674 8448 13720
rect 8588 13674 8687 13720
rect 8785 13801 8888 13847
rect 9028 13801 9040 13847
rect 8337 13434 8383 13455
rect 8641 13595 8687 13614
rect 8641 13388 8687 13455
rect 8785 13595 8831 13801
rect 9089 13720 9135 13920
rect 9374 13886 9385 14033
rect 9431 13886 9442 14033
rect 9569 13966 9615 14052
rect 9569 13903 9615 13920
rect 9873 13966 9919 14006
rect 9374 13875 9442 13886
rect 9569 13801 9672 13847
rect 9812 13801 9824 13847
rect 8882 13674 8896 13720
rect 9036 13674 9135 13720
rect 9374 13715 9442 13726
rect 9374 13669 9385 13715
rect 9431 13669 9442 13715
rect 8785 13434 8831 13455
rect 9089 13595 9135 13614
rect 9089 13388 9135 13455
rect 9374 13587 9442 13669
rect 9374 13541 9385 13587
rect 9431 13541 9442 13587
rect 9374 13459 9442 13541
rect 9374 13413 9385 13459
rect 9431 13413 9442 13459
rect 9569 13595 9615 13801
rect 9873 13720 9919 13920
rect 10017 13966 10063 14052
rect 10017 13903 10063 13920
rect 10321 13966 10367 14006
rect 9666 13674 9680 13720
rect 9820 13674 9919 13720
rect 10017 13801 10120 13847
rect 10260 13801 10272 13847
rect 9569 13434 9615 13455
rect 9873 13595 9919 13614
rect 9374 13388 9442 13413
rect 9873 13388 9919 13455
rect 10017 13595 10063 13801
rect 10321 13720 10367 13920
rect 10465 13966 10511 14052
rect 10465 13903 10511 13920
rect 10769 13966 10815 14006
rect 10114 13674 10128 13720
rect 10268 13674 10367 13720
rect 10465 13801 10568 13847
rect 10708 13801 10720 13847
rect 10017 13434 10063 13455
rect 10321 13595 10367 13614
rect 10321 13388 10367 13455
rect 10465 13595 10511 13801
rect 10769 13720 10815 13920
rect 10913 13966 10959 14052
rect 10913 13903 10959 13920
rect 11217 13966 11263 14006
rect 10562 13674 10576 13720
rect 10716 13674 10815 13720
rect 10913 13801 11016 13847
rect 11156 13801 11168 13847
rect 10465 13434 10511 13455
rect 10769 13595 10815 13614
rect 10769 13388 10815 13455
rect 10913 13595 10959 13801
rect 11217 13720 11263 13920
rect 11361 13966 11407 14052
rect 11361 13903 11407 13920
rect 11665 13966 11711 14006
rect 11010 13674 11024 13720
rect 11164 13674 11263 13720
rect 11361 13801 11464 13847
rect 11604 13801 11616 13847
rect 10913 13434 10959 13455
rect 11217 13595 11263 13614
rect 11217 13388 11263 13455
rect 11361 13595 11407 13801
rect 11665 13720 11711 13920
rect 11809 13966 11855 14052
rect 11809 13903 11855 13920
rect 12113 13966 12159 14006
rect 11458 13674 11472 13720
rect 11612 13674 11711 13720
rect 11809 13801 11912 13847
rect 12052 13801 12064 13847
rect 11361 13434 11407 13455
rect 11665 13595 11711 13614
rect 11665 13388 11711 13455
rect 11809 13595 11855 13801
rect 12113 13720 12159 13920
rect 12257 13966 12303 14052
rect 12257 13903 12303 13920
rect 12561 13966 12607 14006
rect 11906 13674 11920 13720
rect 12060 13674 12159 13720
rect 12257 13801 12360 13847
rect 12500 13801 12512 13847
rect 11809 13434 11855 13455
rect 12113 13595 12159 13614
rect 12113 13388 12159 13455
rect 12257 13595 12303 13801
rect 12561 13720 12607 13920
rect 12705 13966 12751 14052
rect 12705 13903 12751 13920
rect 13009 13966 13055 14006
rect 12354 13674 12368 13720
rect 12508 13674 12607 13720
rect 12705 13801 12808 13847
rect 12948 13801 12960 13847
rect 12257 13434 12303 13455
rect 12561 13595 12607 13614
rect 12561 13388 12607 13455
rect 12705 13595 12751 13801
rect 13009 13720 13055 13920
rect 13153 13966 13199 14052
rect 13153 13898 13199 13920
rect 13457 13966 13503 14006
rect 12802 13674 12816 13720
rect 12956 13674 13055 13720
rect 13153 13801 13256 13847
rect 13396 13801 13408 13847
rect 12705 13434 12751 13455
rect 13009 13595 13055 13614
rect 13009 13388 13055 13455
rect 13153 13595 13199 13801
rect 13457 13720 13503 13920
rect 13601 13966 13647 14052
rect 13601 13898 13647 13920
rect 13905 13966 13951 14006
rect 13250 13674 13264 13720
rect 13404 13674 13503 13720
rect 13601 13801 13704 13847
rect 13844 13801 13856 13847
rect 13153 13434 13199 13455
rect 13457 13595 13503 13614
rect 13457 13388 13503 13455
rect 13601 13595 13647 13801
rect 13905 13720 13951 13920
rect 14049 13966 14095 14052
rect 14049 13898 14095 13920
rect 14353 13966 14399 14006
rect 13698 13674 13712 13720
rect 13852 13674 13951 13720
rect 14049 13801 14152 13847
rect 14292 13801 14304 13847
rect 13601 13434 13647 13455
rect 13905 13595 13951 13614
rect 13905 13388 13951 13455
rect 14049 13595 14095 13801
rect 14353 13720 14399 13920
rect 14497 13966 14543 14052
rect 14497 13898 14543 13920
rect 14801 13966 14847 14006
rect 14146 13674 14160 13720
rect 14300 13674 14399 13720
rect 14497 13801 14600 13847
rect 14740 13801 14752 13847
rect 14049 13434 14095 13455
rect 14353 13595 14399 13614
rect 14353 13388 14399 13455
rect 14497 13595 14543 13801
rect 14801 13720 14847 13920
rect 14945 13966 14991 14052
rect 14945 13895 14991 13920
rect 15249 13966 15295 14006
rect 14594 13674 14608 13720
rect 14748 13674 14847 13720
rect 14945 13801 15048 13847
rect 15188 13801 15200 13847
rect 14497 13434 14543 13455
rect 14801 13595 14847 13614
rect 14801 13388 14847 13455
rect 14945 13595 14991 13801
rect 15249 13720 15295 13920
rect 15393 13966 15439 14052
rect 15393 13895 15439 13920
rect 15697 13966 15743 14006
rect 15042 13674 15056 13720
rect 15196 13674 15295 13720
rect 15393 13801 15496 13847
rect 15636 13801 15648 13847
rect 14945 13434 14991 13455
rect 15249 13595 15295 13614
rect 15249 13388 15295 13455
rect 15393 13595 15439 13801
rect 15697 13720 15743 13920
rect 16065 13966 16111 14052
rect 16065 13880 16111 13920
rect 16269 13966 16335 14006
rect 16269 13920 16289 13966
rect 15490 13674 15504 13720
rect 15644 13674 15743 13720
rect 16158 13829 16223 13872
rect 16158 13746 16173 13829
rect 16158 13689 16173 13694
rect 16219 13689 16223 13829
rect 16158 13672 16223 13689
rect 15393 13434 15439 13455
rect 15697 13595 15743 13614
rect 15697 13388 15743 13455
rect 16085 13587 16131 13606
rect 16085 13388 16131 13447
rect 16269 13587 16335 13920
rect 16737 13966 16783 14052
rect 17326 14033 17394 14052
rect 16737 13880 16783 13920
rect 16941 13966 17007 14006
rect 16941 13920 16961 13966
rect 16830 13829 16895 13872
rect 16830 13746 16845 13829
rect 16830 13689 16845 13694
rect 16891 13689 16895 13829
rect 16830 13672 16895 13689
rect 16269 13522 16289 13587
rect 16269 13470 16270 13522
rect 16269 13447 16289 13470
rect 16269 13434 16335 13447
rect 16757 13587 16803 13606
rect 16757 13388 16803 13447
rect 16941 13587 17007 13920
rect 17326 13886 17337 14033
rect 17383 13886 17394 14033
rect 17326 13875 17394 13886
rect 17633 13966 17679 14052
rect 17633 13880 17679 13920
rect 17837 13966 17903 14006
rect 17837 13920 17857 13966
rect 17726 13829 17791 13872
rect 17726 13746 17741 13829
rect 16941 13522 16961 13587
rect 16941 13470 16942 13522
rect 16941 13447 16961 13470
rect 16941 13434 17007 13447
rect 17326 13715 17394 13726
rect 17326 13669 17337 13715
rect 17383 13669 17394 13715
rect 17726 13689 17741 13694
rect 17787 13689 17791 13829
rect 17726 13672 17791 13689
rect 17326 13587 17394 13669
rect 17326 13541 17337 13587
rect 17383 13541 17394 13587
rect 17326 13459 17394 13541
rect 17326 13413 17337 13459
rect 17383 13413 17394 13459
rect 17326 13388 17394 13413
rect 17653 13587 17699 13606
rect 17653 13388 17699 13447
rect 17837 13587 17903 13920
rect 18305 13966 18351 14052
rect 18305 13880 18351 13920
rect 18509 13966 18575 14006
rect 18509 13920 18529 13966
rect 18398 13829 18463 13872
rect 18398 13746 18413 13829
rect 18398 13689 18413 13694
rect 18459 13689 18463 13829
rect 18398 13672 18463 13689
rect 17837 13522 17857 13587
rect 17837 13470 17838 13522
rect 17837 13447 17857 13470
rect 17837 13434 17903 13447
rect 18325 13587 18371 13606
rect 18325 13388 18371 13447
rect 18509 13587 18575 13920
rect 18753 13966 18799 14052
rect 18753 13903 18799 13920
rect 19057 13966 19103 14006
rect 18509 13522 18529 13587
rect 18509 13470 18510 13522
rect 18509 13447 18529 13470
rect 18509 13434 18575 13447
rect 18753 13801 18856 13847
rect 18996 13801 19008 13847
rect 18753 13595 18799 13801
rect 19057 13720 19103 13920
rect 19201 13966 19247 14052
rect 19201 13903 19247 13920
rect 19505 13966 19551 14006
rect 18850 13674 18864 13720
rect 19004 13674 19103 13720
rect 19201 13801 19304 13847
rect 19444 13801 19456 13847
rect 18753 13434 18799 13455
rect 19057 13595 19103 13614
rect 19057 13388 19103 13455
rect 19201 13595 19247 13801
rect 19505 13720 19551 13920
rect 19649 13966 19695 14052
rect 19649 13903 19695 13920
rect 19953 13966 19999 14006
rect 19298 13674 19312 13720
rect 19452 13674 19551 13720
rect 19649 13801 19752 13847
rect 19892 13801 19904 13847
rect 19201 13434 19247 13455
rect 19505 13595 19551 13614
rect 19505 13388 19551 13455
rect 19649 13595 19695 13801
rect 19953 13720 19999 13920
rect 20097 13966 20143 14052
rect 20097 13903 20143 13920
rect 20401 13966 20447 14006
rect 19746 13674 19760 13720
rect 19900 13674 19999 13720
rect 20097 13801 20200 13847
rect 20340 13801 20352 13847
rect 19649 13434 19695 13455
rect 19953 13595 19999 13614
rect 19953 13388 19999 13455
rect 20097 13595 20143 13801
rect 20401 13720 20447 13920
rect 20545 13966 20591 14052
rect 20545 13903 20591 13920
rect 20849 13966 20895 14006
rect 20194 13674 20208 13720
rect 20348 13674 20447 13720
rect 20545 13801 20648 13847
rect 20788 13801 20800 13847
rect 20097 13434 20143 13455
rect 20401 13595 20447 13614
rect 20401 13388 20447 13455
rect 20545 13595 20591 13801
rect 20849 13720 20895 13920
rect 20993 13966 21039 14052
rect 20993 13903 21039 13920
rect 21297 13966 21343 14006
rect 20642 13674 20656 13720
rect 20796 13674 20895 13720
rect 20993 13801 21096 13847
rect 21236 13801 21248 13847
rect 20545 13434 20591 13455
rect 20849 13595 20895 13614
rect 20849 13388 20895 13455
rect 20993 13595 21039 13801
rect 21297 13720 21343 13920
rect 21441 13966 21487 14052
rect 21441 13903 21487 13920
rect 21745 13966 21791 14006
rect 21090 13674 21104 13720
rect 21244 13674 21343 13720
rect 21441 13801 21544 13847
rect 21684 13801 21696 13847
rect 20993 13434 21039 13455
rect 21297 13595 21343 13614
rect 21297 13388 21343 13455
rect 21441 13595 21487 13801
rect 21745 13720 21791 13920
rect 21889 13966 21935 14052
rect 22482 14033 22550 14052
rect 21889 13903 21935 13920
rect 22193 13966 22239 14006
rect 21538 13674 21552 13720
rect 21692 13674 21791 13720
rect 21889 13801 21992 13847
rect 22132 13801 22144 13847
rect 21441 13434 21487 13455
rect 21745 13595 21791 13614
rect 21745 13388 21791 13455
rect 21889 13595 21935 13801
rect 22193 13720 22239 13920
rect 22482 13886 22493 14033
rect 22539 13886 22550 14033
rect 22482 13874 22550 13886
rect 21986 13674 22000 13720
rect 22140 13674 22239 13720
rect 22482 13715 22550 13728
rect 22482 13669 22493 13715
rect 22539 13669 22550 13715
rect 21889 13434 21935 13455
rect 22193 13595 22239 13614
rect 22193 13388 22239 13455
rect 22482 13587 22550 13669
rect 22482 13541 22493 13587
rect 22539 13541 22550 13587
rect 22482 13459 22550 13541
rect 22482 13413 22493 13459
rect 22539 13413 22550 13459
rect 22482 13388 22550 13413
rect 1344 13354 22624 13388
rect 1344 13302 3874 13354
rect 4134 13302 9194 13354
rect 9454 13302 14514 13354
rect 14774 13302 19834 13354
rect 20094 13302 22624 13354
rect 1344 13268 22624 13302
rect 1418 13243 1486 13268
rect 1418 13197 1429 13243
rect 1475 13197 1486 13243
rect 1418 13115 1486 13197
rect 1418 13069 1429 13115
rect 1475 13069 1486 13115
rect 1418 12987 1486 13069
rect 1418 12941 1429 12987
rect 1475 12941 1486 12987
rect 1418 12928 1486 12941
rect 1617 13201 1663 13222
rect 1617 12855 1663 13061
rect 1921 13201 1967 13268
rect 1921 13042 1967 13061
rect 2065 13201 2111 13222
rect 1714 12936 1728 12982
rect 1868 12936 1967 12982
rect 1617 12809 1720 12855
rect 1860 12809 1872 12855
rect 1418 12770 1486 12782
rect 1418 12623 1429 12770
rect 1475 12623 1486 12770
rect 1418 12604 1486 12623
rect 1617 12736 1663 12753
rect 1617 12604 1663 12690
rect 1921 12736 1967 12936
rect 2065 12855 2111 13061
rect 2369 13201 2415 13268
rect 2369 13042 2415 13061
rect 2513 13201 2559 13222
rect 2162 12936 2176 12982
rect 2316 12936 2415 12982
rect 2065 12809 2168 12855
rect 2308 12809 2320 12855
rect 1921 12650 1967 12690
rect 2065 12736 2111 12753
rect 2065 12604 2111 12690
rect 2369 12736 2415 12936
rect 2513 12855 2559 13061
rect 2817 13201 2863 13268
rect 2817 13042 2863 13061
rect 2961 13201 3007 13222
rect 2610 12936 2624 12982
rect 2764 12936 2863 12982
rect 2513 12809 2616 12855
rect 2756 12809 2768 12855
rect 2369 12650 2415 12690
rect 2513 12736 2559 12753
rect 2513 12604 2559 12690
rect 2817 12736 2863 12936
rect 2961 12855 3007 13061
rect 3265 13201 3311 13268
rect 3265 13042 3311 13061
rect 3409 13201 3455 13222
rect 3058 12936 3072 12982
rect 3212 12936 3311 12982
rect 2961 12809 3064 12855
rect 3204 12809 3216 12855
rect 2817 12650 2863 12690
rect 2961 12736 3007 12753
rect 2961 12604 3007 12690
rect 3265 12736 3311 12936
rect 3409 12855 3455 13061
rect 3713 13201 3759 13268
rect 3713 13042 3759 13061
rect 3857 13201 3903 13222
rect 3506 12936 3520 12982
rect 3660 12936 3759 12982
rect 3409 12809 3512 12855
rect 3652 12809 3664 12855
rect 3265 12650 3311 12690
rect 3409 12736 3455 12753
rect 3409 12604 3455 12690
rect 3713 12736 3759 12936
rect 3857 12855 3903 13061
rect 4161 13201 4207 13268
rect 4161 13042 4207 13061
rect 4305 13201 4351 13222
rect 3954 12936 3968 12982
rect 4108 12936 4207 12982
rect 3857 12809 3960 12855
rect 4100 12809 4112 12855
rect 3713 12650 3759 12690
rect 3857 12736 3903 12753
rect 3857 12604 3903 12690
rect 4161 12736 4207 12936
rect 4305 12855 4351 13061
rect 4609 13201 4655 13268
rect 4609 13042 4655 13061
rect 4753 13201 4799 13222
rect 4402 12936 4416 12982
rect 4556 12936 4655 12982
rect 4305 12809 4408 12855
rect 4548 12809 4560 12855
rect 4161 12650 4207 12690
rect 4305 12736 4351 12753
rect 4305 12604 4351 12690
rect 4609 12736 4655 12936
rect 4753 12855 4799 13061
rect 5057 13201 5103 13268
rect 5057 13042 5103 13061
rect 5342 13243 5410 13268
rect 5342 13197 5353 13243
rect 5399 13197 5410 13243
rect 5342 13115 5410 13197
rect 5342 13069 5353 13115
rect 5399 13069 5410 13115
rect 5342 12987 5410 13069
rect 4850 12936 4864 12982
rect 5004 12936 5103 12982
rect 4753 12809 4856 12855
rect 4996 12809 5008 12855
rect 4609 12650 4655 12690
rect 4753 12736 4799 12753
rect 4753 12604 4799 12690
rect 5057 12736 5103 12936
rect 5342 12941 5353 12987
rect 5399 12941 5410 12987
rect 5342 12930 5410 12941
rect 5537 13201 5583 13222
rect 5537 12855 5583 13061
rect 5841 13201 5887 13268
rect 5841 13042 5887 13061
rect 5985 13201 6031 13222
rect 5634 12936 5648 12982
rect 5788 12936 5887 12982
rect 5537 12809 5640 12855
rect 5780 12809 5792 12855
rect 5057 12650 5103 12690
rect 5342 12770 5410 12781
rect 5342 12623 5353 12770
rect 5399 12623 5410 12770
rect 5342 12604 5410 12623
rect 5537 12736 5583 12755
rect 5537 12604 5583 12690
rect 5841 12736 5887 12936
rect 5985 12855 6031 13061
rect 6289 13201 6335 13268
rect 6289 13042 6335 13061
rect 6433 13201 6479 13222
rect 6082 12936 6096 12982
rect 6236 12936 6335 12982
rect 5985 12809 6088 12855
rect 6228 12809 6240 12855
rect 5841 12650 5887 12690
rect 5985 12736 6031 12755
rect 5985 12604 6031 12690
rect 6289 12736 6335 12936
rect 6433 12855 6479 13061
rect 6737 13201 6783 13268
rect 6737 13042 6783 13061
rect 6881 13201 6927 13222
rect 6530 12936 6544 12982
rect 6684 12936 6783 12982
rect 6433 12809 6536 12855
rect 6676 12809 6688 12855
rect 6289 12650 6335 12690
rect 6433 12736 6479 12755
rect 6433 12604 6479 12690
rect 6737 12736 6783 12936
rect 6881 12855 6927 13061
rect 7185 13201 7231 13268
rect 7185 13042 7231 13061
rect 7329 13201 7375 13222
rect 6978 12936 6992 12982
rect 7132 12936 7231 12982
rect 6881 12809 6984 12855
rect 7124 12809 7136 12855
rect 6737 12650 6783 12690
rect 6881 12736 6927 12755
rect 6881 12604 6927 12690
rect 7185 12736 7231 12936
rect 7329 12855 7375 13061
rect 7633 13201 7679 13268
rect 7633 13042 7679 13061
rect 7777 13201 7823 13222
rect 7426 12936 7440 12982
rect 7580 12936 7679 12982
rect 7329 12809 7432 12855
rect 7572 12809 7584 12855
rect 7185 12650 7231 12690
rect 7329 12736 7375 12755
rect 7329 12604 7375 12690
rect 7633 12736 7679 12936
rect 7777 12855 7823 13061
rect 8081 13201 8127 13268
rect 8081 13042 8127 13061
rect 8225 13201 8271 13222
rect 7874 12936 7888 12982
rect 8028 12936 8127 12982
rect 7777 12809 7880 12855
rect 8020 12809 8032 12855
rect 7633 12650 7679 12690
rect 7777 12736 7823 12755
rect 7777 12604 7823 12690
rect 8081 12736 8127 12936
rect 8225 12855 8271 13061
rect 8529 13201 8575 13268
rect 8529 13042 8575 13061
rect 8673 13201 8719 13222
rect 8322 12936 8336 12982
rect 8476 12936 8575 12982
rect 8225 12809 8328 12855
rect 8468 12809 8480 12855
rect 8081 12650 8127 12690
rect 8225 12736 8271 12755
rect 8225 12604 8271 12690
rect 8529 12736 8575 12936
rect 8673 12855 8719 13061
rect 8977 13201 9023 13268
rect 8977 13042 9023 13061
rect 9121 13201 9167 13222
rect 8770 12936 8784 12982
rect 8924 12936 9023 12982
rect 8673 12809 8776 12855
rect 8916 12809 8928 12855
rect 8529 12650 8575 12690
rect 8673 12736 8719 12755
rect 8673 12604 8719 12690
rect 8977 12736 9023 12936
rect 9121 12855 9167 13061
rect 9425 13201 9471 13268
rect 9425 13042 9471 13061
rect 9569 13201 9615 13222
rect 9218 12936 9232 12982
rect 9372 12936 9471 12982
rect 9121 12809 9224 12855
rect 9364 12809 9376 12855
rect 8977 12650 9023 12690
rect 9121 12736 9167 12755
rect 9121 12604 9167 12690
rect 9425 12736 9471 12936
rect 9569 12855 9615 13061
rect 9873 13201 9919 13268
rect 9873 13042 9919 13061
rect 10017 13201 10063 13222
rect 9666 12936 9680 12982
rect 9820 12936 9919 12982
rect 9569 12809 9672 12855
rect 9812 12809 9824 12855
rect 9425 12650 9471 12690
rect 9569 12736 9615 12755
rect 9569 12604 9615 12690
rect 9873 12736 9919 12936
rect 10017 12855 10063 13061
rect 10321 13201 10367 13268
rect 10321 13042 10367 13061
rect 10465 13201 10511 13222
rect 10114 12936 10128 12982
rect 10268 12936 10367 12982
rect 10017 12809 10120 12855
rect 10260 12809 10272 12855
rect 9873 12650 9919 12690
rect 10017 12736 10063 12755
rect 10017 12604 10063 12690
rect 10321 12736 10367 12936
rect 10465 12855 10511 13061
rect 10769 13201 10815 13268
rect 10769 13042 10815 13061
rect 10913 13201 10959 13222
rect 10562 12936 10576 12982
rect 10716 12936 10815 12982
rect 10465 12809 10568 12855
rect 10708 12809 10720 12855
rect 10321 12650 10367 12690
rect 10465 12736 10511 12755
rect 10465 12604 10511 12690
rect 10769 12736 10815 12936
rect 10913 12855 10959 13061
rect 11217 13201 11263 13268
rect 11217 13042 11263 13061
rect 11361 13201 11407 13222
rect 11010 12936 11024 12982
rect 11164 12936 11263 12982
rect 10913 12809 11016 12855
rect 11156 12809 11168 12855
rect 10769 12650 10815 12690
rect 10913 12736 10959 12755
rect 10913 12604 10959 12690
rect 11217 12736 11263 12936
rect 11361 12855 11407 13061
rect 11665 13201 11711 13268
rect 11665 13042 11711 13061
rect 11809 13201 11855 13222
rect 11458 12936 11472 12982
rect 11612 12936 11711 12982
rect 11361 12809 11464 12855
rect 11604 12809 11616 12855
rect 11217 12650 11263 12690
rect 11361 12736 11407 12755
rect 11361 12604 11407 12690
rect 11665 12736 11711 12936
rect 11809 12855 11855 13061
rect 12113 13201 12159 13268
rect 12113 13042 12159 13061
rect 12257 13201 12303 13222
rect 11906 12936 11920 12982
rect 12060 12936 12159 12982
rect 11809 12809 11912 12855
rect 12052 12809 12064 12855
rect 11665 12650 11711 12690
rect 11809 12736 11855 12755
rect 11809 12604 11855 12690
rect 12113 12736 12159 12936
rect 12257 12855 12303 13061
rect 12561 13201 12607 13268
rect 12561 13042 12607 13061
rect 12705 13201 12751 13222
rect 12354 12936 12368 12982
rect 12508 12936 12607 12982
rect 12257 12809 12360 12855
rect 12500 12809 12512 12855
rect 12113 12650 12159 12690
rect 12257 12736 12303 12755
rect 12257 12604 12303 12690
rect 12561 12736 12607 12936
rect 12705 12855 12751 13061
rect 13009 13201 13055 13268
rect 13009 13042 13055 13061
rect 13294 13243 13362 13268
rect 13294 13197 13305 13243
rect 13351 13197 13362 13243
rect 13294 13115 13362 13197
rect 13294 13069 13305 13115
rect 13351 13069 13362 13115
rect 13294 12987 13362 13069
rect 12802 12936 12816 12982
rect 12956 12936 13055 12982
rect 12705 12809 12808 12855
rect 12948 12809 12960 12855
rect 12561 12650 12607 12690
rect 12705 12736 12751 12763
rect 12705 12604 12751 12690
rect 13009 12736 13055 12936
rect 13294 12941 13305 12987
rect 13351 12941 13362 12987
rect 13294 12930 13362 12941
rect 13489 13201 13535 13222
rect 13489 12855 13535 13061
rect 13793 13201 13839 13268
rect 13793 13042 13839 13061
rect 13937 13201 13983 13222
rect 13586 12936 13600 12982
rect 13740 12936 13839 12982
rect 13489 12809 13592 12855
rect 13732 12809 13744 12855
rect 13009 12650 13055 12690
rect 13294 12770 13362 12781
rect 13294 12623 13305 12770
rect 13351 12623 13362 12770
rect 13294 12604 13362 12623
rect 13489 12736 13535 12761
rect 13489 12604 13535 12690
rect 13793 12736 13839 12936
rect 13937 12855 13983 13061
rect 14241 13201 14287 13268
rect 14241 13042 14287 13061
rect 14741 13209 14787 13268
rect 14741 13050 14787 13069
rect 14925 13209 14991 13222
rect 14925 13186 14945 13209
rect 14925 13134 14926 13186
rect 14925 13069 14945 13134
rect 14034 12936 14048 12982
rect 14188 12936 14287 12982
rect 13937 12809 14040 12855
rect 14180 12809 14192 12855
rect 13793 12650 13839 12690
rect 13937 12736 13983 12761
rect 13937 12604 13983 12690
rect 14241 12736 14287 12936
rect 14814 12967 14879 12984
rect 14814 12850 14829 12967
rect 14875 12827 14879 12967
rect 14866 12798 14879 12827
rect 14814 12784 14879 12798
rect 14241 12650 14287 12690
rect 14721 12736 14767 12776
rect 14721 12604 14767 12690
rect 14925 12736 14991 13069
rect 15413 13209 15459 13268
rect 15413 13050 15459 13069
rect 15597 13209 15663 13222
rect 15597 13069 15617 13209
rect 15486 12967 15551 12984
rect 15486 12850 15501 12967
rect 15547 12827 15551 12967
rect 15538 12798 15551 12827
rect 15486 12784 15551 12798
rect 14925 12690 14945 12736
rect 14925 12650 14991 12690
rect 15393 12736 15439 12776
rect 15393 12604 15439 12690
rect 15597 12738 15663 13069
rect 16085 13209 16131 13268
rect 16085 13050 16131 13069
rect 16269 13209 16335 13222
rect 16269 13069 16289 13209
rect 16158 12967 16223 12984
rect 16158 12850 16173 12967
rect 16219 12827 16223 12967
rect 16210 12798 16223 12827
rect 16158 12784 16223 12798
rect 15597 12686 15598 12738
rect 15650 12736 15663 12738
rect 15650 12686 15663 12690
rect 15597 12650 15663 12686
rect 16065 12736 16111 12776
rect 16065 12604 16111 12690
rect 16269 12738 16335 13069
rect 16757 13209 16803 13268
rect 16757 13050 16803 13069
rect 16941 13209 17007 13222
rect 16941 13069 16961 13209
rect 16830 12967 16895 12984
rect 16830 12850 16845 12967
rect 16891 12827 16895 12967
rect 16882 12798 16895 12827
rect 16830 12784 16895 12798
rect 16269 12686 16270 12738
rect 16322 12736 16335 12738
rect 16322 12686 16335 12690
rect 16269 12650 16335 12686
rect 16737 12736 16783 12776
rect 16737 12604 16783 12690
rect 16941 12738 17007 13069
rect 17429 13209 17475 13268
rect 17429 13050 17475 13069
rect 17613 13209 17679 13222
rect 17613 13069 17633 13209
rect 17502 12967 17567 12984
rect 17502 12962 17517 12967
rect 17502 12827 17517 12910
rect 17563 12827 17567 12967
rect 17502 12784 17567 12827
rect 16941 12686 16942 12738
rect 16994 12736 17007 12738
rect 16994 12686 17007 12690
rect 16941 12650 17007 12686
rect 17409 12736 17455 12776
rect 17409 12604 17455 12690
rect 17613 12738 17679 13069
rect 18101 13209 18147 13268
rect 18101 13050 18147 13069
rect 18285 13209 18351 13222
rect 18285 13186 18305 13209
rect 18285 13134 18286 13186
rect 18285 13069 18305 13134
rect 18174 12967 18239 12984
rect 18174 12850 18189 12967
rect 18235 12827 18239 12967
rect 18226 12798 18239 12827
rect 18174 12784 18239 12798
rect 17613 12686 17614 12738
rect 17666 12736 17679 12738
rect 17666 12686 17679 12690
rect 17613 12650 17679 12686
rect 18081 12736 18127 12776
rect 18081 12604 18127 12690
rect 18285 12736 18351 13069
rect 18773 13209 18819 13268
rect 18773 13050 18819 13069
rect 18957 13209 19023 13222
rect 18957 13186 18977 13209
rect 18957 13134 18958 13186
rect 18957 13069 18977 13134
rect 18846 12967 18911 12984
rect 18846 12962 18861 12967
rect 18846 12827 18861 12910
rect 18907 12827 18911 12967
rect 18846 12784 18911 12827
rect 18285 12690 18305 12736
rect 18285 12650 18351 12690
rect 18753 12736 18799 12776
rect 18753 12604 18799 12690
rect 18957 12736 19023 13069
rect 19445 13209 19491 13268
rect 19445 13050 19491 13069
rect 19629 13209 19695 13222
rect 19629 13069 19649 13209
rect 19518 12967 19583 12984
rect 19518 12850 19533 12967
rect 19579 12827 19583 12967
rect 19570 12798 19583 12827
rect 19518 12784 19583 12798
rect 18957 12690 18977 12736
rect 18957 12650 19023 12690
rect 19425 12736 19471 12776
rect 19425 12604 19471 12690
rect 19629 12738 19695 13069
rect 19873 13201 19919 13222
rect 19873 12855 19919 13061
rect 20177 13201 20223 13268
rect 20177 13042 20223 13061
rect 20321 13201 20367 13222
rect 19970 12936 19984 12982
rect 20124 12936 20223 12982
rect 19873 12809 19976 12855
rect 20116 12809 20128 12855
rect 19629 12686 19630 12738
rect 19682 12736 19695 12738
rect 19682 12686 19695 12690
rect 19629 12650 19695 12686
rect 19873 12736 19919 12761
rect 19873 12604 19919 12690
rect 20177 12736 20223 12936
rect 20321 12855 20367 13061
rect 20625 13201 20671 13268
rect 20625 13042 20671 13061
rect 20769 13201 20815 13222
rect 20418 12936 20432 12982
rect 20572 12936 20671 12982
rect 20321 12809 20424 12855
rect 20564 12809 20576 12855
rect 20177 12650 20223 12690
rect 20321 12736 20367 12761
rect 20321 12604 20367 12690
rect 20625 12736 20671 12936
rect 20769 12855 20815 13061
rect 21073 13201 21119 13268
rect 21073 13042 21119 13061
rect 21246 13243 21314 13268
rect 21246 13197 21257 13243
rect 21303 13197 21314 13243
rect 21246 13115 21314 13197
rect 21246 13069 21257 13115
rect 21303 13069 21314 13115
rect 21246 12987 21314 13069
rect 20866 12936 20880 12982
rect 21020 12936 21119 12982
rect 20769 12809 20872 12855
rect 21012 12809 21024 12855
rect 20625 12650 20671 12690
rect 20769 12736 20815 12763
rect 20769 12604 20815 12690
rect 21073 12736 21119 12936
rect 21246 12941 21257 12987
rect 21303 12941 21314 12987
rect 21246 12930 21314 12941
rect 21441 13201 21487 13222
rect 21441 12855 21487 13061
rect 21745 13201 21791 13268
rect 21745 13042 21791 13061
rect 21889 13201 21935 13222
rect 21538 12936 21552 12982
rect 21692 12936 21791 12982
rect 21441 12809 21544 12855
rect 21684 12809 21696 12855
rect 21073 12650 21119 12690
rect 21246 12770 21314 12781
rect 21246 12623 21257 12770
rect 21303 12623 21314 12770
rect 21246 12604 21314 12623
rect 21441 12736 21487 12761
rect 21441 12604 21487 12690
rect 21745 12736 21791 12936
rect 21889 12855 21935 13061
rect 22193 13201 22239 13268
rect 22193 13042 22239 13061
rect 22482 13243 22550 13268
rect 22482 13197 22493 13243
rect 22539 13197 22550 13243
rect 22482 13115 22550 13197
rect 22482 13069 22493 13115
rect 22539 13069 22550 13115
rect 22482 12987 22550 13069
rect 21986 12936 22000 12982
rect 22140 12936 22239 12982
rect 21889 12809 21992 12855
rect 22132 12809 22144 12855
rect 21745 12650 21791 12690
rect 21889 12736 21935 12761
rect 21889 12604 21935 12690
rect 22193 12736 22239 12936
rect 22482 12941 22493 12987
rect 22539 12941 22550 12987
rect 22482 12928 22550 12941
rect 22193 12650 22239 12690
rect 22482 12770 22550 12782
rect 22482 12623 22493 12770
rect 22539 12623 22550 12770
rect 22482 12604 22550 12623
rect 1344 12570 22784 12604
rect 1344 12518 6534 12570
rect 6794 12518 11854 12570
rect 12114 12518 17174 12570
rect 17434 12518 22494 12570
rect 22754 12518 22784 12570
rect 1344 12484 22784 12518
rect 1418 12465 1486 12484
rect 1418 12318 1429 12465
rect 1475 12318 1486 12465
rect 1617 12398 1663 12484
rect 1617 12333 1663 12352
rect 1921 12398 1967 12438
rect 1418 12306 1486 12318
rect 1617 12233 1720 12279
rect 1860 12233 1872 12279
rect 1418 12147 1486 12160
rect 1418 12101 1429 12147
rect 1475 12101 1486 12147
rect 1418 12019 1486 12101
rect 1418 11973 1429 12019
rect 1475 11973 1486 12019
rect 1418 11891 1486 11973
rect 1418 11845 1429 11891
rect 1475 11845 1486 11891
rect 1617 12027 1663 12233
rect 1921 12152 1967 12352
rect 2065 12398 2111 12484
rect 2065 12333 2111 12352
rect 2369 12398 2415 12438
rect 1714 12106 1728 12152
rect 1868 12106 1967 12152
rect 2065 12233 2168 12279
rect 2308 12233 2320 12279
rect 1617 11866 1663 11887
rect 1921 12027 1967 12046
rect 1418 11820 1486 11845
rect 1921 11820 1967 11887
rect 2065 12027 2111 12233
rect 2369 12152 2415 12352
rect 2513 12398 2559 12484
rect 2513 12333 2559 12352
rect 2817 12398 2863 12438
rect 2162 12106 2176 12152
rect 2316 12106 2415 12152
rect 2513 12233 2616 12279
rect 2756 12233 2768 12279
rect 2065 11866 2111 11887
rect 2369 12027 2415 12046
rect 2369 11820 2415 11887
rect 2513 12027 2559 12233
rect 2817 12152 2863 12352
rect 2961 12398 3007 12484
rect 2961 12333 3007 12352
rect 3265 12398 3311 12438
rect 2610 12106 2624 12152
rect 2764 12106 2863 12152
rect 2961 12233 3064 12279
rect 3204 12233 3216 12279
rect 2513 11866 2559 11887
rect 2817 12027 2863 12046
rect 2817 11820 2863 11887
rect 2961 12027 3007 12233
rect 3265 12152 3311 12352
rect 3409 12398 3455 12484
rect 3409 12333 3455 12352
rect 3713 12398 3759 12438
rect 3058 12106 3072 12152
rect 3212 12106 3311 12152
rect 3409 12233 3512 12279
rect 3652 12233 3664 12279
rect 2961 11866 3007 11887
rect 3265 12027 3311 12046
rect 3265 11820 3311 11887
rect 3409 12027 3455 12233
rect 3713 12152 3759 12352
rect 3857 12398 3903 12484
rect 3857 12333 3903 12352
rect 4161 12398 4207 12438
rect 3506 12106 3520 12152
rect 3660 12106 3759 12152
rect 3857 12233 3960 12279
rect 4100 12233 4112 12279
rect 3409 11866 3455 11887
rect 3713 12027 3759 12046
rect 3713 11820 3759 11887
rect 3857 12027 3903 12233
rect 4161 12152 4207 12352
rect 4305 12398 4351 12484
rect 4305 12333 4351 12352
rect 4609 12398 4655 12438
rect 3954 12106 3968 12152
rect 4108 12106 4207 12152
rect 4305 12233 4408 12279
rect 4548 12233 4560 12279
rect 3857 11866 3903 11887
rect 4161 12027 4207 12046
rect 4161 11820 4207 11887
rect 4305 12027 4351 12233
rect 4609 12152 4655 12352
rect 4753 12398 4799 12484
rect 4753 12333 4799 12352
rect 5057 12398 5103 12438
rect 4402 12106 4416 12152
rect 4556 12106 4655 12152
rect 4753 12233 4856 12279
rect 4996 12233 5008 12279
rect 4305 11866 4351 11887
rect 4609 12027 4655 12046
rect 4609 11820 4655 11887
rect 4753 12027 4799 12233
rect 5057 12152 5103 12352
rect 5201 12398 5247 12484
rect 5201 12333 5247 12352
rect 5505 12398 5551 12438
rect 4850 12106 4864 12152
rect 5004 12106 5103 12152
rect 5201 12233 5304 12279
rect 5444 12233 5456 12279
rect 4753 11866 4799 11887
rect 5057 12027 5103 12046
rect 5057 11820 5103 11887
rect 5201 12027 5247 12233
rect 5505 12152 5551 12352
rect 5649 12398 5695 12484
rect 5649 12333 5695 12352
rect 5953 12398 5999 12438
rect 5298 12106 5312 12152
rect 5452 12106 5551 12152
rect 5649 12233 5752 12279
rect 5892 12233 5904 12279
rect 5201 11866 5247 11887
rect 5505 12027 5551 12046
rect 5505 11820 5551 11887
rect 5649 12027 5695 12233
rect 5953 12152 5999 12352
rect 6097 12398 6143 12484
rect 6097 12333 6143 12352
rect 6401 12398 6447 12438
rect 5746 12106 5760 12152
rect 5900 12106 5999 12152
rect 6097 12233 6200 12279
rect 6340 12233 6352 12279
rect 5649 11866 5695 11887
rect 5953 12027 5999 12046
rect 5953 11820 5999 11887
rect 6097 12027 6143 12233
rect 6401 12152 6447 12352
rect 6545 12398 6591 12484
rect 6545 12333 6591 12352
rect 6849 12398 6895 12438
rect 6194 12106 6208 12152
rect 6348 12106 6447 12152
rect 6545 12233 6648 12279
rect 6788 12233 6800 12279
rect 6097 11866 6143 11887
rect 6401 12027 6447 12046
rect 6401 11820 6447 11887
rect 6545 12027 6591 12233
rect 6849 12152 6895 12352
rect 6993 12398 7039 12484
rect 6993 12333 7039 12352
rect 7297 12398 7343 12438
rect 6642 12106 6656 12152
rect 6796 12106 6895 12152
rect 6993 12233 7096 12279
rect 7236 12233 7248 12279
rect 6545 11866 6591 11887
rect 6849 12027 6895 12046
rect 6849 11820 6895 11887
rect 6993 12027 7039 12233
rect 7297 12152 7343 12352
rect 7441 12398 7487 12484
rect 7441 12333 7487 12352
rect 7745 12398 7791 12438
rect 7090 12106 7104 12152
rect 7244 12106 7343 12152
rect 7441 12233 7544 12279
rect 7684 12233 7696 12279
rect 6993 11866 7039 11887
rect 7297 12027 7343 12046
rect 7297 11820 7343 11887
rect 7441 12027 7487 12233
rect 7745 12152 7791 12352
rect 7889 12398 7935 12484
rect 7889 12333 7935 12352
rect 8193 12398 8239 12438
rect 7538 12106 7552 12152
rect 7692 12106 7791 12152
rect 7889 12233 7992 12279
rect 8132 12233 8144 12279
rect 7441 11866 7487 11887
rect 7745 12027 7791 12046
rect 7745 11820 7791 11887
rect 7889 12027 7935 12233
rect 8193 12152 8239 12352
rect 8337 12398 8383 12484
rect 8337 12333 8383 12352
rect 8641 12398 8687 12438
rect 7986 12106 8000 12152
rect 8140 12106 8239 12152
rect 8337 12233 8440 12279
rect 8580 12233 8592 12279
rect 7889 11866 7935 11887
rect 8193 12027 8239 12046
rect 8193 11820 8239 11887
rect 8337 12027 8383 12233
rect 8641 12152 8687 12352
rect 8785 12398 8831 12484
rect 9374 12465 9442 12484
rect 8785 12325 8831 12352
rect 9089 12398 9135 12438
rect 8434 12106 8448 12152
rect 8588 12106 8687 12152
rect 8785 12233 8888 12279
rect 9028 12233 9040 12279
rect 8337 11866 8383 11887
rect 8641 12027 8687 12046
rect 8641 11820 8687 11887
rect 8785 12027 8831 12233
rect 9089 12152 9135 12352
rect 9374 12318 9385 12465
rect 9431 12318 9442 12465
rect 9569 12398 9615 12484
rect 9569 12335 9615 12352
rect 9873 12398 9919 12438
rect 9374 12307 9442 12318
rect 9569 12233 9672 12279
rect 9812 12233 9824 12279
rect 8882 12106 8896 12152
rect 9036 12106 9135 12152
rect 9374 12147 9442 12158
rect 9374 12101 9385 12147
rect 9431 12101 9442 12147
rect 8785 11866 8831 11887
rect 9089 12027 9135 12046
rect 9089 11820 9135 11887
rect 9374 12019 9442 12101
rect 9374 11973 9385 12019
rect 9431 11973 9442 12019
rect 9374 11891 9442 11973
rect 9374 11845 9385 11891
rect 9431 11845 9442 11891
rect 9569 12027 9615 12233
rect 9873 12152 9919 12352
rect 10017 12398 10063 12484
rect 10017 12335 10063 12352
rect 10321 12398 10367 12438
rect 9666 12106 9680 12152
rect 9820 12106 9919 12152
rect 10017 12233 10120 12279
rect 10260 12233 10272 12279
rect 9569 11866 9615 11887
rect 9873 12027 9919 12046
rect 9374 11820 9442 11845
rect 9873 11820 9919 11887
rect 10017 12027 10063 12233
rect 10321 12152 10367 12352
rect 10465 12398 10511 12484
rect 10465 12335 10511 12352
rect 10769 12398 10815 12438
rect 10114 12106 10128 12152
rect 10268 12106 10367 12152
rect 10465 12233 10568 12279
rect 10708 12233 10720 12279
rect 10017 11866 10063 11887
rect 10321 12027 10367 12046
rect 10321 11820 10367 11887
rect 10465 12027 10511 12233
rect 10769 12152 10815 12352
rect 10913 12398 10959 12484
rect 10913 12335 10959 12352
rect 11217 12398 11263 12438
rect 10562 12106 10576 12152
rect 10716 12106 10815 12152
rect 10913 12233 11016 12279
rect 11156 12233 11168 12279
rect 10465 11866 10511 11887
rect 10769 12027 10815 12046
rect 10769 11820 10815 11887
rect 10913 12027 10959 12233
rect 11217 12152 11263 12352
rect 11361 12398 11407 12484
rect 11361 12335 11407 12352
rect 11665 12398 11711 12438
rect 11010 12106 11024 12152
rect 11164 12106 11263 12152
rect 11361 12233 11464 12279
rect 11604 12233 11616 12279
rect 10913 11866 10959 11887
rect 11217 12027 11263 12046
rect 11217 11820 11263 11887
rect 11361 12027 11407 12233
rect 11665 12152 11711 12352
rect 11809 12398 11855 12484
rect 11809 12335 11855 12352
rect 12113 12398 12159 12438
rect 11458 12106 11472 12152
rect 11612 12106 11711 12152
rect 11809 12233 11912 12279
rect 12052 12233 12064 12279
rect 11361 11866 11407 11887
rect 11665 12027 11711 12046
rect 11665 11820 11711 11887
rect 11809 12027 11855 12233
rect 12113 12152 12159 12352
rect 12257 12398 12303 12484
rect 12257 12335 12303 12352
rect 12561 12398 12607 12438
rect 11906 12106 11920 12152
rect 12060 12106 12159 12152
rect 12257 12233 12360 12279
rect 12500 12233 12512 12279
rect 11809 11866 11855 11887
rect 12113 12027 12159 12046
rect 12113 11820 12159 11887
rect 12257 12027 12303 12233
rect 12561 12152 12607 12352
rect 12705 12398 12751 12484
rect 12705 12335 12751 12352
rect 13009 12398 13055 12438
rect 12354 12106 12368 12152
rect 12508 12106 12607 12152
rect 12705 12233 12808 12279
rect 12948 12233 12960 12279
rect 12257 11866 12303 11887
rect 12561 12027 12607 12046
rect 12561 11820 12607 11887
rect 12705 12027 12751 12233
rect 13009 12152 13055 12352
rect 13153 12398 13199 12484
rect 13153 12327 13199 12352
rect 13457 12398 13503 12438
rect 12802 12106 12816 12152
rect 12956 12106 13055 12152
rect 13153 12233 13256 12279
rect 13396 12233 13408 12279
rect 12705 11866 12751 11887
rect 13009 12027 13055 12046
rect 13009 11820 13055 11887
rect 13153 12027 13199 12233
rect 13457 12152 13503 12352
rect 13601 12398 13647 12484
rect 13601 12327 13647 12352
rect 13905 12398 13951 12438
rect 13250 12106 13264 12152
rect 13404 12106 13503 12152
rect 13601 12233 13704 12279
rect 13844 12233 13856 12279
rect 13153 11866 13199 11887
rect 13457 12027 13503 12046
rect 13457 11820 13503 11887
rect 13601 12027 13647 12233
rect 13905 12152 13951 12352
rect 14049 12398 14095 12484
rect 14049 12312 14095 12352
rect 14253 12398 14319 12438
rect 14253 12352 14273 12398
rect 13698 12106 13712 12152
rect 13852 12106 13951 12152
rect 14142 12261 14207 12304
rect 14142 12178 14157 12261
rect 14142 12121 14157 12126
rect 14203 12121 14207 12261
rect 14142 12104 14207 12121
rect 13601 11866 13647 11887
rect 13905 12027 13951 12046
rect 13905 11820 13951 11887
rect 14069 12019 14115 12038
rect 14069 11820 14115 11879
rect 14253 12019 14319 12352
rect 14721 12398 14767 12484
rect 14721 12312 14767 12352
rect 14925 12398 14991 12438
rect 14925 12352 14945 12398
rect 14814 12261 14879 12304
rect 14814 12178 14829 12261
rect 14814 12121 14829 12126
rect 14875 12121 14879 12261
rect 14814 12104 14879 12121
rect 14253 11954 14273 12019
rect 14253 11902 14254 11954
rect 14253 11879 14273 11902
rect 14253 11866 14319 11879
rect 14741 12019 14787 12038
rect 14741 11820 14787 11879
rect 14925 12019 14991 12352
rect 15393 12398 15439 12484
rect 15393 12312 15439 12352
rect 15597 12398 15663 12438
rect 15597 12352 15617 12398
rect 15486 12261 15551 12304
rect 15486 12178 15501 12261
rect 15486 12121 15501 12126
rect 15547 12121 15551 12261
rect 15486 12104 15551 12121
rect 14925 11954 14945 12019
rect 14925 11902 14926 11954
rect 14925 11879 14945 11902
rect 14925 11866 14991 11879
rect 15413 12019 15459 12038
rect 15413 11820 15459 11879
rect 15597 12019 15663 12352
rect 16065 12398 16111 12484
rect 16065 12312 16111 12352
rect 16269 12398 16335 12438
rect 16269 12352 16289 12398
rect 16158 12261 16223 12304
rect 16158 12178 16173 12261
rect 16158 12121 16173 12126
rect 16219 12121 16223 12261
rect 16158 12104 16223 12121
rect 15597 11954 15617 12019
rect 15597 11902 15598 11954
rect 15597 11879 15617 11902
rect 15597 11866 15663 11879
rect 16085 12019 16131 12038
rect 16085 11820 16131 11879
rect 16269 12019 16335 12352
rect 16737 12398 16783 12484
rect 17326 12465 17394 12484
rect 16737 12312 16783 12352
rect 16941 12398 17007 12438
rect 16941 12352 16961 12398
rect 16830 12261 16895 12304
rect 16830 12178 16845 12261
rect 16830 12121 16845 12126
rect 16891 12121 16895 12261
rect 16830 12104 16895 12121
rect 16269 11954 16289 12019
rect 16269 11902 16270 11954
rect 16269 11879 16289 11902
rect 16269 11866 16335 11879
rect 16757 12019 16803 12038
rect 16757 11820 16803 11879
rect 16941 12019 17007 12352
rect 17326 12318 17337 12465
rect 17383 12318 17394 12465
rect 17326 12307 17394 12318
rect 17633 12398 17679 12484
rect 17633 12312 17679 12352
rect 17837 12398 17903 12438
rect 17837 12352 17857 12398
rect 17726 12290 17791 12304
rect 17778 12261 17791 12290
rect 16941 11954 16961 12019
rect 16941 11902 16942 11954
rect 16941 11879 16961 11902
rect 16941 11866 17007 11879
rect 17326 12147 17394 12158
rect 17326 12101 17337 12147
rect 17383 12101 17394 12147
rect 17726 12121 17741 12238
rect 17787 12121 17791 12261
rect 17726 12104 17791 12121
rect 17837 12290 17903 12352
rect 18305 12398 18351 12484
rect 18305 12312 18351 12352
rect 18509 12398 18575 12438
rect 18509 12352 18529 12398
rect 17837 12238 17838 12290
rect 17890 12238 17903 12290
rect 17326 12019 17394 12101
rect 17326 11973 17337 12019
rect 17383 11973 17394 12019
rect 17326 11891 17394 11973
rect 17326 11845 17337 11891
rect 17383 11845 17394 11891
rect 17326 11820 17394 11845
rect 17653 12019 17699 12038
rect 17653 11820 17699 11879
rect 17837 12019 17903 12238
rect 18398 12290 18463 12304
rect 18450 12261 18463 12290
rect 18398 12121 18413 12238
rect 18459 12121 18463 12261
rect 18398 12104 18463 12121
rect 17837 11879 17857 12019
rect 17837 11866 17903 11879
rect 18325 12019 18371 12038
rect 18325 11820 18371 11879
rect 18509 12019 18575 12352
rect 18977 12398 19023 12484
rect 18977 12312 19023 12352
rect 19181 12402 19247 12438
rect 19181 12350 19182 12402
rect 19234 12398 19247 12402
rect 19234 12350 19247 12352
rect 19070 12290 19135 12304
rect 19122 12261 19135 12290
rect 19070 12121 19085 12238
rect 19131 12121 19135 12261
rect 19070 12104 19135 12121
rect 18509 11954 18529 12019
rect 18509 11902 18510 11954
rect 18509 11879 18529 11902
rect 18509 11866 18575 11879
rect 18997 12019 19043 12038
rect 18997 11820 19043 11879
rect 19181 12019 19247 12350
rect 19649 12398 19695 12484
rect 19649 12312 19695 12352
rect 19853 12402 19919 12438
rect 19853 12350 19854 12402
rect 19906 12398 19919 12402
rect 19906 12350 19919 12352
rect 19742 12290 19807 12304
rect 19794 12261 19807 12290
rect 19742 12121 19757 12238
rect 19803 12121 19807 12261
rect 19742 12104 19807 12121
rect 19181 11879 19201 12019
rect 19181 11866 19247 11879
rect 19669 12019 19715 12038
rect 19669 11820 19715 11879
rect 19853 12019 19919 12350
rect 20321 12398 20367 12484
rect 20321 12312 20367 12352
rect 20525 12398 20591 12438
rect 20525 12352 20545 12398
rect 20414 12290 20479 12304
rect 20466 12261 20479 12290
rect 20414 12121 20429 12238
rect 20475 12121 20479 12261
rect 20414 12104 20479 12121
rect 20525 12290 20591 12352
rect 20769 12398 20815 12484
rect 20769 12327 20815 12352
rect 21073 12398 21119 12438
rect 20525 12238 20526 12290
rect 20578 12238 20591 12290
rect 19853 11879 19873 12019
rect 19853 11866 19919 11879
rect 20341 12019 20387 12038
rect 20341 11820 20387 11879
rect 20525 12019 20591 12238
rect 20525 11879 20545 12019
rect 20525 11866 20591 11879
rect 20769 12233 20872 12279
rect 21012 12233 21024 12279
rect 20769 12027 20815 12233
rect 21073 12152 21119 12352
rect 21217 12398 21263 12484
rect 21217 12327 21263 12352
rect 21521 12398 21567 12438
rect 20866 12106 20880 12152
rect 21020 12106 21119 12152
rect 21217 12233 21320 12279
rect 21460 12233 21472 12279
rect 20769 11866 20815 11887
rect 21073 12027 21119 12046
rect 21073 11820 21119 11887
rect 21217 12027 21263 12233
rect 21521 12152 21567 12352
rect 21665 12398 21711 12484
rect 22482 12465 22550 12484
rect 21665 12325 21711 12352
rect 21969 12398 22015 12438
rect 21314 12106 21328 12152
rect 21468 12106 21567 12152
rect 21665 12233 21768 12279
rect 21908 12233 21920 12279
rect 21217 11866 21263 11887
rect 21521 12027 21567 12046
rect 21521 11820 21567 11887
rect 21665 12027 21711 12233
rect 21969 12152 22015 12352
rect 22482 12318 22493 12465
rect 22539 12318 22550 12465
rect 22482 12306 22550 12318
rect 21762 12106 21776 12152
rect 21916 12106 22015 12152
rect 22482 12147 22550 12160
rect 22482 12101 22493 12147
rect 22539 12101 22550 12147
rect 21665 11866 21711 11887
rect 21969 12027 22015 12046
rect 21969 11820 22015 11887
rect 22482 12019 22550 12101
rect 22482 11973 22493 12019
rect 22539 11973 22550 12019
rect 22482 11891 22550 11973
rect 22482 11845 22493 11891
rect 22539 11845 22550 11891
rect 22482 11820 22550 11845
rect 1344 11786 22624 11820
rect 1344 11734 3874 11786
rect 4134 11734 9194 11786
rect 9454 11734 14514 11786
rect 14774 11734 19834 11786
rect 20094 11734 22624 11786
rect 1344 11700 22624 11734
rect 1418 11675 1486 11700
rect 1418 11629 1429 11675
rect 1475 11629 1486 11675
rect 1418 11547 1486 11629
rect 1418 11501 1429 11547
rect 1475 11501 1486 11547
rect 1418 11419 1486 11501
rect 1418 11373 1429 11419
rect 1475 11373 1486 11419
rect 1418 11360 1486 11373
rect 1617 11633 1663 11654
rect 1617 11287 1663 11493
rect 1921 11633 1967 11700
rect 1921 11474 1967 11493
rect 2065 11633 2111 11654
rect 1714 11368 1728 11414
rect 1868 11368 1967 11414
rect 1617 11241 1720 11287
rect 1860 11241 1872 11287
rect 1418 11202 1486 11214
rect 1418 11055 1429 11202
rect 1475 11055 1486 11202
rect 1418 11036 1486 11055
rect 1617 11168 1663 11185
rect 1617 11036 1663 11122
rect 1921 11168 1967 11368
rect 2065 11287 2111 11493
rect 2369 11633 2415 11700
rect 2369 11474 2415 11493
rect 2513 11633 2559 11654
rect 2162 11368 2176 11414
rect 2316 11368 2415 11414
rect 2065 11241 2168 11287
rect 2308 11241 2320 11287
rect 1921 11082 1967 11122
rect 2065 11168 2111 11185
rect 2065 11036 2111 11122
rect 2369 11168 2415 11368
rect 2513 11287 2559 11493
rect 2817 11633 2863 11700
rect 2817 11474 2863 11493
rect 2961 11633 3007 11654
rect 2610 11368 2624 11414
rect 2764 11368 2863 11414
rect 2513 11241 2616 11287
rect 2756 11241 2768 11287
rect 2369 11082 2415 11122
rect 2513 11168 2559 11185
rect 2513 11036 2559 11122
rect 2817 11168 2863 11368
rect 2961 11287 3007 11493
rect 3265 11633 3311 11700
rect 3265 11474 3311 11493
rect 3409 11633 3455 11654
rect 3058 11368 3072 11414
rect 3212 11368 3311 11414
rect 2961 11241 3064 11287
rect 3204 11241 3216 11287
rect 2817 11082 2863 11122
rect 2961 11168 3007 11185
rect 2961 11036 3007 11122
rect 3265 11168 3311 11368
rect 3409 11287 3455 11493
rect 3713 11633 3759 11700
rect 3713 11474 3759 11493
rect 3857 11633 3903 11654
rect 3506 11368 3520 11414
rect 3660 11368 3759 11414
rect 3409 11241 3512 11287
rect 3652 11241 3664 11287
rect 3265 11082 3311 11122
rect 3409 11168 3455 11185
rect 3409 11036 3455 11122
rect 3713 11168 3759 11368
rect 3857 11287 3903 11493
rect 4161 11633 4207 11700
rect 4161 11474 4207 11493
rect 4305 11633 4351 11654
rect 3954 11368 3968 11414
rect 4108 11368 4207 11414
rect 3857 11241 3960 11287
rect 4100 11241 4112 11287
rect 3713 11082 3759 11122
rect 3857 11168 3903 11185
rect 3857 11036 3903 11122
rect 4161 11168 4207 11368
rect 4305 11287 4351 11493
rect 4609 11633 4655 11700
rect 4609 11474 4655 11493
rect 4753 11633 4799 11654
rect 4402 11368 4416 11414
rect 4556 11368 4655 11414
rect 4305 11241 4408 11287
rect 4548 11241 4560 11287
rect 4161 11082 4207 11122
rect 4305 11168 4351 11185
rect 4305 11036 4351 11122
rect 4609 11168 4655 11368
rect 4753 11287 4799 11493
rect 5057 11633 5103 11700
rect 5057 11474 5103 11493
rect 5342 11675 5410 11700
rect 5342 11629 5353 11675
rect 5399 11629 5410 11675
rect 5342 11547 5410 11629
rect 5342 11501 5353 11547
rect 5399 11501 5410 11547
rect 5342 11419 5410 11501
rect 4850 11368 4864 11414
rect 5004 11368 5103 11414
rect 4753 11241 4856 11287
rect 4996 11241 5008 11287
rect 4609 11082 4655 11122
rect 4753 11168 4799 11185
rect 4753 11036 4799 11122
rect 5057 11168 5103 11368
rect 5342 11373 5353 11419
rect 5399 11373 5410 11419
rect 5342 11362 5410 11373
rect 5537 11633 5583 11654
rect 5537 11287 5583 11493
rect 5841 11633 5887 11700
rect 5841 11474 5887 11493
rect 6065 11641 6131 11654
rect 6111 11501 6131 11641
rect 5634 11368 5648 11414
rect 5788 11368 5887 11414
rect 5537 11241 5640 11287
rect 5780 11241 5792 11287
rect 5057 11082 5103 11122
rect 5342 11202 5410 11213
rect 5342 11055 5353 11202
rect 5399 11055 5410 11202
rect 5342 11036 5410 11055
rect 5537 11168 5583 11195
rect 5537 11036 5583 11122
rect 5841 11168 5887 11368
rect 5841 11082 5887 11122
rect 6065 11282 6131 11501
rect 6269 11641 6315 11700
rect 6269 11482 6315 11501
rect 6849 11641 6915 11654
rect 6895 11501 6915 11641
rect 6065 11230 6078 11282
rect 6130 11230 6131 11282
rect 6065 11168 6131 11230
rect 6177 11399 6242 11416
rect 6177 11259 6181 11399
rect 6227 11282 6242 11399
rect 6177 11230 6190 11259
rect 6177 11216 6242 11230
rect 6111 11122 6131 11168
rect 6065 11082 6131 11122
rect 6289 11168 6335 11208
rect 6289 11036 6335 11122
rect 6849 11170 6915 11501
rect 7053 11641 7099 11700
rect 7053 11482 7099 11501
rect 7521 11641 7587 11654
rect 7567 11501 7587 11641
rect 6961 11399 7026 11416
rect 6961 11259 6965 11399
rect 7011 11282 7026 11399
rect 6961 11230 6974 11259
rect 6961 11216 7026 11230
rect 6849 11168 6862 11170
rect 6849 11118 6862 11122
rect 6914 11118 6915 11170
rect 6849 11082 6915 11118
rect 7073 11168 7119 11208
rect 7073 11036 7119 11122
rect 7521 11170 7587 11501
rect 7725 11641 7771 11700
rect 7725 11482 7771 11501
rect 8193 11641 8259 11654
rect 8239 11501 8259 11641
rect 7633 11399 7698 11416
rect 7633 11259 7637 11399
rect 7683 11282 7698 11399
rect 7633 11230 7646 11259
rect 7633 11216 7698 11230
rect 7521 11168 7534 11170
rect 7521 11118 7534 11122
rect 7586 11118 7587 11170
rect 7521 11082 7587 11118
rect 7745 11168 7791 11208
rect 7745 11036 7791 11122
rect 8193 11170 8259 11501
rect 8397 11641 8443 11700
rect 8397 11482 8443 11501
rect 8561 11633 8607 11654
rect 8305 11399 8370 11416
rect 8305 11259 8309 11399
rect 8355 11282 8370 11399
rect 8305 11230 8318 11259
rect 8561 11287 8607 11493
rect 8865 11633 8911 11700
rect 8865 11474 8911 11493
rect 9141 11641 9187 11700
rect 9141 11482 9187 11501
rect 9325 11641 9391 11654
rect 9325 11501 9345 11641
rect 8658 11368 8672 11414
rect 8812 11368 8911 11414
rect 8561 11241 8664 11287
rect 8804 11241 8816 11287
rect 8305 11216 8370 11230
rect 8193 11168 8206 11170
rect 8193 11118 8206 11122
rect 8258 11118 8259 11170
rect 8193 11082 8259 11118
rect 8417 11168 8463 11208
rect 8417 11036 8463 11122
rect 8561 11168 8607 11195
rect 8561 11036 8607 11122
rect 8865 11168 8911 11368
rect 9214 11399 9279 11416
rect 9214 11282 9229 11399
rect 9275 11259 9279 11399
rect 9266 11230 9279 11259
rect 9214 11216 9279 11230
rect 8865 11082 8911 11122
rect 9121 11168 9167 11208
rect 9121 11036 9167 11122
rect 9325 11170 9391 11501
rect 9813 11641 9859 11700
rect 9813 11482 9859 11501
rect 9997 11641 10063 11654
rect 9997 11501 10017 11641
rect 9886 11399 9951 11416
rect 9886 11282 9901 11399
rect 9947 11259 9951 11399
rect 9938 11230 9951 11259
rect 9886 11216 9951 11230
rect 9325 11118 9326 11170
rect 9378 11168 9391 11170
rect 9378 11118 9391 11122
rect 9325 11082 9391 11118
rect 9793 11168 9839 11208
rect 9793 11036 9839 11122
rect 9997 11170 10063 11501
rect 10485 11641 10531 11700
rect 10485 11482 10531 11501
rect 10669 11641 10735 11654
rect 10669 11506 10689 11641
rect 10669 11454 10670 11506
rect 10722 11454 10735 11501
rect 10558 11399 10623 11416
rect 10558 11282 10573 11399
rect 10619 11259 10623 11399
rect 10610 11230 10623 11259
rect 10558 11216 10623 11230
rect 9997 11118 9998 11170
rect 10050 11168 10063 11170
rect 10050 11118 10063 11122
rect 9997 11082 10063 11118
rect 10465 11168 10511 11208
rect 10465 11036 10511 11122
rect 10669 11168 10735 11454
rect 10913 11633 10959 11654
rect 10913 11287 10959 11493
rect 11217 11633 11263 11700
rect 11217 11474 11263 11493
rect 11361 11633 11407 11654
rect 11010 11368 11024 11414
rect 11164 11368 11263 11414
rect 10913 11241 11016 11287
rect 11156 11241 11168 11287
rect 10669 11122 10689 11168
rect 10669 11082 10735 11122
rect 10913 11168 10959 11193
rect 10913 11036 10959 11122
rect 11217 11168 11263 11368
rect 11361 11287 11407 11493
rect 11665 11633 11711 11700
rect 11665 11474 11711 11493
rect 12053 11641 12099 11700
rect 12053 11482 12099 11501
rect 12237 11641 12303 11654
rect 12237 11501 12257 11641
rect 11458 11368 11472 11414
rect 11612 11368 11711 11414
rect 11361 11241 11464 11287
rect 11604 11241 11616 11287
rect 11217 11082 11263 11122
rect 11361 11168 11407 11193
rect 11361 11036 11407 11122
rect 11665 11168 11711 11368
rect 12126 11399 12191 11416
rect 12126 11282 12141 11399
rect 12187 11259 12191 11399
rect 12178 11230 12191 11259
rect 12126 11216 12191 11230
rect 12237 11282 12303 11501
rect 12725 11641 12771 11700
rect 13294 11675 13362 11700
rect 12725 11482 12771 11501
rect 12909 11641 12975 11654
rect 12909 11501 12929 11641
rect 12237 11230 12238 11282
rect 12290 11230 12303 11282
rect 11665 11082 11711 11122
rect 12033 11168 12079 11208
rect 12033 11036 12079 11122
rect 12237 11168 12303 11230
rect 12798 11399 12863 11416
rect 12798 11282 12813 11399
rect 12859 11259 12863 11399
rect 12850 11230 12863 11259
rect 12798 11216 12863 11230
rect 12237 11122 12257 11168
rect 12237 11082 12303 11122
rect 12705 11168 12751 11208
rect 12705 11036 12751 11122
rect 12909 11170 12975 11501
rect 13294 11629 13305 11675
rect 13351 11629 13362 11675
rect 13294 11547 13362 11629
rect 13294 11501 13305 11547
rect 13351 11501 13362 11547
rect 13294 11419 13362 11501
rect 13621 11641 13667 11700
rect 13621 11482 13667 11501
rect 13805 11641 13871 11654
rect 13805 11501 13825 11641
rect 13294 11373 13305 11419
rect 13351 11373 13362 11419
rect 13294 11362 13362 11373
rect 13694 11399 13759 11416
rect 13694 11282 13709 11399
rect 13755 11259 13759 11399
rect 13746 11230 13759 11259
rect 13694 11216 13759 11230
rect 12909 11118 12910 11170
rect 12962 11168 12975 11170
rect 12962 11118 12975 11122
rect 12909 11082 12975 11118
rect 13294 11202 13362 11213
rect 13294 11055 13305 11202
rect 13351 11055 13362 11202
rect 13294 11036 13362 11055
rect 13601 11168 13647 11208
rect 13601 11036 13647 11122
rect 13805 11170 13871 11501
rect 14049 11633 14095 11654
rect 14049 11287 14095 11493
rect 14353 11633 14399 11700
rect 14353 11474 14399 11493
rect 14741 11641 14787 11700
rect 14741 11482 14787 11501
rect 14925 11641 14991 11654
rect 14925 11501 14945 11641
rect 14146 11368 14160 11414
rect 14300 11368 14399 11414
rect 14049 11241 14152 11287
rect 14292 11241 14304 11287
rect 13805 11118 13806 11170
rect 13858 11168 13871 11170
rect 13858 11118 13871 11122
rect 13805 11082 13871 11118
rect 14049 11168 14095 11195
rect 14049 11036 14095 11122
rect 14353 11168 14399 11368
rect 14814 11399 14879 11416
rect 14814 11282 14829 11399
rect 14875 11259 14879 11399
rect 14866 11230 14879 11259
rect 14814 11216 14879 11230
rect 14925 11394 14991 11501
rect 15413 11641 15459 11700
rect 15413 11482 15459 11501
rect 15597 11641 15663 11654
rect 15597 11501 15617 11641
rect 14925 11342 14926 11394
rect 14978 11342 14991 11394
rect 14353 11082 14399 11122
rect 14721 11168 14767 11208
rect 14721 11036 14767 11122
rect 14925 11168 14991 11342
rect 15486 11399 15551 11416
rect 15486 11282 15501 11399
rect 15547 11259 15551 11399
rect 15538 11230 15551 11259
rect 15486 11216 15551 11230
rect 15597 11394 15663 11501
rect 16085 11641 16131 11700
rect 16085 11482 16131 11501
rect 16269 11641 16335 11654
rect 16269 11501 16289 11641
rect 15597 11342 15598 11394
rect 15650 11342 15663 11394
rect 14925 11122 14945 11168
rect 14925 11082 14991 11122
rect 15393 11168 15439 11208
rect 15393 11036 15439 11122
rect 15597 11168 15663 11342
rect 16158 11399 16223 11416
rect 16158 11282 16173 11399
rect 16219 11259 16223 11399
rect 16210 11230 16223 11259
rect 16158 11216 16223 11230
rect 16269 11394 16335 11501
rect 16757 11641 16803 11700
rect 16757 11482 16803 11501
rect 16941 11641 17007 11654
rect 16941 11501 16961 11641
rect 16269 11342 16270 11394
rect 16322 11342 16335 11394
rect 15597 11122 15617 11168
rect 15597 11082 15663 11122
rect 16065 11168 16111 11208
rect 16065 11036 16111 11122
rect 16269 11168 16335 11342
rect 16830 11399 16895 11416
rect 16830 11394 16845 11399
rect 16830 11259 16845 11342
rect 16891 11259 16895 11399
rect 16830 11216 16895 11259
rect 16941 11394 17007 11501
rect 17429 11641 17475 11700
rect 17429 11482 17475 11501
rect 17613 11641 17679 11654
rect 17613 11618 17633 11641
rect 17613 11566 17614 11618
rect 17613 11501 17633 11566
rect 16941 11342 16942 11394
rect 16994 11342 17007 11394
rect 16269 11122 16289 11168
rect 16269 11082 16335 11122
rect 16737 11168 16783 11208
rect 16737 11036 16783 11122
rect 16941 11168 17007 11342
rect 17502 11399 17567 11416
rect 17502 11394 17517 11399
rect 17502 11259 17517 11342
rect 17563 11259 17567 11399
rect 17502 11216 17567 11259
rect 16941 11122 16961 11168
rect 16941 11082 17007 11122
rect 17409 11168 17455 11208
rect 17409 11036 17455 11122
rect 17613 11168 17679 11501
rect 18101 11641 18147 11700
rect 18101 11482 18147 11501
rect 18285 11641 18351 11654
rect 18285 11501 18305 11641
rect 18174 11399 18239 11416
rect 18174 11394 18189 11399
rect 18174 11259 18189 11342
rect 18235 11259 18239 11399
rect 18174 11216 18239 11259
rect 17613 11122 17633 11168
rect 17613 11082 17679 11122
rect 18081 11168 18127 11208
rect 18081 11036 18127 11122
rect 18285 11170 18351 11501
rect 18773 11641 18819 11700
rect 18773 11482 18819 11501
rect 18957 11641 19023 11654
rect 18957 11501 18977 11641
rect 18846 11399 18911 11416
rect 18846 11394 18861 11399
rect 18846 11259 18861 11342
rect 18907 11259 18911 11399
rect 18846 11216 18911 11259
rect 18285 11118 18286 11170
rect 18338 11168 18351 11170
rect 18338 11118 18351 11122
rect 18285 11082 18351 11118
rect 18753 11168 18799 11208
rect 18753 11036 18799 11122
rect 18957 11170 19023 11501
rect 19445 11641 19491 11700
rect 19445 11482 19491 11501
rect 19629 11641 19695 11654
rect 19629 11618 19649 11641
rect 19629 11566 19630 11618
rect 19629 11501 19649 11566
rect 19518 11399 19583 11416
rect 19518 11394 19533 11399
rect 19518 11259 19533 11342
rect 19579 11259 19583 11399
rect 19518 11216 19583 11259
rect 18957 11118 18958 11170
rect 19010 11168 19023 11170
rect 19010 11118 19023 11122
rect 18957 11082 19023 11118
rect 19425 11168 19471 11208
rect 19425 11036 19471 11122
rect 19629 11168 19695 11501
rect 20117 11641 20163 11700
rect 20117 11482 20163 11501
rect 20301 11641 20367 11654
rect 20301 11501 20321 11641
rect 20190 11399 20255 11416
rect 20190 11282 20205 11399
rect 20251 11259 20255 11399
rect 20242 11230 20255 11259
rect 20190 11216 20255 11230
rect 19629 11122 19649 11168
rect 19629 11082 19695 11122
rect 20097 11168 20143 11208
rect 20097 11036 20143 11122
rect 20301 11170 20367 11501
rect 20545 11633 20591 11654
rect 20545 11287 20591 11493
rect 20849 11633 20895 11700
rect 20849 11474 20895 11493
rect 21246 11675 21314 11700
rect 21246 11629 21257 11675
rect 21303 11629 21314 11675
rect 21246 11547 21314 11629
rect 21246 11501 21257 11547
rect 21303 11501 21314 11547
rect 21246 11419 21314 11501
rect 20642 11368 20656 11414
rect 20796 11368 20895 11414
rect 20545 11241 20648 11287
rect 20788 11241 20800 11287
rect 20301 11118 20302 11170
rect 20354 11168 20367 11170
rect 20354 11118 20367 11122
rect 20301 11082 20367 11118
rect 20545 11168 20591 11195
rect 20545 11036 20591 11122
rect 20849 11168 20895 11368
rect 21246 11373 21257 11419
rect 21303 11373 21314 11419
rect 21246 11362 21314 11373
rect 21441 11633 21487 11654
rect 21441 11287 21487 11493
rect 21745 11633 21791 11700
rect 21745 11474 21791 11493
rect 21889 11633 21935 11654
rect 21538 11368 21552 11414
rect 21692 11368 21791 11414
rect 21441 11241 21544 11287
rect 21684 11241 21696 11287
rect 20849 11082 20895 11122
rect 21246 11202 21314 11213
rect 21246 11055 21257 11202
rect 21303 11055 21314 11202
rect 21246 11036 21314 11055
rect 21441 11168 21487 11193
rect 21441 11036 21487 11122
rect 21745 11168 21791 11368
rect 21889 11287 21935 11493
rect 22193 11633 22239 11700
rect 22193 11474 22239 11493
rect 22482 11675 22550 11700
rect 22482 11629 22493 11675
rect 22539 11629 22550 11675
rect 22482 11547 22550 11629
rect 22482 11501 22493 11547
rect 22539 11501 22550 11547
rect 22482 11419 22550 11501
rect 21986 11368 22000 11414
rect 22140 11368 22239 11414
rect 21889 11241 21992 11287
rect 22132 11241 22144 11287
rect 21745 11082 21791 11122
rect 21889 11168 21935 11193
rect 21889 11036 21935 11122
rect 22193 11168 22239 11368
rect 22482 11373 22493 11419
rect 22539 11373 22550 11419
rect 22482 11360 22550 11373
rect 22193 11082 22239 11122
rect 22482 11202 22550 11214
rect 22482 11055 22493 11202
rect 22539 11055 22550 11202
rect 22482 11036 22550 11055
rect 1344 11002 22784 11036
rect 1344 10950 6534 11002
rect 6794 10950 11854 11002
rect 12114 10950 17174 11002
rect 17434 10950 22494 11002
rect 22754 10950 22784 11002
rect 1344 10916 22784 10950
rect 1418 10897 1486 10916
rect 1418 10750 1429 10897
rect 1475 10750 1486 10897
rect 1617 10830 1663 10916
rect 1617 10767 1663 10784
rect 1921 10830 1967 10870
rect 1418 10738 1486 10750
rect 1617 10665 1720 10711
rect 1860 10665 1872 10711
rect 1418 10579 1486 10592
rect 1418 10533 1429 10579
rect 1475 10533 1486 10579
rect 1418 10451 1486 10533
rect 1418 10405 1429 10451
rect 1475 10405 1486 10451
rect 1418 10323 1486 10405
rect 1418 10277 1429 10323
rect 1475 10277 1486 10323
rect 1617 10459 1663 10665
rect 1921 10584 1967 10784
rect 2065 10830 2111 10916
rect 2065 10767 2111 10784
rect 2369 10830 2415 10870
rect 1714 10538 1728 10584
rect 1868 10538 1967 10584
rect 2065 10665 2168 10711
rect 2308 10665 2320 10711
rect 1617 10298 1663 10319
rect 1921 10459 1967 10478
rect 1418 10252 1486 10277
rect 1921 10252 1967 10319
rect 2065 10459 2111 10665
rect 2369 10584 2415 10784
rect 2513 10830 2559 10916
rect 2513 10767 2559 10784
rect 2817 10830 2863 10870
rect 2162 10538 2176 10584
rect 2316 10538 2415 10584
rect 2513 10665 2616 10711
rect 2756 10665 2768 10711
rect 2065 10298 2111 10319
rect 2369 10459 2415 10478
rect 2369 10252 2415 10319
rect 2513 10459 2559 10665
rect 2817 10584 2863 10784
rect 2961 10830 3007 10916
rect 2961 10767 3007 10784
rect 3265 10830 3311 10870
rect 2610 10538 2624 10584
rect 2764 10538 2863 10584
rect 2961 10665 3064 10711
rect 3204 10665 3216 10711
rect 2513 10298 2559 10319
rect 2817 10459 2863 10478
rect 2817 10252 2863 10319
rect 2961 10459 3007 10665
rect 3265 10584 3311 10784
rect 3409 10830 3455 10916
rect 3409 10767 3455 10784
rect 3713 10830 3759 10870
rect 3058 10538 3072 10584
rect 3212 10538 3311 10584
rect 3409 10665 3512 10711
rect 3652 10665 3664 10711
rect 2961 10298 3007 10319
rect 3265 10459 3311 10478
rect 3265 10252 3311 10319
rect 3409 10459 3455 10665
rect 3713 10584 3759 10784
rect 3857 10830 3903 10916
rect 3857 10767 3903 10784
rect 4161 10830 4207 10870
rect 3506 10538 3520 10584
rect 3660 10538 3759 10584
rect 3857 10665 3960 10711
rect 4100 10665 4112 10711
rect 3409 10298 3455 10319
rect 3713 10459 3759 10478
rect 3713 10252 3759 10319
rect 3857 10459 3903 10665
rect 4161 10584 4207 10784
rect 4305 10830 4351 10916
rect 4305 10767 4351 10784
rect 4609 10830 4655 10870
rect 3954 10538 3968 10584
rect 4108 10538 4207 10584
rect 4305 10665 4408 10711
rect 4548 10665 4560 10711
rect 3857 10298 3903 10319
rect 4161 10459 4207 10478
rect 4161 10252 4207 10319
rect 4305 10459 4351 10665
rect 4609 10584 4655 10784
rect 4753 10830 4799 10916
rect 4753 10767 4799 10784
rect 5057 10830 5103 10870
rect 4402 10538 4416 10584
rect 4556 10538 4655 10584
rect 4753 10665 4856 10711
rect 4996 10665 5008 10711
rect 4305 10298 4351 10319
rect 4609 10459 4655 10478
rect 4609 10252 4655 10319
rect 4753 10459 4799 10665
rect 5057 10584 5103 10784
rect 5313 10830 5359 10916
rect 5313 10744 5359 10784
rect 5517 10830 5583 10870
rect 5517 10784 5537 10830
rect 4850 10538 4864 10584
rect 5004 10538 5103 10584
rect 5406 10722 5471 10736
rect 5458 10693 5471 10722
rect 5406 10553 5421 10670
rect 5467 10553 5471 10693
rect 5406 10536 5471 10553
rect 5517 10722 5583 10784
rect 5985 10830 6031 10916
rect 5985 10744 6031 10784
rect 6189 10830 6255 10870
rect 6189 10784 6209 10830
rect 5517 10670 5518 10722
rect 5570 10670 5583 10722
rect 4753 10298 4799 10319
rect 5057 10459 5103 10478
rect 5057 10252 5103 10319
rect 5333 10451 5379 10470
rect 5333 10252 5379 10311
rect 5517 10451 5583 10670
rect 6078 10722 6143 10736
rect 6130 10693 6143 10722
rect 6078 10553 6093 10670
rect 6139 10553 6143 10693
rect 6078 10536 6143 10553
rect 5517 10311 5537 10451
rect 5517 10298 5583 10311
rect 6005 10451 6051 10470
rect 6005 10252 6051 10311
rect 6189 10451 6255 10784
rect 6657 10830 6703 10916
rect 6657 10744 6703 10784
rect 6861 10834 6927 10870
rect 6861 10782 6862 10834
rect 6914 10830 6927 10834
rect 6914 10782 6927 10784
rect 6750 10693 6815 10736
rect 6750 10610 6765 10693
rect 6750 10553 6765 10558
rect 6811 10553 6815 10693
rect 6750 10536 6815 10553
rect 6189 10386 6209 10451
rect 6189 10334 6190 10386
rect 6189 10311 6209 10334
rect 6189 10298 6255 10311
rect 6677 10451 6723 10470
rect 6677 10252 6723 10311
rect 6861 10451 6927 10782
rect 7329 10830 7375 10916
rect 7329 10744 7375 10784
rect 7533 10830 7599 10870
rect 7533 10784 7553 10830
rect 7422 10693 7487 10736
rect 7422 10610 7437 10693
rect 7422 10553 7437 10558
rect 7483 10553 7487 10693
rect 7422 10536 7487 10553
rect 7533 10610 7599 10784
rect 8001 10830 8047 10916
rect 8001 10744 8047 10784
rect 8205 10830 8271 10870
rect 8205 10784 8225 10830
rect 7533 10558 7534 10610
rect 7586 10558 7599 10610
rect 6861 10311 6881 10451
rect 6861 10298 6927 10311
rect 7349 10451 7395 10470
rect 7349 10252 7395 10311
rect 7533 10451 7599 10558
rect 8094 10722 8159 10736
rect 8146 10693 8159 10722
rect 8094 10553 8109 10670
rect 8155 10553 8159 10693
rect 8094 10536 8159 10553
rect 7533 10311 7553 10451
rect 7533 10298 7599 10311
rect 8021 10451 8067 10470
rect 8021 10252 8067 10311
rect 8205 10451 8271 10784
rect 8785 10830 8831 10916
rect 9374 10897 9442 10916
rect 8785 10744 8831 10784
rect 8989 10830 9055 10870
rect 8989 10784 9009 10830
rect 8878 10693 8943 10736
rect 8878 10610 8893 10693
rect 8878 10553 8893 10558
rect 8939 10553 8943 10693
rect 8878 10536 8943 10553
rect 8205 10386 8225 10451
rect 8205 10334 8206 10386
rect 8205 10311 8225 10334
rect 8205 10298 8271 10311
rect 8805 10451 8851 10470
rect 8805 10252 8851 10311
rect 8989 10451 9055 10784
rect 9374 10750 9385 10897
rect 9431 10750 9442 10897
rect 9374 10739 9442 10750
rect 9793 10830 9839 10916
rect 9793 10744 9839 10784
rect 9997 10830 10063 10870
rect 9997 10784 10017 10830
rect 9886 10693 9951 10736
rect 9886 10610 9901 10693
rect 8989 10386 9009 10451
rect 8989 10334 8990 10386
rect 8989 10311 9009 10334
rect 8989 10298 9055 10311
rect 9374 10579 9442 10590
rect 9374 10533 9385 10579
rect 9431 10533 9442 10579
rect 9886 10553 9901 10558
rect 9947 10553 9951 10693
rect 9886 10536 9951 10553
rect 9374 10451 9442 10533
rect 9374 10405 9385 10451
rect 9431 10405 9442 10451
rect 9374 10323 9442 10405
rect 9374 10277 9385 10323
rect 9431 10277 9442 10323
rect 9374 10252 9442 10277
rect 9813 10451 9859 10470
rect 9813 10252 9859 10311
rect 9997 10451 10063 10784
rect 10465 10830 10511 10916
rect 10465 10744 10511 10784
rect 10669 10830 10735 10870
rect 10669 10784 10689 10830
rect 10558 10693 10623 10736
rect 10558 10610 10573 10693
rect 10558 10553 10573 10558
rect 10619 10553 10623 10693
rect 10558 10536 10623 10553
rect 9997 10386 10017 10451
rect 9997 10334 9998 10386
rect 9997 10311 10017 10334
rect 9997 10298 10063 10311
rect 10485 10451 10531 10470
rect 10485 10252 10531 10311
rect 10669 10451 10735 10784
rect 11137 10830 11183 10916
rect 11137 10744 11183 10784
rect 11341 10830 11407 10870
rect 11341 10784 11361 10830
rect 11230 10693 11295 10736
rect 11230 10610 11245 10693
rect 11230 10553 11245 10558
rect 11291 10553 11295 10693
rect 11230 10536 11295 10553
rect 10669 10386 10689 10451
rect 10669 10334 10670 10386
rect 10669 10311 10689 10334
rect 10669 10298 10735 10311
rect 11157 10451 11203 10470
rect 11157 10252 11203 10311
rect 11341 10451 11407 10784
rect 11921 10830 11967 10916
rect 11921 10744 11967 10784
rect 12125 10830 12191 10870
rect 12125 10784 12145 10830
rect 12014 10693 12079 10736
rect 12014 10610 12029 10693
rect 12014 10553 12029 10558
rect 12075 10553 12079 10693
rect 12014 10536 12079 10553
rect 11341 10386 11361 10451
rect 11341 10334 11342 10386
rect 11341 10311 11361 10334
rect 11341 10298 11407 10311
rect 11941 10451 11987 10470
rect 11941 10252 11987 10311
rect 12125 10451 12191 10784
rect 12593 10830 12639 10916
rect 12593 10744 12639 10784
rect 12797 10830 12863 10870
rect 12797 10784 12817 10830
rect 12686 10693 12751 10736
rect 12686 10610 12701 10693
rect 12686 10553 12701 10558
rect 12747 10553 12751 10693
rect 12686 10536 12751 10553
rect 12797 10610 12863 10784
rect 13265 10830 13311 10916
rect 13265 10744 13311 10784
rect 13469 10830 13535 10870
rect 13469 10784 13489 10830
rect 12797 10558 12798 10610
rect 12850 10558 12863 10610
rect 12125 10386 12145 10451
rect 12125 10334 12126 10386
rect 12125 10311 12145 10334
rect 12125 10298 12191 10311
rect 12613 10451 12659 10470
rect 12613 10252 12659 10311
rect 12797 10451 12863 10558
rect 13358 10693 13423 10736
rect 13358 10610 13373 10693
rect 13358 10553 13373 10558
rect 13419 10553 13423 10693
rect 13358 10536 13423 10553
rect 13469 10610 13535 10784
rect 13937 10830 13983 10916
rect 13937 10744 13983 10784
rect 14141 10830 14207 10870
rect 14141 10784 14161 10830
rect 13469 10558 13470 10610
rect 13522 10558 13535 10610
rect 12797 10311 12817 10451
rect 12797 10298 12863 10311
rect 13285 10451 13331 10470
rect 13285 10252 13331 10311
rect 13469 10451 13535 10558
rect 14030 10693 14095 10736
rect 14030 10610 14045 10693
rect 14030 10553 14045 10558
rect 14091 10553 14095 10693
rect 14030 10536 14095 10553
rect 14141 10610 14207 10784
rect 14609 10830 14655 10916
rect 14609 10744 14655 10784
rect 14813 10830 14879 10870
rect 14813 10784 14833 10830
rect 14141 10558 14142 10610
rect 14194 10558 14207 10610
rect 13469 10311 13489 10451
rect 13469 10298 13535 10311
rect 13957 10451 14003 10470
rect 13957 10252 14003 10311
rect 14141 10451 14207 10558
rect 14702 10693 14767 10736
rect 14702 10610 14717 10693
rect 14702 10553 14717 10558
rect 14763 10553 14767 10693
rect 14702 10536 14767 10553
rect 14813 10610 14879 10784
rect 15281 10830 15327 10916
rect 15281 10744 15327 10784
rect 15485 10830 15551 10870
rect 15485 10784 15505 10830
rect 14813 10558 14814 10610
rect 14866 10558 14879 10610
rect 14141 10311 14161 10451
rect 14141 10298 14207 10311
rect 14629 10451 14675 10470
rect 14629 10252 14675 10311
rect 14813 10451 14879 10558
rect 15374 10693 15439 10736
rect 15374 10610 15389 10693
rect 15374 10553 15389 10558
rect 15435 10553 15439 10693
rect 15374 10536 15439 10553
rect 15485 10610 15551 10784
rect 15953 10830 15999 10916
rect 15953 10744 15999 10784
rect 16157 10830 16223 10870
rect 16157 10784 16177 10830
rect 15485 10558 15486 10610
rect 15538 10558 15551 10610
rect 14813 10311 14833 10451
rect 14813 10298 14879 10311
rect 15301 10451 15347 10470
rect 15301 10252 15347 10311
rect 15485 10451 15551 10558
rect 16046 10693 16111 10736
rect 16046 10610 16061 10693
rect 16046 10553 16061 10558
rect 16107 10553 16111 10693
rect 16046 10536 16111 10553
rect 15485 10311 15505 10451
rect 15485 10298 15551 10311
rect 15973 10451 16019 10470
rect 15973 10252 16019 10311
rect 16157 10451 16223 10784
rect 16625 10830 16671 10916
rect 17326 10897 17394 10916
rect 16625 10744 16671 10784
rect 16829 10830 16895 10870
rect 16829 10784 16849 10830
rect 16718 10722 16783 10736
rect 16770 10693 16783 10722
rect 16718 10553 16733 10670
rect 16779 10553 16783 10693
rect 16718 10536 16783 10553
rect 16157 10386 16177 10451
rect 16157 10334 16158 10386
rect 16157 10311 16177 10334
rect 16157 10298 16223 10311
rect 16645 10451 16691 10470
rect 16645 10252 16691 10311
rect 16829 10451 16895 10784
rect 17326 10750 17337 10897
rect 17383 10750 17394 10897
rect 17326 10739 17394 10750
rect 17633 10830 17679 10916
rect 17633 10744 17679 10784
rect 17837 10830 17903 10870
rect 17837 10784 17857 10830
rect 17726 10722 17791 10736
rect 17778 10693 17791 10722
rect 16829 10386 16849 10451
rect 16829 10334 16830 10386
rect 16829 10311 16849 10334
rect 16829 10298 16895 10311
rect 17326 10579 17394 10590
rect 17326 10533 17337 10579
rect 17383 10533 17394 10579
rect 17726 10553 17741 10670
rect 17787 10553 17791 10693
rect 17726 10536 17791 10553
rect 17326 10451 17394 10533
rect 17326 10405 17337 10451
rect 17383 10405 17394 10451
rect 17326 10323 17394 10405
rect 17326 10277 17337 10323
rect 17383 10277 17394 10323
rect 17326 10252 17394 10277
rect 17653 10451 17699 10470
rect 17653 10252 17699 10311
rect 17837 10451 17903 10784
rect 18305 10830 18351 10916
rect 18305 10744 18351 10784
rect 18509 10830 18575 10870
rect 18509 10784 18529 10830
rect 18398 10722 18463 10736
rect 18450 10693 18463 10722
rect 18398 10553 18413 10670
rect 18459 10553 18463 10693
rect 18398 10536 18463 10553
rect 17837 10386 17857 10451
rect 17837 10334 17838 10386
rect 17837 10311 17857 10334
rect 17837 10298 17903 10311
rect 18325 10451 18371 10470
rect 18325 10252 18371 10311
rect 18509 10451 18575 10784
rect 18977 10830 19023 10916
rect 18977 10744 19023 10784
rect 19181 10834 19247 10870
rect 19181 10782 19182 10834
rect 19234 10830 19247 10834
rect 19234 10782 19247 10784
rect 19070 10722 19135 10736
rect 19122 10693 19135 10722
rect 19070 10553 19085 10670
rect 19131 10553 19135 10693
rect 19070 10536 19135 10553
rect 18509 10386 18529 10451
rect 18509 10334 18510 10386
rect 18509 10311 18529 10334
rect 18509 10298 18575 10311
rect 18997 10451 19043 10470
rect 18997 10252 19043 10311
rect 19181 10451 19247 10782
rect 19649 10830 19695 10916
rect 19649 10744 19695 10784
rect 19853 10834 19919 10870
rect 19853 10782 19854 10834
rect 19906 10830 19919 10834
rect 19906 10782 19919 10784
rect 19742 10722 19807 10736
rect 19794 10693 19807 10722
rect 19742 10553 19757 10670
rect 19803 10553 19807 10693
rect 19742 10536 19807 10553
rect 19181 10311 19201 10451
rect 19181 10298 19247 10311
rect 19669 10451 19715 10470
rect 19669 10252 19715 10311
rect 19853 10451 19919 10782
rect 20321 10830 20367 10916
rect 20321 10744 20367 10784
rect 20525 10830 20591 10870
rect 20525 10784 20545 10830
rect 20414 10722 20479 10736
rect 20466 10693 20479 10722
rect 20414 10553 20429 10670
rect 20475 10553 20479 10693
rect 20414 10536 20479 10553
rect 19853 10311 19873 10451
rect 19853 10298 19919 10311
rect 20341 10451 20387 10470
rect 20341 10252 20387 10311
rect 20525 10451 20591 10784
rect 20993 10830 21039 10916
rect 20993 10744 21039 10784
rect 21197 10830 21263 10870
rect 21197 10784 21217 10830
rect 21086 10722 21151 10736
rect 21138 10693 21151 10722
rect 21086 10553 21101 10670
rect 21147 10553 21151 10693
rect 21086 10536 21151 10553
rect 20525 10386 20545 10451
rect 20525 10334 20526 10386
rect 20525 10311 20545 10334
rect 20525 10298 20591 10311
rect 21013 10451 21059 10470
rect 21013 10252 21059 10311
rect 21197 10451 21263 10784
rect 21665 10830 21711 10916
rect 22482 10897 22550 10916
rect 21665 10744 21711 10784
rect 21869 10830 21935 10870
rect 21869 10784 21889 10830
rect 21758 10722 21823 10736
rect 21810 10693 21823 10722
rect 21758 10553 21773 10670
rect 21819 10553 21823 10693
rect 21758 10536 21823 10553
rect 21869 10722 21935 10784
rect 22482 10750 22493 10897
rect 22539 10750 22550 10897
rect 22482 10738 22550 10750
rect 21869 10670 21870 10722
rect 21922 10670 21935 10722
rect 21197 10386 21217 10451
rect 21197 10334 21198 10386
rect 21197 10311 21217 10334
rect 21197 10298 21263 10311
rect 21685 10451 21731 10470
rect 21685 10252 21731 10311
rect 21869 10451 21935 10670
rect 21869 10311 21889 10451
rect 21869 10298 21935 10311
rect 22482 10579 22550 10592
rect 22482 10533 22493 10579
rect 22539 10533 22550 10579
rect 22482 10451 22550 10533
rect 22482 10405 22493 10451
rect 22539 10405 22550 10451
rect 22482 10323 22550 10405
rect 22482 10277 22493 10323
rect 22539 10277 22550 10323
rect 22482 10252 22550 10277
rect 1344 10218 22624 10252
rect 1344 10166 3874 10218
rect 4134 10166 9194 10218
rect 9454 10166 14514 10218
rect 14774 10166 19834 10218
rect 20094 10166 22624 10218
rect 1344 10132 22624 10166
rect 1418 10107 1486 10132
rect 1418 10061 1429 10107
rect 1475 10061 1486 10107
rect 1418 9979 1486 10061
rect 1418 9933 1429 9979
rect 1475 9933 1486 9979
rect 1418 9851 1486 9933
rect 1418 9805 1429 9851
rect 1475 9805 1486 9851
rect 1418 9792 1486 9805
rect 1617 10065 1663 10086
rect 1617 9719 1663 9925
rect 1921 10065 1967 10132
rect 1921 9906 1967 9925
rect 2065 10065 2111 10086
rect 1714 9800 1728 9846
rect 1868 9800 1967 9846
rect 1617 9673 1720 9719
rect 1860 9673 1872 9719
rect 1418 9634 1486 9646
rect 1418 9487 1429 9634
rect 1475 9487 1486 9634
rect 1418 9468 1486 9487
rect 1617 9600 1663 9622
rect 1617 9468 1663 9554
rect 1921 9600 1967 9800
rect 2065 9719 2111 9925
rect 2369 10065 2415 10132
rect 2369 9906 2415 9925
rect 2513 10065 2559 10086
rect 2162 9800 2176 9846
rect 2316 9800 2415 9846
rect 2065 9673 2168 9719
rect 2308 9673 2320 9719
rect 1921 9514 1967 9554
rect 2065 9600 2111 9622
rect 2065 9468 2111 9554
rect 2369 9600 2415 9800
rect 2513 9719 2559 9925
rect 2817 10065 2863 10132
rect 2817 9906 2863 9925
rect 2961 10065 3007 10086
rect 2610 9800 2624 9846
rect 2764 9800 2863 9846
rect 2513 9673 2616 9719
rect 2756 9673 2768 9719
rect 2369 9514 2415 9554
rect 2513 9600 2559 9622
rect 2513 9468 2559 9554
rect 2817 9600 2863 9800
rect 2961 9719 3007 9925
rect 3265 10065 3311 10132
rect 3265 9906 3311 9925
rect 3409 10065 3455 10086
rect 3058 9800 3072 9846
rect 3212 9800 3311 9846
rect 2961 9673 3064 9719
rect 3204 9673 3216 9719
rect 2817 9514 2863 9554
rect 2961 9600 3007 9622
rect 2961 9468 3007 9554
rect 3265 9600 3311 9800
rect 3409 9719 3455 9925
rect 3713 10065 3759 10132
rect 3713 9906 3759 9925
rect 4101 10073 4147 10132
rect 4101 9914 4147 9933
rect 4285 10073 4351 10086
rect 4285 9933 4305 10073
rect 3506 9800 3520 9846
rect 3660 9800 3759 9846
rect 3409 9673 3512 9719
rect 3652 9673 3664 9719
rect 3265 9514 3311 9554
rect 3409 9600 3455 9627
rect 3409 9468 3455 9554
rect 3713 9600 3759 9800
rect 4174 9831 4239 9848
rect 4174 9826 4189 9831
rect 4174 9691 4189 9774
rect 4235 9691 4239 9831
rect 4174 9648 4239 9691
rect 4285 9826 4351 9933
rect 4773 10073 4819 10132
rect 5342 10107 5410 10132
rect 4773 9914 4819 9933
rect 4957 10073 5023 10086
rect 4957 9933 4977 10073
rect 4285 9774 4286 9826
rect 4338 9774 4351 9826
rect 3713 9514 3759 9554
rect 4081 9600 4127 9640
rect 4081 9468 4127 9554
rect 4285 9600 4351 9774
rect 4846 9831 4911 9848
rect 4846 9826 4861 9831
rect 4846 9691 4861 9774
rect 4907 9691 4911 9831
rect 4846 9648 4911 9691
rect 4285 9554 4305 9600
rect 4285 9514 4351 9554
rect 4753 9600 4799 9640
rect 4753 9468 4799 9554
rect 4957 9602 5023 9933
rect 5342 10061 5353 10107
rect 5399 10061 5410 10107
rect 5342 9979 5410 10061
rect 5342 9933 5353 9979
rect 5399 9933 5410 9979
rect 5342 9851 5410 9933
rect 5781 10073 5827 10132
rect 5781 9914 5827 9933
rect 5965 10073 6031 10086
rect 5965 9933 5985 10073
rect 5342 9805 5353 9851
rect 5399 9805 5410 9851
rect 5342 9794 5410 9805
rect 5854 9831 5919 9848
rect 5854 9714 5869 9831
rect 5915 9691 5919 9831
rect 5906 9662 5919 9691
rect 5854 9648 5919 9662
rect 4957 9550 4958 9602
rect 5010 9600 5023 9602
rect 5010 9550 5023 9554
rect 4957 9514 5023 9550
rect 5342 9634 5410 9645
rect 5342 9487 5353 9634
rect 5399 9487 5410 9634
rect 5342 9468 5410 9487
rect 5761 9600 5807 9640
rect 5761 9468 5807 9554
rect 5965 9602 6031 9933
rect 6453 10073 6499 10132
rect 6453 9914 6499 9933
rect 6637 10073 6703 10086
rect 6637 9933 6657 10073
rect 6526 9831 6591 9848
rect 6526 9714 6541 9831
rect 6587 9691 6591 9831
rect 6578 9662 6591 9691
rect 6526 9648 6591 9662
rect 6637 9714 6703 9933
rect 7125 10073 7171 10132
rect 7125 9914 7171 9933
rect 7309 10073 7375 10086
rect 7309 9933 7329 10073
rect 6637 9662 6638 9714
rect 6690 9662 6703 9714
rect 5965 9550 5966 9602
rect 6018 9600 6031 9602
rect 6018 9550 6031 9554
rect 5965 9514 6031 9550
rect 6433 9600 6479 9640
rect 6433 9468 6479 9554
rect 6637 9600 6703 9662
rect 7198 9831 7263 9848
rect 7198 9714 7213 9831
rect 7259 9691 7263 9831
rect 7250 9662 7263 9691
rect 7198 9648 7263 9662
rect 7309 9714 7375 9933
rect 7797 10073 7843 10132
rect 7797 9914 7843 9933
rect 7981 10073 8047 10086
rect 7981 9933 8001 10073
rect 7309 9662 7310 9714
rect 7362 9662 7375 9714
rect 6637 9554 6657 9600
rect 6637 9514 6703 9554
rect 7105 9600 7151 9640
rect 7105 9468 7151 9554
rect 7309 9600 7375 9662
rect 7870 9831 7935 9848
rect 7870 9826 7885 9831
rect 7870 9691 7885 9774
rect 7931 9691 7935 9831
rect 7870 9648 7935 9691
rect 7309 9554 7329 9600
rect 7309 9514 7375 9554
rect 7777 9600 7823 9640
rect 7777 9468 7823 9554
rect 7981 9602 8047 9933
rect 8469 10073 8515 10132
rect 8469 9914 8515 9933
rect 8653 10073 8719 10086
rect 8653 9933 8673 10073
rect 8542 9831 8607 9848
rect 8542 9826 8557 9831
rect 8542 9691 8557 9774
rect 8603 9691 8607 9831
rect 8542 9648 8607 9691
rect 7981 9550 7982 9602
rect 8034 9600 8047 9602
rect 8034 9550 8047 9554
rect 7981 9514 8047 9550
rect 8449 9600 8495 9640
rect 8449 9468 8495 9554
rect 8653 9602 8719 9933
rect 9141 10073 9187 10132
rect 9141 9914 9187 9933
rect 9325 10073 9391 10086
rect 9325 9933 9345 10073
rect 9214 9831 9279 9848
rect 9214 9826 9229 9831
rect 9214 9691 9229 9774
rect 9275 9691 9279 9831
rect 9214 9648 9279 9691
rect 8653 9550 8654 9602
rect 8706 9600 8719 9602
rect 8706 9550 8719 9554
rect 8653 9514 8719 9550
rect 9121 9600 9167 9640
rect 9121 9468 9167 9554
rect 9325 9602 9391 9933
rect 9813 10073 9859 10132
rect 9813 9914 9859 9933
rect 9997 10073 10063 10086
rect 9997 9933 10017 10073
rect 9886 9831 9951 9848
rect 9886 9714 9901 9831
rect 9947 9691 9951 9831
rect 9938 9662 9951 9691
rect 9886 9648 9951 9662
rect 9325 9550 9326 9602
rect 9378 9600 9391 9602
rect 9378 9550 9391 9554
rect 9325 9514 9391 9550
rect 9793 9600 9839 9640
rect 9793 9468 9839 9554
rect 9997 9602 10063 9933
rect 10485 10073 10531 10132
rect 10485 9914 10531 9933
rect 10669 10073 10735 10086
rect 10669 9933 10689 10073
rect 10558 9831 10623 9848
rect 10558 9826 10573 9831
rect 10558 9691 10573 9774
rect 10619 9691 10623 9831
rect 10558 9648 10623 9691
rect 9997 9550 9998 9602
rect 10050 9600 10063 9602
rect 10050 9550 10063 9554
rect 9997 9514 10063 9550
rect 10465 9600 10511 9640
rect 10465 9468 10511 9554
rect 10669 9602 10735 9933
rect 10913 10065 10959 10086
rect 10913 9719 10959 9925
rect 11217 10065 11263 10132
rect 11217 9906 11263 9925
rect 11381 10073 11427 10132
rect 11381 9914 11427 9933
rect 11565 10073 11631 10086
rect 11565 10050 11585 10073
rect 11565 9998 11566 10050
rect 11565 9933 11585 9998
rect 11010 9800 11024 9846
rect 11164 9800 11263 9846
rect 10913 9673 11016 9719
rect 11156 9673 11168 9719
rect 10669 9550 10670 9602
rect 10722 9600 10735 9602
rect 10722 9550 10735 9554
rect 10669 9514 10735 9550
rect 10913 9600 10959 9627
rect 10913 9468 10959 9554
rect 11217 9600 11263 9800
rect 11454 9831 11519 9848
rect 11454 9714 11469 9831
rect 11515 9691 11519 9831
rect 11506 9662 11519 9691
rect 11454 9648 11519 9662
rect 11217 9514 11263 9554
rect 11361 9600 11407 9640
rect 11361 9468 11407 9554
rect 11565 9600 11631 9933
rect 12053 10073 12099 10132
rect 12053 9914 12099 9933
rect 12237 10073 12303 10086
rect 12237 9933 12257 10073
rect 12126 9831 12191 9848
rect 12126 9826 12141 9831
rect 12126 9691 12141 9774
rect 12187 9691 12191 9831
rect 12126 9648 12191 9691
rect 12237 9826 12303 9933
rect 12725 10073 12771 10132
rect 13294 10107 13362 10132
rect 12725 9914 12771 9933
rect 12909 10073 12975 10086
rect 12909 9933 12929 10073
rect 12237 9774 12238 9826
rect 12290 9774 12303 9826
rect 11565 9554 11585 9600
rect 11565 9514 11631 9554
rect 12033 9600 12079 9640
rect 12033 9468 12079 9554
rect 12237 9600 12303 9774
rect 12798 9831 12863 9848
rect 12798 9714 12813 9831
rect 12859 9691 12863 9831
rect 12850 9662 12863 9691
rect 12798 9648 12863 9662
rect 12909 9714 12975 9933
rect 13294 10061 13305 10107
rect 13351 10061 13362 10107
rect 13294 9979 13362 10061
rect 13294 9933 13305 9979
rect 13351 9933 13362 9979
rect 13294 9851 13362 9933
rect 13621 10073 13667 10132
rect 13621 9914 13667 9933
rect 13805 10073 13871 10086
rect 13805 9933 13825 10073
rect 13294 9805 13305 9851
rect 13351 9805 13362 9851
rect 13294 9794 13362 9805
rect 13694 9831 13759 9848
rect 12909 9662 12910 9714
rect 12962 9662 12975 9714
rect 12237 9554 12257 9600
rect 12237 9514 12303 9554
rect 12705 9600 12751 9640
rect 12705 9468 12751 9554
rect 12909 9600 12975 9662
rect 13694 9714 13709 9831
rect 13755 9691 13759 9831
rect 13746 9662 13759 9691
rect 13694 9648 13759 9662
rect 13805 9714 13871 9933
rect 14293 10073 14339 10132
rect 14293 9914 14339 9933
rect 14477 10073 14543 10086
rect 14477 9933 14497 10073
rect 13805 9662 13806 9714
rect 13858 9662 13871 9714
rect 12909 9554 12929 9600
rect 12909 9514 12975 9554
rect 13294 9634 13362 9645
rect 13294 9487 13305 9634
rect 13351 9487 13362 9634
rect 13294 9468 13362 9487
rect 13601 9600 13647 9640
rect 13601 9468 13647 9554
rect 13805 9600 13871 9662
rect 14366 9831 14431 9848
rect 14366 9714 14381 9831
rect 14427 9691 14431 9831
rect 14418 9662 14431 9691
rect 14366 9648 14431 9662
rect 14477 9826 14543 9933
rect 14965 10073 15011 10132
rect 14965 9914 15011 9933
rect 15149 10073 15215 10086
rect 15149 9933 15169 10073
rect 14477 9774 14478 9826
rect 14530 9774 14543 9826
rect 13805 9554 13825 9600
rect 13805 9514 13871 9554
rect 14273 9600 14319 9640
rect 14273 9468 14319 9554
rect 14477 9600 14543 9774
rect 15038 9831 15103 9848
rect 15038 9826 15053 9831
rect 15038 9691 15053 9774
rect 15099 9691 15103 9831
rect 15038 9648 15103 9691
rect 14477 9554 14497 9600
rect 14477 9514 14543 9554
rect 14945 9600 14991 9640
rect 14945 9468 14991 9554
rect 15149 9602 15215 9933
rect 15637 10073 15683 10132
rect 15637 9914 15683 9933
rect 15821 10073 15887 10086
rect 15821 9933 15841 10073
rect 15710 9831 15775 9848
rect 15710 9826 15725 9831
rect 15710 9691 15725 9774
rect 15771 9691 15775 9831
rect 15710 9648 15775 9691
rect 15149 9550 15150 9602
rect 15202 9600 15215 9602
rect 15202 9550 15215 9554
rect 15149 9514 15215 9550
rect 15617 9600 15663 9640
rect 15617 9468 15663 9554
rect 15821 9602 15887 9933
rect 16309 10073 16355 10132
rect 16309 9914 16355 9933
rect 16493 10073 16559 10086
rect 16493 9933 16513 10073
rect 16382 9831 16447 9848
rect 16382 9714 16397 9831
rect 16443 9691 16447 9831
rect 16434 9662 16447 9691
rect 16382 9648 16447 9662
rect 15821 9550 15822 9602
rect 15874 9600 15887 9602
rect 15874 9550 15887 9554
rect 15821 9514 15887 9550
rect 16289 9600 16335 9640
rect 16289 9468 16335 9554
rect 16493 9602 16559 9933
rect 16981 10073 17027 10132
rect 16981 9914 17027 9933
rect 17165 10073 17231 10086
rect 17165 9933 17185 10073
rect 17054 9831 17119 9848
rect 17054 9714 17069 9831
rect 17115 9691 17119 9831
rect 17106 9662 17119 9691
rect 17054 9648 17119 9662
rect 16493 9550 16494 9602
rect 16546 9600 16559 9602
rect 16546 9550 16559 9554
rect 16493 9514 16559 9550
rect 16961 9600 17007 9640
rect 16961 9468 17007 9554
rect 17165 9602 17231 9933
rect 17165 9550 17166 9602
rect 17218 9600 17231 9602
rect 17218 9550 17231 9554
rect 17165 9514 17231 9550
rect 17713 10073 17779 10086
rect 17759 9933 17779 10073
rect 17713 9602 17779 9933
rect 17917 10073 17963 10132
rect 17917 9914 17963 9933
rect 18325 10073 18371 10132
rect 18325 9914 18371 9933
rect 18509 10073 18575 10086
rect 18509 10050 18529 10073
rect 18509 9998 18510 10050
rect 18509 9933 18529 9998
rect 17825 9831 17890 9848
rect 17825 9691 17829 9831
rect 17875 9826 17890 9831
rect 17875 9691 17890 9774
rect 17825 9648 17890 9691
rect 18398 9831 18463 9848
rect 18398 9714 18413 9831
rect 18459 9691 18463 9831
rect 18450 9662 18463 9691
rect 18398 9648 18463 9662
rect 17713 9600 17726 9602
rect 17713 9550 17726 9554
rect 17778 9550 17779 9602
rect 17713 9514 17779 9550
rect 17937 9600 17983 9640
rect 17937 9468 17983 9554
rect 18305 9600 18351 9640
rect 18305 9468 18351 9554
rect 18509 9600 18575 9933
rect 18997 10073 19043 10132
rect 18997 9914 19043 9933
rect 19181 10073 19247 10086
rect 19181 9933 19201 10073
rect 19070 9831 19135 9848
rect 19070 9826 19085 9831
rect 19070 9691 19085 9774
rect 19131 9691 19135 9831
rect 19070 9648 19135 9691
rect 18509 9554 18529 9600
rect 18509 9514 18575 9554
rect 18977 9600 19023 9640
rect 18977 9468 19023 9554
rect 19181 9602 19247 9933
rect 19669 10073 19715 10132
rect 19669 9914 19715 9933
rect 19853 10073 19919 10086
rect 19853 9933 19873 10073
rect 19742 9831 19807 9848
rect 19742 9826 19757 9831
rect 19742 9691 19757 9774
rect 19803 9691 19807 9831
rect 19742 9648 19807 9691
rect 19181 9550 19182 9602
rect 19234 9600 19247 9602
rect 19234 9550 19247 9554
rect 19181 9514 19247 9550
rect 19649 9600 19695 9640
rect 19649 9468 19695 9554
rect 19853 9602 19919 9933
rect 20341 10073 20387 10132
rect 20341 9914 20387 9933
rect 20525 10073 20591 10086
rect 20525 10050 20545 10073
rect 20525 9998 20526 10050
rect 20525 9933 20545 9998
rect 20414 9831 20479 9848
rect 20414 9826 20429 9831
rect 20414 9691 20429 9774
rect 20475 9691 20479 9831
rect 20414 9648 20479 9691
rect 19853 9550 19854 9602
rect 19906 9600 19919 9602
rect 19906 9550 19919 9554
rect 19853 9514 19919 9550
rect 20321 9600 20367 9640
rect 20321 9468 20367 9554
rect 20525 9600 20591 9933
rect 20769 10065 20815 10086
rect 20769 9719 20815 9925
rect 21073 10065 21119 10132
rect 21073 9906 21119 9925
rect 21246 10107 21314 10132
rect 21246 10061 21257 10107
rect 21303 10061 21314 10107
rect 21246 9979 21314 10061
rect 21246 9933 21257 9979
rect 21303 9933 21314 9979
rect 21246 9851 21314 9933
rect 21573 10073 21619 10132
rect 21573 9914 21619 9933
rect 21757 10073 21823 10086
rect 21757 10050 21777 10073
rect 21757 9998 21758 10050
rect 21757 9933 21777 9998
rect 20866 9800 20880 9846
rect 21020 9800 21119 9846
rect 20769 9673 20872 9719
rect 21012 9673 21024 9719
rect 20525 9554 20545 9600
rect 20525 9514 20591 9554
rect 20769 9600 20815 9627
rect 20769 9468 20815 9554
rect 21073 9600 21119 9800
rect 21246 9805 21257 9851
rect 21303 9805 21314 9851
rect 21246 9794 21314 9805
rect 21646 9831 21711 9848
rect 21646 9826 21661 9831
rect 21646 9691 21661 9774
rect 21707 9691 21711 9831
rect 21646 9648 21711 9691
rect 21073 9514 21119 9554
rect 21246 9634 21314 9645
rect 21246 9487 21257 9634
rect 21303 9487 21314 9634
rect 21246 9468 21314 9487
rect 21553 9600 21599 9640
rect 21553 9468 21599 9554
rect 21757 9600 21823 9933
rect 22001 10065 22047 10086
rect 22001 9719 22047 9925
rect 22305 10065 22351 10132
rect 22305 9906 22351 9925
rect 22482 10107 22550 10132
rect 22482 10061 22493 10107
rect 22539 10061 22550 10107
rect 22482 9979 22550 10061
rect 22482 9933 22493 9979
rect 22539 9933 22550 9979
rect 22482 9851 22550 9933
rect 22098 9800 22112 9846
rect 22252 9800 22351 9846
rect 22001 9673 22104 9719
rect 22244 9673 22256 9719
rect 21757 9554 21777 9600
rect 21757 9514 21823 9554
rect 22001 9600 22047 9627
rect 22001 9468 22047 9554
rect 22305 9600 22351 9800
rect 22482 9805 22493 9851
rect 22539 9805 22550 9851
rect 22482 9792 22550 9805
rect 22305 9514 22351 9554
rect 22482 9634 22550 9646
rect 22482 9487 22493 9634
rect 22539 9487 22550 9634
rect 22482 9468 22550 9487
rect 1344 9434 22784 9468
rect 1344 9382 6534 9434
rect 6794 9382 11854 9434
rect 12114 9382 17174 9434
rect 17434 9382 22494 9434
rect 22754 9382 22784 9434
rect 1344 9348 22784 9382
rect 1418 9329 1486 9348
rect 1418 9182 1429 9329
rect 1475 9182 1486 9329
rect 1617 9262 1663 9348
rect 1617 9191 1663 9216
rect 1921 9262 1967 9302
rect 1418 9170 1486 9182
rect 1617 9097 1720 9143
rect 1860 9097 1872 9143
rect 1418 9011 1486 9024
rect 1418 8965 1429 9011
rect 1475 8965 1486 9011
rect 1418 8883 1486 8965
rect 1418 8837 1429 8883
rect 1475 8837 1486 8883
rect 1418 8755 1486 8837
rect 1418 8709 1429 8755
rect 1475 8709 1486 8755
rect 1617 8891 1663 9097
rect 1921 9016 1967 9216
rect 2065 9262 2111 9348
rect 2065 9191 2111 9216
rect 2369 9262 2415 9302
rect 1714 8970 1728 9016
rect 1868 8970 1967 9016
rect 2065 9097 2168 9143
rect 2308 9097 2320 9143
rect 1617 8730 1663 8751
rect 1921 8891 1967 8910
rect 1418 8684 1486 8709
rect 1921 8684 1967 8751
rect 2065 8891 2111 9097
rect 2369 9016 2415 9216
rect 2513 9262 2559 9348
rect 2513 9189 2559 9216
rect 2817 9262 2863 9302
rect 2162 8970 2176 9016
rect 2316 8970 2415 9016
rect 2513 9097 2616 9143
rect 2756 9097 2768 9143
rect 2065 8730 2111 8751
rect 2369 8891 2415 8910
rect 2369 8684 2415 8751
rect 2513 8891 2559 9097
rect 2817 9016 2863 9216
rect 3297 9262 3343 9348
rect 3297 9176 3343 9216
rect 3501 9262 3567 9302
rect 3501 9216 3521 9262
rect 2610 8970 2624 9016
rect 2764 8970 2863 9016
rect 3390 9154 3455 9168
rect 3442 9125 3455 9154
rect 3390 8985 3405 9102
rect 3451 8985 3455 9125
rect 3390 8968 3455 8985
rect 3501 9154 3567 9216
rect 3969 9262 4015 9348
rect 3969 9176 4015 9216
rect 4173 9262 4239 9302
rect 4173 9216 4193 9262
rect 3501 9102 3502 9154
rect 3554 9102 3567 9154
rect 2513 8730 2559 8751
rect 2817 8891 2863 8910
rect 2817 8684 2863 8751
rect 3317 8883 3363 8902
rect 3317 8684 3363 8743
rect 3501 8883 3567 9102
rect 4062 9154 4127 9168
rect 4114 9125 4127 9154
rect 4062 8985 4077 9102
rect 4123 8985 4127 9125
rect 4062 8968 4127 8985
rect 3501 8743 3521 8883
rect 3501 8730 3567 8743
rect 3989 8883 4035 8902
rect 3989 8684 4035 8743
rect 4173 8883 4239 9216
rect 4641 9262 4687 9348
rect 4641 9176 4687 9216
rect 4845 9266 4911 9302
rect 4845 9214 4846 9266
rect 4898 9262 4911 9266
rect 4898 9214 4911 9216
rect 4734 9125 4799 9168
rect 4734 9042 4749 9125
rect 4734 8985 4749 8990
rect 4795 8985 4799 9125
rect 4734 8968 4799 8985
rect 4173 8818 4193 8883
rect 4173 8766 4174 8818
rect 4173 8743 4193 8766
rect 4173 8730 4239 8743
rect 4661 8883 4707 8902
rect 4661 8684 4707 8743
rect 4845 8883 4911 9214
rect 5313 9262 5359 9348
rect 5313 9176 5359 9216
rect 5517 9262 5583 9302
rect 5517 9216 5537 9262
rect 5406 9125 5471 9168
rect 5406 9042 5421 9125
rect 5406 8985 5421 8990
rect 5467 8985 5471 9125
rect 5406 8968 5471 8985
rect 4845 8743 4865 8883
rect 4845 8730 4911 8743
rect 5333 8883 5379 8902
rect 5333 8684 5379 8743
rect 5517 8883 5583 9216
rect 5985 9262 6031 9348
rect 5985 9176 6031 9216
rect 6189 9262 6255 9302
rect 6189 9216 6209 9262
rect 6078 9125 6143 9168
rect 6078 9042 6093 9125
rect 6078 8985 6093 8990
rect 6139 8985 6143 9125
rect 6078 8968 6143 8985
rect 6189 9042 6255 9216
rect 6657 9262 6703 9348
rect 6657 9176 6703 9216
rect 6861 9262 6927 9302
rect 6861 9216 6881 9262
rect 6189 8990 6190 9042
rect 6242 8990 6255 9042
rect 5517 8818 5537 8883
rect 5517 8766 5518 8818
rect 5517 8743 5537 8766
rect 5517 8730 5583 8743
rect 6005 8883 6051 8902
rect 6005 8684 6051 8743
rect 6189 8883 6255 8990
rect 6750 9125 6815 9168
rect 6750 9042 6765 9125
rect 6750 8985 6765 8990
rect 6811 8985 6815 9125
rect 6750 8968 6815 8985
rect 6861 9042 6927 9216
rect 7329 9262 7375 9348
rect 7329 9176 7375 9216
rect 7533 9262 7599 9302
rect 7533 9216 7553 9262
rect 6861 8990 6862 9042
rect 6914 8990 6927 9042
rect 6189 8743 6209 8883
rect 6189 8730 6255 8743
rect 6677 8883 6723 8902
rect 6677 8684 6723 8743
rect 6861 8883 6927 8990
rect 7422 9154 7487 9168
rect 7474 9125 7487 9154
rect 7422 8985 7437 9102
rect 7483 8985 7487 9125
rect 7422 8968 7487 8985
rect 7533 9154 7599 9216
rect 8113 9262 8159 9348
rect 8113 9176 8159 9216
rect 8317 9262 8383 9302
rect 8317 9216 8337 9262
rect 7533 9102 7534 9154
rect 7586 9102 7599 9154
rect 6861 8743 6881 8883
rect 6861 8730 6927 8743
rect 7349 8883 7395 8902
rect 7349 8684 7395 8743
rect 7533 8883 7599 9102
rect 8206 9154 8271 9168
rect 8258 9125 8271 9154
rect 8206 8985 8221 9102
rect 8267 8985 8271 9125
rect 8206 8968 8271 8985
rect 7533 8743 7553 8883
rect 7533 8730 7599 8743
rect 8133 8883 8179 8902
rect 8133 8684 8179 8743
rect 8317 8883 8383 9216
rect 8785 9262 8831 9348
rect 9374 9329 9442 9348
rect 8785 9176 8831 9216
rect 8989 9266 9055 9302
rect 8989 9214 8990 9266
rect 9042 9262 9055 9266
rect 9042 9214 9055 9216
rect 8878 9125 8943 9168
rect 8878 9042 8893 9125
rect 8878 8985 8893 8990
rect 8939 8985 8943 9125
rect 8878 8968 8943 8985
rect 8317 8818 8337 8883
rect 8317 8766 8318 8818
rect 8317 8743 8337 8766
rect 8317 8730 8383 8743
rect 8805 8883 8851 8902
rect 8805 8684 8851 8743
rect 8989 8883 9055 9214
rect 9374 9182 9385 9329
rect 9431 9182 9442 9329
rect 9569 9262 9615 9348
rect 9569 9189 9615 9216
rect 9873 9262 9919 9302
rect 9374 9171 9442 9182
rect 9569 9097 9672 9143
rect 9812 9097 9824 9143
rect 8989 8743 9009 8883
rect 8989 8730 9055 8743
rect 9374 9011 9442 9022
rect 9374 8965 9385 9011
rect 9431 8965 9442 9011
rect 9374 8883 9442 8965
rect 9374 8837 9385 8883
rect 9431 8837 9442 8883
rect 9374 8755 9442 8837
rect 9374 8709 9385 8755
rect 9431 8709 9442 8755
rect 9569 8891 9615 9097
rect 9873 9016 9919 9216
rect 10241 9262 10287 9348
rect 10241 9176 10287 9216
rect 10445 9262 10511 9302
rect 10445 9216 10465 9262
rect 9666 8970 9680 9016
rect 9820 8970 9919 9016
rect 10334 9154 10399 9168
rect 10386 9125 10399 9154
rect 10334 8985 10349 9102
rect 10395 8985 10399 9125
rect 10334 8968 10399 8985
rect 10445 8930 10511 9216
rect 10913 9262 10959 9348
rect 10913 9176 10959 9216
rect 11117 9262 11183 9302
rect 11117 9216 11137 9262
rect 11006 9125 11071 9168
rect 11006 9042 11021 9125
rect 11006 8985 11021 8990
rect 11067 8985 11071 9125
rect 11006 8968 11071 8985
rect 9569 8730 9615 8751
rect 9873 8891 9919 8910
rect 9374 8684 9442 8709
rect 9873 8684 9919 8751
rect 10261 8883 10307 8902
rect 10261 8684 10307 8743
rect 10445 8878 10446 8930
rect 10498 8883 10511 8930
rect 10445 8743 10465 8878
rect 10445 8730 10511 8743
rect 10933 8883 10979 8902
rect 10933 8684 10979 8743
rect 11117 8883 11183 9216
rect 11585 9262 11631 9348
rect 11585 9176 11631 9216
rect 11789 9262 11855 9302
rect 11789 9216 11809 9262
rect 11678 9125 11743 9168
rect 11678 9042 11693 9125
rect 11678 8985 11693 8990
rect 11739 8985 11743 9125
rect 11678 8968 11743 8985
rect 11117 8818 11137 8883
rect 11117 8766 11118 8818
rect 11117 8743 11137 8766
rect 11117 8730 11183 8743
rect 11605 8883 11651 8902
rect 11605 8684 11651 8743
rect 11789 8883 11855 9216
rect 12257 9262 12303 9348
rect 12257 9176 12303 9216
rect 12461 9262 12527 9302
rect 12461 9216 12481 9262
rect 12350 9154 12415 9168
rect 12402 9125 12415 9154
rect 12350 8985 12365 9102
rect 12411 8985 12415 9125
rect 12350 8968 12415 8985
rect 11789 8818 11809 8883
rect 11789 8766 11790 8818
rect 11789 8743 11809 8766
rect 11789 8730 11855 8743
rect 12277 8883 12323 8902
rect 12277 8684 12323 8743
rect 12461 8883 12527 9216
rect 12929 9262 12975 9348
rect 12929 9176 12975 9216
rect 13133 9262 13199 9302
rect 13133 9216 13153 9262
rect 13022 9154 13087 9168
rect 13074 9125 13087 9154
rect 13022 8985 13037 9102
rect 13083 8985 13087 9125
rect 13022 8968 13087 8985
rect 12461 8818 12481 8883
rect 12461 8766 12462 8818
rect 12461 8743 12481 8766
rect 12461 8730 12527 8743
rect 12949 8883 12995 8902
rect 12949 8684 12995 8743
rect 13133 8883 13199 9216
rect 13601 9262 13647 9348
rect 13601 9176 13647 9216
rect 13805 9262 13871 9302
rect 13805 9216 13825 9262
rect 13694 9125 13759 9168
rect 13694 9042 13709 9125
rect 13694 8985 13709 8990
rect 13755 8985 13759 9125
rect 13694 8968 13759 8985
rect 13133 8818 13153 8883
rect 13133 8766 13134 8818
rect 13133 8743 13153 8766
rect 13133 8730 13199 8743
rect 13621 8883 13667 8902
rect 13621 8684 13667 8743
rect 13805 8883 13871 9216
rect 14273 9262 14319 9348
rect 14273 9176 14319 9216
rect 14477 9266 14543 9302
rect 14477 9214 14478 9266
rect 14530 9262 14543 9266
rect 14530 9214 14543 9216
rect 14366 9125 14431 9168
rect 14366 9042 14381 9125
rect 14366 8985 14381 8990
rect 14427 8985 14431 9125
rect 14366 8968 14431 8985
rect 13805 8818 13825 8883
rect 13805 8766 13806 8818
rect 13805 8743 13825 8766
rect 13805 8730 13871 8743
rect 14293 8883 14339 8902
rect 14293 8684 14339 8743
rect 14477 8883 14543 9214
rect 14945 9262 14991 9348
rect 14945 9176 14991 9216
rect 15149 9266 15215 9302
rect 15149 9214 15150 9266
rect 15202 9262 15215 9266
rect 15202 9214 15215 9216
rect 15038 9125 15103 9168
rect 15038 9042 15053 9125
rect 15038 8985 15053 8990
rect 15099 8985 15103 9125
rect 15038 8968 15103 8985
rect 14477 8743 14497 8883
rect 14477 8730 14543 8743
rect 14965 8883 15011 8902
rect 14965 8684 15011 8743
rect 15149 8883 15215 9214
rect 15617 9262 15663 9348
rect 15617 9176 15663 9216
rect 15821 9262 15887 9302
rect 15821 9216 15841 9262
rect 15710 9154 15775 9168
rect 15762 9125 15775 9154
rect 15710 8985 15725 9102
rect 15771 8985 15775 9125
rect 15710 8968 15775 8985
rect 15149 8743 15169 8883
rect 15149 8730 15215 8743
rect 15637 8883 15683 8902
rect 15637 8684 15683 8743
rect 15821 8883 15887 9216
rect 16289 9262 16335 9348
rect 16289 9176 16335 9216
rect 16493 9262 16559 9302
rect 16493 9216 16513 9262
rect 16382 9125 16447 9168
rect 16382 9042 16397 9125
rect 16382 8985 16397 8990
rect 16443 8985 16447 9125
rect 16382 8968 16447 8985
rect 15821 8818 15841 8883
rect 15821 8766 15822 8818
rect 15821 8743 15841 8766
rect 15821 8730 15887 8743
rect 16309 8883 16355 8902
rect 16309 8684 16355 8743
rect 16493 8883 16559 9216
rect 16737 9262 16783 9348
rect 17326 9329 17394 9348
rect 16737 9189 16783 9216
rect 17041 9262 17087 9302
rect 16493 8818 16513 8883
rect 16493 8766 16494 8818
rect 16493 8743 16513 8766
rect 16493 8730 16559 8743
rect 16737 9097 16840 9143
rect 16980 9097 16992 9143
rect 16737 8891 16783 9097
rect 17041 9016 17087 9216
rect 17326 9182 17337 9329
rect 17383 9182 17394 9329
rect 17326 9171 17394 9182
rect 17633 9262 17679 9348
rect 17633 9176 17679 9216
rect 17837 9262 17903 9302
rect 17837 9216 17857 9262
rect 17726 9154 17791 9168
rect 17778 9125 17791 9154
rect 16834 8970 16848 9016
rect 16988 8970 17087 9016
rect 17326 9011 17394 9022
rect 17326 8965 17337 9011
rect 17383 8965 17394 9011
rect 17726 8985 17741 9102
rect 17787 8985 17791 9125
rect 17726 8968 17791 8985
rect 16737 8730 16783 8751
rect 17041 8891 17087 8910
rect 17041 8684 17087 8751
rect 17326 8883 17394 8965
rect 17326 8837 17337 8883
rect 17383 8837 17394 8883
rect 17326 8755 17394 8837
rect 17326 8709 17337 8755
rect 17383 8709 17394 8755
rect 17326 8684 17394 8709
rect 17653 8883 17699 8902
rect 17653 8684 17699 8743
rect 17837 8883 17903 9216
rect 18305 9262 18351 9348
rect 18305 9176 18351 9216
rect 18509 9262 18575 9302
rect 18509 9216 18529 9262
rect 18398 9125 18463 9168
rect 18398 9042 18413 9125
rect 18398 8985 18413 8990
rect 18459 8985 18463 9125
rect 18398 8968 18463 8985
rect 17837 8818 17857 8883
rect 17837 8766 17838 8818
rect 17837 8743 17857 8766
rect 17837 8730 17903 8743
rect 18325 8883 18371 8902
rect 18325 8684 18371 8743
rect 18509 8883 18575 9216
rect 18977 9262 19023 9348
rect 18977 9176 19023 9216
rect 19181 9262 19247 9302
rect 19181 9216 19201 9262
rect 19070 9154 19135 9168
rect 19122 9125 19135 9154
rect 19070 8985 19085 9102
rect 19131 8985 19135 9125
rect 19070 8968 19135 8985
rect 18509 8818 18529 8883
rect 18509 8766 18510 8818
rect 18509 8743 18529 8766
rect 18509 8730 18575 8743
rect 18997 8883 19043 8902
rect 18997 8684 19043 8743
rect 19181 8883 19247 9216
rect 19649 9262 19695 9348
rect 19649 9176 19695 9216
rect 19853 9266 19919 9302
rect 19853 9214 19854 9266
rect 19906 9262 19919 9266
rect 19906 9214 19919 9216
rect 19742 9125 19807 9168
rect 19742 9042 19757 9125
rect 19742 8985 19757 8990
rect 19803 8985 19807 9125
rect 19742 8968 19807 8985
rect 19181 8818 19201 8883
rect 19181 8766 19182 8818
rect 19181 8743 19201 8766
rect 19181 8730 19247 8743
rect 19669 8883 19715 8902
rect 19669 8684 19715 8743
rect 19853 8883 19919 9214
rect 20321 9262 20367 9348
rect 20321 9176 20367 9216
rect 20525 9266 20591 9302
rect 20525 9214 20526 9266
rect 20578 9262 20591 9266
rect 20578 9214 20591 9216
rect 20414 9154 20479 9168
rect 20466 9125 20479 9154
rect 20414 8985 20429 9102
rect 20475 8985 20479 9125
rect 20414 8968 20479 8985
rect 19853 8743 19873 8883
rect 19853 8730 19919 8743
rect 20341 8883 20387 8902
rect 20341 8684 20387 8743
rect 20525 8883 20591 9214
rect 20769 9262 20815 9348
rect 20769 9191 20815 9216
rect 21073 9262 21119 9302
rect 20525 8743 20545 8883
rect 20525 8730 20591 8743
rect 20769 9097 20872 9143
rect 21012 9097 21024 9143
rect 20769 8891 20815 9097
rect 21073 9016 21119 9216
rect 21217 9262 21263 9348
rect 21217 9191 21263 9216
rect 21521 9262 21567 9302
rect 20866 8970 20880 9016
rect 21020 8970 21119 9016
rect 21217 9097 21320 9143
rect 21460 9097 21472 9143
rect 20769 8730 20815 8751
rect 21073 8891 21119 8910
rect 21073 8684 21119 8751
rect 21217 8891 21263 9097
rect 21521 9016 21567 9216
rect 21665 9262 21711 9348
rect 22482 9329 22550 9348
rect 21665 9189 21711 9216
rect 21969 9262 22015 9302
rect 21314 8970 21328 9016
rect 21468 8970 21567 9016
rect 21665 9097 21768 9143
rect 21908 9097 21920 9143
rect 21217 8730 21263 8751
rect 21521 8891 21567 8910
rect 21521 8684 21567 8751
rect 21665 8891 21711 9097
rect 21969 9016 22015 9216
rect 22482 9182 22493 9329
rect 22539 9182 22550 9329
rect 22482 9170 22550 9182
rect 21762 8970 21776 9016
rect 21916 8970 22015 9016
rect 22482 9011 22550 9024
rect 22482 8965 22493 9011
rect 22539 8965 22550 9011
rect 21665 8730 21711 8751
rect 21969 8891 22015 8910
rect 21969 8684 22015 8751
rect 22482 8883 22550 8965
rect 22482 8837 22493 8883
rect 22539 8837 22550 8883
rect 22482 8755 22550 8837
rect 22482 8709 22493 8755
rect 22539 8709 22550 8755
rect 22482 8684 22550 8709
rect 1344 8650 22624 8684
rect 1344 8598 3874 8650
rect 4134 8598 9194 8650
rect 9454 8598 14514 8650
rect 14774 8598 19834 8650
rect 20094 8598 22624 8650
rect 1344 8564 22624 8598
rect 1418 8539 1486 8564
rect 1418 8493 1429 8539
rect 1475 8493 1486 8539
rect 1418 8411 1486 8493
rect 1418 8365 1429 8411
rect 1475 8365 1486 8411
rect 1418 8283 1486 8365
rect 1418 8237 1429 8283
rect 1475 8237 1486 8283
rect 1418 8224 1486 8237
rect 1617 8497 1663 8518
rect 1617 8151 1663 8357
rect 1921 8497 1967 8564
rect 1921 8338 1967 8357
rect 2065 8497 2111 8518
rect 1714 8232 1728 8278
rect 1868 8232 1967 8278
rect 1617 8105 1720 8151
rect 1860 8105 1872 8151
rect 1418 8066 1486 8078
rect 1418 7919 1429 8066
rect 1475 7919 1486 8066
rect 1418 7900 1486 7919
rect 1617 8032 1663 8057
rect 1617 7900 1663 7986
rect 1921 8032 1967 8232
rect 2065 8151 2111 8357
rect 2369 8497 2415 8564
rect 2369 8338 2415 8357
rect 2817 8505 2883 8518
rect 2863 8365 2883 8505
rect 2162 8232 2176 8278
rect 2316 8232 2415 8278
rect 2065 8105 2168 8151
rect 2308 8105 2320 8151
rect 1921 7946 1967 7986
rect 2065 8032 2111 8057
rect 2065 7900 2111 7986
rect 2369 8032 2415 8232
rect 2369 7946 2415 7986
rect 2817 8034 2883 8365
rect 3021 8505 3067 8564
rect 3021 8346 3067 8365
rect 3429 8505 3475 8564
rect 3429 8346 3475 8365
rect 3613 8505 3679 8518
rect 3613 8365 3633 8505
rect 2929 8263 2994 8280
rect 2929 8123 2933 8263
rect 2979 8146 2994 8263
rect 2929 8094 2942 8123
rect 2929 8080 2994 8094
rect 3502 8263 3567 8280
rect 3502 8146 3517 8263
rect 3563 8123 3567 8263
rect 3554 8094 3567 8123
rect 3502 8080 3567 8094
rect 2817 8032 2830 8034
rect 2817 7982 2830 7986
rect 2882 7982 2883 8034
rect 2817 7946 2883 7982
rect 3041 8032 3087 8072
rect 3041 7900 3087 7986
rect 3409 8032 3455 8072
rect 3409 7900 3455 7986
rect 3613 8034 3679 8365
rect 4101 8505 4147 8564
rect 4101 8346 4147 8365
rect 4285 8505 4351 8518
rect 4285 8365 4305 8505
rect 4174 8263 4239 8280
rect 4174 8146 4189 8263
rect 4235 8123 4239 8263
rect 4226 8094 4239 8123
rect 4174 8080 4239 8094
rect 3613 7982 3614 8034
rect 3666 8032 3679 8034
rect 3666 7982 3679 7986
rect 3613 7946 3679 7982
rect 4081 8032 4127 8072
rect 4081 7900 4127 7986
rect 4285 8034 4351 8365
rect 4773 8505 4819 8564
rect 5342 8539 5410 8564
rect 4773 8346 4819 8365
rect 4957 8505 5023 8518
rect 4957 8482 4977 8505
rect 4957 8430 4958 8482
rect 4957 8365 4977 8430
rect 4846 8263 4911 8280
rect 4846 8146 4861 8263
rect 4907 8123 4911 8263
rect 4898 8094 4911 8123
rect 4846 8080 4911 8094
rect 4285 7982 4286 8034
rect 4338 8032 4351 8034
rect 4338 7982 4351 7986
rect 4285 7946 4351 7982
rect 4753 8032 4799 8072
rect 4753 7900 4799 7986
rect 4957 8032 5023 8365
rect 5342 8493 5353 8539
rect 5399 8493 5410 8539
rect 5342 8411 5410 8493
rect 5342 8365 5353 8411
rect 5399 8365 5410 8411
rect 5342 8283 5410 8365
rect 5781 8505 5827 8564
rect 5781 8346 5827 8365
rect 5965 8505 6031 8518
rect 5965 8482 5985 8505
rect 5965 8430 5966 8482
rect 5965 8365 5985 8430
rect 5342 8237 5353 8283
rect 5399 8237 5410 8283
rect 5342 8226 5410 8237
rect 5854 8263 5919 8280
rect 5854 8146 5869 8263
rect 5915 8123 5919 8263
rect 5906 8094 5919 8123
rect 5854 8080 5919 8094
rect 4957 7986 4977 8032
rect 4957 7946 5023 7986
rect 5342 8066 5410 8077
rect 5342 7919 5353 8066
rect 5399 7919 5410 8066
rect 5342 7900 5410 7919
rect 5761 8032 5807 8072
rect 5761 7900 5807 7986
rect 5965 8032 6031 8365
rect 6453 8505 6499 8564
rect 6453 8346 6499 8365
rect 6637 8505 6703 8518
rect 6637 8482 6657 8505
rect 6637 8430 6638 8482
rect 6637 8365 6657 8430
rect 6526 8263 6591 8280
rect 6526 8258 6541 8263
rect 6526 8123 6541 8206
rect 6587 8123 6591 8263
rect 6526 8080 6591 8123
rect 5965 7986 5985 8032
rect 5965 7946 6031 7986
rect 6433 8032 6479 8072
rect 6433 7900 6479 7986
rect 6637 8032 6703 8365
rect 7125 8505 7171 8564
rect 7125 8346 7171 8365
rect 7309 8505 7375 8518
rect 7309 8365 7329 8505
rect 7198 8263 7263 8280
rect 7198 8258 7213 8263
rect 7198 8123 7213 8206
rect 7259 8123 7263 8263
rect 7198 8080 7263 8123
rect 6637 7986 6657 8032
rect 6637 7946 6703 7986
rect 7105 8032 7151 8072
rect 7105 7900 7151 7986
rect 7309 8034 7375 8365
rect 7797 8505 7843 8564
rect 7797 8346 7843 8365
rect 7981 8505 8047 8518
rect 7981 8365 8001 8505
rect 7870 8263 7935 8280
rect 7870 8258 7885 8263
rect 7870 8123 7885 8206
rect 7931 8123 7935 8263
rect 7870 8080 7935 8123
rect 7309 7982 7310 8034
rect 7362 8032 7375 8034
rect 7362 7982 7375 7986
rect 7309 7946 7375 7982
rect 7777 8032 7823 8072
rect 7777 7900 7823 7986
rect 7981 8034 8047 8365
rect 8469 8505 8515 8564
rect 8469 8346 8515 8365
rect 8653 8505 8719 8518
rect 8653 8365 8673 8505
rect 8542 8263 8607 8280
rect 8542 8146 8557 8263
rect 8603 8123 8607 8263
rect 8594 8094 8607 8123
rect 8542 8080 8607 8094
rect 7981 7982 7982 8034
rect 8034 8032 8047 8034
rect 8034 7982 8047 7986
rect 7981 7946 8047 7982
rect 8449 8032 8495 8072
rect 8449 7900 8495 7986
rect 8653 8034 8719 8365
rect 9141 8505 9187 8564
rect 9141 8346 9187 8365
rect 9325 8505 9391 8518
rect 9325 8482 9345 8505
rect 9325 8430 9326 8482
rect 9325 8365 9345 8430
rect 9214 8263 9279 8280
rect 9214 8258 9229 8263
rect 9214 8123 9229 8206
rect 9275 8123 9279 8263
rect 9214 8080 9279 8123
rect 8653 7982 8654 8034
rect 8706 8032 8719 8034
rect 8706 7982 8719 7986
rect 8653 7946 8719 7982
rect 9121 8032 9167 8072
rect 9121 7900 9167 7986
rect 9325 8032 9391 8365
rect 9813 8505 9859 8564
rect 9813 8346 9859 8365
rect 9997 8505 10063 8518
rect 9997 8482 10017 8505
rect 9997 8430 9998 8482
rect 9997 8365 10017 8430
rect 9886 8263 9951 8280
rect 9886 8258 9901 8263
rect 9886 8123 9901 8206
rect 9947 8123 9951 8263
rect 9886 8080 9951 8123
rect 9325 7986 9345 8032
rect 9325 7946 9391 7986
rect 9793 8032 9839 8072
rect 9793 7900 9839 7986
rect 9997 8032 10063 8365
rect 10485 8505 10531 8564
rect 10485 8346 10531 8365
rect 10669 8505 10735 8518
rect 10669 8482 10689 8505
rect 10669 8430 10670 8482
rect 10669 8365 10689 8430
rect 10558 8263 10623 8280
rect 10558 8258 10573 8263
rect 10558 8123 10573 8206
rect 10619 8123 10623 8263
rect 10558 8080 10623 8123
rect 9997 7986 10017 8032
rect 9997 7946 10063 7986
rect 10465 8032 10511 8072
rect 10465 7900 10511 7986
rect 10669 8032 10735 8365
rect 10669 7986 10689 8032
rect 10669 7946 10735 7986
rect 11217 8505 11283 8518
rect 11263 8370 11283 8505
rect 11217 8318 11230 8365
rect 11282 8318 11283 8370
rect 11421 8505 11467 8564
rect 11421 8346 11467 8365
rect 11585 8497 11631 8518
rect 11217 8032 11283 8318
rect 11329 8263 11394 8280
rect 11329 8123 11333 8263
rect 11379 8146 11394 8263
rect 11329 8094 11342 8123
rect 11585 8151 11631 8357
rect 11889 8497 11935 8564
rect 11889 8338 11935 8357
rect 12053 8505 12099 8564
rect 12053 8346 12099 8365
rect 12237 8505 12303 8518
rect 12237 8365 12257 8505
rect 11682 8232 11696 8278
rect 11836 8232 11935 8278
rect 11585 8105 11688 8151
rect 11828 8105 11840 8151
rect 11329 8080 11394 8094
rect 11263 7986 11283 8032
rect 11217 7946 11283 7986
rect 11441 8032 11487 8072
rect 11441 7900 11487 7986
rect 11585 8032 11631 8059
rect 11585 7900 11631 7986
rect 11889 8032 11935 8232
rect 12126 8263 12191 8280
rect 12126 8258 12141 8263
rect 12126 8123 12141 8206
rect 12187 8123 12191 8263
rect 12126 8080 12191 8123
rect 12237 8258 12303 8365
rect 12725 8505 12771 8564
rect 13294 8539 13362 8564
rect 12725 8346 12771 8365
rect 12909 8505 12975 8518
rect 12909 8365 12929 8505
rect 12237 8206 12238 8258
rect 12290 8206 12303 8258
rect 11889 7946 11935 7986
rect 12033 8032 12079 8072
rect 12033 7900 12079 7986
rect 12237 8032 12303 8206
rect 12798 8263 12863 8280
rect 12798 8146 12813 8263
rect 12859 8123 12863 8263
rect 12850 8094 12863 8123
rect 12798 8080 12863 8094
rect 12909 8258 12975 8365
rect 12909 8206 12910 8258
rect 12962 8206 12975 8258
rect 13294 8493 13305 8539
rect 13351 8493 13362 8539
rect 13294 8411 13362 8493
rect 13294 8365 13305 8411
rect 13351 8365 13362 8411
rect 13294 8283 13362 8365
rect 13621 8505 13667 8564
rect 13621 8346 13667 8365
rect 13805 8505 13871 8518
rect 13805 8365 13825 8505
rect 13294 8237 13305 8283
rect 13351 8237 13362 8283
rect 13294 8226 13362 8237
rect 13694 8263 13759 8280
rect 13694 8258 13709 8263
rect 12237 7986 12257 8032
rect 12237 7946 12303 7986
rect 12705 8032 12751 8072
rect 12705 7900 12751 7986
rect 12909 8032 12975 8206
rect 13694 8123 13709 8206
rect 13755 8123 13759 8263
rect 13694 8080 13759 8123
rect 13805 8258 13871 8365
rect 14293 8505 14339 8564
rect 14293 8346 14339 8365
rect 14477 8505 14543 8518
rect 14477 8365 14497 8505
rect 13805 8206 13806 8258
rect 13858 8206 13871 8258
rect 12909 7986 12929 8032
rect 12909 7946 12975 7986
rect 13294 8066 13362 8077
rect 13294 7919 13305 8066
rect 13351 7919 13362 8066
rect 13294 7900 13362 7919
rect 13601 8032 13647 8072
rect 13601 7900 13647 7986
rect 13805 8032 13871 8206
rect 14366 8263 14431 8280
rect 14366 8258 14381 8263
rect 14366 8123 14381 8206
rect 14427 8123 14431 8263
rect 14366 8080 14431 8123
rect 14477 8258 14543 8365
rect 14965 8505 15011 8564
rect 14965 8346 15011 8365
rect 15149 8505 15215 8518
rect 15149 8482 15169 8505
rect 15149 8430 15150 8482
rect 15149 8365 15169 8430
rect 14477 8206 14478 8258
rect 14530 8206 14543 8258
rect 13805 7986 13825 8032
rect 13805 7946 13871 7986
rect 14273 8032 14319 8072
rect 14273 7900 14319 7986
rect 14477 8032 14543 8206
rect 15038 8263 15103 8280
rect 15038 8258 15053 8263
rect 15038 8123 15053 8206
rect 15099 8123 15103 8263
rect 15038 8080 15103 8123
rect 14477 7986 14497 8032
rect 14477 7946 14543 7986
rect 14945 8032 14991 8072
rect 14945 7900 14991 7986
rect 15149 8032 15215 8365
rect 15637 8505 15683 8564
rect 15637 8346 15683 8365
rect 15821 8505 15887 8518
rect 15821 8365 15841 8505
rect 15710 8263 15775 8280
rect 15710 8146 15725 8263
rect 15771 8123 15775 8263
rect 15762 8094 15775 8123
rect 15710 8080 15775 8094
rect 15821 8258 15887 8365
rect 16309 8505 16355 8564
rect 16309 8346 16355 8365
rect 16493 8505 16559 8518
rect 16493 8365 16513 8505
rect 15821 8206 15822 8258
rect 15874 8206 15887 8258
rect 15149 7986 15169 8032
rect 15149 7946 15215 7986
rect 15617 8032 15663 8072
rect 15617 7900 15663 7986
rect 15821 8032 15887 8206
rect 16382 8263 16447 8280
rect 16382 8146 16397 8263
rect 16443 8123 16447 8263
rect 16434 8094 16447 8123
rect 16382 8080 16447 8094
rect 16493 8258 16559 8365
rect 16981 8505 17027 8564
rect 16981 8346 17027 8365
rect 17165 8505 17231 8518
rect 17165 8482 17185 8505
rect 17165 8430 17166 8482
rect 17165 8365 17185 8430
rect 16493 8206 16494 8258
rect 16546 8206 16559 8258
rect 15821 7986 15841 8032
rect 15821 7946 15887 7986
rect 16289 8032 16335 8072
rect 16289 7900 16335 7986
rect 16493 8032 16559 8206
rect 17054 8263 17119 8280
rect 17054 8258 17069 8263
rect 17054 8123 17069 8206
rect 17115 8123 17119 8263
rect 17054 8080 17119 8123
rect 16493 7986 16513 8032
rect 16493 7946 16559 7986
rect 16961 8032 17007 8072
rect 16961 7900 17007 7986
rect 17165 8032 17231 8365
rect 17653 8505 17699 8564
rect 17653 8346 17699 8365
rect 17837 8505 17903 8518
rect 17837 8482 17857 8505
rect 17837 8430 17838 8482
rect 17837 8365 17857 8430
rect 17726 8263 17791 8280
rect 17726 8146 17741 8263
rect 17787 8123 17791 8263
rect 17778 8094 17791 8123
rect 17726 8080 17791 8094
rect 17165 7986 17185 8032
rect 17165 7946 17231 7986
rect 17633 8032 17679 8072
rect 17633 7900 17679 7986
rect 17837 8032 17903 8365
rect 18325 8505 18371 8564
rect 18325 8346 18371 8365
rect 18509 8505 18575 8518
rect 18509 8482 18529 8505
rect 18509 8430 18510 8482
rect 18509 8365 18529 8430
rect 18398 8263 18463 8280
rect 18398 8258 18413 8263
rect 18398 8123 18413 8206
rect 18459 8123 18463 8263
rect 18398 8080 18463 8123
rect 17837 7986 17857 8032
rect 17837 7946 17903 7986
rect 18305 8032 18351 8072
rect 18305 7900 18351 7986
rect 18509 8032 18575 8365
rect 18997 8505 19043 8564
rect 18997 8346 19043 8365
rect 19181 8505 19247 8518
rect 19181 8482 19201 8505
rect 19181 8430 19182 8482
rect 19181 8365 19201 8430
rect 19070 8263 19135 8280
rect 19070 8258 19085 8263
rect 19070 8123 19085 8206
rect 19131 8123 19135 8263
rect 19070 8080 19135 8123
rect 18509 7986 18529 8032
rect 18509 7946 18575 7986
rect 18977 8032 19023 8072
rect 18977 7900 19023 7986
rect 19181 8032 19247 8365
rect 19669 8505 19715 8564
rect 19669 8346 19715 8365
rect 19853 8505 19919 8518
rect 19853 8365 19873 8505
rect 19742 8263 19807 8280
rect 19742 8258 19757 8263
rect 19742 8123 19757 8206
rect 19803 8123 19807 8263
rect 19742 8080 19807 8123
rect 19853 8258 19919 8365
rect 19853 8206 19854 8258
rect 19906 8206 19919 8258
rect 19181 7986 19201 8032
rect 19181 7946 19247 7986
rect 19649 8032 19695 8072
rect 19649 7900 19695 7986
rect 19853 8032 19919 8206
rect 19853 7986 19873 8032
rect 19853 7946 19919 7986
rect 20401 8505 20467 8518
rect 20447 8365 20467 8505
rect 20401 8034 20467 8365
rect 20605 8505 20651 8564
rect 20605 8346 20651 8365
rect 20769 8497 20815 8518
rect 20513 8263 20578 8280
rect 20513 8123 20517 8263
rect 20563 8146 20578 8263
rect 20513 8094 20526 8123
rect 20769 8151 20815 8357
rect 21073 8497 21119 8564
rect 21073 8338 21119 8357
rect 21246 8539 21314 8564
rect 21246 8493 21257 8539
rect 21303 8493 21314 8539
rect 21246 8411 21314 8493
rect 21246 8365 21257 8411
rect 21303 8365 21314 8411
rect 21246 8283 21314 8365
rect 20866 8232 20880 8278
rect 21020 8232 21119 8278
rect 20769 8105 20872 8151
rect 21012 8105 21024 8151
rect 20513 8080 20578 8094
rect 20401 8032 20414 8034
rect 20401 7982 20414 7986
rect 20466 7982 20467 8034
rect 20401 7946 20467 7982
rect 20625 8032 20671 8072
rect 20625 7900 20671 7986
rect 20769 8032 20815 8059
rect 20769 7900 20815 7986
rect 21073 8032 21119 8232
rect 21246 8237 21257 8283
rect 21303 8237 21314 8283
rect 21246 8226 21314 8237
rect 21441 8497 21487 8518
rect 21441 8151 21487 8357
rect 21745 8497 21791 8564
rect 21745 8338 21791 8357
rect 21889 8497 21935 8518
rect 21538 8232 21552 8278
rect 21692 8232 21791 8278
rect 21441 8105 21544 8151
rect 21684 8105 21696 8151
rect 21073 7946 21119 7986
rect 21246 8066 21314 8077
rect 21246 7919 21257 8066
rect 21303 7919 21314 8066
rect 21246 7900 21314 7919
rect 21441 8032 21487 8057
rect 21441 7900 21487 7986
rect 21745 8032 21791 8232
rect 21889 8151 21935 8357
rect 22193 8497 22239 8564
rect 22193 8338 22239 8357
rect 22482 8539 22550 8564
rect 22482 8493 22493 8539
rect 22539 8493 22550 8539
rect 22482 8411 22550 8493
rect 22482 8365 22493 8411
rect 22539 8365 22550 8411
rect 22482 8283 22550 8365
rect 21986 8232 22000 8278
rect 22140 8232 22239 8278
rect 21889 8105 21992 8151
rect 22132 8105 22144 8151
rect 21745 7946 21791 7986
rect 21889 8032 21935 8057
rect 21889 7900 21935 7986
rect 22193 8032 22239 8232
rect 22482 8237 22493 8283
rect 22539 8237 22550 8283
rect 22482 8224 22550 8237
rect 22193 7946 22239 7986
rect 22482 8066 22550 8078
rect 22482 7919 22493 8066
rect 22539 7919 22550 8066
rect 22482 7900 22550 7919
rect 1344 7866 22784 7900
rect 1344 7814 6534 7866
rect 6794 7814 11854 7866
rect 12114 7814 17174 7866
rect 17434 7814 22494 7866
rect 22754 7814 22784 7866
rect 1344 7780 22784 7814
rect 1418 7761 1486 7780
rect 1418 7614 1429 7761
rect 1475 7614 1486 7761
rect 1418 7602 1486 7614
rect 2033 7694 2099 7734
rect 2079 7648 2099 7694
rect 1418 7443 1486 7456
rect 1418 7397 1429 7443
rect 1475 7397 1486 7443
rect 1418 7315 1486 7397
rect 1418 7269 1429 7315
rect 1475 7269 1486 7315
rect 1418 7187 1486 7269
rect 1418 7141 1429 7187
rect 1475 7141 1486 7187
rect 2033 7315 2099 7648
rect 2257 7694 2303 7780
rect 2257 7608 2303 7648
rect 2625 7694 2671 7780
rect 2625 7608 2671 7648
rect 2829 7694 2895 7734
rect 2829 7648 2849 7694
rect 2145 7557 2210 7600
rect 2145 7417 2149 7557
rect 2195 7474 2210 7557
rect 2195 7417 2210 7422
rect 2145 7400 2210 7417
rect 2718 7557 2783 7600
rect 2718 7474 2733 7557
rect 2718 7417 2733 7422
rect 2779 7417 2783 7557
rect 2718 7400 2783 7417
rect 2079 7250 2099 7315
rect 2098 7198 2099 7250
rect 2079 7175 2099 7198
rect 2033 7162 2099 7175
rect 2237 7315 2283 7334
rect 1418 7116 1486 7141
rect 2237 7116 2283 7175
rect 2645 7315 2691 7334
rect 2645 7116 2691 7175
rect 2829 7315 2895 7648
rect 3297 7694 3343 7780
rect 3297 7608 3343 7648
rect 3501 7694 3567 7734
rect 3501 7648 3521 7694
rect 3390 7557 3455 7600
rect 3390 7474 3405 7557
rect 3390 7417 3405 7422
rect 3451 7417 3455 7557
rect 3390 7400 3455 7417
rect 2829 7250 2849 7315
rect 2829 7198 2830 7250
rect 2829 7175 2849 7198
rect 2829 7162 2895 7175
rect 3317 7315 3363 7334
rect 3317 7116 3363 7175
rect 3501 7315 3567 7648
rect 3969 7694 4015 7780
rect 3969 7608 4015 7648
rect 4173 7694 4239 7734
rect 4173 7648 4193 7694
rect 4062 7557 4127 7600
rect 4062 7474 4077 7557
rect 4062 7417 4077 7422
rect 4123 7417 4127 7557
rect 4062 7400 4127 7417
rect 3501 7250 3521 7315
rect 3501 7198 3502 7250
rect 3501 7175 3521 7198
rect 3501 7162 3567 7175
rect 3989 7315 4035 7334
rect 3989 7116 4035 7175
rect 4173 7315 4239 7648
rect 4641 7694 4687 7780
rect 4641 7608 4687 7648
rect 4845 7694 4911 7734
rect 4845 7648 4865 7694
rect 4734 7586 4799 7600
rect 4786 7557 4799 7586
rect 4734 7417 4749 7534
rect 4795 7417 4799 7557
rect 4734 7400 4799 7417
rect 4845 7474 4911 7648
rect 5313 7694 5359 7780
rect 5313 7608 5359 7648
rect 5517 7694 5583 7734
rect 5517 7648 5537 7694
rect 4845 7422 4846 7474
rect 4898 7422 4911 7474
rect 4173 7250 4193 7315
rect 4173 7198 4174 7250
rect 4173 7175 4193 7198
rect 4173 7162 4239 7175
rect 4661 7315 4707 7334
rect 4661 7116 4707 7175
rect 4845 7315 4911 7422
rect 5406 7557 5471 7600
rect 5406 7474 5421 7557
rect 5406 7417 5421 7422
rect 5467 7417 5471 7557
rect 5406 7400 5471 7417
rect 4845 7175 4865 7315
rect 4845 7162 4911 7175
rect 5333 7315 5379 7334
rect 5333 7116 5379 7175
rect 5517 7315 5583 7648
rect 5985 7694 6031 7780
rect 5985 7608 6031 7648
rect 6189 7698 6255 7734
rect 6189 7646 6190 7698
rect 6242 7694 6255 7698
rect 6242 7646 6255 7648
rect 6078 7557 6143 7600
rect 6078 7474 6093 7557
rect 6078 7417 6093 7422
rect 6139 7417 6143 7557
rect 6078 7400 6143 7417
rect 5517 7250 5537 7315
rect 5517 7198 5518 7250
rect 5517 7175 5537 7198
rect 5517 7162 5583 7175
rect 6005 7315 6051 7334
rect 6005 7116 6051 7175
rect 6189 7315 6255 7646
rect 6657 7694 6703 7780
rect 6657 7608 6703 7648
rect 6861 7698 6927 7734
rect 6861 7646 6862 7698
rect 6914 7694 6927 7698
rect 6914 7646 6927 7648
rect 6750 7557 6815 7600
rect 6750 7474 6765 7557
rect 6750 7417 6765 7422
rect 6811 7417 6815 7557
rect 6750 7400 6815 7417
rect 6189 7175 6209 7315
rect 6189 7162 6255 7175
rect 6677 7315 6723 7334
rect 6677 7116 6723 7175
rect 6861 7315 6927 7646
rect 7329 7694 7375 7780
rect 7329 7608 7375 7648
rect 7533 7694 7599 7734
rect 7533 7648 7553 7694
rect 7422 7557 7487 7600
rect 7422 7474 7437 7557
rect 7422 7417 7437 7422
rect 7483 7417 7487 7557
rect 7422 7400 7487 7417
rect 6861 7175 6881 7315
rect 6861 7162 6927 7175
rect 7349 7315 7395 7334
rect 7349 7116 7395 7175
rect 7533 7315 7599 7648
rect 8113 7694 8159 7780
rect 8113 7608 8159 7648
rect 8317 7694 8383 7734
rect 8317 7648 8337 7694
rect 8206 7557 8271 7600
rect 8206 7474 8221 7557
rect 8206 7417 8221 7422
rect 8267 7417 8271 7557
rect 8206 7400 8271 7417
rect 7533 7250 7553 7315
rect 7533 7198 7534 7250
rect 7533 7175 7553 7198
rect 7533 7162 7599 7175
rect 8133 7315 8179 7334
rect 8133 7116 8179 7175
rect 8317 7315 8383 7648
rect 8785 7694 8831 7780
rect 9374 7761 9442 7780
rect 8785 7608 8831 7648
rect 8989 7698 9055 7734
rect 8989 7646 8990 7698
rect 9042 7694 9055 7698
rect 9042 7646 9055 7648
rect 8878 7557 8943 7600
rect 8878 7474 8893 7557
rect 8878 7417 8893 7422
rect 8939 7417 8943 7557
rect 8878 7400 8943 7417
rect 8317 7250 8337 7315
rect 8317 7198 8318 7250
rect 8317 7175 8337 7198
rect 8317 7162 8383 7175
rect 8805 7315 8851 7334
rect 8805 7116 8851 7175
rect 8989 7315 9055 7646
rect 9374 7614 9385 7761
rect 9431 7614 9442 7761
rect 9374 7603 9442 7614
rect 9793 7694 9839 7780
rect 9793 7608 9839 7648
rect 9997 7698 10063 7734
rect 9997 7646 9998 7698
rect 10050 7694 10063 7698
rect 10050 7646 10063 7648
rect 9886 7557 9951 7600
rect 9886 7474 9901 7557
rect 8989 7175 9009 7315
rect 8989 7162 9055 7175
rect 9374 7443 9442 7454
rect 9374 7397 9385 7443
rect 9431 7397 9442 7443
rect 9886 7417 9901 7422
rect 9947 7417 9951 7557
rect 9886 7400 9951 7417
rect 9374 7315 9442 7397
rect 9374 7269 9385 7315
rect 9431 7269 9442 7315
rect 9374 7187 9442 7269
rect 9374 7141 9385 7187
rect 9431 7141 9442 7187
rect 9374 7116 9442 7141
rect 9813 7315 9859 7334
rect 9813 7116 9859 7175
rect 9997 7315 10063 7646
rect 10465 7694 10511 7780
rect 10465 7608 10511 7648
rect 10669 7698 10735 7734
rect 10669 7646 10670 7698
rect 10722 7694 10735 7698
rect 10722 7646 10735 7648
rect 10558 7586 10623 7600
rect 10610 7557 10623 7586
rect 10558 7417 10573 7534
rect 10619 7417 10623 7557
rect 10558 7400 10623 7417
rect 9997 7175 10017 7315
rect 9997 7162 10063 7175
rect 10485 7315 10531 7334
rect 10485 7116 10531 7175
rect 10669 7315 10735 7646
rect 10669 7175 10689 7315
rect 10669 7162 10735 7175
rect 11217 7698 11283 7734
rect 11217 7694 11230 7698
rect 11217 7646 11230 7648
rect 11282 7646 11283 7698
rect 11217 7315 11283 7646
rect 11441 7694 11487 7780
rect 11441 7608 11487 7648
rect 11809 7694 11855 7780
rect 11809 7608 11855 7648
rect 12013 7694 12079 7734
rect 12013 7648 12033 7694
rect 11329 7557 11394 7600
rect 11329 7417 11333 7557
rect 11379 7474 11394 7557
rect 11379 7417 11394 7422
rect 11329 7400 11394 7417
rect 11902 7557 11967 7600
rect 11902 7474 11917 7557
rect 11902 7417 11917 7422
rect 11963 7417 11967 7557
rect 11902 7400 11967 7417
rect 11263 7175 11283 7315
rect 11217 7162 11283 7175
rect 11421 7315 11467 7334
rect 11421 7116 11467 7175
rect 11829 7315 11875 7334
rect 11829 7116 11875 7175
rect 12013 7315 12079 7648
rect 12481 7694 12527 7780
rect 12481 7608 12527 7648
rect 12685 7694 12751 7734
rect 12685 7648 12705 7694
rect 12574 7557 12639 7600
rect 12574 7474 12589 7557
rect 12574 7417 12589 7422
rect 12635 7417 12639 7557
rect 12574 7400 12639 7417
rect 12013 7250 12033 7315
rect 12013 7198 12014 7250
rect 12013 7175 12033 7198
rect 12013 7162 12079 7175
rect 12501 7315 12547 7334
rect 12501 7116 12547 7175
rect 12685 7315 12751 7648
rect 13153 7694 13199 7780
rect 13153 7608 13199 7648
rect 13357 7698 13423 7734
rect 13357 7646 13358 7698
rect 13410 7694 13423 7698
rect 13410 7646 13423 7648
rect 13246 7557 13311 7600
rect 13246 7474 13261 7557
rect 13246 7417 13261 7422
rect 13307 7417 13311 7557
rect 13246 7400 13311 7417
rect 12685 7250 12705 7315
rect 12685 7198 12686 7250
rect 12685 7175 12705 7198
rect 12685 7162 12751 7175
rect 13173 7315 13219 7334
rect 13173 7116 13219 7175
rect 13357 7315 13423 7646
rect 13825 7694 13871 7780
rect 13825 7608 13871 7648
rect 14029 7694 14095 7734
rect 14029 7648 14049 7694
rect 13918 7586 13983 7600
rect 13970 7557 13983 7586
rect 13918 7417 13933 7534
rect 13979 7417 13983 7557
rect 13918 7400 13983 7417
rect 14029 7362 14095 7648
rect 14497 7694 14543 7780
rect 14497 7608 14543 7648
rect 14701 7698 14767 7734
rect 14701 7646 14702 7698
rect 14754 7694 14767 7698
rect 14754 7646 14767 7648
rect 14590 7557 14655 7600
rect 14590 7474 14605 7557
rect 14590 7417 14605 7422
rect 14651 7417 14655 7557
rect 14590 7400 14655 7417
rect 13357 7175 13377 7315
rect 13357 7162 13423 7175
rect 13845 7315 13891 7334
rect 13845 7116 13891 7175
rect 14029 7310 14030 7362
rect 14082 7315 14095 7362
rect 14029 7175 14049 7310
rect 14029 7162 14095 7175
rect 14517 7315 14563 7334
rect 14517 7116 14563 7175
rect 14701 7315 14767 7646
rect 15169 7694 15215 7780
rect 15169 7608 15215 7648
rect 15373 7694 15439 7734
rect 15373 7648 15393 7694
rect 15262 7586 15327 7600
rect 15314 7557 15327 7586
rect 15262 7417 15277 7534
rect 15323 7417 15327 7557
rect 15262 7400 15327 7417
rect 14701 7175 14721 7315
rect 14701 7162 14767 7175
rect 15189 7315 15235 7334
rect 15189 7116 15235 7175
rect 15373 7315 15439 7648
rect 15841 7694 15887 7780
rect 15841 7608 15887 7648
rect 16045 7694 16111 7734
rect 16045 7648 16065 7694
rect 15934 7586 15999 7600
rect 15986 7557 15999 7586
rect 15934 7417 15949 7534
rect 15995 7417 15999 7557
rect 15934 7400 15999 7417
rect 15373 7250 15393 7315
rect 15373 7198 15374 7250
rect 15373 7175 15393 7198
rect 15373 7162 15439 7175
rect 15861 7315 15907 7334
rect 15861 7116 15907 7175
rect 16045 7315 16111 7648
rect 16513 7694 16559 7780
rect 17326 7761 17394 7780
rect 16513 7608 16559 7648
rect 16717 7698 16783 7734
rect 16717 7646 16718 7698
rect 16770 7694 16783 7698
rect 16770 7646 16783 7648
rect 16606 7557 16671 7600
rect 16606 7474 16621 7557
rect 16606 7417 16621 7422
rect 16667 7417 16671 7557
rect 16606 7400 16671 7417
rect 16045 7250 16065 7315
rect 16045 7198 16046 7250
rect 16045 7175 16065 7198
rect 16045 7162 16111 7175
rect 16533 7315 16579 7334
rect 16533 7116 16579 7175
rect 16717 7315 16783 7646
rect 17326 7614 17337 7761
rect 17383 7614 17394 7761
rect 17326 7603 17394 7614
rect 17633 7694 17679 7780
rect 17633 7608 17679 7648
rect 17837 7698 17903 7734
rect 17837 7646 17838 7698
rect 17890 7694 17903 7698
rect 17890 7646 17903 7648
rect 17726 7557 17791 7600
rect 17726 7474 17741 7557
rect 16717 7175 16737 7315
rect 16717 7162 16783 7175
rect 17326 7443 17394 7454
rect 17326 7397 17337 7443
rect 17383 7397 17394 7443
rect 17726 7417 17741 7422
rect 17787 7417 17791 7557
rect 17726 7400 17791 7417
rect 17326 7315 17394 7397
rect 17326 7269 17337 7315
rect 17383 7269 17394 7315
rect 17326 7187 17394 7269
rect 17326 7141 17337 7187
rect 17383 7141 17394 7187
rect 17326 7116 17394 7141
rect 17653 7315 17699 7334
rect 17653 7116 17699 7175
rect 17837 7315 17903 7646
rect 18305 7694 18351 7780
rect 18305 7608 18351 7648
rect 18509 7698 18575 7734
rect 18509 7646 18510 7698
rect 18562 7694 18575 7698
rect 18562 7646 18575 7648
rect 18398 7557 18463 7600
rect 18398 7474 18413 7557
rect 18398 7417 18413 7422
rect 18459 7417 18463 7557
rect 18398 7400 18463 7417
rect 17837 7175 17857 7315
rect 17837 7162 17903 7175
rect 18325 7315 18371 7334
rect 18325 7116 18371 7175
rect 18509 7315 18575 7646
rect 18977 7694 19023 7780
rect 18977 7608 19023 7648
rect 19181 7694 19247 7734
rect 19181 7648 19201 7694
rect 19070 7557 19135 7600
rect 19070 7474 19085 7557
rect 19070 7417 19085 7422
rect 19131 7417 19135 7557
rect 19070 7400 19135 7417
rect 18509 7175 18529 7315
rect 18509 7162 18575 7175
rect 18997 7315 19043 7334
rect 18997 7116 19043 7175
rect 19181 7315 19247 7648
rect 19649 7694 19695 7780
rect 19649 7608 19695 7648
rect 19853 7694 19919 7734
rect 19853 7648 19873 7694
rect 19742 7557 19807 7600
rect 19742 7474 19757 7557
rect 19742 7417 19757 7422
rect 19803 7417 19807 7557
rect 19742 7400 19807 7417
rect 19181 7250 19201 7315
rect 19181 7198 19182 7250
rect 19181 7175 19201 7198
rect 19181 7162 19247 7175
rect 19669 7315 19715 7334
rect 19669 7116 19715 7175
rect 19853 7315 19919 7648
rect 20321 7694 20367 7780
rect 20321 7608 20367 7648
rect 20525 7694 20591 7734
rect 20525 7648 20545 7694
rect 20414 7557 20479 7600
rect 20414 7474 20429 7557
rect 20414 7417 20429 7422
rect 20475 7417 20479 7557
rect 20414 7400 20479 7417
rect 19853 7250 19873 7315
rect 19853 7198 19854 7250
rect 19853 7175 19873 7198
rect 19853 7162 19919 7175
rect 20341 7315 20387 7334
rect 20341 7116 20387 7175
rect 20525 7315 20591 7648
rect 20993 7694 21039 7780
rect 20993 7608 21039 7648
rect 21197 7694 21263 7734
rect 21197 7648 21217 7694
rect 21086 7557 21151 7600
rect 21086 7474 21101 7557
rect 21086 7417 21101 7422
rect 21147 7417 21151 7557
rect 21086 7400 21151 7417
rect 20525 7250 20545 7315
rect 20525 7198 20526 7250
rect 20525 7175 20545 7198
rect 20525 7162 20591 7175
rect 21013 7315 21059 7334
rect 21013 7116 21059 7175
rect 21197 7315 21263 7648
rect 21441 7694 21487 7780
rect 21441 7623 21487 7648
rect 21745 7694 21791 7734
rect 21197 7250 21217 7315
rect 21197 7198 21198 7250
rect 21197 7175 21217 7198
rect 21197 7162 21263 7175
rect 21441 7529 21544 7575
rect 21684 7529 21696 7575
rect 21441 7323 21487 7529
rect 21745 7448 21791 7648
rect 21889 7694 21935 7780
rect 22482 7761 22550 7780
rect 21889 7623 21935 7648
rect 22193 7694 22239 7734
rect 21538 7402 21552 7448
rect 21692 7402 21791 7448
rect 21889 7529 21992 7575
rect 22132 7529 22144 7575
rect 21441 7162 21487 7183
rect 21745 7323 21791 7342
rect 21745 7116 21791 7183
rect 21889 7323 21935 7529
rect 22193 7448 22239 7648
rect 22482 7614 22493 7761
rect 22539 7614 22550 7761
rect 22482 7602 22550 7614
rect 21986 7402 22000 7448
rect 22140 7402 22239 7448
rect 22482 7443 22550 7456
rect 22482 7397 22493 7443
rect 22539 7397 22550 7443
rect 21889 7162 21935 7183
rect 22193 7323 22239 7342
rect 22193 7116 22239 7183
rect 22482 7315 22550 7397
rect 22482 7269 22493 7315
rect 22539 7269 22550 7315
rect 22482 7187 22550 7269
rect 22482 7141 22493 7187
rect 22539 7141 22550 7187
rect 22482 7116 22550 7141
rect 1344 7082 22624 7116
rect 1344 7030 3874 7082
rect 4134 7030 9194 7082
rect 9454 7030 14514 7082
rect 14774 7030 19834 7082
rect 20094 7030 22624 7082
rect 1344 6996 22624 7030
rect 1418 6971 1486 6996
rect 1418 6925 1429 6971
rect 1475 6925 1486 6971
rect 1418 6843 1486 6925
rect 1418 6797 1429 6843
rect 1475 6797 1486 6843
rect 1418 6715 1486 6797
rect 1418 6669 1429 6715
rect 1475 6669 1486 6715
rect 1418 6656 1486 6669
rect 1617 6929 1663 6950
rect 1617 6583 1663 6789
rect 1921 6929 1967 6996
rect 1921 6770 1967 6789
rect 2085 6937 2131 6996
rect 2085 6778 2131 6797
rect 2269 6937 2335 6950
rect 2269 6797 2289 6937
rect 1714 6664 1728 6710
rect 1868 6664 1967 6710
rect 1617 6537 1720 6583
rect 1860 6537 1872 6583
rect 1418 6498 1486 6510
rect 1418 6351 1429 6498
rect 1475 6351 1486 6498
rect 1418 6332 1486 6351
rect 1617 6464 1663 6491
rect 1617 6332 1663 6418
rect 1921 6464 1967 6664
rect 2158 6695 2223 6712
rect 2158 6578 2173 6695
rect 2219 6555 2223 6695
rect 2210 6526 2223 6555
rect 2158 6512 2223 6526
rect 1921 6378 1967 6418
rect 2065 6464 2111 6504
rect 2065 6332 2111 6418
rect 2269 6466 2335 6797
rect 2757 6937 2803 6996
rect 2757 6778 2803 6797
rect 2941 6937 3007 6950
rect 2941 6797 2961 6937
rect 2830 6695 2895 6712
rect 2830 6578 2845 6695
rect 2891 6555 2895 6695
rect 2882 6526 2895 6555
rect 2830 6512 2895 6526
rect 2269 6414 2270 6466
rect 2322 6464 2335 6466
rect 2322 6414 2335 6418
rect 2269 6378 2335 6414
rect 2737 6464 2783 6504
rect 2737 6332 2783 6418
rect 2941 6466 3007 6797
rect 3429 6937 3475 6996
rect 3429 6778 3475 6797
rect 3613 6937 3679 6950
rect 3613 6797 3633 6937
rect 3502 6695 3567 6712
rect 3502 6578 3517 6695
rect 3563 6555 3567 6695
rect 3554 6526 3567 6555
rect 3502 6512 3567 6526
rect 2941 6414 2942 6466
rect 2994 6464 3007 6466
rect 2994 6414 3007 6418
rect 2941 6378 3007 6414
rect 3409 6464 3455 6504
rect 3409 6332 3455 6418
rect 3613 6466 3679 6797
rect 4101 6937 4147 6996
rect 4101 6778 4147 6797
rect 4285 6937 4351 6950
rect 4285 6914 4305 6937
rect 4285 6862 4286 6914
rect 4285 6797 4305 6862
rect 4174 6695 4239 6712
rect 4174 6578 4189 6695
rect 4235 6555 4239 6695
rect 4226 6526 4239 6555
rect 4174 6512 4239 6526
rect 3613 6414 3614 6466
rect 3666 6464 3679 6466
rect 3666 6414 3679 6418
rect 3613 6378 3679 6414
rect 4081 6464 4127 6504
rect 4081 6332 4127 6418
rect 4285 6464 4351 6797
rect 4773 6937 4819 6996
rect 5342 6971 5410 6996
rect 4773 6778 4819 6797
rect 4957 6937 5023 6950
rect 4957 6914 4977 6937
rect 4957 6862 4958 6914
rect 4957 6797 4977 6862
rect 4846 6695 4911 6712
rect 4846 6578 4861 6695
rect 4907 6555 4911 6695
rect 4898 6526 4911 6555
rect 4846 6512 4911 6526
rect 4285 6418 4305 6464
rect 4285 6378 4351 6418
rect 4753 6464 4799 6504
rect 4753 6332 4799 6418
rect 4957 6464 5023 6797
rect 5342 6925 5353 6971
rect 5399 6925 5410 6971
rect 5342 6843 5410 6925
rect 5342 6797 5353 6843
rect 5399 6797 5410 6843
rect 5342 6715 5410 6797
rect 5669 6937 5715 6996
rect 5669 6778 5715 6797
rect 5853 6937 5919 6950
rect 5853 6797 5873 6937
rect 5342 6669 5353 6715
rect 5399 6669 5410 6715
rect 5342 6658 5410 6669
rect 5742 6695 5807 6712
rect 5742 6690 5757 6695
rect 5742 6555 5757 6638
rect 5803 6555 5807 6695
rect 5742 6512 5807 6555
rect 5853 6690 5919 6797
rect 6341 6937 6387 6996
rect 6341 6778 6387 6797
rect 6525 6937 6591 6950
rect 6525 6797 6545 6937
rect 5853 6638 5854 6690
rect 5906 6638 5919 6690
rect 4957 6418 4977 6464
rect 4957 6378 5023 6418
rect 5342 6498 5410 6509
rect 5342 6351 5353 6498
rect 5399 6351 5410 6498
rect 5342 6332 5410 6351
rect 5649 6464 5695 6504
rect 5649 6332 5695 6418
rect 5853 6464 5919 6638
rect 6414 6695 6479 6712
rect 6414 6690 6429 6695
rect 6414 6555 6429 6638
rect 6475 6555 6479 6695
rect 6414 6512 6479 6555
rect 6525 6690 6591 6797
rect 7013 6937 7059 6996
rect 7013 6778 7059 6797
rect 7197 6937 7263 6950
rect 7197 6797 7217 6937
rect 6525 6638 6526 6690
rect 6578 6638 6591 6690
rect 5853 6418 5873 6464
rect 5853 6378 5919 6418
rect 6321 6464 6367 6504
rect 6321 6332 6367 6418
rect 6525 6464 6591 6638
rect 7086 6695 7151 6712
rect 7086 6578 7101 6695
rect 7147 6555 7151 6695
rect 7138 6526 7151 6555
rect 7086 6512 7151 6526
rect 6525 6418 6545 6464
rect 6525 6378 6591 6418
rect 6993 6464 7039 6504
rect 6993 6332 7039 6418
rect 7197 6466 7263 6797
rect 7685 6937 7731 6996
rect 7685 6778 7731 6797
rect 7869 6937 7935 6950
rect 7869 6797 7889 6937
rect 7758 6695 7823 6712
rect 7758 6578 7773 6695
rect 7819 6555 7823 6695
rect 7810 6526 7823 6555
rect 7758 6512 7823 6526
rect 7197 6414 7198 6466
rect 7250 6464 7263 6466
rect 7250 6414 7263 6418
rect 7197 6378 7263 6414
rect 7665 6464 7711 6504
rect 7665 6332 7711 6418
rect 7869 6466 7935 6797
rect 8357 6937 8403 6996
rect 8357 6778 8403 6797
rect 8541 6937 8607 6950
rect 8541 6797 8561 6937
rect 8430 6695 8495 6712
rect 8430 6578 8445 6695
rect 8491 6555 8495 6695
rect 8482 6526 8495 6555
rect 8430 6512 8495 6526
rect 8541 6690 8607 6797
rect 9029 6937 9075 6996
rect 9029 6778 9075 6797
rect 9213 6937 9279 6950
rect 9213 6797 9233 6937
rect 8541 6638 8542 6690
rect 8594 6638 8607 6690
rect 7869 6414 7870 6466
rect 7922 6464 7935 6466
rect 7922 6414 7935 6418
rect 7869 6378 7935 6414
rect 8337 6464 8383 6504
rect 8337 6332 8383 6418
rect 8541 6464 8607 6638
rect 9102 6695 9167 6712
rect 9102 6578 9117 6695
rect 9163 6555 9167 6695
rect 9154 6526 9167 6555
rect 9102 6512 9167 6526
rect 9213 6690 9279 6797
rect 9701 6937 9747 6996
rect 9701 6778 9747 6797
rect 9885 6937 9951 6950
rect 9885 6797 9905 6937
rect 9213 6638 9214 6690
rect 9266 6638 9279 6690
rect 8541 6418 8561 6464
rect 8541 6378 8607 6418
rect 9009 6464 9055 6504
rect 9009 6332 9055 6418
rect 9213 6464 9279 6638
rect 9774 6695 9839 6712
rect 9774 6690 9789 6695
rect 9774 6555 9789 6638
rect 9835 6555 9839 6695
rect 9774 6512 9839 6555
rect 9213 6418 9233 6464
rect 9213 6378 9279 6418
rect 9681 6464 9727 6504
rect 9681 6332 9727 6418
rect 9885 6466 9951 6797
rect 10373 6937 10419 6996
rect 10373 6778 10419 6797
rect 10557 6937 10623 6950
rect 10557 6914 10577 6937
rect 10557 6862 10558 6914
rect 10557 6797 10577 6862
rect 10446 6695 10511 6712
rect 10446 6690 10461 6695
rect 10446 6555 10461 6638
rect 10507 6555 10511 6695
rect 10446 6512 10511 6555
rect 9885 6414 9886 6466
rect 9938 6464 9951 6466
rect 9938 6414 9951 6418
rect 9885 6378 9951 6414
rect 10353 6464 10399 6504
rect 10353 6332 10399 6418
rect 10557 6464 10623 6797
rect 11045 6937 11091 6996
rect 11045 6778 11091 6797
rect 11229 6937 11295 6950
rect 11229 6914 11249 6937
rect 11229 6862 11230 6914
rect 11229 6797 11249 6862
rect 11118 6695 11183 6712
rect 11118 6690 11133 6695
rect 11118 6555 11133 6638
rect 11179 6555 11183 6695
rect 11118 6512 11183 6555
rect 10557 6418 10577 6464
rect 10557 6378 10623 6418
rect 11025 6464 11071 6504
rect 11025 6332 11071 6418
rect 11229 6464 11295 6797
rect 11717 6937 11763 6996
rect 11717 6778 11763 6797
rect 11901 6937 11967 6950
rect 11901 6797 11921 6937
rect 11790 6695 11855 6712
rect 11790 6690 11805 6695
rect 11790 6555 11805 6638
rect 11851 6555 11855 6695
rect 11790 6512 11855 6555
rect 11229 6418 11249 6464
rect 11229 6378 11295 6418
rect 11697 6464 11743 6504
rect 11697 6332 11743 6418
rect 11901 6466 11967 6797
rect 12389 6937 12435 6996
rect 12389 6778 12435 6797
rect 12573 6937 12639 6950
rect 12573 6797 12593 6937
rect 12462 6695 12527 6712
rect 12462 6690 12477 6695
rect 12462 6555 12477 6638
rect 12523 6555 12527 6695
rect 12462 6512 12527 6555
rect 11901 6414 11902 6466
rect 11954 6464 11967 6466
rect 11954 6414 11967 6418
rect 11901 6378 11967 6414
rect 12369 6464 12415 6504
rect 12369 6332 12415 6418
rect 12573 6466 12639 6797
rect 12817 6929 12863 6950
rect 12817 6583 12863 6789
rect 13121 6929 13167 6996
rect 13121 6770 13167 6789
rect 13294 6971 13362 6996
rect 13294 6925 13305 6971
rect 13351 6925 13362 6971
rect 13294 6843 13362 6925
rect 13294 6797 13305 6843
rect 13351 6797 13362 6843
rect 13294 6715 13362 6797
rect 12914 6664 12928 6710
rect 13068 6664 13167 6710
rect 12817 6537 12920 6583
rect 13060 6537 13072 6583
rect 12573 6414 12574 6466
rect 12626 6464 12639 6466
rect 12626 6414 12639 6418
rect 12573 6378 12639 6414
rect 12817 6464 12863 6491
rect 12817 6332 12863 6418
rect 13121 6464 13167 6664
rect 13294 6669 13305 6715
rect 13351 6669 13362 6715
rect 13294 6658 13362 6669
rect 13489 6929 13535 6950
rect 13489 6583 13535 6789
rect 13793 6929 13839 6996
rect 13793 6770 13839 6789
rect 14069 6937 14115 6996
rect 14069 6778 14115 6797
rect 14253 6937 14319 6950
rect 14253 6914 14273 6937
rect 14253 6862 14254 6914
rect 14253 6797 14273 6862
rect 13586 6664 13600 6710
rect 13740 6664 13839 6710
rect 13489 6537 13592 6583
rect 13732 6537 13744 6583
rect 13121 6378 13167 6418
rect 13294 6498 13362 6509
rect 13294 6351 13305 6498
rect 13351 6351 13362 6498
rect 13294 6332 13362 6351
rect 13489 6464 13535 6491
rect 13489 6332 13535 6418
rect 13793 6464 13839 6664
rect 14142 6695 14207 6712
rect 14142 6690 14157 6695
rect 14142 6555 14157 6638
rect 14203 6555 14207 6695
rect 14142 6512 14207 6555
rect 13793 6378 13839 6418
rect 14049 6464 14095 6504
rect 14049 6332 14095 6418
rect 14253 6464 14319 6797
rect 14741 6937 14787 6996
rect 14741 6778 14787 6797
rect 14925 6937 14991 6950
rect 14925 6914 14945 6937
rect 14925 6862 14926 6914
rect 14925 6797 14945 6862
rect 14814 6695 14879 6712
rect 14814 6690 14829 6695
rect 14814 6555 14829 6638
rect 14875 6555 14879 6695
rect 14814 6512 14879 6555
rect 14253 6418 14273 6464
rect 14253 6378 14319 6418
rect 14721 6464 14767 6504
rect 14721 6332 14767 6418
rect 14925 6464 14991 6797
rect 15413 6937 15459 6996
rect 15413 6778 15459 6797
rect 15597 6937 15663 6950
rect 15597 6914 15617 6937
rect 15597 6862 15598 6914
rect 15597 6797 15617 6862
rect 15486 6695 15551 6712
rect 15486 6690 15501 6695
rect 15486 6555 15501 6638
rect 15547 6555 15551 6695
rect 15486 6512 15551 6555
rect 14925 6418 14945 6464
rect 14925 6378 14991 6418
rect 15393 6464 15439 6504
rect 15393 6332 15439 6418
rect 15597 6464 15663 6797
rect 16085 6937 16131 6996
rect 16085 6778 16131 6797
rect 16269 6937 16335 6950
rect 16269 6797 16289 6937
rect 16158 6695 16223 6712
rect 16158 6578 16173 6695
rect 16219 6555 16223 6695
rect 16210 6526 16223 6555
rect 16158 6512 16223 6526
rect 16269 6578 16335 6797
rect 16757 6937 16803 6996
rect 16757 6778 16803 6797
rect 16941 6937 17007 6950
rect 16941 6797 16961 6937
rect 16269 6526 16270 6578
rect 16322 6526 16335 6578
rect 15597 6418 15617 6464
rect 15597 6378 15663 6418
rect 16065 6464 16111 6504
rect 16065 6332 16111 6418
rect 16269 6464 16335 6526
rect 16830 6695 16895 6712
rect 16830 6578 16845 6695
rect 16891 6555 16895 6695
rect 16882 6526 16895 6555
rect 16830 6512 16895 6526
rect 16941 6578 17007 6797
rect 17429 6937 17475 6996
rect 17429 6778 17475 6797
rect 17613 6937 17679 6950
rect 17613 6914 17633 6937
rect 17613 6862 17614 6914
rect 17613 6797 17633 6862
rect 16941 6526 16942 6578
rect 16994 6526 17007 6578
rect 16269 6418 16289 6464
rect 16269 6378 16335 6418
rect 16737 6464 16783 6504
rect 16737 6332 16783 6418
rect 16941 6464 17007 6526
rect 17502 6695 17567 6712
rect 17502 6578 17517 6695
rect 17563 6555 17567 6695
rect 17554 6526 17567 6555
rect 17502 6512 17567 6526
rect 16941 6418 16961 6464
rect 16941 6378 17007 6418
rect 17409 6464 17455 6504
rect 17409 6332 17455 6418
rect 17613 6464 17679 6797
rect 18101 6937 18147 6996
rect 18101 6778 18147 6797
rect 18285 6937 18351 6950
rect 18285 6797 18305 6937
rect 18174 6695 18239 6712
rect 18174 6578 18189 6695
rect 18235 6555 18239 6695
rect 18226 6526 18239 6555
rect 18174 6512 18239 6526
rect 17613 6418 17633 6464
rect 17613 6378 17679 6418
rect 18081 6464 18127 6504
rect 18081 6332 18127 6418
rect 18285 6466 18351 6797
rect 18773 6937 18819 6996
rect 18773 6778 18819 6797
rect 18957 6937 19023 6950
rect 18957 6797 18977 6937
rect 18846 6695 18911 6712
rect 18846 6578 18861 6695
rect 18907 6555 18911 6695
rect 18898 6526 18911 6555
rect 18846 6512 18911 6526
rect 18957 6690 19023 6797
rect 19445 6937 19491 6996
rect 19445 6778 19491 6797
rect 19629 6937 19695 6950
rect 19629 6914 19649 6937
rect 19629 6862 19630 6914
rect 19629 6797 19649 6862
rect 18957 6638 18958 6690
rect 19010 6638 19023 6690
rect 18285 6414 18286 6466
rect 18338 6464 18351 6466
rect 18338 6414 18351 6418
rect 18285 6378 18351 6414
rect 18753 6464 18799 6504
rect 18753 6332 18799 6418
rect 18957 6464 19023 6638
rect 19518 6695 19583 6712
rect 19518 6578 19533 6695
rect 19579 6555 19583 6695
rect 19570 6526 19583 6555
rect 19518 6512 19583 6526
rect 18957 6418 18977 6464
rect 18957 6378 19023 6418
rect 19425 6464 19471 6504
rect 19425 6332 19471 6418
rect 19629 6464 19695 6797
rect 19629 6418 19649 6464
rect 19629 6378 19695 6418
rect 20177 6937 20243 6950
rect 20223 6797 20243 6937
rect 20177 6466 20243 6797
rect 20381 6937 20427 6996
rect 20381 6778 20427 6797
rect 20545 6929 20591 6950
rect 20289 6695 20354 6712
rect 20289 6555 20293 6695
rect 20339 6578 20354 6695
rect 20289 6526 20302 6555
rect 20545 6583 20591 6789
rect 20849 6929 20895 6996
rect 20849 6770 20895 6789
rect 21246 6971 21314 6996
rect 21246 6925 21257 6971
rect 21303 6925 21314 6971
rect 21246 6843 21314 6925
rect 21246 6797 21257 6843
rect 21303 6797 21314 6843
rect 21246 6715 21314 6797
rect 21573 6937 21619 6996
rect 21573 6778 21619 6797
rect 21757 6937 21823 6950
rect 21757 6797 21777 6937
rect 20642 6664 20656 6710
rect 20796 6664 20895 6710
rect 20545 6537 20648 6583
rect 20788 6537 20800 6583
rect 20289 6512 20354 6526
rect 20177 6464 20190 6466
rect 20177 6414 20190 6418
rect 20242 6414 20243 6466
rect 20177 6378 20243 6414
rect 20401 6464 20447 6504
rect 20401 6332 20447 6418
rect 20545 6464 20591 6491
rect 20545 6332 20591 6418
rect 20849 6464 20895 6664
rect 21246 6669 21257 6715
rect 21303 6669 21314 6715
rect 21246 6658 21314 6669
rect 21646 6695 21711 6712
rect 21646 6690 21661 6695
rect 21646 6555 21661 6638
rect 21707 6555 21711 6695
rect 21646 6512 21711 6555
rect 20849 6378 20895 6418
rect 21246 6498 21314 6509
rect 21246 6351 21257 6498
rect 21303 6351 21314 6498
rect 21246 6332 21314 6351
rect 21553 6464 21599 6504
rect 21553 6332 21599 6418
rect 21757 6466 21823 6797
rect 22001 6929 22047 6950
rect 22001 6583 22047 6789
rect 22305 6929 22351 6996
rect 22305 6770 22351 6789
rect 22482 6971 22550 6996
rect 22482 6925 22493 6971
rect 22539 6925 22550 6971
rect 22482 6843 22550 6925
rect 22482 6797 22493 6843
rect 22539 6797 22550 6843
rect 22482 6715 22550 6797
rect 22098 6664 22112 6710
rect 22252 6664 22351 6710
rect 22001 6537 22104 6583
rect 22244 6537 22256 6583
rect 21757 6414 21758 6466
rect 21810 6464 21823 6466
rect 21810 6414 21823 6418
rect 21757 6378 21823 6414
rect 22001 6464 22047 6491
rect 22001 6332 22047 6418
rect 22305 6464 22351 6664
rect 22482 6669 22493 6715
rect 22539 6669 22550 6715
rect 22482 6656 22550 6669
rect 22305 6378 22351 6418
rect 22482 6498 22550 6510
rect 22482 6351 22493 6498
rect 22539 6351 22550 6498
rect 22482 6332 22550 6351
rect 1344 6298 22784 6332
rect 1344 6246 6534 6298
rect 6794 6246 11854 6298
rect 12114 6246 17174 6298
rect 17434 6246 22494 6298
rect 22754 6246 22784 6298
rect 1344 6212 22784 6246
rect 1418 6193 1486 6212
rect 1418 6046 1429 6193
rect 1475 6046 1486 6193
rect 1418 6034 1486 6046
rect 1953 6126 1999 6212
rect 1953 6040 1999 6080
rect 2157 6126 2223 6166
rect 2157 6080 2177 6126
rect 2046 5989 2111 6032
rect 2046 5906 2061 5989
rect 1418 5875 1486 5888
rect 1418 5829 1429 5875
rect 1475 5829 1486 5875
rect 2046 5849 2061 5854
rect 2107 5849 2111 5989
rect 2046 5832 2111 5849
rect 1418 5747 1486 5829
rect 1418 5701 1429 5747
rect 1475 5701 1486 5747
rect 1418 5619 1486 5701
rect 1418 5573 1429 5619
rect 1475 5573 1486 5619
rect 1418 5548 1486 5573
rect 1973 5747 2019 5766
rect 1973 5548 2019 5607
rect 2157 5747 2223 6080
rect 2625 6126 2671 6212
rect 2625 6040 2671 6080
rect 2829 6126 2895 6166
rect 2829 6080 2849 6126
rect 2718 5989 2783 6032
rect 2718 5906 2733 5989
rect 2718 5849 2733 5854
rect 2779 5849 2783 5989
rect 2718 5832 2783 5849
rect 2157 5682 2177 5747
rect 2157 5630 2158 5682
rect 2157 5607 2177 5630
rect 2157 5594 2223 5607
rect 2645 5747 2691 5766
rect 2645 5548 2691 5607
rect 2829 5747 2895 6080
rect 3297 6126 3343 6212
rect 3297 6040 3343 6080
rect 3501 6126 3567 6166
rect 3501 6080 3521 6126
rect 3390 5989 3455 6032
rect 3390 5906 3405 5989
rect 3390 5849 3405 5854
rect 3451 5849 3455 5989
rect 3390 5832 3455 5849
rect 2829 5682 2849 5747
rect 2829 5630 2830 5682
rect 2829 5607 2849 5630
rect 2829 5594 2895 5607
rect 3317 5747 3363 5766
rect 3317 5548 3363 5607
rect 3501 5747 3567 6080
rect 3969 6126 4015 6212
rect 3969 6040 4015 6080
rect 4173 6126 4239 6166
rect 4173 6080 4193 6126
rect 4062 5989 4127 6032
rect 4062 5906 4077 5989
rect 4062 5849 4077 5854
rect 4123 5849 4127 5989
rect 4062 5832 4127 5849
rect 3501 5682 3521 5747
rect 3501 5630 3502 5682
rect 3501 5607 3521 5630
rect 3501 5594 3567 5607
rect 3989 5747 4035 5766
rect 3989 5548 4035 5607
rect 4173 5747 4239 6080
rect 4641 6126 4687 6212
rect 4641 6040 4687 6080
rect 4845 6126 4911 6166
rect 4845 6080 4865 6126
rect 4734 5989 4799 6032
rect 4734 5906 4749 5989
rect 4734 5849 4749 5854
rect 4795 5849 4799 5989
rect 4734 5832 4799 5849
rect 4173 5682 4193 5747
rect 4173 5630 4174 5682
rect 4173 5607 4193 5630
rect 4173 5594 4239 5607
rect 4661 5747 4707 5766
rect 4661 5548 4707 5607
rect 4845 5747 4911 6080
rect 5313 6126 5359 6212
rect 5313 6040 5359 6080
rect 5517 6130 5583 6166
rect 5517 6078 5518 6130
rect 5570 6126 5583 6130
rect 5570 6078 5583 6080
rect 5406 5989 5471 6032
rect 5406 5906 5421 5989
rect 5406 5849 5421 5854
rect 5467 5849 5471 5989
rect 5406 5832 5471 5849
rect 4845 5682 4865 5747
rect 4845 5630 4846 5682
rect 4845 5607 4865 5630
rect 4845 5594 4911 5607
rect 5333 5747 5379 5766
rect 5333 5548 5379 5607
rect 5517 5747 5583 6078
rect 5985 6126 6031 6212
rect 5985 6040 6031 6080
rect 6189 6130 6255 6166
rect 6189 6078 6190 6130
rect 6242 6126 6255 6130
rect 6242 6078 6255 6080
rect 6078 5989 6143 6032
rect 6078 5906 6093 5989
rect 6078 5849 6093 5854
rect 6139 5849 6143 5989
rect 6078 5832 6143 5849
rect 5517 5607 5537 5747
rect 5517 5594 5583 5607
rect 6005 5747 6051 5766
rect 6005 5548 6051 5607
rect 6189 5747 6255 6078
rect 6657 6126 6703 6212
rect 6657 6040 6703 6080
rect 6861 6126 6927 6166
rect 6861 6080 6881 6126
rect 6750 6018 6815 6032
rect 6802 5989 6815 6018
rect 6750 5849 6765 5966
rect 6811 5849 6815 5989
rect 6750 5832 6815 5849
rect 6861 6018 6927 6080
rect 7329 6126 7375 6212
rect 7329 6040 7375 6080
rect 7533 6126 7599 6166
rect 7533 6080 7553 6126
rect 6861 5966 6862 6018
rect 6914 5966 6927 6018
rect 6189 5607 6209 5747
rect 6189 5594 6255 5607
rect 6677 5747 6723 5766
rect 6677 5548 6723 5607
rect 6861 5747 6927 5966
rect 7422 6018 7487 6032
rect 7474 5989 7487 6018
rect 7422 5849 7437 5966
rect 7483 5849 7487 5989
rect 7422 5832 7487 5849
rect 6861 5607 6881 5747
rect 6861 5594 6927 5607
rect 7349 5747 7395 5766
rect 7349 5548 7395 5607
rect 7533 5747 7599 6080
rect 8001 6126 8047 6212
rect 8001 6040 8047 6080
rect 8205 6126 8271 6166
rect 8205 6080 8225 6126
rect 8094 6018 8159 6032
rect 8146 5989 8159 6018
rect 8094 5849 8109 5966
rect 8155 5849 8159 5989
rect 8094 5832 8159 5849
rect 7533 5682 7553 5747
rect 7533 5630 7534 5682
rect 7533 5607 7553 5630
rect 7533 5594 7599 5607
rect 8021 5747 8067 5766
rect 8021 5548 8067 5607
rect 8205 5747 8271 6080
rect 8673 6126 8719 6212
rect 9374 6193 9442 6212
rect 8673 6040 8719 6080
rect 8877 6130 8943 6166
rect 8877 6078 8878 6130
rect 8930 6126 8943 6130
rect 8930 6078 8943 6080
rect 8766 6018 8831 6032
rect 8818 5989 8831 6018
rect 8766 5849 8781 5966
rect 8827 5849 8831 5989
rect 8766 5832 8831 5849
rect 8205 5682 8225 5747
rect 8205 5630 8206 5682
rect 8205 5607 8225 5630
rect 8205 5594 8271 5607
rect 8693 5747 8739 5766
rect 8693 5548 8739 5607
rect 8877 5747 8943 6078
rect 9374 6046 9385 6193
rect 9431 6046 9442 6193
rect 9374 6035 9442 6046
rect 9681 6126 9727 6212
rect 9681 6040 9727 6080
rect 9885 6130 9951 6166
rect 9885 6078 9886 6130
rect 9938 6126 9951 6130
rect 9938 6078 9951 6080
rect 9774 5989 9839 6032
rect 9774 5906 9789 5989
rect 8877 5607 8897 5747
rect 8877 5594 8943 5607
rect 9374 5875 9442 5886
rect 9374 5829 9385 5875
rect 9431 5829 9442 5875
rect 9774 5849 9789 5854
rect 9835 5849 9839 5989
rect 9774 5832 9839 5849
rect 9374 5747 9442 5829
rect 9374 5701 9385 5747
rect 9431 5701 9442 5747
rect 9374 5619 9442 5701
rect 9374 5573 9385 5619
rect 9431 5573 9442 5619
rect 9374 5548 9442 5573
rect 9701 5747 9747 5766
rect 9701 5548 9747 5607
rect 9885 5747 9951 6078
rect 10353 6126 10399 6212
rect 10353 6040 10399 6080
rect 10557 6130 10623 6166
rect 10557 6078 10558 6130
rect 10610 6126 10623 6130
rect 10610 6078 10623 6080
rect 10446 5989 10511 6032
rect 10446 5906 10461 5989
rect 10446 5849 10461 5854
rect 10507 5849 10511 5989
rect 10446 5832 10511 5849
rect 9885 5607 9905 5747
rect 9885 5594 9951 5607
rect 10373 5747 10419 5766
rect 10373 5548 10419 5607
rect 10557 5747 10623 6078
rect 11025 6126 11071 6212
rect 11025 6040 11071 6080
rect 11229 6130 11295 6166
rect 11229 6078 11230 6130
rect 11282 6126 11295 6130
rect 11282 6078 11295 6080
rect 11118 6018 11183 6032
rect 11170 5989 11183 6018
rect 11118 5849 11133 5966
rect 11179 5849 11183 5989
rect 11118 5832 11183 5849
rect 10557 5607 10577 5747
rect 10557 5594 10623 5607
rect 11045 5747 11091 5766
rect 11045 5548 11091 5607
rect 11229 5747 11295 6078
rect 11697 6126 11743 6212
rect 11697 6040 11743 6080
rect 11901 6130 11967 6166
rect 11901 6078 11902 6130
rect 11954 6126 11967 6130
rect 11954 6078 11967 6080
rect 11790 6018 11855 6032
rect 11842 5989 11855 6018
rect 11790 5849 11805 5966
rect 11851 5849 11855 5989
rect 11790 5832 11855 5849
rect 11229 5607 11249 5747
rect 11229 5594 11295 5607
rect 11717 5747 11763 5766
rect 11717 5548 11763 5607
rect 11901 5747 11967 6078
rect 12481 6126 12527 6212
rect 12481 6040 12527 6080
rect 12685 6126 12751 6166
rect 12685 6080 12705 6126
rect 12574 6018 12639 6032
rect 12626 5989 12639 6018
rect 12574 5849 12589 5966
rect 12635 5849 12639 5989
rect 12574 5832 12639 5849
rect 11901 5607 11921 5747
rect 11901 5594 11967 5607
rect 12501 5747 12547 5766
rect 12501 5548 12547 5607
rect 12685 5747 12751 6080
rect 13153 6126 13199 6212
rect 13153 6040 13199 6080
rect 13357 6130 13423 6166
rect 13357 6078 13358 6130
rect 13410 6126 13423 6130
rect 13410 6078 13423 6080
rect 13246 5989 13311 6032
rect 13246 5906 13261 5989
rect 13246 5849 13261 5854
rect 13307 5849 13311 5989
rect 13246 5832 13311 5849
rect 12685 5682 12705 5747
rect 12685 5630 12686 5682
rect 12685 5607 12705 5630
rect 12685 5594 12751 5607
rect 13173 5747 13219 5766
rect 13173 5548 13219 5607
rect 13357 5747 13423 6078
rect 13825 6126 13871 6212
rect 13825 6040 13871 6080
rect 14029 6130 14095 6166
rect 14029 6078 14030 6130
rect 14082 6126 14095 6130
rect 14082 6078 14095 6080
rect 13918 5989 13983 6032
rect 13918 5906 13933 5989
rect 13918 5849 13933 5854
rect 13979 5849 13983 5989
rect 13918 5832 13983 5849
rect 13357 5607 13377 5747
rect 13357 5594 13423 5607
rect 13845 5747 13891 5766
rect 13845 5548 13891 5607
rect 14029 5747 14095 6078
rect 14497 6126 14543 6212
rect 14497 6040 14543 6080
rect 14701 6130 14767 6166
rect 14701 6078 14702 6130
rect 14754 6126 14767 6130
rect 14754 6078 14767 6080
rect 14590 6018 14655 6032
rect 14642 5989 14655 6018
rect 14590 5849 14605 5966
rect 14651 5849 14655 5989
rect 14590 5832 14655 5849
rect 14029 5607 14049 5747
rect 14029 5594 14095 5607
rect 14517 5747 14563 5766
rect 14517 5548 14563 5607
rect 14701 5747 14767 6078
rect 15169 6126 15215 6212
rect 15169 6040 15215 6080
rect 15373 6130 15439 6166
rect 15373 6078 15374 6130
rect 15426 6126 15439 6130
rect 15426 6078 15439 6080
rect 15262 6018 15327 6032
rect 15314 5989 15327 6018
rect 15262 5849 15277 5966
rect 15323 5849 15327 5989
rect 15262 5832 15327 5849
rect 14701 5607 14721 5747
rect 14701 5594 14767 5607
rect 15189 5747 15235 5766
rect 15189 5548 15235 5607
rect 15373 5747 15439 6078
rect 15841 6126 15887 6212
rect 15841 6040 15887 6080
rect 16045 6130 16111 6166
rect 16045 6078 16046 6130
rect 16098 6126 16111 6130
rect 16098 6078 16111 6080
rect 15934 6018 15999 6032
rect 15986 5989 15999 6018
rect 15934 5849 15949 5966
rect 15995 5849 15999 5989
rect 15934 5832 15999 5849
rect 15373 5607 15393 5747
rect 15373 5594 15439 5607
rect 15861 5747 15907 5766
rect 15861 5548 15907 5607
rect 16045 5747 16111 6078
rect 16513 6126 16559 6212
rect 17326 6193 17394 6212
rect 16513 6040 16559 6080
rect 16717 6130 16783 6166
rect 16717 6078 16718 6130
rect 16770 6126 16783 6130
rect 16770 6078 16783 6080
rect 16606 6018 16671 6032
rect 16658 5989 16671 6018
rect 16606 5849 16621 5966
rect 16667 5849 16671 5989
rect 16606 5832 16671 5849
rect 16045 5607 16065 5747
rect 16045 5594 16111 5607
rect 16533 5747 16579 5766
rect 16533 5548 16579 5607
rect 16717 5747 16783 6078
rect 17326 6046 17337 6193
rect 17383 6046 17394 6193
rect 17326 6035 17394 6046
rect 17633 6126 17679 6212
rect 17633 6040 17679 6080
rect 17837 6126 17903 6166
rect 17837 6080 17857 6126
rect 17726 5989 17791 6032
rect 17726 5906 17741 5989
rect 16717 5607 16737 5747
rect 16717 5594 16783 5607
rect 17326 5875 17394 5886
rect 17326 5829 17337 5875
rect 17383 5829 17394 5875
rect 17726 5849 17741 5854
rect 17787 5849 17791 5989
rect 17726 5832 17791 5849
rect 17326 5747 17394 5829
rect 17326 5701 17337 5747
rect 17383 5701 17394 5747
rect 17326 5619 17394 5701
rect 17326 5573 17337 5619
rect 17383 5573 17394 5619
rect 17326 5548 17394 5573
rect 17653 5747 17699 5766
rect 17653 5548 17699 5607
rect 17837 5747 17903 6080
rect 18305 6126 18351 6212
rect 18305 6040 18351 6080
rect 18509 6126 18575 6166
rect 18509 6080 18529 6126
rect 18398 5989 18463 6032
rect 18398 5906 18413 5989
rect 18398 5849 18413 5854
rect 18459 5849 18463 5989
rect 18398 5832 18463 5849
rect 18509 5794 18575 6080
rect 18977 6126 19023 6212
rect 18977 6040 19023 6080
rect 19181 6126 19247 6166
rect 19181 6080 19201 6126
rect 19070 6018 19135 6032
rect 19122 5989 19135 6018
rect 19070 5849 19085 5966
rect 19131 5849 19135 5989
rect 19070 5832 19135 5849
rect 17837 5682 17857 5747
rect 17837 5630 17838 5682
rect 17837 5607 17857 5630
rect 17837 5594 17903 5607
rect 18325 5747 18371 5766
rect 18325 5548 18371 5607
rect 18509 5742 18510 5794
rect 18562 5747 18575 5794
rect 19181 5794 19247 6080
rect 19649 6126 19695 6212
rect 19649 6040 19695 6080
rect 19853 6126 19919 6166
rect 19853 6080 19873 6126
rect 19742 6018 19807 6032
rect 19794 5989 19807 6018
rect 19742 5849 19757 5966
rect 19803 5849 19807 5989
rect 19742 5832 19807 5849
rect 18509 5607 18529 5742
rect 18509 5594 18575 5607
rect 18997 5747 19043 5766
rect 18997 5548 19043 5607
rect 19181 5742 19182 5794
rect 19234 5747 19247 5794
rect 19181 5607 19201 5742
rect 19181 5594 19247 5607
rect 19669 5747 19715 5766
rect 19669 5548 19715 5607
rect 19853 5747 19919 6080
rect 20321 6126 20367 6212
rect 20321 6040 20367 6080
rect 20525 6126 20591 6166
rect 20525 6080 20545 6126
rect 20414 5989 20479 6032
rect 20414 5906 20429 5989
rect 20414 5849 20429 5854
rect 20475 5849 20479 5989
rect 20414 5832 20479 5849
rect 19853 5682 19873 5747
rect 19853 5630 19854 5682
rect 19853 5607 19873 5630
rect 19853 5594 19919 5607
rect 20341 5747 20387 5766
rect 20341 5548 20387 5607
rect 20525 5747 20591 6080
rect 20993 6126 21039 6212
rect 20993 6040 21039 6080
rect 21197 6126 21263 6166
rect 21197 6080 21217 6126
rect 21086 5989 21151 6032
rect 21086 5906 21101 5989
rect 21086 5849 21101 5854
rect 21147 5849 21151 5989
rect 21086 5832 21151 5849
rect 20525 5682 20545 5747
rect 20525 5630 20526 5682
rect 20525 5607 20545 5630
rect 20525 5594 20591 5607
rect 21013 5747 21059 5766
rect 21013 5548 21059 5607
rect 21197 5747 21263 6080
rect 21197 5682 21217 5747
rect 21197 5630 21198 5682
rect 21197 5607 21217 5630
rect 21197 5594 21263 5607
rect 21745 6126 21811 6166
rect 21791 6080 21811 6126
rect 21745 5747 21811 6080
rect 21969 6126 22015 6212
rect 21969 6040 22015 6080
rect 22482 6193 22550 6212
rect 22482 6046 22493 6193
rect 22539 6046 22550 6193
rect 22482 6034 22550 6046
rect 21857 5989 21922 6032
rect 21857 5849 21861 5989
rect 21907 5906 21922 5989
rect 21907 5849 21922 5854
rect 21857 5832 21922 5849
rect 22482 5875 22550 5888
rect 22482 5829 22493 5875
rect 22539 5829 22550 5875
rect 21791 5682 21811 5747
rect 21810 5630 21811 5682
rect 21791 5607 21811 5630
rect 21745 5594 21811 5607
rect 21949 5747 21995 5766
rect 21949 5548 21995 5607
rect 22482 5747 22550 5829
rect 22482 5701 22493 5747
rect 22539 5701 22550 5747
rect 22482 5619 22550 5701
rect 22482 5573 22493 5619
rect 22539 5573 22550 5619
rect 22482 5548 22550 5573
rect 1344 5514 22624 5548
rect 1344 5462 3874 5514
rect 4134 5462 9194 5514
rect 9454 5462 14514 5514
rect 14774 5462 19834 5514
rect 20094 5462 22624 5514
rect 1344 5428 22624 5462
rect 1418 5403 1486 5428
rect 1418 5357 1429 5403
rect 1475 5357 1486 5403
rect 1418 5275 1486 5357
rect 1418 5229 1429 5275
rect 1475 5229 1486 5275
rect 1418 5147 1486 5229
rect 1418 5101 1429 5147
rect 1475 5101 1486 5147
rect 1418 5088 1486 5101
rect 1617 5361 1663 5382
rect 1617 5015 1663 5221
rect 1921 5361 1967 5428
rect 1921 5202 1967 5221
rect 2085 5369 2131 5428
rect 2085 5210 2131 5229
rect 2269 5369 2335 5382
rect 2269 5229 2289 5369
rect 1714 5096 1728 5142
rect 1868 5096 1967 5142
rect 1617 4969 1720 5015
rect 1860 4969 1872 5015
rect 1418 4930 1486 4942
rect 1418 4783 1429 4930
rect 1475 4783 1486 4930
rect 1418 4764 1486 4783
rect 1617 4896 1663 4923
rect 1617 4764 1663 4850
rect 1921 4896 1967 5096
rect 2158 5127 2223 5144
rect 2158 5010 2173 5127
rect 2219 4987 2223 5127
rect 2210 4958 2223 4987
rect 2158 4944 2223 4958
rect 1921 4810 1967 4850
rect 2065 4896 2111 4936
rect 2065 4764 2111 4850
rect 2269 4898 2335 5229
rect 2757 5369 2803 5428
rect 2757 5210 2803 5229
rect 2941 5369 3007 5382
rect 2941 5229 2961 5369
rect 2830 5127 2895 5144
rect 2830 5010 2845 5127
rect 2891 4987 2895 5127
rect 2882 4958 2895 4987
rect 2830 4944 2895 4958
rect 2269 4846 2270 4898
rect 2322 4896 2335 4898
rect 2322 4846 2335 4850
rect 2269 4810 2335 4846
rect 2737 4896 2783 4936
rect 2737 4764 2783 4850
rect 2941 4898 3007 5229
rect 3429 5369 3475 5428
rect 3429 5210 3475 5229
rect 3613 5369 3679 5382
rect 3613 5229 3633 5369
rect 3502 5127 3567 5144
rect 3502 5010 3517 5127
rect 3563 4987 3567 5127
rect 3554 4958 3567 4987
rect 3502 4944 3567 4958
rect 3613 5010 3679 5229
rect 4101 5369 4147 5428
rect 4101 5210 4147 5229
rect 4285 5369 4351 5382
rect 4285 5229 4305 5369
rect 3613 4958 3614 5010
rect 3666 4958 3679 5010
rect 2941 4846 2942 4898
rect 2994 4896 3007 4898
rect 2994 4846 3007 4850
rect 2941 4810 3007 4846
rect 3409 4896 3455 4936
rect 3409 4764 3455 4850
rect 3613 4896 3679 4958
rect 4174 5127 4239 5144
rect 4174 5122 4189 5127
rect 4174 4987 4189 5070
rect 4235 4987 4239 5127
rect 4174 4944 4239 4987
rect 3613 4850 3633 4896
rect 3613 4810 3679 4850
rect 4081 4896 4127 4936
rect 4081 4764 4127 4850
rect 4285 4898 4351 5229
rect 4773 5369 4819 5428
rect 5342 5403 5410 5428
rect 4773 5210 4819 5229
rect 4957 5369 5023 5382
rect 4957 5229 4977 5369
rect 4846 5127 4911 5144
rect 4846 5122 4861 5127
rect 4846 4987 4861 5070
rect 4907 4987 4911 5127
rect 4846 4944 4911 4987
rect 4285 4846 4286 4898
rect 4338 4896 4351 4898
rect 4338 4846 4351 4850
rect 4285 4810 4351 4846
rect 4753 4896 4799 4936
rect 4753 4764 4799 4850
rect 4957 4898 5023 5229
rect 5342 5357 5353 5403
rect 5399 5357 5410 5403
rect 5342 5275 5410 5357
rect 5342 5229 5353 5275
rect 5399 5229 5410 5275
rect 5342 5147 5410 5229
rect 5669 5369 5715 5428
rect 5669 5210 5715 5229
rect 5853 5369 5919 5382
rect 5853 5346 5873 5369
rect 5853 5294 5854 5346
rect 5853 5229 5873 5294
rect 5342 5101 5353 5147
rect 5399 5101 5410 5147
rect 5342 5090 5410 5101
rect 5742 5127 5807 5144
rect 5742 5010 5757 5127
rect 5803 4987 5807 5127
rect 5794 4958 5807 4987
rect 5742 4944 5807 4958
rect 4957 4846 4958 4898
rect 5010 4896 5023 4898
rect 5010 4846 5023 4850
rect 4957 4810 5023 4846
rect 5342 4930 5410 4941
rect 5342 4783 5353 4930
rect 5399 4783 5410 4930
rect 5342 4764 5410 4783
rect 5649 4896 5695 4936
rect 5649 4764 5695 4850
rect 5853 4896 5919 5229
rect 6341 5369 6387 5428
rect 6341 5210 6387 5229
rect 6525 5369 6591 5382
rect 6525 5346 6545 5369
rect 6525 5294 6526 5346
rect 6525 5229 6545 5294
rect 6414 5127 6479 5144
rect 6414 5010 6429 5127
rect 6475 4987 6479 5127
rect 6466 4958 6479 4987
rect 6414 4944 6479 4958
rect 5853 4850 5873 4896
rect 5853 4810 5919 4850
rect 6321 4896 6367 4936
rect 6321 4764 6367 4850
rect 6525 4896 6591 5229
rect 7013 5369 7059 5428
rect 7013 5210 7059 5229
rect 7197 5369 7263 5382
rect 7197 5346 7217 5369
rect 7197 5294 7198 5346
rect 7197 5229 7217 5294
rect 7086 5127 7151 5144
rect 7086 5122 7101 5127
rect 7086 4987 7101 5070
rect 7147 4987 7151 5127
rect 7086 4944 7151 4987
rect 6525 4850 6545 4896
rect 6525 4810 6591 4850
rect 6993 4896 7039 4936
rect 6993 4764 7039 4850
rect 7197 4896 7263 5229
rect 7685 5369 7731 5428
rect 7685 5210 7731 5229
rect 7869 5369 7935 5382
rect 7869 5229 7889 5369
rect 7758 5127 7823 5144
rect 7758 5122 7773 5127
rect 7758 4987 7773 5070
rect 7819 4987 7823 5127
rect 7758 4944 7823 4987
rect 7869 5122 7935 5229
rect 8357 5369 8403 5428
rect 8357 5210 8403 5229
rect 8541 5369 8607 5382
rect 8541 5346 8561 5369
rect 8541 5294 8542 5346
rect 8541 5229 8561 5294
rect 7869 5070 7870 5122
rect 7922 5070 7935 5122
rect 7197 4850 7217 4896
rect 7197 4810 7263 4850
rect 7665 4896 7711 4936
rect 7665 4764 7711 4850
rect 7869 4896 7935 5070
rect 8430 5127 8495 5144
rect 8430 5122 8445 5127
rect 8430 4987 8445 5070
rect 8491 4987 8495 5127
rect 8430 4944 8495 4987
rect 7869 4850 7889 4896
rect 7869 4810 7935 4850
rect 8337 4896 8383 4936
rect 8337 4764 8383 4850
rect 8541 4896 8607 5229
rect 9029 5369 9075 5428
rect 9029 5210 9075 5229
rect 9213 5369 9279 5382
rect 9213 5229 9233 5369
rect 9102 5127 9167 5144
rect 9102 5122 9117 5127
rect 9102 4987 9117 5070
rect 9163 4987 9167 5127
rect 9102 4944 9167 4987
rect 9213 5122 9279 5229
rect 9701 5369 9747 5428
rect 9701 5210 9747 5229
rect 9885 5369 9951 5382
rect 9885 5346 9905 5369
rect 9885 5294 9886 5346
rect 9885 5229 9905 5294
rect 9213 5070 9214 5122
rect 9266 5070 9279 5122
rect 8541 4850 8561 4896
rect 8541 4810 8607 4850
rect 9009 4896 9055 4936
rect 9009 4764 9055 4850
rect 9213 4896 9279 5070
rect 9774 5127 9839 5144
rect 9774 5010 9789 5127
rect 9835 4987 9839 5127
rect 9826 4958 9839 4987
rect 9774 4944 9839 4958
rect 9213 4850 9233 4896
rect 9213 4810 9279 4850
rect 9681 4896 9727 4936
rect 9681 4764 9727 4850
rect 9885 4896 9951 5229
rect 10373 5369 10419 5428
rect 10373 5210 10419 5229
rect 10557 5369 10623 5382
rect 10557 5346 10577 5369
rect 10557 5294 10558 5346
rect 10557 5229 10577 5294
rect 10446 5127 10511 5144
rect 10446 5122 10461 5127
rect 10446 4987 10461 5070
rect 10507 4987 10511 5127
rect 10446 4944 10511 4987
rect 9885 4850 9905 4896
rect 9885 4810 9951 4850
rect 10353 4896 10399 4936
rect 10353 4764 10399 4850
rect 10557 4896 10623 5229
rect 10801 5361 10847 5382
rect 10801 5015 10847 5221
rect 11105 5361 11151 5428
rect 11105 5202 11151 5221
rect 11381 5369 11427 5428
rect 11381 5210 11427 5229
rect 11565 5369 11631 5382
rect 11565 5229 11585 5369
rect 10898 5096 10912 5142
rect 11052 5096 11151 5142
rect 10801 4969 10904 5015
rect 11044 4969 11056 5015
rect 10557 4850 10577 4896
rect 10557 4810 10623 4850
rect 10801 4896 10847 4923
rect 10801 4764 10847 4850
rect 11105 4896 11151 5096
rect 11454 5127 11519 5144
rect 11454 5122 11469 5127
rect 11454 4987 11469 5070
rect 11515 4987 11519 5127
rect 11454 4944 11519 4987
rect 11565 5122 11631 5229
rect 12053 5369 12099 5428
rect 12053 5210 12099 5229
rect 12237 5369 12303 5382
rect 12237 5229 12257 5369
rect 11565 5070 11566 5122
rect 11618 5070 11631 5122
rect 11105 4810 11151 4850
rect 11361 4896 11407 4936
rect 11361 4764 11407 4850
rect 11565 4896 11631 5070
rect 12126 5127 12191 5144
rect 12126 5010 12141 5127
rect 12187 4987 12191 5127
rect 12178 4958 12191 4987
rect 12126 4944 12191 4958
rect 11565 4850 11585 4896
rect 11565 4810 11631 4850
rect 12033 4896 12079 4936
rect 12033 4764 12079 4850
rect 12237 4898 12303 5229
rect 12725 5369 12771 5428
rect 13294 5403 13362 5428
rect 12725 5210 12771 5229
rect 12909 5369 12975 5382
rect 12909 5229 12929 5369
rect 12798 5127 12863 5144
rect 12798 5010 12813 5127
rect 12859 4987 12863 5127
rect 12850 4958 12863 4987
rect 12798 4944 12863 4958
rect 12237 4846 12238 4898
rect 12290 4896 12303 4898
rect 12290 4846 12303 4850
rect 12237 4810 12303 4846
rect 12705 4896 12751 4936
rect 12705 4764 12751 4850
rect 12909 4898 12975 5229
rect 13294 5357 13305 5403
rect 13351 5357 13362 5403
rect 13294 5275 13362 5357
rect 13294 5229 13305 5275
rect 13351 5229 13362 5275
rect 13294 5147 13362 5229
rect 13294 5101 13305 5147
rect 13351 5101 13362 5147
rect 13294 5090 13362 5101
rect 13489 5361 13535 5382
rect 13489 5015 13535 5221
rect 13793 5361 13839 5428
rect 13793 5202 13839 5221
rect 13957 5369 14003 5428
rect 13957 5210 14003 5229
rect 14141 5369 14207 5382
rect 14141 5346 14161 5369
rect 14141 5294 14142 5346
rect 14141 5229 14161 5294
rect 13586 5096 13600 5142
rect 13740 5096 13839 5142
rect 13489 4969 13592 5015
rect 13732 4969 13744 5015
rect 12909 4846 12910 4898
rect 12962 4896 12975 4898
rect 12962 4846 12975 4850
rect 12909 4810 12975 4846
rect 13294 4930 13362 4941
rect 13294 4783 13305 4930
rect 13351 4783 13362 4930
rect 13294 4764 13362 4783
rect 13489 4896 13535 4923
rect 13489 4764 13535 4850
rect 13793 4896 13839 5096
rect 14030 5127 14095 5144
rect 14030 5010 14045 5127
rect 14091 4987 14095 5127
rect 14082 4958 14095 4987
rect 14030 4944 14095 4958
rect 13793 4810 13839 4850
rect 13937 4896 13983 4936
rect 13937 4764 13983 4850
rect 14141 4896 14207 5229
rect 14629 5369 14675 5428
rect 14629 5210 14675 5229
rect 14813 5369 14879 5382
rect 14813 5346 14833 5369
rect 14813 5294 14814 5346
rect 14813 5229 14833 5294
rect 14702 5127 14767 5144
rect 14702 5010 14717 5127
rect 14763 4987 14767 5127
rect 14754 4958 14767 4987
rect 14702 4944 14767 4958
rect 14141 4850 14161 4896
rect 14141 4810 14207 4850
rect 14609 4896 14655 4936
rect 14609 4764 14655 4850
rect 14813 4896 14879 5229
rect 15301 5369 15347 5428
rect 15301 5210 15347 5229
rect 15485 5369 15551 5382
rect 15485 5346 15505 5369
rect 15485 5294 15486 5346
rect 15485 5229 15505 5294
rect 15374 5127 15439 5144
rect 15374 5122 15389 5127
rect 15374 4987 15389 5070
rect 15435 4987 15439 5127
rect 15374 4944 15439 4987
rect 14813 4850 14833 4896
rect 14813 4810 14879 4850
rect 15281 4896 15327 4936
rect 15281 4764 15327 4850
rect 15485 4896 15551 5229
rect 15973 5369 16019 5428
rect 15973 5210 16019 5229
rect 16157 5369 16223 5382
rect 16157 5229 16177 5369
rect 16046 5127 16111 5144
rect 16046 5010 16061 5127
rect 16107 4987 16111 5127
rect 16098 4958 16111 4987
rect 16046 4944 16111 4958
rect 15485 4850 15505 4896
rect 15485 4810 15551 4850
rect 15953 4896 15999 4936
rect 15953 4764 15999 4850
rect 16157 4898 16223 5229
rect 16645 5369 16691 5428
rect 16645 5210 16691 5229
rect 16829 5369 16895 5382
rect 16829 5229 16849 5369
rect 16718 5127 16783 5144
rect 16718 5010 16733 5127
rect 16779 4987 16783 5127
rect 16770 4958 16783 4987
rect 16718 4944 16783 4958
rect 16829 5122 16895 5229
rect 17317 5369 17363 5428
rect 17317 5210 17363 5229
rect 17501 5369 17567 5382
rect 17501 5229 17521 5369
rect 16829 5070 16830 5122
rect 16882 5070 16895 5122
rect 16157 4846 16158 4898
rect 16210 4896 16223 4898
rect 16210 4846 16223 4850
rect 16157 4810 16223 4846
rect 16625 4896 16671 4936
rect 16625 4764 16671 4850
rect 16829 4896 16895 5070
rect 17390 5127 17455 5144
rect 17390 5122 17405 5127
rect 17390 4987 17405 5070
rect 17451 4987 17455 5127
rect 17390 4944 17455 4987
rect 16829 4850 16849 4896
rect 16829 4810 16895 4850
rect 17297 4896 17343 4936
rect 17297 4764 17343 4850
rect 17501 4898 17567 5229
rect 17989 5369 18035 5428
rect 17989 5210 18035 5229
rect 18173 5369 18239 5382
rect 18173 5346 18193 5369
rect 18173 5294 18174 5346
rect 18173 5229 18193 5294
rect 18062 5127 18127 5144
rect 18062 5122 18077 5127
rect 18062 4987 18077 5070
rect 18123 4987 18127 5127
rect 18062 4944 18127 4987
rect 17501 4846 17502 4898
rect 17554 4896 17567 4898
rect 17554 4846 17567 4850
rect 17501 4810 17567 4846
rect 17969 4896 18015 4936
rect 17969 4764 18015 4850
rect 18173 4896 18239 5229
rect 18661 5369 18707 5428
rect 18661 5210 18707 5229
rect 18845 5369 18911 5382
rect 18845 5229 18865 5369
rect 18734 5127 18799 5144
rect 18734 5122 18749 5127
rect 18734 4987 18749 5070
rect 18795 4987 18799 5127
rect 18734 4944 18799 4987
rect 18845 5122 18911 5229
rect 19333 5369 19379 5428
rect 19333 5210 19379 5229
rect 19517 5369 19583 5382
rect 19517 5234 19537 5369
rect 19517 5182 19518 5234
rect 19570 5182 19583 5229
rect 20005 5369 20051 5428
rect 20005 5210 20051 5229
rect 20189 5369 20255 5382
rect 20189 5346 20209 5369
rect 20189 5294 20190 5346
rect 20189 5229 20209 5294
rect 18845 5070 18846 5122
rect 18898 5070 18911 5122
rect 18173 4850 18193 4896
rect 18173 4810 18239 4850
rect 18641 4896 18687 4936
rect 18641 4764 18687 4850
rect 18845 4896 18911 5070
rect 19406 5127 19471 5144
rect 19406 5122 19421 5127
rect 19406 4987 19421 5070
rect 19467 4987 19471 5127
rect 19406 4944 19471 4987
rect 18845 4850 18865 4896
rect 18845 4810 18911 4850
rect 19313 4896 19359 4936
rect 19313 4764 19359 4850
rect 19517 4896 19583 5182
rect 20078 5127 20143 5144
rect 20078 5122 20093 5127
rect 20078 4987 20093 5070
rect 20139 4987 20143 5127
rect 20078 4944 20143 4987
rect 19517 4850 19537 4896
rect 19517 4810 19583 4850
rect 19985 4896 20031 4936
rect 19985 4764 20031 4850
rect 20189 4896 20255 5229
rect 20677 5369 20723 5428
rect 21246 5403 21314 5428
rect 20677 5210 20723 5229
rect 20861 5369 20927 5382
rect 20861 5229 20881 5369
rect 20750 5127 20815 5144
rect 20750 5010 20765 5127
rect 20811 4987 20815 5127
rect 20802 4958 20815 4987
rect 20750 4944 20815 4958
rect 20189 4850 20209 4896
rect 20189 4810 20255 4850
rect 20657 4896 20703 4936
rect 20657 4764 20703 4850
rect 20861 4898 20927 5229
rect 21246 5357 21257 5403
rect 21303 5357 21314 5403
rect 21246 5275 21314 5357
rect 21246 5229 21257 5275
rect 21303 5229 21314 5275
rect 21246 5147 21314 5229
rect 21573 5369 21619 5428
rect 21573 5210 21619 5229
rect 21757 5369 21823 5382
rect 21757 5229 21777 5369
rect 21246 5101 21257 5147
rect 21303 5101 21314 5147
rect 21246 5090 21314 5101
rect 21646 5127 21711 5144
rect 21646 5010 21661 5127
rect 21707 4987 21711 5127
rect 21698 4958 21711 4987
rect 21646 4944 21711 4958
rect 20861 4846 20862 4898
rect 20914 4896 20927 4898
rect 20914 4846 20927 4850
rect 20861 4810 20927 4846
rect 21246 4930 21314 4941
rect 21246 4783 21257 4930
rect 21303 4783 21314 4930
rect 21246 4764 21314 4783
rect 21553 4896 21599 4936
rect 21553 4764 21599 4850
rect 21757 4898 21823 5229
rect 22001 5361 22047 5382
rect 22001 5015 22047 5221
rect 22305 5361 22351 5428
rect 22305 5202 22351 5221
rect 22482 5403 22550 5428
rect 22482 5357 22493 5403
rect 22539 5357 22550 5403
rect 22482 5275 22550 5357
rect 22482 5229 22493 5275
rect 22539 5229 22550 5275
rect 22482 5147 22550 5229
rect 22098 5096 22112 5142
rect 22252 5096 22351 5142
rect 22001 4969 22104 5015
rect 22244 4969 22256 5015
rect 21757 4846 21758 4898
rect 21810 4896 21823 4898
rect 21810 4846 21823 4850
rect 21757 4810 21823 4846
rect 22001 4896 22047 4923
rect 22001 4764 22047 4850
rect 22305 4896 22351 5096
rect 22482 5101 22493 5147
rect 22539 5101 22550 5147
rect 22482 5088 22550 5101
rect 22305 4810 22351 4850
rect 22482 4930 22550 4942
rect 22482 4783 22493 4930
rect 22539 4783 22550 4930
rect 22482 4764 22550 4783
rect 1344 4730 22784 4764
rect 1344 4678 6534 4730
rect 6794 4678 11854 4730
rect 12114 4678 17174 4730
rect 17434 4678 22494 4730
rect 22754 4678 22784 4730
rect 1344 4644 22784 4678
rect 1418 4625 1486 4644
rect 1418 4478 1429 4625
rect 1475 4478 1486 4625
rect 1617 4558 1663 4644
rect 1617 4485 1663 4512
rect 1921 4558 1967 4598
rect 1418 4466 1486 4478
rect 1617 4393 1720 4439
rect 1860 4393 1872 4439
rect 1418 4307 1486 4320
rect 1418 4261 1429 4307
rect 1475 4261 1486 4307
rect 1418 4179 1486 4261
rect 1418 4133 1429 4179
rect 1475 4133 1486 4179
rect 1418 4051 1486 4133
rect 1418 4005 1429 4051
rect 1475 4005 1486 4051
rect 1617 4187 1663 4393
rect 1921 4312 1967 4512
rect 2289 4558 2335 4644
rect 2289 4472 2335 4512
rect 2493 4558 2559 4598
rect 2493 4512 2513 4558
rect 1714 4266 1728 4312
rect 1868 4266 1967 4312
rect 2382 4450 2447 4464
rect 2434 4421 2447 4450
rect 2382 4281 2397 4398
rect 2443 4281 2447 4421
rect 2382 4264 2447 4281
rect 2493 4338 2559 4512
rect 2961 4558 3007 4644
rect 2961 4472 3007 4512
rect 3165 4558 3231 4598
rect 3165 4512 3185 4558
rect 2493 4286 2494 4338
rect 2546 4286 2559 4338
rect 1617 4026 1663 4047
rect 1921 4187 1967 4206
rect 1418 3980 1486 4005
rect 1921 3980 1967 4047
rect 2309 4179 2355 4198
rect 2309 3980 2355 4039
rect 2493 4179 2559 4286
rect 3054 4421 3119 4464
rect 3054 4338 3069 4421
rect 3054 4281 3069 4286
rect 3115 4281 3119 4421
rect 3054 4264 3119 4281
rect 3165 4338 3231 4512
rect 3633 4558 3679 4644
rect 3633 4472 3679 4512
rect 3837 4562 3903 4598
rect 3837 4510 3838 4562
rect 3890 4558 3903 4562
rect 3890 4510 3903 4512
rect 3165 4286 3166 4338
rect 3218 4286 3231 4338
rect 2493 4039 2513 4179
rect 2493 4026 2559 4039
rect 2981 4179 3027 4198
rect 2981 3980 3027 4039
rect 3165 4179 3231 4286
rect 3726 4421 3791 4464
rect 3726 4338 3741 4421
rect 3726 4281 3741 4286
rect 3787 4281 3791 4421
rect 3726 4264 3791 4281
rect 3165 4039 3185 4179
rect 3165 4026 3231 4039
rect 3653 4179 3699 4198
rect 3653 3980 3699 4039
rect 3837 4179 3903 4510
rect 4305 4558 4351 4644
rect 4305 4472 4351 4512
rect 4509 4562 4575 4598
rect 4509 4510 4510 4562
rect 4562 4558 4575 4562
rect 4562 4510 4575 4512
rect 4398 4421 4463 4464
rect 4398 4338 4413 4421
rect 4398 4281 4413 4286
rect 4459 4281 4463 4421
rect 4398 4264 4463 4281
rect 3837 4039 3857 4179
rect 3837 4026 3903 4039
rect 4325 4179 4371 4198
rect 4325 3980 4371 4039
rect 4509 4179 4575 4510
rect 4977 4558 5023 4644
rect 4977 4472 5023 4512
rect 5181 4558 5247 4598
rect 5181 4512 5201 4558
rect 5070 4450 5135 4464
rect 5122 4421 5135 4450
rect 5070 4281 5085 4398
rect 5131 4281 5135 4421
rect 5070 4264 5135 4281
rect 4509 4039 4529 4179
rect 4509 4026 4575 4039
rect 4997 4179 5043 4198
rect 4997 3980 5043 4039
rect 5181 4179 5247 4512
rect 5649 4558 5695 4644
rect 5649 4472 5695 4512
rect 5853 4558 5919 4598
rect 5853 4512 5873 4558
rect 5742 4450 5807 4464
rect 5794 4421 5807 4450
rect 5742 4281 5757 4398
rect 5803 4281 5807 4421
rect 5742 4264 5807 4281
rect 5181 4114 5201 4179
rect 5181 4062 5182 4114
rect 5181 4039 5201 4062
rect 5181 4026 5247 4039
rect 5669 4179 5715 4198
rect 5669 3980 5715 4039
rect 5853 4179 5919 4512
rect 6321 4558 6367 4644
rect 6321 4472 6367 4512
rect 6525 4558 6591 4598
rect 6525 4512 6545 4558
rect 6414 4421 6479 4464
rect 6414 4338 6429 4421
rect 6414 4281 6429 4286
rect 6475 4281 6479 4421
rect 6414 4264 6479 4281
rect 5853 4114 5873 4179
rect 5853 4062 5854 4114
rect 5853 4039 5873 4062
rect 5853 4026 5919 4039
rect 6341 4179 6387 4198
rect 6341 3980 6387 4039
rect 6525 4179 6591 4512
rect 6993 4558 7039 4644
rect 6993 4472 7039 4512
rect 7197 4562 7263 4598
rect 7197 4510 7198 4562
rect 7250 4558 7263 4562
rect 7250 4510 7263 4512
rect 7086 4421 7151 4464
rect 7086 4338 7101 4421
rect 7086 4281 7101 4286
rect 7147 4281 7151 4421
rect 7086 4264 7151 4281
rect 6525 4114 6545 4179
rect 6525 4062 6526 4114
rect 6525 4039 6545 4062
rect 6525 4026 6591 4039
rect 7013 4179 7059 4198
rect 7013 3980 7059 4039
rect 7197 4179 7263 4510
rect 7665 4558 7711 4644
rect 7665 4472 7711 4512
rect 7869 4558 7935 4598
rect 7869 4512 7889 4558
rect 7758 4421 7823 4464
rect 7758 4338 7773 4421
rect 7758 4281 7773 4286
rect 7819 4281 7823 4421
rect 7758 4264 7823 4281
rect 7197 4039 7217 4179
rect 7197 4026 7263 4039
rect 7685 4179 7731 4198
rect 7685 3980 7731 4039
rect 7869 4179 7935 4512
rect 8337 4558 8383 4644
rect 8337 4472 8383 4512
rect 8541 4562 8607 4598
rect 8541 4510 8542 4562
rect 8594 4558 8607 4562
rect 8594 4510 8607 4512
rect 8430 4450 8495 4464
rect 8482 4421 8495 4450
rect 8430 4281 8445 4398
rect 8491 4281 8495 4421
rect 8430 4264 8495 4281
rect 7869 4114 7889 4179
rect 7869 4062 7870 4114
rect 7869 4039 7889 4062
rect 7869 4026 7935 4039
rect 8357 4179 8403 4198
rect 8357 3980 8403 4039
rect 8541 4179 8607 4510
rect 8785 4558 8831 4644
rect 9374 4625 9442 4644
rect 8785 4485 8831 4512
rect 9089 4558 9135 4598
rect 8541 4039 8561 4179
rect 8541 4026 8607 4039
rect 8785 4393 8888 4439
rect 9028 4393 9040 4439
rect 8785 4187 8831 4393
rect 9089 4312 9135 4512
rect 9374 4478 9385 4625
rect 9431 4478 9442 4625
rect 9374 4467 9442 4478
rect 9681 4558 9727 4644
rect 9681 4472 9727 4512
rect 9885 4558 9951 4598
rect 9885 4512 9905 4558
rect 9774 4450 9839 4464
rect 9826 4421 9839 4450
rect 8882 4266 8896 4312
rect 9036 4266 9135 4312
rect 9374 4307 9442 4318
rect 9374 4261 9385 4307
rect 9431 4261 9442 4307
rect 9774 4281 9789 4398
rect 9835 4281 9839 4421
rect 9774 4264 9839 4281
rect 8785 4026 8831 4047
rect 9089 4187 9135 4206
rect 9089 3980 9135 4047
rect 9374 4179 9442 4261
rect 9374 4133 9385 4179
rect 9431 4133 9442 4179
rect 9374 4051 9442 4133
rect 9374 4005 9385 4051
rect 9431 4005 9442 4051
rect 9374 3980 9442 4005
rect 9701 4179 9747 4198
rect 9701 3980 9747 4039
rect 9885 4179 9951 4512
rect 10353 4558 10399 4644
rect 10353 4472 10399 4512
rect 10557 4558 10623 4598
rect 10557 4512 10577 4558
rect 10446 4450 10511 4464
rect 10498 4421 10511 4450
rect 10446 4281 10461 4398
rect 10507 4281 10511 4421
rect 10446 4264 10511 4281
rect 9885 4114 9905 4179
rect 9885 4062 9886 4114
rect 9885 4039 9905 4062
rect 9885 4026 9951 4039
rect 10373 4179 10419 4198
rect 10373 3980 10419 4039
rect 10557 4179 10623 4512
rect 11025 4558 11071 4644
rect 11025 4472 11071 4512
rect 11229 4558 11295 4598
rect 11229 4512 11249 4558
rect 11118 4421 11183 4464
rect 11118 4338 11133 4421
rect 11118 4281 11133 4286
rect 11179 4281 11183 4421
rect 11118 4264 11183 4281
rect 10557 4114 10577 4179
rect 10557 4062 10558 4114
rect 10557 4039 10577 4062
rect 10557 4026 10623 4039
rect 11045 4179 11091 4198
rect 11045 3980 11091 4039
rect 11229 4179 11295 4512
rect 11473 4558 11519 4644
rect 11473 4485 11519 4512
rect 11777 4558 11823 4598
rect 11229 4114 11249 4179
rect 11229 4062 11230 4114
rect 11229 4039 11249 4062
rect 11229 4026 11295 4039
rect 11473 4393 11576 4439
rect 11716 4393 11728 4439
rect 11473 4187 11519 4393
rect 11777 4312 11823 4512
rect 12257 4558 12303 4644
rect 12257 4472 12303 4512
rect 12461 4558 12527 4598
rect 12461 4512 12481 4558
rect 11570 4266 11584 4312
rect 11724 4266 11823 4312
rect 12350 4421 12415 4464
rect 12350 4338 12365 4421
rect 12350 4281 12365 4286
rect 12411 4281 12415 4421
rect 12350 4264 12415 4281
rect 11473 4026 11519 4047
rect 11777 4187 11823 4206
rect 11777 3980 11823 4047
rect 12277 4179 12323 4198
rect 12277 3980 12323 4039
rect 12461 4179 12527 4512
rect 12929 4558 12975 4644
rect 12929 4472 12975 4512
rect 13133 4558 13199 4598
rect 13133 4512 13153 4558
rect 13022 4421 13087 4464
rect 13022 4338 13037 4421
rect 13022 4281 13037 4286
rect 13083 4281 13087 4421
rect 13022 4264 13087 4281
rect 12461 4114 12481 4179
rect 12461 4062 12462 4114
rect 12461 4039 12481 4062
rect 12461 4026 12527 4039
rect 12949 4179 12995 4198
rect 12949 3980 12995 4039
rect 13133 4179 13199 4512
rect 13601 4558 13647 4644
rect 13601 4472 13647 4512
rect 13805 4558 13871 4598
rect 13805 4512 13825 4558
rect 13694 4421 13759 4464
rect 13694 4338 13709 4421
rect 13694 4281 13709 4286
rect 13755 4281 13759 4421
rect 13694 4264 13759 4281
rect 13133 4114 13153 4179
rect 13133 4062 13134 4114
rect 13133 4039 13153 4062
rect 13133 4026 13199 4039
rect 13621 4179 13667 4198
rect 13621 3980 13667 4039
rect 13805 4179 13871 4512
rect 14273 4558 14319 4644
rect 14273 4472 14319 4512
rect 14477 4558 14543 4598
rect 14477 4512 14497 4558
rect 14366 4450 14431 4464
rect 14418 4421 14431 4450
rect 14366 4281 14381 4398
rect 14427 4281 14431 4421
rect 14366 4264 14431 4281
rect 14477 4338 14543 4512
rect 14945 4558 14991 4644
rect 14945 4472 14991 4512
rect 15149 4562 15215 4598
rect 15149 4510 15150 4562
rect 15202 4558 15215 4562
rect 15202 4510 15215 4512
rect 14477 4286 14478 4338
rect 14530 4286 14543 4338
rect 13805 4114 13825 4179
rect 13805 4062 13806 4114
rect 13805 4039 13825 4062
rect 13805 4026 13871 4039
rect 14293 4179 14339 4198
rect 14293 3980 14339 4039
rect 14477 4179 14543 4286
rect 15038 4421 15103 4464
rect 15038 4338 15053 4421
rect 15038 4281 15053 4286
rect 15099 4281 15103 4421
rect 15038 4264 15103 4281
rect 14477 4039 14497 4179
rect 14477 4026 14543 4039
rect 14965 4179 15011 4198
rect 14965 3980 15011 4039
rect 15149 4179 15215 4510
rect 15617 4558 15663 4644
rect 15617 4472 15663 4512
rect 15821 4562 15887 4598
rect 15821 4510 15822 4562
rect 15874 4558 15887 4562
rect 15874 4510 15887 4512
rect 15710 4421 15775 4464
rect 15710 4338 15725 4421
rect 15710 4281 15725 4286
rect 15771 4281 15775 4421
rect 15710 4264 15775 4281
rect 15149 4039 15169 4179
rect 15149 4026 15215 4039
rect 15637 4179 15683 4198
rect 15637 3980 15683 4039
rect 15821 4179 15887 4510
rect 16289 4558 16335 4644
rect 16289 4472 16335 4512
rect 16493 4558 16559 4598
rect 16493 4512 16513 4558
rect 16382 4450 16447 4464
rect 16434 4421 16447 4450
rect 16382 4281 16397 4398
rect 16443 4281 16447 4421
rect 16382 4264 16447 4281
rect 16493 4450 16559 4512
rect 16737 4558 16783 4644
rect 17326 4625 17394 4644
rect 16737 4485 16783 4512
rect 17041 4558 17087 4598
rect 16493 4398 16494 4450
rect 16546 4398 16559 4450
rect 15821 4039 15841 4179
rect 15821 4026 15887 4039
rect 16309 4179 16355 4198
rect 16309 3980 16355 4039
rect 16493 4179 16559 4398
rect 16493 4039 16513 4179
rect 16493 4026 16559 4039
rect 16737 4393 16840 4439
rect 16980 4393 16992 4439
rect 16737 4187 16783 4393
rect 17041 4312 17087 4512
rect 17326 4478 17337 4625
rect 17383 4478 17394 4625
rect 17326 4467 17394 4478
rect 17633 4558 17679 4644
rect 17633 4472 17679 4512
rect 17837 4562 17903 4598
rect 17837 4510 17838 4562
rect 17890 4558 17903 4562
rect 17890 4510 17903 4512
rect 17726 4450 17791 4464
rect 17778 4421 17791 4450
rect 16834 4266 16848 4312
rect 16988 4266 17087 4312
rect 17326 4307 17394 4318
rect 17326 4261 17337 4307
rect 17383 4261 17394 4307
rect 17726 4281 17741 4398
rect 17787 4281 17791 4421
rect 17726 4264 17791 4281
rect 16737 4026 16783 4047
rect 17041 4187 17087 4206
rect 17041 3980 17087 4047
rect 17326 4179 17394 4261
rect 17326 4133 17337 4179
rect 17383 4133 17394 4179
rect 17326 4051 17394 4133
rect 17326 4005 17337 4051
rect 17383 4005 17394 4051
rect 17326 3980 17394 4005
rect 17653 4179 17699 4198
rect 17653 3980 17699 4039
rect 17837 4179 17903 4510
rect 18305 4558 18351 4644
rect 18305 4472 18351 4512
rect 18509 4562 18575 4598
rect 18509 4510 18510 4562
rect 18562 4558 18575 4562
rect 18562 4510 18575 4512
rect 18398 4450 18463 4464
rect 18450 4421 18463 4450
rect 18398 4281 18413 4398
rect 18459 4281 18463 4421
rect 18398 4264 18463 4281
rect 17837 4039 17857 4179
rect 17837 4026 17903 4039
rect 18325 4179 18371 4198
rect 18325 3980 18371 4039
rect 18509 4179 18575 4510
rect 18977 4558 19023 4644
rect 18977 4472 19023 4512
rect 19181 4558 19247 4598
rect 19181 4512 19201 4558
rect 19070 4450 19135 4464
rect 19122 4421 19135 4450
rect 19070 4281 19085 4398
rect 19131 4281 19135 4421
rect 19070 4264 19135 4281
rect 18509 4039 18529 4179
rect 18509 4026 18575 4039
rect 18997 4179 19043 4198
rect 18997 3980 19043 4039
rect 19181 4179 19247 4512
rect 19649 4558 19695 4644
rect 19649 4472 19695 4512
rect 19853 4562 19919 4598
rect 19853 4510 19854 4562
rect 19906 4558 19919 4562
rect 19906 4510 19919 4512
rect 19742 4421 19807 4464
rect 19742 4338 19757 4421
rect 19742 4281 19757 4286
rect 19803 4281 19807 4421
rect 19742 4264 19807 4281
rect 19181 4114 19201 4179
rect 19181 4062 19182 4114
rect 19181 4039 19201 4062
rect 19181 4026 19247 4039
rect 19669 4179 19715 4198
rect 19669 3980 19715 4039
rect 19853 4179 19919 4510
rect 20321 4558 20367 4644
rect 20321 4472 20367 4512
rect 20525 4562 20591 4598
rect 20525 4510 20526 4562
rect 20578 4558 20591 4562
rect 20578 4510 20591 4512
rect 20414 4450 20479 4464
rect 20466 4421 20479 4450
rect 20414 4281 20429 4398
rect 20475 4281 20479 4421
rect 20414 4264 20479 4281
rect 19853 4039 19873 4179
rect 19853 4026 19919 4039
rect 20341 4179 20387 4198
rect 20341 3980 20387 4039
rect 20525 4179 20591 4510
rect 20993 4558 21039 4644
rect 20993 4472 21039 4512
rect 21197 4562 21263 4598
rect 21197 4510 21198 4562
rect 21250 4558 21263 4562
rect 21250 4510 21263 4512
rect 21086 4450 21151 4464
rect 21138 4421 21151 4450
rect 21086 4281 21101 4398
rect 21147 4281 21151 4421
rect 21086 4264 21151 4281
rect 20525 4039 20545 4179
rect 20525 4026 20591 4039
rect 21013 4179 21059 4198
rect 21013 3980 21059 4039
rect 21197 4179 21263 4510
rect 21197 4039 21217 4179
rect 21197 4026 21263 4039
rect 21745 4558 21811 4598
rect 21791 4512 21811 4558
rect 21745 4179 21811 4512
rect 21969 4558 22015 4644
rect 21969 4472 22015 4512
rect 22482 4625 22550 4644
rect 22482 4478 22493 4625
rect 22539 4478 22550 4625
rect 22482 4466 22550 4478
rect 21857 4421 21922 4464
rect 21857 4281 21861 4421
rect 21907 4338 21922 4421
rect 21907 4281 21922 4286
rect 21857 4264 21922 4281
rect 22482 4307 22550 4320
rect 22482 4261 22493 4307
rect 22539 4261 22550 4307
rect 21791 4114 21811 4179
rect 21810 4062 21811 4114
rect 21791 4039 21811 4062
rect 21745 4026 21811 4039
rect 21949 4179 21995 4198
rect 21949 3980 21995 4039
rect 22482 4179 22550 4261
rect 22482 4133 22493 4179
rect 22539 4133 22550 4179
rect 22482 4051 22550 4133
rect 22482 4005 22493 4051
rect 22539 4005 22550 4051
rect 22482 3980 22550 4005
rect 1344 3946 22624 3980
rect 1344 3894 3874 3946
rect 4134 3894 9194 3946
rect 9454 3894 14514 3946
rect 14774 3894 19834 3946
rect 20094 3894 22624 3946
rect 1344 3860 22624 3894
rect 1418 3835 1486 3860
rect 1418 3789 1429 3835
rect 1475 3789 1486 3835
rect 1418 3707 1486 3789
rect 1418 3661 1429 3707
rect 1475 3661 1486 3707
rect 1418 3579 1486 3661
rect 1418 3533 1429 3579
rect 1475 3533 1486 3579
rect 1418 3520 1486 3533
rect 1617 3793 1663 3814
rect 1617 3447 1663 3653
rect 1921 3793 1967 3860
rect 1921 3634 1967 3653
rect 2065 3793 2111 3814
rect 1714 3528 1728 3574
rect 1868 3528 1967 3574
rect 1617 3401 1720 3447
rect 1860 3401 1872 3447
rect 1418 3362 1486 3374
rect 1418 3215 1429 3362
rect 1475 3215 1486 3362
rect 1418 3196 1486 3215
rect 1617 3328 1663 3353
rect 1617 3196 1663 3282
rect 1921 3328 1967 3528
rect 2065 3447 2111 3653
rect 2369 3793 2415 3860
rect 2369 3634 2415 3653
rect 2757 3801 2803 3860
rect 2757 3642 2803 3661
rect 2941 3801 3007 3814
rect 2941 3778 2961 3801
rect 2941 3726 2942 3778
rect 2941 3661 2961 3726
rect 2162 3528 2176 3574
rect 2316 3528 2415 3574
rect 2065 3401 2168 3447
rect 2308 3401 2320 3447
rect 1921 3242 1967 3282
rect 2065 3328 2111 3353
rect 2065 3196 2111 3282
rect 2369 3328 2415 3528
rect 2830 3559 2895 3576
rect 2830 3554 2845 3559
rect 2830 3419 2845 3502
rect 2891 3419 2895 3559
rect 2830 3376 2895 3419
rect 2369 3242 2415 3282
rect 2737 3328 2783 3368
rect 2737 3196 2783 3282
rect 2941 3328 3007 3661
rect 3429 3801 3475 3860
rect 3429 3642 3475 3661
rect 3613 3801 3679 3814
rect 3613 3778 3633 3801
rect 3613 3726 3614 3778
rect 3613 3661 3633 3726
rect 3502 3559 3567 3576
rect 3502 3554 3517 3559
rect 3502 3419 3517 3502
rect 3563 3419 3567 3559
rect 3502 3376 3567 3419
rect 2941 3282 2961 3328
rect 2941 3242 3007 3282
rect 3409 3328 3455 3368
rect 3409 3196 3455 3282
rect 3613 3328 3679 3661
rect 4101 3801 4147 3860
rect 4101 3642 4147 3661
rect 4285 3801 4351 3814
rect 4285 3778 4305 3801
rect 4285 3726 4286 3778
rect 4285 3661 4305 3726
rect 4174 3559 4239 3576
rect 4174 3554 4189 3559
rect 4174 3419 4189 3502
rect 4235 3419 4239 3559
rect 4174 3376 4239 3419
rect 3613 3282 3633 3328
rect 3613 3242 3679 3282
rect 4081 3328 4127 3368
rect 4081 3196 4127 3282
rect 4285 3328 4351 3661
rect 4773 3801 4819 3860
rect 5342 3835 5410 3860
rect 4773 3642 4819 3661
rect 4957 3801 5023 3814
rect 4957 3778 4977 3801
rect 4957 3726 4958 3778
rect 4957 3661 4977 3726
rect 4846 3559 4911 3576
rect 4846 3442 4861 3559
rect 4907 3419 4911 3559
rect 4898 3390 4911 3419
rect 4846 3376 4911 3390
rect 4285 3282 4305 3328
rect 4285 3242 4351 3282
rect 4753 3328 4799 3368
rect 4753 3196 4799 3282
rect 4957 3328 5023 3661
rect 5342 3789 5353 3835
rect 5399 3789 5410 3835
rect 5342 3707 5410 3789
rect 5342 3661 5353 3707
rect 5399 3661 5410 3707
rect 5342 3579 5410 3661
rect 5342 3533 5353 3579
rect 5399 3533 5410 3579
rect 5342 3522 5410 3533
rect 5729 3801 5795 3814
rect 5775 3661 5795 3801
rect 5729 3442 5795 3661
rect 5933 3801 5979 3860
rect 5933 3642 5979 3661
rect 6401 3801 6467 3814
rect 6447 3778 6467 3801
rect 6466 3726 6467 3778
rect 6447 3661 6467 3726
rect 5729 3390 5742 3442
rect 5794 3390 5795 3442
rect 4957 3282 4977 3328
rect 4957 3242 5023 3282
rect 5342 3362 5410 3373
rect 5342 3215 5353 3362
rect 5399 3215 5410 3362
rect 5729 3328 5795 3390
rect 5841 3559 5906 3576
rect 5841 3419 5845 3559
rect 5891 3554 5906 3559
rect 5891 3419 5906 3502
rect 5841 3376 5906 3419
rect 5775 3282 5795 3328
rect 5729 3242 5795 3282
rect 5953 3328 5999 3368
rect 5342 3196 5410 3215
rect 5953 3196 5999 3282
rect 6401 3328 6467 3661
rect 6605 3801 6651 3860
rect 6605 3642 6651 3661
rect 7073 3801 7139 3814
rect 7119 3778 7139 3801
rect 7138 3726 7139 3778
rect 7119 3661 7139 3726
rect 6513 3559 6578 3576
rect 6513 3419 6517 3559
rect 6563 3554 6578 3559
rect 6563 3419 6578 3502
rect 6513 3376 6578 3419
rect 6447 3282 6467 3328
rect 6401 3242 6467 3282
rect 6625 3328 6671 3368
rect 6625 3196 6671 3282
rect 7073 3328 7139 3661
rect 7277 3801 7323 3860
rect 7277 3642 7323 3661
rect 7685 3801 7731 3860
rect 7685 3642 7731 3661
rect 7869 3801 7935 3814
rect 7869 3778 7889 3801
rect 7869 3726 7870 3778
rect 7869 3661 7889 3726
rect 7185 3559 7250 3576
rect 7185 3419 7189 3559
rect 7235 3554 7250 3559
rect 7235 3419 7250 3502
rect 7185 3376 7250 3419
rect 7758 3559 7823 3576
rect 7758 3554 7773 3559
rect 7758 3419 7773 3502
rect 7819 3419 7823 3559
rect 7758 3376 7823 3419
rect 7119 3282 7139 3328
rect 7073 3242 7139 3282
rect 7297 3328 7343 3368
rect 7297 3196 7343 3282
rect 7665 3328 7711 3368
rect 7665 3196 7711 3282
rect 7869 3328 7935 3661
rect 7869 3282 7889 3328
rect 7869 3242 7935 3282
rect 8417 3801 8483 3814
rect 8463 3661 8483 3801
rect 8417 3554 8483 3661
rect 8621 3801 8667 3860
rect 8621 3642 8667 3661
rect 8785 3793 8831 3814
rect 8417 3502 8430 3554
rect 8482 3502 8483 3554
rect 8417 3328 8483 3502
rect 8529 3559 8594 3576
rect 8529 3419 8533 3559
rect 8579 3554 8594 3559
rect 8579 3419 8594 3502
rect 8529 3376 8594 3419
rect 8785 3447 8831 3653
rect 9089 3793 9135 3860
rect 9089 3634 9135 3653
rect 9262 3835 9330 3860
rect 9262 3789 9273 3835
rect 9319 3789 9330 3835
rect 9262 3707 9330 3789
rect 9262 3661 9273 3707
rect 9319 3661 9330 3707
rect 9262 3579 9330 3661
rect 8882 3528 8896 3574
rect 9036 3528 9135 3574
rect 8785 3401 8888 3447
rect 9028 3401 9040 3447
rect 8463 3282 8483 3328
rect 8417 3242 8483 3282
rect 8641 3328 8687 3368
rect 8641 3196 8687 3282
rect 8785 3328 8831 3355
rect 8785 3196 8831 3282
rect 9089 3328 9135 3528
rect 9262 3533 9273 3579
rect 9319 3533 9330 3579
rect 9262 3522 9330 3533
rect 9649 3801 9715 3814
rect 9695 3661 9715 3801
rect 9649 3554 9715 3661
rect 9853 3801 9899 3860
rect 9853 3642 9899 3661
rect 10261 3801 10307 3860
rect 10261 3642 10307 3661
rect 10445 3801 10511 3814
rect 10445 3661 10465 3801
rect 9649 3502 9662 3554
rect 9714 3502 9715 3554
rect 9089 3242 9135 3282
rect 9262 3362 9330 3373
rect 9262 3215 9273 3362
rect 9319 3215 9330 3362
rect 9649 3328 9715 3502
rect 9761 3559 9826 3576
rect 9761 3419 9765 3559
rect 9811 3554 9826 3559
rect 9811 3419 9826 3502
rect 9761 3376 9826 3419
rect 10334 3559 10399 3576
rect 10334 3554 10349 3559
rect 10334 3419 10349 3502
rect 10395 3419 10399 3559
rect 10334 3376 10399 3419
rect 10445 3554 10511 3661
rect 10933 3801 10979 3860
rect 10933 3642 10979 3661
rect 11117 3801 11183 3814
rect 11117 3661 11137 3801
rect 10445 3502 10446 3554
rect 10498 3502 10511 3554
rect 9695 3282 9715 3328
rect 9649 3242 9715 3282
rect 9873 3328 9919 3368
rect 9262 3196 9330 3215
rect 9873 3196 9919 3282
rect 10241 3328 10287 3368
rect 10241 3196 10287 3282
rect 10445 3328 10511 3502
rect 11006 3559 11071 3576
rect 11006 3442 11021 3559
rect 11067 3419 11071 3559
rect 11058 3390 11071 3419
rect 11006 3376 11071 3390
rect 11117 3554 11183 3661
rect 11117 3502 11118 3554
rect 11170 3502 11183 3554
rect 10445 3282 10465 3328
rect 10445 3242 10511 3282
rect 10913 3328 10959 3368
rect 10913 3196 10959 3282
rect 11117 3328 11183 3502
rect 11117 3282 11137 3328
rect 11117 3242 11183 3282
rect 11665 3801 11731 3814
rect 11711 3661 11731 3801
rect 11665 3554 11731 3661
rect 11869 3801 11915 3860
rect 11869 3642 11915 3661
rect 12033 3793 12079 3814
rect 11665 3502 11678 3554
rect 11730 3502 11731 3554
rect 11665 3328 11731 3502
rect 11777 3559 11842 3576
rect 11777 3419 11781 3559
rect 11827 3442 11842 3559
rect 11777 3390 11790 3419
rect 12033 3447 12079 3653
rect 12337 3793 12383 3860
rect 12337 3634 12383 3653
rect 12481 3793 12527 3814
rect 12130 3528 12144 3574
rect 12284 3528 12383 3574
rect 12033 3401 12136 3447
rect 12276 3401 12288 3447
rect 11777 3376 11842 3390
rect 11711 3282 11731 3328
rect 11665 3242 11731 3282
rect 11889 3328 11935 3368
rect 11889 3196 11935 3282
rect 12033 3328 12079 3353
rect 12033 3196 12079 3282
rect 12337 3328 12383 3528
rect 12481 3447 12527 3653
rect 12785 3793 12831 3860
rect 12785 3634 12831 3653
rect 13182 3835 13250 3860
rect 13182 3789 13193 3835
rect 13239 3789 13250 3835
rect 13182 3707 13250 3789
rect 13182 3661 13193 3707
rect 13239 3661 13250 3707
rect 13182 3579 13250 3661
rect 12578 3528 12592 3574
rect 12732 3528 12831 3574
rect 12481 3401 12584 3447
rect 12724 3401 12736 3447
rect 12337 3242 12383 3282
rect 12481 3328 12527 3353
rect 12481 3196 12527 3282
rect 12785 3328 12831 3528
rect 13182 3533 13193 3579
rect 13239 3533 13250 3579
rect 13182 3522 13250 3533
rect 13377 3793 13423 3814
rect 13377 3447 13423 3653
rect 13681 3793 13727 3860
rect 13681 3634 13727 3653
rect 13845 3801 13891 3860
rect 13845 3642 13891 3661
rect 14029 3801 14095 3814
rect 14029 3661 14049 3801
rect 13474 3528 13488 3574
rect 13628 3528 13727 3574
rect 13377 3401 13480 3447
rect 13620 3401 13632 3447
rect 12785 3242 12831 3282
rect 13182 3362 13250 3373
rect 13182 3215 13193 3362
rect 13239 3215 13250 3362
rect 13182 3196 13250 3215
rect 13377 3328 13423 3355
rect 13377 3196 13423 3282
rect 13681 3328 13727 3528
rect 13918 3559 13983 3576
rect 13918 3442 13933 3559
rect 13979 3419 13983 3559
rect 13970 3390 13983 3419
rect 13918 3376 13983 3390
rect 14029 3442 14095 3661
rect 14517 3801 14563 3860
rect 14517 3642 14563 3661
rect 14701 3801 14767 3814
rect 14701 3661 14721 3801
rect 14029 3390 14030 3442
rect 14082 3390 14095 3442
rect 13681 3242 13727 3282
rect 13825 3328 13871 3368
rect 13825 3196 13871 3282
rect 14029 3328 14095 3390
rect 14590 3559 14655 3576
rect 14590 3554 14605 3559
rect 14590 3419 14605 3502
rect 14651 3419 14655 3559
rect 14590 3376 14655 3419
rect 14701 3442 14767 3661
rect 15189 3801 15235 3860
rect 15189 3642 15235 3661
rect 15373 3801 15439 3814
rect 15373 3661 15393 3801
rect 14701 3390 14702 3442
rect 14754 3390 14767 3442
rect 14029 3282 14049 3328
rect 14029 3242 14095 3282
rect 14497 3328 14543 3368
rect 14497 3196 14543 3282
rect 14701 3328 14767 3390
rect 15262 3559 15327 3576
rect 15262 3554 15277 3559
rect 15262 3419 15277 3502
rect 15323 3419 15327 3559
rect 15262 3376 15327 3419
rect 15373 3442 15439 3661
rect 15861 3801 15907 3860
rect 15861 3642 15907 3661
rect 16045 3801 16111 3814
rect 16045 3661 16065 3801
rect 15934 3559 15999 3576
rect 15586 3502 15598 3554
rect 15650 3551 15662 3554
rect 15810 3551 15822 3554
rect 15650 3505 15822 3551
rect 15650 3502 15662 3505
rect 15810 3502 15822 3505
rect 15874 3502 15886 3554
rect 15373 3390 15374 3442
rect 15426 3390 15439 3442
rect 14701 3282 14721 3328
rect 14701 3242 14767 3282
rect 15169 3328 15215 3368
rect 15169 3196 15215 3282
rect 15373 3328 15439 3390
rect 15934 3442 15949 3559
rect 15995 3419 15999 3559
rect 15986 3390 15999 3419
rect 15934 3376 15999 3390
rect 16045 3442 16111 3661
rect 16533 3801 16579 3860
rect 17102 3835 17170 3860
rect 16533 3642 16579 3661
rect 16717 3801 16783 3814
rect 16717 3661 16737 3801
rect 16045 3390 16046 3442
rect 16098 3390 16111 3442
rect 15373 3282 15393 3328
rect 15373 3242 15439 3282
rect 15841 3328 15887 3368
rect 15841 3196 15887 3282
rect 16045 3328 16111 3390
rect 16606 3559 16671 3576
rect 16606 3554 16621 3559
rect 16606 3419 16621 3502
rect 16667 3419 16671 3559
rect 16606 3376 16671 3419
rect 16717 3442 16783 3661
rect 17102 3789 17113 3835
rect 17159 3789 17170 3835
rect 17102 3707 17170 3789
rect 17102 3661 17113 3707
rect 17159 3661 17170 3707
rect 17102 3579 17170 3661
rect 17429 3801 17475 3860
rect 17429 3642 17475 3661
rect 17613 3801 17679 3814
rect 17613 3778 17633 3801
rect 17613 3726 17614 3778
rect 17613 3661 17633 3726
rect 17102 3533 17113 3579
rect 17159 3533 17170 3579
rect 17102 3522 17170 3533
rect 17502 3559 17567 3576
rect 17502 3554 17517 3559
rect 16717 3390 16718 3442
rect 16770 3390 16783 3442
rect 16045 3282 16065 3328
rect 16045 3242 16111 3282
rect 16513 3328 16559 3368
rect 16513 3196 16559 3282
rect 16717 3328 16783 3390
rect 17502 3419 17517 3502
rect 17563 3419 17567 3559
rect 17502 3376 17567 3419
rect 16717 3282 16737 3328
rect 16717 3242 16783 3282
rect 17102 3362 17170 3373
rect 17102 3215 17113 3362
rect 17159 3215 17170 3362
rect 17102 3196 17170 3215
rect 17409 3328 17455 3368
rect 17409 3196 17455 3282
rect 17613 3328 17679 3661
rect 18101 3801 18147 3860
rect 18101 3642 18147 3661
rect 18285 3801 18351 3814
rect 18285 3661 18305 3801
rect 18174 3559 18239 3576
rect 18174 3554 18189 3559
rect 18174 3419 18189 3502
rect 18235 3419 18239 3559
rect 18174 3376 18239 3419
rect 18285 3442 18351 3661
rect 18773 3801 18819 3860
rect 18773 3642 18819 3661
rect 18957 3801 19023 3814
rect 18957 3661 18977 3801
rect 18285 3390 18286 3442
rect 18338 3390 18351 3442
rect 17613 3282 17633 3328
rect 17613 3242 17679 3282
rect 18081 3328 18127 3368
rect 18081 3196 18127 3282
rect 18285 3328 18351 3390
rect 18846 3559 18911 3576
rect 18846 3554 18861 3559
rect 18846 3419 18861 3502
rect 18907 3419 18911 3559
rect 18846 3376 18911 3419
rect 18957 3442 19023 3661
rect 19445 3801 19491 3860
rect 19445 3642 19491 3661
rect 19629 3801 19695 3814
rect 19629 3778 19649 3801
rect 19629 3726 19630 3778
rect 19629 3661 19649 3726
rect 18957 3390 18958 3442
rect 19010 3390 19023 3442
rect 18285 3282 18305 3328
rect 18285 3242 18351 3282
rect 18753 3328 18799 3368
rect 18753 3196 18799 3282
rect 18957 3328 19023 3390
rect 19518 3559 19583 3576
rect 19518 3442 19533 3559
rect 19579 3419 19583 3559
rect 19570 3390 19583 3419
rect 19518 3376 19583 3390
rect 18957 3282 18977 3328
rect 18957 3242 19023 3282
rect 19425 3328 19471 3368
rect 19425 3196 19471 3282
rect 19629 3328 19695 3661
rect 20117 3801 20163 3860
rect 20117 3642 20163 3661
rect 20301 3801 20367 3814
rect 20301 3778 20321 3801
rect 20301 3726 20302 3778
rect 20301 3661 20321 3726
rect 20190 3559 20255 3576
rect 20190 3554 20205 3559
rect 20190 3419 20205 3502
rect 20251 3419 20255 3559
rect 20190 3376 20255 3419
rect 19629 3282 19649 3328
rect 19629 3242 19695 3282
rect 20097 3328 20143 3368
rect 20097 3196 20143 3282
rect 20301 3328 20367 3661
rect 20545 3793 20591 3814
rect 20545 3447 20591 3653
rect 20849 3793 20895 3860
rect 20849 3634 20895 3653
rect 21022 3835 21090 3860
rect 21022 3789 21033 3835
rect 21079 3789 21090 3835
rect 21022 3707 21090 3789
rect 21022 3661 21033 3707
rect 21079 3661 21090 3707
rect 21022 3579 21090 3661
rect 20642 3528 20656 3574
rect 20796 3528 20895 3574
rect 20545 3401 20648 3447
rect 20788 3401 20800 3447
rect 20301 3282 20321 3328
rect 20301 3242 20367 3282
rect 20545 3328 20591 3355
rect 20545 3196 20591 3282
rect 20849 3328 20895 3528
rect 21022 3533 21033 3579
rect 21079 3533 21090 3579
rect 21022 3522 21090 3533
rect 21217 3793 21263 3814
rect 21217 3447 21263 3653
rect 21521 3793 21567 3860
rect 21521 3634 21567 3653
rect 21665 3793 21711 3814
rect 21314 3528 21328 3574
rect 21468 3528 21567 3574
rect 21217 3401 21320 3447
rect 21460 3401 21472 3447
rect 20849 3242 20895 3282
rect 21022 3362 21090 3373
rect 21022 3215 21033 3362
rect 21079 3215 21090 3362
rect 21022 3196 21090 3215
rect 21217 3328 21263 3353
rect 21217 3196 21263 3282
rect 21521 3328 21567 3528
rect 21665 3447 21711 3653
rect 21969 3793 22015 3860
rect 21969 3634 22015 3653
rect 22482 3835 22550 3860
rect 22482 3789 22493 3835
rect 22539 3789 22550 3835
rect 22482 3707 22550 3789
rect 22482 3661 22493 3707
rect 22539 3661 22550 3707
rect 22482 3579 22550 3661
rect 21762 3528 21776 3574
rect 21916 3528 22015 3574
rect 21665 3401 21768 3447
rect 21908 3401 21920 3447
rect 21521 3242 21567 3282
rect 21665 3328 21711 3353
rect 21665 3196 21711 3282
rect 21969 3328 22015 3528
rect 22482 3533 22493 3579
rect 22539 3533 22550 3579
rect 22482 3520 22550 3533
rect 21969 3242 22015 3282
rect 22482 3362 22550 3374
rect 22482 3215 22493 3362
rect 22539 3215 22550 3362
rect 22482 3196 22550 3215
rect 1344 3162 22784 3196
rect 1344 3110 6534 3162
rect 6794 3110 11854 3162
rect 12114 3110 17174 3162
rect 17434 3110 22494 3162
rect 22754 3110 22784 3162
rect 1344 3076 22784 3110
<< via1 >>
rect 3874 16438 4134 16490
rect 9194 16438 9454 16490
rect 14514 16438 14774 16490
rect 19834 16438 20094 16490
rect 6534 15654 6794 15706
rect 11854 15654 12114 15706
rect 17174 15654 17434 15706
rect 22494 15654 22754 15706
rect 3874 14870 4134 14922
rect 9194 14870 9454 14922
rect 14514 14870 14774 14922
rect 19834 14870 20094 14922
rect 16830 14637 16863 14642
rect 16863 14637 16882 14642
rect 16830 14590 16882 14637
rect 16942 14395 16979 14418
rect 16979 14395 16994 14418
rect 16942 14366 16994 14395
rect 17614 14395 17651 14418
rect 17651 14395 17666 14418
rect 17614 14366 17666 14395
rect 17502 14304 17554 14306
rect 17502 14258 17535 14304
rect 17535 14258 17554 14304
rect 17502 14254 17554 14258
rect 6534 14086 6794 14138
rect 11854 14086 12114 14138
rect 17174 14086 17434 14138
rect 22494 14086 22754 14138
rect 16158 13694 16173 13746
rect 16173 13694 16210 13746
rect 16830 13694 16845 13746
rect 16845 13694 16882 13746
rect 16270 13470 16289 13522
rect 16289 13470 16322 13522
rect 16942 13470 16961 13522
rect 16961 13470 16994 13522
rect 17726 13694 17741 13746
rect 17741 13694 17778 13746
rect 18398 13694 18413 13746
rect 18413 13694 18450 13746
rect 17838 13470 17857 13522
rect 17857 13470 17890 13522
rect 18510 13470 18529 13522
rect 18529 13470 18562 13522
rect 3874 13302 4134 13354
rect 9194 13302 9454 13354
rect 14514 13302 14774 13354
rect 19834 13302 20094 13354
rect 14926 13134 14945 13186
rect 14945 13134 14978 13186
rect 14814 12827 14829 12850
rect 14829 12827 14866 12850
rect 14814 12798 14866 12827
rect 15486 12827 15501 12850
rect 15501 12827 15538 12850
rect 15486 12798 15538 12827
rect 16158 12827 16173 12850
rect 16173 12827 16210 12850
rect 16158 12798 16210 12827
rect 15598 12736 15650 12738
rect 15598 12690 15617 12736
rect 15617 12690 15650 12736
rect 15598 12686 15650 12690
rect 16830 12827 16845 12850
rect 16845 12827 16882 12850
rect 16830 12798 16882 12827
rect 16270 12736 16322 12738
rect 16270 12690 16289 12736
rect 16289 12690 16322 12736
rect 16270 12686 16322 12690
rect 17502 12910 17517 12962
rect 17517 12910 17554 12962
rect 16942 12736 16994 12738
rect 16942 12690 16961 12736
rect 16961 12690 16994 12736
rect 16942 12686 16994 12690
rect 18286 13134 18305 13186
rect 18305 13134 18338 13186
rect 18174 12827 18189 12850
rect 18189 12827 18226 12850
rect 18174 12798 18226 12827
rect 17614 12736 17666 12738
rect 17614 12690 17633 12736
rect 17633 12690 17666 12736
rect 17614 12686 17666 12690
rect 18958 13134 18977 13186
rect 18977 13134 19010 13186
rect 18846 12910 18861 12962
rect 18861 12910 18898 12962
rect 19518 12827 19533 12850
rect 19533 12827 19570 12850
rect 19518 12798 19570 12827
rect 19630 12736 19682 12738
rect 19630 12690 19649 12736
rect 19649 12690 19682 12736
rect 19630 12686 19682 12690
rect 6534 12518 6794 12570
rect 11854 12518 12114 12570
rect 17174 12518 17434 12570
rect 22494 12518 22754 12570
rect 14142 12126 14157 12178
rect 14157 12126 14194 12178
rect 14814 12126 14829 12178
rect 14829 12126 14866 12178
rect 14254 11902 14273 11954
rect 14273 11902 14306 11954
rect 15486 12126 15501 12178
rect 15501 12126 15538 12178
rect 14926 11902 14945 11954
rect 14945 11902 14978 11954
rect 16158 12126 16173 12178
rect 16173 12126 16210 12178
rect 15598 11902 15617 11954
rect 15617 11902 15650 11954
rect 16830 12126 16845 12178
rect 16845 12126 16882 12178
rect 16270 11902 16289 11954
rect 16289 11902 16322 11954
rect 17726 12261 17778 12290
rect 17726 12238 17741 12261
rect 17741 12238 17778 12261
rect 16942 11902 16961 11954
rect 16961 11902 16994 11954
rect 17838 12238 17890 12290
rect 18398 12261 18450 12290
rect 18398 12238 18413 12261
rect 18413 12238 18450 12261
rect 19182 12398 19234 12402
rect 19182 12352 19201 12398
rect 19201 12352 19234 12398
rect 19182 12350 19234 12352
rect 19070 12261 19122 12290
rect 19070 12238 19085 12261
rect 19085 12238 19122 12261
rect 18510 11902 18529 11954
rect 18529 11902 18562 11954
rect 19854 12398 19906 12402
rect 19854 12352 19873 12398
rect 19873 12352 19906 12398
rect 19854 12350 19906 12352
rect 19742 12261 19794 12290
rect 19742 12238 19757 12261
rect 19757 12238 19794 12261
rect 20414 12261 20466 12290
rect 20414 12238 20429 12261
rect 20429 12238 20466 12261
rect 20526 12238 20578 12290
rect 3874 11734 4134 11786
rect 9194 11734 9454 11786
rect 14514 11734 14774 11786
rect 19834 11734 20094 11786
rect 6078 11230 6130 11282
rect 6190 11259 6227 11282
rect 6227 11259 6242 11282
rect 6190 11230 6242 11259
rect 6974 11259 7011 11282
rect 7011 11259 7026 11282
rect 6974 11230 7026 11259
rect 6862 11168 6914 11170
rect 6862 11122 6895 11168
rect 6895 11122 6914 11168
rect 6862 11118 6914 11122
rect 7646 11259 7683 11282
rect 7683 11259 7698 11282
rect 7646 11230 7698 11259
rect 7534 11168 7586 11170
rect 7534 11122 7567 11168
rect 7567 11122 7586 11168
rect 7534 11118 7586 11122
rect 8318 11259 8355 11282
rect 8355 11259 8370 11282
rect 8318 11230 8370 11259
rect 8206 11168 8258 11170
rect 8206 11122 8239 11168
rect 8239 11122 8258 11168
rect 8206 11118 8258 11122
rect 9214 11259 9229 11282
rect 9229 11259 9266 11282
rect 9214 11230 9266 11259
rect 9886 11259 9901 11282
rect 9901 11259 9938 11282
rect 9886 11230 9938 11259
rect 9326 11168 9378 11170
rect 9326 11122 9345 11168
rect 9345 11122 9378 11168
rect 9326 11118 9378 11122
rect 10670 11501 10689 11506
rect 10689 11501 10722 11506
rect 10670 11454 10722 11501
rect 10558 11259 10573 11282
rect 10573 11259 10610 11282
rect 10558 11230 10610 11259
rect 9998 11168 10050 11170
rect 9998 11122 10017 11168
rect 10017 11122 10050 11168
rect 9998 11118 10050 11122
rect 12126 11259 12141 11282
rect 12141 11259 12178 11282
rect 12126 11230 12178 11259
rect 12238 11230 12290 11282
rect 12798 11259 12813 11282
rect 12813 11259 12850 11282
rect 12798 11230 12850 11259
rect 13694 11259 13709 11282
rect 13709 11259 13746 11282
rect 13694 11230 13746 11259
rect 12910 11168 12962 11170
rect 12910 11122 12929 11168
rect 12929 11122 12962 11168
rect 12910 11118 12962 11122
rect 13806 11168 13858 11170
rect 13806 11122 13825 11168
rect 13825 11122 13858 11168
rect 13806 11118 13858 11122
rect 14814 11259 14829 11282
rect 14829 11259 14866 11282
rect 14814 11230 14866 11259
rect 14926 11342 14978 11394
rect 15486 11259 15501 11282
rect 15501 11259 15538 11282
rect 15486 11230 15538 11259
rect 15598 11342 15650 11394
rect 16158 11259 16173 11282
rect 16173 11259 16210 11282
rect 16158 11230 16210 11259
rect 16270 11342 16322 11394
rect 16830 11342 16845 11394
rect 16845 11342 16882 11394
rect 17614 11566 17633 11618
rect 17633 11566 17666 11618
rect 16942 11342 16994 11394
rect 17502 11342 17517 11394
rect 17517 11342 17554 11394
rect 18174 11342 18189 11394
rect 18189 11342 18226 11394
rect 18846 11342 18861 11394
rect 18861 11342 18898 11394
rect 18286 11168 18338 11170
rect 18286 11122 18305 11168
rect 18305 11122 18338 11168
rect 18286 11118 18338 11122
rect 19630 11566 19649 11618
rect 19649 11566 19682 11618
rect 19518 11342 19533 11394
rect 19533 11342 19570 11394
rect 18958 11168 19010 11170
rect 18958 11122 18977 11168
rect 18977 11122 19010 11168
rect 18958 11118 19010 11122
rect 20190 11259 20205 11282
rect 20205 11259 20242 11282
rect 20190 11230 20242 11259
rect 20302 11168 20354 11170
rect 20302 11122 20321 11168
rect 20321 11122 20354 11168
rect 20302 11118 20354 11122
rect 6534 10950 6794 11002
rect 11854 10950 12114 11002
rect 17174 10950 17434 11002
rect 22494 10950 22754 11002
rect 5406 10693 5458 10722
rect 5406 10670 5421 10693
rect 5421 10670 5458 10693
rect 5518 10670 5570 10722
rect 6078 10693 6130 10722
rect 6078 10670 6093 10693
rect 6093 10670 6130 10693
rect 6862 10830 6914 10834
rect 6862 10784 6881 10830
rect 6881 10784 6914 10830
rect 6862 10782 6914 10784
rect 6750 10558 6765 10610
rect 6765 10558 6802 10610
rect 6190 10334 6209 10386
rect 6209 10334 6242 10386
rect 7422 10558 7437 10610
rect 7437 10558 7474 10610
rect 7534 10558 7586 10610
rect 8094 10693 8146 10722
rect 8094 10670 8109 10693
rect 8109 10670 8146 10693
rect 8878 10558 8893 10610
rect 8893 10558 8930 10610
rect 8206 10334 8225 10386
rect 8225 10334 8258 10386
rect 8990 10334 9009 10386
rect 9009 10334 9042 10386
rect 9886 10558 9901 10610
rect 9901 10558 9938 10610
rect 10558 10558 10573 10610
rect 10573 10558 10610 10610
rect 9998 10334 10017 10386
rect 10017 10334 10050 10386
rect 11230 10558 11245 10610
rect 11245 10558 11282 10610
rect 10670 10334 10689 10386
rect 10689 10334 10722 10386
rect 12014 10558 12029 10610
rect 12029 10558 12066 10610
rect 11342 10334 11361 10386
rect 11361 10334 11394 10386
rect 12686 10558 12701 10610
rect 12701 10558 12738 10610
rect 12798 10558 12850 10610
rect 12126 10334 12145 10386
rect 12145 10334 12178 10386
rect 13358 10558 13373 10610
rect 13373 10558 13410 10610
rect 13470 10558 13522 10610
rect 14030 10558 14045 10610
rect 14045 10558 14082 10610
rect 14142 10558 14194 10610
rect 14702 10558 14717 10610
rect 14717 10558 14754 10610
rect 14814 10558 14866 10610
rect 15374 10558 15389 10610
rect 15389 10558 15426 10610
rect 15486 10558 15538 10610
rect 16046 10558 16061 10610
rect 16061 10558 16098 10610
rect 16718 10693 16770 10722
rect 16718 10670 16733 10693
rect 16733 10670 16770 10693
rect 16158 10334 16177 10386
rect 16177 10334 16210 10386
rect 17726 10693 17778 10722
rect 17726 10670 17741 10693
rect 17741 10670 17778 10693
rect 16830 10334 16849 10386
rect 16849 10334 16882 10386
rect 18398 10693 18450 10722
rect 18398 10670 18413 10693
rect 18413 10670 18450 10693
rect 17838 10334 17857 10386
rect 17857 10334 17890 10386
rect 19182 10830 19234 10834
rect 19182 10784 19201 10830
rect 19201 10784 19234 10830
rect 19182 10782 19234 10784
rect 19070 10693 19122 10722
rect 19070 10670 19085 10693
rect 19085 10670 19122 10693
rect 18510 10334 18529 10386
rect 18529 10334 18562 10386
rect 19854 10830 19906 10834
rect 19854 10784 19873 10830
rect 19873 10784 19906 10830
rect 19854 10782 19906 10784
rect 19742 10693 19794 10722
rect 19742 10670 19757 10693
rect 19757 10670 19794 10693
rect 20414 10693 20466 10722
rect 20414 10670 20429 10693
rect 20429 10670 20466 10693
rect 21086 10693 21138 10722
rect 21086 10670 21101 10693
rect 21101 10670 21138 10693
rect 20526 10334 20545 10386
rect 20545 10334 20578 10386
rect 21758 10693 21810 10722
rect 21758 10670 21773 10693
rect 21773 10670 21810 10693
rect 21870 10670 21922 10722
rect 21198 10334 21217 10386
rect 21217 10334 21250 10386
rect 3874 10166 4134 10218
rect 9194 10166 9454 10218
rect 14514 10166 14774 10218
rect 19834 10166 20094 10218
rect 4174 9774 4189 9826
rect 4189 9774 4226 9826
rect 4286 9774 4338 9826
rect 4846 9774 4861 9826
rect 4861 9774 4898 9826
rect 5854 9691 5869 9714
rect 5869 9691 5906 9714
rect 5854 9662 5906 9691
rect 4958 9600 5010 9602
rect 4958 9554 4977 9600
rect 4977 9554 5010 9600
rect 4958 9550 5010 9554
rect 6526 9691 6541 9714
rect 6541 9691 6578 9714
rect 6526 9662 6578 9691
rect 6638 9662 6690 9714
rect 5966 9600 6018 9602
rect 5966 9554 5985 9600
rect 5985 9554 6018 9600
rect 5966 9550 6018 9554
rect 7198 9691 7213 9714
rect 7213 9691 7250 9714
rect 7198 9662 7250 9691
rect 7310 9662 7362 9714
rect 7870 9774 7885 9826
rect 7885 9774 7922 9826
rect 8542 9774 8557 9826
rect 8557 9774 8594 9826
rect 7982 9600 8034 9602
rect 7982 9554 8001 9600
rect 8001 9554 8034 9600
rect 7982 9550 8034 9554
rect 9214 9774 9229 9826
rect 9229 9774 9266 9826
rect 8654 9600 8706 9602
rect 8654 9554 8673 9600
rect 8673 9554 8706 9600
rect 8654 9550 8706 9554
rect 9886 9691 9901 9714
rect 9901 9691 9938 9714
rect 9886 9662 9938 9691
rect 9326 9600 9378 9602
rect 9326 9554 9345 9600
rect 9345 9554 9378 9600
rect 9326 9550 9378 9554
rect 10558 9774 10573 9826
rect 10573 9774 10610 9826
rect 9998 9600 10050 9602
rect 9998 9554 10017 9600
rect 10017 9554 10050 9600
rect 9998 9550 10050 9554
rect 11566 9998 11585 10050
rect 11585 9998 11618 10050
rect 10670 9600 10722 9602
rect 10670 9554 10689 9600
rect 10689 9554 10722 9600
rect 10670 9550 10722 9554
rect 11454 9691 11469 9714
rect 11469 9691 11506 9714
rect 11454 9662 11506 9691
rect 12126 9774 12141 9826
rect 12141 9774 12178 9826
rect 12238 9774 12290 9826
rect 12798 9691 12813 9714
rect 12813 9691 12850 9714
rect 12798 9662 12850 9691
rect 12910 9662 12962 9714
rect 13694 9691 13709 9714
rect 13709 9691 13746 9714
rect 13694 9662 13746 9691
rect 13806 9662 13858 9714
rect 14366 9691 14381 9714
rect 14381 9691 14418 9714
rect 14366 9662 14418 9691
rect 14478 9774 14530 9826
rect 15038 9774 15053 9826
rect 15053 9774 15090 9826
rect 15710 9774 15725 9826
rect 15725 9774 15762 9826
rect 15150 9600 15202 9602
rect 15150 9554 15169 9600
rect 15169 9554 15202 9600
rect 15150 9550 15202 9554
rect 16382 9691 16397 9714
rect 16397 9691 16434 9714
rect 16382 9662 16434 9691
rect 15822 9600 15874 9602
rect 15822 9554 15841 9600
rect 15841 9554 15874 9600
rect 15822 9550 15874 9554
rect 17054 9691 17069 9714
rect 17069 9691 17106 9714
rect 17054 9662 17106 9691
rect 16494 9600 16546 9602
rect 16494 9554 16513 9600
rect 16513 9554 16546 9600
rect 16494 9550 16546 9554
rect 17166 9600 17218 9602
rect 17166 9554 17185 9600
rect 17185 9554 17218 9600
rect 17166 9550 17218 9554
rect 18510 9998 18529 10050
rect 18529 9998 18562 10050
rect 17838 9774 17875 9826
rect 17875 9774 17890 9826
rect 18398 9691 18413 9714
rect 18413 9691 18450 9714
rect 18398 9662 18450 9691
rect 17726 9600 17778 9602
rect 17726 9554 17759 9600
rect 17759 9554 17778 9600
rect 17726 9550 17778 9554
rect 19070 9774 19085 9826
rect 19085 9774 19122 9826
rect 19742 9774 19757 9826
rect 19757 9774 19794 9826
rect 19182 9600 19234 9602
rect 19182 9554 19201 9600
rect 19201 9554 19234 9600
rect 19182 9550 19234 9554
rect 20526 9998 20545 10050
rect 20545 9998 20578 10050
rect 20414 9774 20429 9826
rect 20429 9774 20466 9826
rect 19854 9600 19906 9602
rect 19854 9554 19873 9600
rect 19873 9554 19906 9600
rect 19854 9550 19906 9554
rect 21758 9998 21777 10050
rect 21777 9998 21810 10050
rect 21646 9774 21661 9826
rect 21661 9774 21698 9826
rect 6534 9382 6794 9434
rect 11854 9382 12114 9434
rect 17174 9382 17434 9434
rect 22494 9382 22754 9434
rect 3390 9125 3442 9154
rect 3390 9102 3405 9125
rect 3405 9102 3442 9125
rect 3502 9102 3554 9154
rect 4062 9125 4114 9154
rect 4062 9102 4077 9125
rect 4077 9102 4114 9125
rect 4846 9262 4898 9266
rect 4846 9216 4865 9262
rect 4865 9216 4898 9262
rect 4846 9214 4898 9216
rect 4734 8990 4749 9042
rect 4749 8990 4786 9042
rect 4174 8766 4193 8818
rect 4193 8766 4226 8818
rect 5406 8990 5421 9042
rect 5421 8990 5458 9042
rect 6078 8990 6093 9042
rect 6093 8990 6130 9042
rect 6190 8990 6242 9042
rect 5518 8766 5537 8818
rect 5537 8766 5570 8818
rect 6750 8990 6765 9042
rect 6765 8990 6802 9042
rect 6862 8990 6914 9042
rect 7422 9125 7474 9154
rect 7422 9102 7437 9125
rect 7437 9102 7474 9125
rect 7534 9102 7586 9154
rect 8206 9125 8258 9154
rect 8206 9102 8221 9125
rect 8221 9102 8258 9125
rect 8990 9262 9042 9266
rect 8990 9216 9009 9262
rect 9009 9216 9042 9262
rect 8990 9214 9042 9216
rect 8878 8990 8893 9042
rect 8893 8990 8930 9042
rect 8318 8766 8337 8818
rect 8337 8766 8370 8818
rect 10334 9125 10386 9154
rect 10334 9102 10349 9125
rect 10349 9102 10386 9125
rect 11006 8990 11021 9042
rect 11021 8990 11058 9042
rect 10446 8883 10498 8930
rect 10446 8878 10465 8883
rect 10465 8878 10498 8883
rect 11678 8990 11693 9042
rect 11693 8990 11730 9042
rect 11118 8766 11137 8818
rect 11137 8766 11170 8818
rect 12350 9125 12402 9154
rect 12350 9102 12365 9125
rect 12365 9102 12402 9125
rect 11790 8766 11809 8818
rect 11809 8766 11842 8818
rect 13022 9125 13074 9154
rect 13022 9102 13037 9125
rect 13037 9102 13074 9125
rect 12462 8766 12481 8818
rect 12481 8766 12514 8818
rect 13694 8990 13709 9042
rect 13709 8990 13746 9042
rect 13134 8766 13153 8818
rect 13153 8766 13186 8818
rect 14478 9262 14530 9266
rect 14478 9216 14497 9262
rect 14497 9216 14530 9262
rect 14478 9214 14530 9216
rect 14366 8990 14381 9042
rect 14381 8990 14418 9042
rect 13806 8766 13825 8818
rect 13825 8766 13858 8818
rect 15150 9262 15202 9266
rect 15150 9216 15169 9262
rect 15169 9216 15202 9262
rect 15150 9214 15202 9216
rect 15038 8990 15053 9042
rect 15053 8990 15090 9042
rect 15710 9125 15762 9154
rect 15710 9102 15725 9125
rect 15725 9102 15762 9125
rect 16382 8990 16397 9042
rect 16397 8990 16434 9042
rect 15822 8766 15841 8818
rect 15841 8766 15874 8818
rect 16494 8766 16513 8818
rect 16513 8766 16546 8818
rect 17726 9125 17778 9154
rect 17726 9102 17741 9125
rect 17741 9102 17778 9125
rect 18398 8990 18413 9042
rect 18413 8990 18450 9042
rect 17838 8766 17857 8818
rect 17857 8766 17890 8818
rect 19070 9125 19122 9154
rect 19070 9102 19085 9125
rect 19085 9102 19122 9125
rect 18510 8766 18529 8818
rect 18529 8766 18562 8818
rect 19854 9262 19906 9266
rect 19854 9216 19873 9262
rect 19873 9216 19906 9262
rect 19854 9214 19906 9216
rect 19742 8990 19757 9042
rect 19757 8990 19794 9042
rect 19182 8766 19201 8818
rect 19201 8766 19234 8818
rect 20526 9262 20578 9266
rect 20526 9216 20545 9262
rect 20545 9216 20578 9262
rect 20526 9214 20578 9216
rect 20414 9125 20466 9154
rect 20414 9102 20429 9125
rect 20429 9102 20466 9125
rect 3874 8598 4134 8650
rect 9194 8598 9454 8650
rect 14514 8598 14774 8650
rect 19834 8598 20094 8650
rect 2942 8123 2979 8146
rect 2979 8123 2994 8146
rect 2942 8094 2994 8123
rect 3502 8123 3517 8146
rect 3517 8123 3554 8146
rect 3502 8094 3554 8123
rect 2830 8032 2882 8034
rect 2830 7986 2863 8032
rect 2863 7986 2882 8032
rect 2830 7982 2882 7986
rect 4174 8123 4189 8146
rect 4189 8123 4226 8146
rect 4174 8094 4226 8123
rect 3614 8032 3666 8034
rect 3614 7986 3633 8032
rect 3633 7986 3666 8032
rect 3614 7982 3666 7986
rect 4958 8430 4977 8482
rect 4977 8430 5010 8482
rect 4846 8123 4861 8146
rect 4861 8123 4898 8146
rect 4846 8094 4898 8123
rect 4286 8032 4338 8034
rect 4286 7986 4305 8032
rect 4305 7986 4338 8032
rect 4286 7982 4338 7986
rect 5966 8430 5985 8482
rect 5985 8430 6018 8482
rect 5854 8123 5869 8146
rect 5869 8123 5906 8146
rect 5854 8094 5906 8123
rect 6638 8430 6657 8482
rect 6657 8430 6690 8482
rect 6526 8206 6541 8258
rect 6541 8206 6578 8258
rect 7198 8206 7213 8258
rect 7213 8206 7250 8258
rect 7870 8206 7885 8258
rect 7885 8206 7922 8258
rect 7310 8032 7362 8034
rect 7310 7986 7329 8032
rect 7329 7986 7362 8032
rect 7310 7982 7362 7986
rect 8542 8123 8557 8146
rect 8557 8123 8594 8146
rect 8542 8094 8594 8123
rect 7982 8032 8034 8034
rect 7982 7986 8001 8032
rect 8001 7986 8034 8032
rect 7982 7982 8034 7986
rect 9326 8430 9345 8482
rect 9345 8430 9378 8482
rect 9214 8206 9229 8258
rect 9229 8206 9266 8258
rect 8654 8032 8706 8034
rect 8654 7986 8673 8032
rect 8673 7986 8706 8032
rect 8654 7982 8706 7986
rect 9998 8430 10017 8482
rect 10017 8430 10050 8482
rect 9886 8206 9901 8258
rect 9901 8206 9938 8258
rect 10670 8430 10689 8482
rect 10689 8430 10722 8482
rect 10558 8206 10573 8258
rect 10573 8206 10610 8258
rect 11230 8365 11263 8370
rect 11263 8365 11282 8370
rect 11230 8318 11282 8365
rect 11342 8123 11379 8146
rect 11379 8123 11394 8146
rect 11342 8094 11394 8123
rect 12126 8206 12141 8258
rect 12141 8206 12178 8258
rect 12238 8206 12290 8258
rect 12798 8123 12813 8146
rect 12813 8123 12850 8146
rect 12798 8094 12850 8123
rect 12910 8206 12962 8258
rect 13694 8206 13709 8258
rect 13709 8206 13746 8258
rect 13806 8206 13858 8258
rect 14366 8206 14381 8258
rect 14381 8206 14418 8258
rect 15150 8430 15169 8482
rect 15169 8430 15202 8482
rect 14478 8206 14530 8258
rect 15038 8206 15053 8258
rect 15053 8206 15090 8258
rect 15710 8123 15725 8146
rect 15725 8123 15762 8146
rect 15710 8094 15762 8123
rect 15822 8206 15874 8258
rect 16382 8123 16397 8146
rect 16397 8123 16434 8146
rect 16382 8094 16434 8123
rect 17166 8430 17185 8482
rect 17185 8430 17218 8482
rect 16494 8206 16546 8258
rect 17054 8206 17069 8258
rect 17069 8206 17106 8258
rect 17838 8430 17857 8482
rect 17857 8430 17890 8482
rect 17726 8123 17741 8146
rect 17741 8123 17778 8146
rect 17726 8094 17778 8123
rect 18510 8430 18529 8482
rect 18529 8430 18562 8482
rect 18398 8206 18413 8258
rect 18413 8206 18450 8258
rect 19182 8430 19201 8482
rect 19201 8430 19234 8482
rect 19070 8206 19085 8258
rect 19085 8206 19122 8258
rect 19742 8206 19757 8258
rect 19757 8206 19794 8258
rect 19854 8206 19906 8258
rect 20526 8123 20563 8146
rect 20563 8123 20578 8146
rect 20526 8094 20578 8123
rect 20414 8032 20466 8034
rect 20414 7986 20447 8032
rect 20447 7986 20466 8032
rect 20414 7982 20466 7986
rect 6534 7814 6794 7866
rect 11854 7814 12114 7866
rect 17174 7814 17434 7866
rect 22494 7814 22754 7866
rect 2158 7422 2195 7474
rect 2195 7422 2210 7474
rect 2718 7422 2733 7474
rect 2733 7422 2770 7474
rect 2046 7198 2079 7250
rect 2079 7198 2098 7250
rect 3390 7422 3405 7474
rect 3405 7422 3442 7474
rect 2830 7198 2849 7250
rect 2849 7198 2882 7250
rect 4062 7422 4077 7474
rect 4077 7422 4114 7474
rect 3502 7198 3521 7250
rect 3521 7198 3554 7250
rect 4734 7557 4786 7586
rect 4734 7534 4749 7557
rect 4749 7534 4786 7557
rect 4846 7422 4898 7474
rect 4174 7198 4193 7250
rect 4193 7198 4226 7250
rect 5406 7422 5421 7474
rect 5421 7422 5458 7474
rect 6190 7694 6242 7698
rect 6190 7648 6209 7694
rect 6209 7648 6242 7694
rect 6190 7646 6242 7648
rect 6078 7422 6093 7474
rect 6093 7422 6130 7474
rect 5518 7198 5537 7250
rect 5537 7198 5570 7250
rect 6862 7694 6914 7698
rect 6862 7648 6881 7694
rect 6881 7648 6914 7694
rect 6862 7646 6914 7648
rect 6750 7422 6765 7474
rect 6765 7422 6802 7474
rect 7422 7422 7437 7474
rect 7437 7422 7474 7474
rect 8206 7422 8221 7474
rect 8221 7422 8258 7474
rect 7534 7198 7553 7250
rect 7553 7198 7586 7250
rect 8990 7694 9042 7698
rect 8990 7648 9009 7694
rect 9009 7648 9042 7694
rect 8990 7646 9042 7648
rect 8878 7422 8893 7474
rect 8893 7422 8930 7474
rect 8318 7198 8337 7250
rect 8337 7198 8370 7250
rect 9998 7694 10050 7698
rect 9998 7648 10017 7694
rect 10017 7648 10050 7694
rect 9998 7646 10050 7648
rect 9886 7422 9901 7474
rect 9901 7422 9938 7474
rect 10670 7694 10722 7698
rect 10670 7648 10689 7694
rect 10689 7648 10722 7694
rect 10670 7646 10722 7648
rect 10558 7557 10610 7586
rect 10558 7534 10573 7557
rect 10573 7534 10610 7557
rect 11230 7694 11282 7698
rect 11230 7648 11263 7694
rect 11263 7648 11282 7694
rect 11230 7646 11282 7648
rect 11342 7422 11379 7474
rect 11379 7422 11394 7474
rect 11902 7422 11917 7474
rect 11917 7422 11954 7474
rect 12574 7422 12589 7474
rect 12589 7422 12626 7474
rect 12014 7198 12033 7250
rect 12033 7198 12066 7250
rect 13358 7694 13410 7698
rect 13358 7648 13377 7694
rect 13377 7648 13410 7694
rect 13358 7646 13410 7648
rect 13246 7422 13261 7474
rect 13261 7422 13298 7474
rect 12686 7198 12705 7250
rect 12705 7198 12738 7250
rect 13918 7557 13970 7586
rect 13918 7534 13933 7557
rect 13933 7534 13970 7557
rect 14702 7694 14754 7698
rect 14702 7648 14721 7694
rect 14721 7648 14754 7694
rect 14702 7646 14754 7648
rect 14590 7422 14605 7474
rect 14605 7422 14642 7474
rect 14030 7315 14082 7362
rect 14030 7310 14049 7315
rect 14049 7310 14082 7315
rect 15262 7557 15314 7586
rect 15262 7534 15277 7557
rect 15277 7534 15314 7557
rect 15934 7557 15986 7586
rect 15934 7534 15949 7557
rect 15949 7534 15986 7557
rect 15374 7198 15393 7250
rect 15393 7198 15426 7250
rect 16718 7694 16770 7698
rect 16718 7648 16737 7694
rect 16737 7648 16770 7694
rect 16718 7646 16770 7648
rect 16606 7422 16621 7474
rect 16621 7422 16658 7474
rect 16046 7198 16065 7250
rect 16065 7198 16098 7250
rect 17838 7694 17890 7698
rect 17838 7648 17857 7694
rect 17857 7648 17890 7694
rect 17838 7646 17890 7648
rect 17726 7422 17741 7474
rect 17741 7422 17778 7474
rect 18510 7694 18562 7698
rect 18510 7648 18529 7694
rect 18529 7648 18562 7694
rect 18510 7646 18562 7648
rect 18398 7422 18413 7474
rect 18413 7422 18450 7474
rect 19070 7422 19085 7474
rect 19085 7422 19122 7474
rect 19742 7422 19757 7474
rect 19757 7422 19794 7474
rect 19182 7198 19201 7250
rect 19201 7198 19234 7250
rect 20414 7422 20429 7474
rect 20429 7422 20466 7474
rect 19854 7198 19873 7250
rect 19873 7198 19906 7250
rect 21086 7422 21101 7474
rect 21101 7422 21138 7474
rect 20526 7198 20545 7250
rect 20545 7198 20578 7250
rect 21198 7198 21217 7250
rect 21217 7198 21250 7250
rect 3874 7030 4134 7082
rect 9194 7030 9454 7082
rect 14514 7030 14774 7082
rect 19834 7030 20094 7082
rect 2158 6555 2173 6578
rect 2173 6555 2210 6578
rect 2158 6526 2210 6555
rect 2830 6555 2845 6578
rect 2845 6555 2882 6578
rect 2830 6526 2882 6555
rect 2270 6464 2322 6466
rect 2270 6418 2289 6464
rect 2289 6418 2322 6464
rect 2270 6414 2322 6418
rect 3502 6555 3517 6578
rect 3517 6555 3554 6578
rect 3502 6526 3554 6555
rect 2942 6464 2994 6466
rect 2942 6418 2961 6464
rect 2961 6418 2994 6464
rect 2942 6414 2994 6418
rect 4286 6862 4305 6914
rect 4305 6862 4338 6914
rect 4174 6555 4189 6578
rect 4189 6555 4226 6578
rect 4174 6526 4226 6555
rect 3614 6464 3666 6466
rect 3614 6418 3633 6464
rect 3633 6418 3666 6464
rect 3614 6414 3666 6418
rect 4958 6862 4977 6914
rect 4977 6862 5010 6914
rect 4846 6555 4861 6578
rect 4861 6555 4898 6578
rect 4846 6526 4898 6555
rect 5742 6638 5757 6690
rect 5757 6638 5794 6690
rect 5854 6638 5906 6690
rect 6414 6638 6429 6690
rect 6429 6638 6466 6690
rect 6526 6638 6578 6690
rect 7086 6555 7101 6578
rect 7101 6555 7138 6578
rect 7086 6526 7138 6555
rect 7758 6555 7773 6578
rect 7773 6555 7810 6578
rect 7758 6526 7810 6555
rect 7198 6464 7250 6466
rect 7198 6418 7217 6464
rect 7217 6418 7250 6464
rect 7198 6414 7250 6418
rect 8430 6555 8445 6578
rect 8445 6555 8482 6578
rect 8430 6526 8482 6555
rect 8542 6638 8594 6690
rect 7870 6464 7922 6466
rect 7870 6418 7889 6464
rect 7889 6418 7922 6464
rect 7870 6414 7922 6418
rect 9102 6555 9117 6578
rect 9117 6555 9154 6578
rect 9102 6526 9154 6555
rect 9214 6638 9266 6690
rect 9774 6638 9789 6690
rect 9789 6638 9826 6690
rect 10558 6862 10577 6914
rect 10577 6862 10610 6914
rect 10446 6638 10461 6690
rect 10461 6638 10498 6690
rect 9886 6464 9938 6466
rect 9886 6418 9905 6464
rect 9905 6418 9938 6464
rect 9886 6414 9938 6418
rect 11230 6862 11249 6914
rect 11249 6862 11282 6914
rect 11118 6638 11133 6690
rect 11133 6638 11170 6690
rect 11790 6638 11805 6690
rect 11805 6638 11842 6690
rect 12462 6638 12477 6690
rect 12477 6638 12514 6690
rect 11902 6464 11954 6466
rect 11902 6418 11921 6464
rect 11921 6418 11954 6464
rect 11902 6414 11954 6418
rect 12574 6464 12626 6466
rect 12574 6418 12593 6464
rect 12593 6418 12626 6464
rect 12574 6414 12626 6418
rect 14254 6862 14273 6914
rect 14273 6862 14306 6914
rect 14142 6638 14157 6690
rect 14157 6638 14194 6690
rect 14926 6862 14945 6914
rect 14945 6862 14978 6914
rect 14814 6638 14829 6690
rect 14829 6638 14866 6690
rect 15598 6862 15617 6914
rect 15617 6862 15650 6914
rect 15486 6638 15501 6690
rect 15501 6638 15538 6690
rect 16158 6555 16173 6578
rect 16173 6555 16210 6578
rect 16158 6526 16210 6555
rect 16270 6526 16322 6578
rect 16830 6555 16845 6578
rect 16845 6555 16882 6578
rect 16830 6526 16882 6555
rect 17614 6862 17633 6914
rect 17633 6862 17666 6914
rect 16942 6526 16994 6578
rect 17502 6555 17517 6578
rect 17517 6555 17554 6578
rect 17502 6526 17554 6555
rect 18174 6555 18189 6578
rect 18189 6555 18226 6578
rect 18174 6526 18226 6555
rect 18846 6555 18861 6578
rect 18861 6555 18898 6578
rect 18846 6526 18898 6555
rect 19630 6862 19649 6914
rect 19649 6862 19682 6914
rect 18958 6638 19010 6690
rect 18286 6464 18338 6466
rect 18286 6418 18305 6464
rect 18305 6418 18338 6464
rect 18286 6414 18338 6418
rect 19518 6555 19533 6578
rect 19533 6555 19570 6578
rect 19518 6526 19570 6555
rect 20302 6555 20339 6578
rect 20339 6555 20354 6578
rect 20302 6526 20354 6555
rect 20190 6464 20242 6466
rect 20190 6418 20223 6464
rect 20223 6418 20242 6464
rect 20190 6414 20242 6418
rect 21646 6638 21661 6690
rect 21661 6638 21698 6690
rect 21758 6464 21810 6466
rect 21758 6418 21777 6464
rect 21777 6418 21810 6464
rect 21758 6414 21810 6418
rect 6534 6246 6794 6298
rect 11854 6246 12114 6298
rect 17174 6246 17434 6298
rect 22494 6246 22754 6298
rect 2046 5854 2061 5906
rect 2061 5854 2098 5906
rect 2718 5854 2733 5906
rect 2733 5854 2770 5906
rect 2158 5630 2177 5682
rect 2177 5630 2210 5682
rect 3390 5854 3405 5906
rect 3405 5854 3442 5906
rect 2830 5630 2849 5682
rect 2849 5630 2882 5682
rect 4062 5854 4077 5906
rect 4077 5854 4114 5906
rect 3502 5630 3521 5682
rect 3521 5630 3554 5682
rect 4734 5854 4749 5906
rect 4749 5854 4786 5906
rect 4174 5630 4193 5682
rect 4193 5630 4226 5682
rect 5518 6126 5570 6130
rect 5518 6080 5537 6126
rect 5537 6080 5570 6126
rect 5518 6078 5570 6080
rect 5406 5854 5421 5906
rect 5421 5854 5458 5906
rect 4846 5630 4865 5682
rect 4865 5630 4898 5682
rect 6190 6126 6242 6130
rect 6190 6080 6209 6126
rect 6209 6080 6242 6126
rect 6190 6078 6242 6080
rect 6078 5854 6093 5906
rect 6093 5854 6130 5906
rect 6750 5989 6802 6018
rect 6750 5966 6765 5989
rect 6765 5966 6802 5989
rect 6862 5966 6914 6018
rect 7422 5989 7474 6018
rect 7422 5966 7437 5989
rect 7437 5966 7474 5989
rect 8094 5989 8146 6018
rect 8094 5966 8109 5989
rect 8109 5966 8146 5989
rect 7534 5630 7553 5682
rect 7553 5630 7586 5682
rect 8878 6126 8930 6130
rect 8878 6080 8897 6126
rect 8897 6080 8930 6126
rect 8878 6078 8930 6080
rect 8766 5989 8818 6018
rect 8766 5966 8781 5989
rect 8781 5966 8818 5989
rect 8206 5630 8225 5682
rect 8225 5630 8258 5682
rect 9886 6126 9938 6130
rect 9886 6080 9905 6126
rect 9905 6080 9938 6126
rect 9886 6078 9938 6080
rect 9774 5854 9789 5906
rect 9789 5854 9826 5906
rect 10558 6126 10610 6130
rect 10558 6080 10577 6126
rect 10577 6080 10610 6126
rect 10558 6078 10610 6080
rect 10446 5854 10461 5906
rect 10461 5854 10498 5906
rect 11230 6126 11282 6130
rect 11230 6080 11249 6126
rect 11249 6080 11282 6126
rect 11230 6078 11282 6080
rect 11118 5989 11170 6018
rect 11118 5966 11133 5989
rect 11133 5966 11170 5989
rect 11902 6126 11954 6130
rect 11902 6080 11921 6126
rect 11921 6080 11954 6126
rect 11902 6078 11954 6080
rect 11790 5989 11842 6018
rect 11790 5966 11805 5989
rect 11805 5966 11842 5989
rect 12574 5989 12626 6018
rect 12574 5966 12589 5989
rect 12589 5966 12626 5989
rect 13358 6126 13410 6130
rect 13358 6080 13377 6126
rect 13377 6080 13410 6126
rect 13358 6078 13410 6080
rect 13246 5854 13261 5906
rect 13261 5854 13298 5906
rect 12686 5630 12705 5682
rect 12705 5630 12738 5682
rect 14030 6126 14082 6130
rect 14030 6080 14049 6126
rect 14049 6080 14082 6126
rect 14030 6078 14082 6080
rect 13918 5854 13933 5906
rect 13933 5854 13970 5906
rect 14702 6126 14754 6130
rect 14702 6080 14721 6126
rect 14721 6080 14754 6126
rect 14702 6078 14754 6080
rect 14590 5989 14642 6018
rect 14590 5966 14605 5989
rect 14605 5966 14642 5989
rect 15374 6126 15426 6130
rect 15374 6080 15393 6126
rect 15393 6080 15426 6126
rect 15374 6078 15426 6080
rect 15262 5989 15314 6018
rect 15262 5966 15277 5989
rect 15277 5966 15314 5989
rect 16046 6126 16098 6130
rect 16046 6080 16065 6126
rect 16065 6080 16098 6126
rect 16046 6078 16098 6080
rect 15934 5989 15986 6018
rect 15934 5966 15949 5989
rect 15949 5966 15986 5989
rect 16718 6126 16770 6130
rect 16718 6080 16737 6126
rect 16737 6080 16770 6126
rect 16718 6078 16770 6080
rect 16606 5989 16658 6018
rect 16606 5966 16621 5989
rect 16621 5966 16658 5989
rect 17726 5854 17741 5906
rect 17741 5854 17778 5906
rect 18398 5854 18413 5906
rect 18413 5854 18450 5906
rect 19070 5989 19122 6018
rect 19070 5966 19085 5989
rect 19085 5966 19122 5989
rect 17838 5630 17857 5682
rect 17857 5630 17890 5682
rect 18510 5747 18562 5794
rect 19742 5989 19794 6018
rect 19742 5966 19757 5989
rect 19757 5966 19794 5989
rect 18510 5742 18529 5747
rect 18529 5742 18562 5747
rect 19182 5747 19234 5794
rect 19182 5742 19201 5747
rect 19201 5742 19234 5747
rect 20414 5854 20429 5906
rect 20429 5854 20466 5906
rect 19854 5630 19873 5682
rect 19873 5630 19906 5682
rect 21086 5854 21101 5906
rect 21101 5854 21138 5906
rect 20526 5630 20545 5682
rect 20545 5630 20578 5682
rect 21198 5630 21217 5682
rect 21217 5630 21250 5682
rect 21870 5854 21907 5906
rect 21907 5854 21922 5906
rect 21758 5630 21791 5682
rect 21791 5630 21810 5682
rect 3874 5462 4134 5514
rect 9194 5462 9454 5514
rect 14514 5462 14774 5514
rect 19834 5462 20094 5514
rect 2158 4987 2173 5010
rect 2173 4987 2210 5010
rect 2158 4958 2210 4987
rect 2830 4987 2845 5010
rect 2845 4987 2882 5010
rect 2830 4958 2882 4987
rect 2270 4896 2322 4898
rect 2270 4850 2289 4896
rect 2289 4850 2322 4896
rect 2270 4846 2322 4850
rect 3502 4987 3517 5010
rect 3517 4987 3554 5010
rect 3502 4958 3554 4987
rect 3614 4958 3666 5010
rect 2942 4896 2994 4898
rect 2942 4850 2961 4896
rect 2961 4850 2994 4896
rect 2942 4846 2994 4850
rect 4174 5070 4189 5122
rect 4189 5070 4226 5122
rect 4846 5070 4861 5122
rect 4861 5070 4898 5122
rect 4286 4896 4338 4898
rect 4286 4850 4305 4896
rect 4305 4850 4338 4896
rect 4286 4846 4338 4850
rect 5854 5294 5873 5346
rect 5873 5294 5906 5346
rect 5742 4987 5757 5010
rect 5757 4987 5794 5010
rect 5742 4958 5794 4987
rect 4958 4896 5010 4898
rect 4958 4850 4977 4896
rect 4977 4850 5010 4896
rect 4958 4846 5010 4850
rect 6526 5294 6545 5346
rect 6545 5294 6578 5346
rect 6414 4987 6429 5010
rect 6429 4987 6466 5010
rect 6414 4958 6466 4987
rect 7198 5294 7217 5346
rect 7217 5294 7250 5346
rect 7086 5070 7101 5122
rect 7101 5070 7138 5122
rect 7758 5070 7773 5122
rect 7773 5070 7810 5122
rect 8542 5294 8561 5346
rect 8561 5294 8594 5346
rect 7870 5070 7922 5122
rect 8430 5070 8445 5122
rect 8445 5070 8482 5122
rect 9102 5070 9117 5122
rect 9117 5070 9154 5122
rect 9886 5294 9905 5346
rect 9905 5294 9938 5346
rect 9214 5070 9266 5122
rect 9774 4987 9789 5010
rect 9789 4987 9826 5010
rect 9774 4958 9826 4987
rect 10558 5294 10577 5346
rect 10577 5294 10610 5346
rect 10446 5070 10461 5122
rect 10461 5070 10498 5122
rect 11454 5070 11469 5122
rect 11469 5070 11506 5122
rect 11566 5070 11618 5122
rect 12126 4987 12141 5010
rect 12141 4987 12178 5010
rect 12126 4958 12178 4987
rect 12798 4987 12813 5010
rect 12813 4987 12850 5010
rect 12798 4958 12850 4987
rect 12238 4896 12290 4898
rect 12238 4850 12257 4896
rect 12257 4850 12290 4896
rect 12238 4846 12290 4850
rect 14142 5294 14161 5346
rect 14161 5294 14194 5346
rect 12910 4896 12962 4898
rect 12910 4850 12929 4896
rect 12929 4850 12962 4896
rect 12910 4846 12962 4850
rect 14030 4987 14045 5010
rect 14045 4987 14082 5010
rect 14030 4958 14082 4987
rect 14814 5294 14833 5346
rect 14833 5294 14866 5346
rect 14702 4987 14717 5010
rect 14717 4987 14754 5010
rect 14702 4958 14754 4987
rect 15486 5294 15505 5346
rect 15505 5294 15538 5346
rect 15374 5070 15389 5122
rect 15389 5070 15426 5122
rect 16046 4987 16061 5010
rect 16061 4987 16098 5010
rect 16046 4958 16098 4987
rect 16718 4987 16733 5010
rect 16733 4987 16770 5010
rect 16718 4958 16770 4987
rect 16830 5070 16882 5122
rect 16158 4896 16210 4898
rect 16158 4850 16177 4896
rect 16177 4850 16210 4896
rect 16158 4846 16210 4850
rect 17390 5070 17405 5122
rect 17405 5070 17442 5122
rect 18174 5294 18193 5346
rect 18193 5294 18226 5346
rect 18062 5070 18077 5122
rect 18077 5070 18114 5122
rect 17502 4896 17554 4898
rect 17502 4850 17521 4896
rect 17521 4850 17554 4896
rect 17502 4846 17554 4850
rect 18734 5070 18749 5122
rect 18749 5070 18786 5122
rect 19518 5229 19537 5234
rect 19537 5229 19570 5234
rect 19518 5182 19570 5229
rect 20190 5294 20209 5346
rect 20209 5294 20242 5346
rect 18846 5070 18898 5122
rect 19406 5070 19421 5122
rect 19421 5070 19458 5122
rect 20078 5070 20093 5122
rect 20093 5070 20130 5122
rect 20750 4987 20765 5010
rect 20765 4987 20802 5010
rect 20750 4958 20802 4987
rect 21646 4987 21661 5010
rect 21661 4987 21698 5010
rect 21646 4958 21698 4987
rect 20862 4896 20914 4898
rect 20862 4850 20881 4896
rect 20881 4850 20914 4896
rect 20862 4846 20914 4850
rect 21758 4896 21810 4898
rect 21758 4850 21777 4896
rect 21777 4850 21810 4896
rect 21758 4846 21810 4850
rect 6534 4678 6794 4730
rect 11854 4678 12114 4730
rect 17174 4678 17434 4730
rect 22494 4678 22754 4730
rect 2382 4421 2434 4450
rect 2382 4398 2397 4421
rect 2397 4398 2434 4421
rect 2494 4286 2546 4338
rect 3054 4286 3069 4338
rect 3069 4286 3106 4338
rect 3838 4558 3890 4562
rect 3838 4512 3857 4558
rect 3857 4512 3890 4558
rect 3838 4510 3890 4512
rect 3166 4286 3218 4338
rect 3726 4286 3741 4338
rect 3741 4286 3778 4338
rect 4510 4558 4562 4562
rect 4510 4512 4529 4558
rect 4529 4512 4562 4558
rect 4510 4510 4562 4512
rect 4398 4286 4413 4338
rect 4413 4286 4450 4338
rect 5070 4421 5122 4450
rect 5070 4398 5085 4421
rect 5085 4398 5122 4421
rect 5742 4421 5794 4450
rect 5742 4398 5757 4421
rect 5757 4398 5794 4421
rect 5182 4062 5201 4114
rect 5201 4062 5234 4114
rect 6414 4286 6429 4338
rect 6429 4286 6466 4338
rect 5854 4062 5873 4114
rect 5873 4062 5906 4114
rect 7198 4558 7250 4562
rect 7198 4512 7217 4558
rect 7217 4512 7250 4558
rect 7198 4510 7250 4512
rect 7086 4286 7101 4338
rect 7101 4286 7138 4338
rect 6526 4062 6545 4114
rect 6545 4062 6578 4114
rect 7758 4286 7773 4338
rect 7773 4286 7810 4338
rect 8542 4558 8594 4562
rect 8542 4512 8561 4558
rect 8561 4512 8594 4558
rect 8542 4510 8594 4512
rect 8430 4421 8482 4450
rect 8430 4398 8445 4421
rect 8445 4398 8482 4421
rect 7870 4062 7889 4114
rect 7889 4062 7922 4114
rect 9774 4421 9826 4450
rect 9774 4398 9789 4421
rect 9789 4398 9826 4421
rect 10446 4421 10498 4450
rect 10446 4398 10461 4421
rect 10461 4398 10498 4421
rect 9886 4062 9905 4114
rect 9905 4062 9938 4114
rect 11118 4286 11133 4338
rect 11133 4286 11170 4338
rect 10558 4062 10577 4114
rect 10577 4062 10610 4114
rect 11230 4062 11249 4114
rect 11249 4062 11282 4114
rect 12350 4286 12365 4338
rect 12365 4286 12402 4338
rect 13022 4286 13037 4338
rect 13037 4286 13074 4338
rect 12462 4062 12481 4114
rect 12481 4062 12514 4114
rect 13694 4286 13709 4338
rect 13709 4286 13746 4338
rect 13134 4062 13153 4114
rect 13153 4062 13186 4114
rect 14366 4421 14418 4450
rect 14366 4398 14381 4421
rect 14381 4398 14418 4421
rect 15150 4558 15202 4562
rect 15150 4512 15169 4558
rect 15169 4512 15202 4558
rect 15150 4510 15202 4512
rect 14478 4286 14530 4338
rect 13806 4062 13825 4114
rect 13825 4062 13858 4114
rect 15038 4286 15053 4338
rect 15053 4286 15090 4338
rect 15822 4558 15874 4562
rect 15822 4512 15841 4558
rect 15841 4512 15874 4558
rect 15822 4510 15874 4512
rect 15710 4286 15725 4338
rect 15725 4286 15762 4338
rect 16382 4421 16434 4450
rect 16382 4398 16397 4421
rect 16397 4398 16434 4421
rect 16494 4398 16546 4450
rect 17838 4558 17890 4562
rect 17838 4512 17857 4558
rect 17857 4512 17890 4558
rect 17838 4510 17890 4512
rect 17726 4421 17778 4450
rect 17726 4398 17741 4421
rect 17741 4398 17778 4421
rect 18510 4558 18562 4562
rect 18510 4512 18529 4558
rect 18529 4512 18562 4558
rect 18510 4510 18562 4512
rect 18398 4421 18450 4450
rect 18398 4398 18413 4421
rect 18413 4398 18450 4421
rect 19070 4421 19122 4450
rect 19070 4398 19085 4421
rect 19085 4398 19122 4421
rect 19854 4558 19906 4562
rect 19854 4512 19873 4558
rect 19873 4512 19906 4558
rect 19854 4510 19906 4512
rect 19742 4286 19757 4338
rect 19757 4286 19794 4338
rect 19182 4062 19201 4114
rect 19201 4062 19234 4114
rect 20526 4558 20578 4562
rect 20526 4512 20545 4558
rect 20545 4512 20578 4558
rect 20526 4510 20578 4512
rect 20414 4421 20466 4450
rect 20414 4398 20429 4421
rect 20429 4398 20466 4421
rect 21198 4558 21250 4562
rect 21198 4512 21217 4558
rect 21217 4512 21250 4558
rect 21198 4510 21250 4512
rect 21086 4421 21138 4450
rect 21086 4398 21101 4421
rect 21101 4398 21138 4421
rect 21870 4286 21907 4338
rect 21907 4286 21922 4338
rect 21758 4062 21791 4114
rect 21791 4062 21810 4114
rect 3874 3894 4134 3946
rect 9194 3894 9454 3946
rect 14514 3894 14774 3946
rect 19834 3894 20094 3946
rect 2942 3726 2961 3778
rect 2961 3726 2994 3778
rect 2830 3502 2845 3554
rect 2845 3502 2882 3554
rect 3614 3726 3633 3778
rect 3633 3726 3666 3778
rect 3502 3502 3517 3554
rect 3517 3502 3554 3554
rect 4286 3726 4305 3778
rect 4305 3726 4338 3778
rect 4174 3502 4189 3554
rect 4189 3502 4226 3554
rect 4958 3726 4977 3778
rect 4977 3726 5010 3778
rect 4846 3419 4861 3442
rect 4861 3419 4898 3442
rect 4846 3390 4898 3419
rect 6414 3726 6447 3778
rect 6447 3726 6466 3778
rect 5742 3390 5794 3442
rect 5854 3502 5891 3554
rect 5891 3502 5906 3554
rect 7086 3726 7119 3778
rect 7119 3726 7138 3778
rect 6526 3502 6563 3554
rect 6563 3502 6578 3554
rect 7870 3726 7889 3778
rect 7889 3726 7922 3778
rect 7198 3502 7235 3554
rect 7235 3502 7250 3554
rect 7758 3502 7773 3554
rect 7773 3502 7810 3554
rect 8430 3502 8482 3554
rect 8542 3502 8579 3554
rect 8579 3502 8594 3554
rect 9662 3502 9714 3554
rect 9774 3502 9811 3554
rect 9811 3502 9826 3554
rect 10334 3502 10349 3554
rect 10349 3502 10386 3554
rect 10446 3502 10498 3554
rect 11006 3419 11021 3442
rect 11021 3419 11058 3442
rect 11006 3390 11058 3419
rect 11118 3502 11170 3554
rect 11678 3502 11730 3554
rect 11790 3419 11827 3442
rect 11827 3419 11842 3442
rect 11790 3390 11842 3419
rect 13918 3419 13933 3442
rect 13933 3419 13970 3442
rect 13918 3390 13970 3419
rect 14030 3390 14082 3442
rect 14590 3502 14605 3554
rect 14605 3502 14642 3554
rect 14702 3390 14754 3442
rect 15262 3502 15277 3554
rect 15277 3502 15314 3554
rect 15598 3502 15650 3554
rect 15822 3502 15874 3554
rect 15374 3390 15426 3442
rect 15934 3419 15949 3442
rect 15949 3419 15986 3442
rect 15934 3390 15986 3419
rect 16046 3390 16098 3442
rect 16606 3502 16621 3554
rect 16621 3502 16658 3554
rect 17614 3726 17633 3778
rect 17633 3726 17666 3778
rect 16718 3390 16770 3442
rect 17502 3502 17517 3554
rect 17517 3502 17554 3554
rect 18174 3502 18189 3554
rect 18189 3502 18226 3554
rect 18286 3390 18338 3442
rect 18846 3502 18861 3554
rect 18861 3502 18898 3554
rect 19630 3726 19649 3778
rect 19649 3726 19682 3778
rect 18958 3390 19010 3442
rect 19518 3419 19533 3442
rect 19533 3419 19570 3442
rect 19518 3390 19570 3419
rect 20302 3726 20321 3778
rect 20321 3726 20354 3778
rect 20190 3502 20205 3554
rect 20205 3502 20242 3554
rect 6534 3110 6794 3162
rect 11854 3110 12114 3162
rect 17174 3110 17434 3162
rect 22494 3110 22754 3162
<< metal2 >>
rect 3872 16492 4136 16502
rect 3872 16426 4136 16436
rect 9192 16492 9456 16502
rect 9192 16426 9456 16436
rect 14512 16492 14776 16502
rect 14512 16426 14776 16436
rect 19832 16492 20096 16502
rect 19832 16426 20096 16436
rect 6532 15708 6796 15718
rect 6532 15642 6796 15652
rect 11852 15708 12116 15718
rect 11852 15642 12116 15652
rect 17172 15708 17436 15718
rect 17172 15642 17436 15652
rect 22492 15708 22756 15718
rect 22492 15642 22756 15652
rect 3612 14980 3668 14990
rect 3388 9156 3444 9166
rect 3500 9156 3556 9166
rect 3388 9154 3500 9156
rect 3388 9102 3390 9154
rect 3442 9102 3500 9154
rect 3388 9100 3500 9102
rect 2940 8148 2996 8158
rect 3388 8148 3444 9100
rect 3500 9062 3556 9100
rect 3612 8484 3668 14924
rect 3872 14924 4136 14934
rect 3872 14858 4136 14868
rect 9192 14924 9456 14934
rect 9192 14858 9456 14868
rect 14512 14924 14776 14934
rect 14512 14858 14776 14868
rect 19832 14924 20096 14934
rect 19832 14858 20096 14868
rect 19628 14756 19684 14766
rect 16828 14644 16884 14654
rect 16828 14642 17108 14644
rect 16828 14590 16830 14642
rect 16882 14590 17108 14642
rect 16828 14588 17108 14590
rect 16828 14578 16884 14588
rect 16940 14418 16996 14430
rect 16940 14366 16942 14418
rect 16994 14366 16996 14418
rect 6532 14140 6796 14150
rect 6532 14074 6796 14084
rect 11852 14140 12116 14150
rect 11852 14074 12116 14084
rect 16156 13746 16212 13758
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 3872 13356 4136 13366
rect 3872 13290 4136 13300
rect 9192 13356 9456 13366
rect 9192 13290 9456 13300
rect 14512 13356 14776 13366
rect 14512 13290 14776 13300
rect 14924 13188 14980 13198
rect 14924 13094 14980 13132
rect 16156 13076 16212 13694
rect 16828 13746 16884 13758
rect 16828 13694 16830 13746
rect 16882 13694 16884 13746
rect 16268 13524 16324 13534
rect 16268 13430 16324 13468
rect 16156 13020 16324 13076
rect 14812 12852 14868 12862
rect 14812 12850 15092 12852
rect 14812 12798 14814 12850
rect 14866 12798 15092 12850
rect 14812 12796 15092 12798
rect 14812 12786 14868 12796
rect 6532 12572 6796 12582
rect 6532 12506 6796 12516
rect 11852 12572 12116 12582
rect 11852 12506 12116 12516
rect 14140 12178 14196 12190
rect 14140 12126 14142 12178
rect 14194 12126 14196 12178
rect 3872 11788 4136 11798
rect 3872 11722 4136 11732
rect 9192 11788 9456 11798
rect 9192 11722 9456 11732
rect 10668 11508 10724 11518
rect 7532 11452 8148 11508
rect 6076 11284 6132 11294
rect 6188 11284 6244 11294
rect 6076 11282 6188 11284
rect 6076 11230 6078 11282
rect 6130 11230 6188 11282
rect 6076 11228 6188 11230
rect 5404 10724 5460 10734
rect 5516 10724 5572 10734
rect 5404 10722 5516 10724
rect 5404 10670 5406 10722
rect 5458 10670 5516 10722
rect 5404 10668 5516 10670
rect 3872 10220 4136 10230
rect 3872 10154 4136 10164
rect 4172 9828 4228 9838
rect 4284 9828 4340 9838
rect 4172 9826 4284 9828
rect 4172 9774 4174 9826
rect 4226 9774 4284 9826
rect 4172 9772 4284 9774
rect 4060 9156 4116 9166
rect 4172 9156 4228 9772
rect 4284 9734 4340 9772
rect 4844 9828 4900 9838
rect 4844 9734 4900 9772
rect 5404 9828 5460 10668
rect 5516 10630 5572 10668
rect 6076 10724 6132 11228
rect 6188 11190 6244 11228
rect 6972 11284 7028 11294
rect 6972 11190 7028 11228
rect 6860 11170 6916 11182
rect 7532 11172 7588 11452
rect 7644 11284 7700 11294
rect 7644 11282 7812 11284
rect 7644 11230 7646 11282
rect 7698 11230 7812 11282
rect 7644 11228 7812 11230
rect 7644 11218 7700 11228
rect 6860 11118 6862 11170
rect 6914 11118 6916 11170
rect 6860 11060 6916 11118
rect 7420 11170 7588 11172
rect 7420 11118 7534 11170
rect 7586 11118 7588 11170
rect 7420 11116 7588 11118
rect 7756 11172 7812 11228
rect 8092 11172 8148 11452
rect 10444 11506 10724 11508
rect 10444 11454 10670 11506
rect 10722 11454 10724 11506
rect 10444 11452 10724 11454
rect 8316 11282 8372 11294
rect 8316 11230 8318 11282
rect 8370 11230 8372 11282
rect 8204 11172 8260 11182
rect 7756 11116 7924 11172
rect 7420 11060 7476 11116
rect 7532 11106 7588 11116
rect 6532 11004 6796 11014
rect 6532 10938 6796 10948
rect 6860 11004 7476 11060
rect 6860 10836 6916 11004
rect 6076 10592 6132 10668
rect 6188 10834 6916 10836
rect 6188 10782 6862 10834
rect 6914 10782 6916 10834
rect 6188 10780 6916 10782
rect 5404 9762 5460 9772
rect 6188 10386 6244 10780
rect 6860 10770 6916 10780
rect 6748 10612 6804 10622
rect 7420 10612 7476 10622
rect 7532 10612 7588 10622
rect 7868 10612 7924 11116
rect 8092 11170 8260 11172
rect 8092 11118 8206 11170
rect 8258 11118 8260 11170
rect 8092 11116 8260 11118
rect 8092 10722 8148 11116
rect 8204 11106 8260 11116
rect 8092 10670 8094 10722
rect 8146 10670 8148 10722
rect 8092 10658 8148 10670
rect 6636 10610 6804 10612
rect 6636 10558 6750 10610
rect 6802 10558 6804 10610
rect 6636 10556 6804 10558
rect 6636 10500 6692 10556
rect 6748 10546 6804 10556
rect 7308 10610 7924 10612
rect 7308 10558 7422 10610
rect 7474 10558 7534 10610
rect 7586 10558 7924 10610
rect 7308 10556 7924 10558
rect 6188 10334 6190 10386
rect 6242 10334 6244 10386
rect 5852 9716 5908 9726
rect 5740 9660 5852 9716
rect 4956 9602 5012 9614
rect 4956 9550 4958 9602
rect 5010 9550 5012 9602
rect 4116 9100 4228 9156
rect 4844 9268 4900 9278
rect 4956 9268 5012 9550
rect 4844 9266 5012 9268
rect 4844 9214 4846 9266
rect 4898 9214 5012 9266
rect 4844 9212 5012 9214
rect 4060 9024 4116 9100
rect 4732 9042 4788 9054
rect 4732 8990 4734 9042
rect 4786 8990 4788 9042
rect 4172 8820 4228 8830
rect 4172 8818 4340 8820
rect 4172 8766 4174 8818
rect 4226 8766 4340 8818
rect 4172 8764 4340 8766
rect 4172 8754 4228 8764
rect 3872 8652 4136 8662
rect 3872 8586 4136 8596
rect 2940 8146 3444 8148
rect 2940 8094 2942 8146
rect 2994 8094 3444 8146
rect 2940 8092 3444 8094
rect 3500 8372 3668 8428
rect 4172 8484 4228 8494
rect 3500 8146 3556 8372
rect 3500 8094 3502 8146
rect 3554 8094 3556 8146
rect 2828 8034 2884 8046
rect 2828 7982 2830 8034
rect 2882 7982 2884 8034
rect 2828 7700 2884 7982
rect 2604 7644 2884 7700
rect 2156 7476 2212 7486
rect 2156 7382 2212 7420
rect 2044 7252 2100 7262
rect 2604 7252 2660 7644
rect 2044 7250 2660 7252
rect 2044 7198 2046 7250
rect 2098 7198 2660 7250
rect 2044 7196 2660 7198
rect 2716 7476 2772 7486
rect 2940 7476 2996 8092
rect 2772 7420 2996 7476
rect 3388 7476 3444 7486
rect 3500 7476 3556 8094
rect 4172 8146 4228 8428
rect 4172 8094 4174 8146
rect 4226 8094 4228 8146
rect 3612 8036 3668 8046
rect 3612 8034 3780 8036
rect 3612 7982 3614 8034
rect 3666 7982 3780 8034
rect 3612 7980 3780 7982
rect 3612 7970 3668 7980
rect 3388 7474 3556 7476
rect 3388 7422 3390 7474
rect 3442 7422 3556 7474
rect 3388 7420 3556 7422
rect 2044 5906 2100 7196
rect 2156 6580 2212 6590
rect 2156 6486 2212 6524
rect 2044 5854 2046 5906
rect 2098 5854 2100 5906
rect 2044 5012 2100 5854
rect 2268 6466 2324 6478
rect 2268 6414 2270 6466
rect 2322 6414 2324 6466
rect 2156 5684 2212 5694
rect 2268 5684 2324 6414
rect 2716 5908 2772 7420
rect 2828 7250 2884 7262
rect 2828 7198 2830 7250
rect 2882 7198 2884 7250
rect 2828 6804 2884 7198
rect 2828 6738 2884 6748
rect 2828 6580 2884 6590
rect 2828 6486 2884 6524
rect 3388 6580 3444 7420
rect 3500 7252 3556 7262
rect 3612 7252 3668 7262
rect 3500 7250 3612 7252
rect 3500 7198 3502 7250
rect 3554 7198 3612 7250
rect 3500 7196 3612 7198
rect 3500 7186 3556 7196
rect 3500 6580 3556 6590
rect 3444 6578 3556 6580
rect 3444 6526 3502 6578
rect 3554 6526 3556 6578
rect 3444 6524 3556 6526
rect 2940 6466 2996 6478
rect 2940 6414 2942 6466
rect 2994 6414 2996 6466
rect 2940 5908 2996 6414
rect 2716 5906 2996 5908
rect 2716 5854 2718 5906
rect 2770 5854 2996 5906
rect 2716 5852 2996 5854
rect 3388 5906 3444 6524
rect 3500 6514 3556 6524
rect 3388 5854 3390 5906
rect 3442 5854 3444 5906
rect 2716 5684 2772 5852
rect 2156 5682 2772 5684
rect 2156 5630 2158 5682
rect 2210 5630 2772 5682
rect 2156 5628 2772 5630
rect 2828 5682 2884 5694
rect 2828 5630 2830 5682
rect 2882 5630 2884 5682
rect 2156 5618 2212 5628
rect 2156 5012 2212 5022
rect 2044 5010 2212 5012
rect 2044 4958 2158 5010
rect 2210 4958 2212 5010
rect 2044 4956 2212 4958
rect 2156 4452 2212 4956
rect 2268 4898 2324 5628
rect 2828 5572 2884 5630
rect 2716 5516 2884 5572
rect 2716 5124 2772 5516
rect 2716 5058 2772 5068
rect 3388 5124 3444 5854
rect 3612 6466 3668 7196
rect 3724 6804 3780 7980
rect 4060 7476 4116 7486
rect 4172 7476 4228 8094
rect 4284 8036 4340 8764
rect 4284 7942 4340 7980
rect 4732 8484 4788 8990
rect 4732 7586 4788 8428
rect 4732 7534 4734 7586
rect 4786 7534 4788 7586
rect 4060 7474 4340 7476
rect 4060 7422 4062 7474
rect 4114 7422 4340 7474
rect 4060 7420 4340 7422
rect 4060 7410 4116 7420
rect 4172 7252 4228 7290
rect 4172 7186 4228 7196
rect 3872 7084 4136 7094
rect 3872 7018 4136 7028
rect 4284 6914 4340 7420
rect 4284 6862 4286 6914
rect 4338 6862 4340 6914
rect 4284 6850 4340 6862
rect 4732 6916 4788 7534
rect 4844 8146 4900 9212
rect 5404 9044 5460 9054
rect 5740 9044 5796 9660
rect 5852 9584 5908 9660
rect 5964 9604 6020 9614
rect 6188 9604 6244 10334
rect 6524 10444 6692 10500
rect 6524 9716 6580 10444
rect 6636 9716 6692 9726
rect 6580 9714 6692 9716
rect 6580 9662 6638 9714
rect 6690 9662 6692 9714
rect 6580 9660 6692 9662
rect 6524 9622 6580 9660
rect 6636 9650 6692 9660
rect 7196 9716 7252 9726
rect 7308 9716 7364 10556
rect 7420 10546 7476 10556
rect 7532 10546 7588 10556
rect 7868 10388 7924 10556
rect 8204 10388 8260 10398
rect 8316 10388 8372 11230
rect 9212 11282 9268 11294
rect 9212 11230 9214 11282
rect 9266 11230 9268 11282
rect 7868 10386 8372 10388
rect 7868 10334 8206 10386
rect 8258 10334 8372 10386
rect 7868 10332 8372 10334
rect 7868 9826 7924 10332
rect 8204 10322 8260 10332
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9762 7924 9774
rect 8316 9828 8372 10332
rect 8876 10612 8932 10622
rect 9212 10612 9268 11230
rect 9884 11282 9940 11294
rect 9884 11230 9886 11282
rect 9938 11230 9940 11282
rect 8876 10610 9268 10612
rect 8876 10558 8878 10610
rect 8930 10558 9268 10610
rect 8876 10556 9268 10558
rect 9324 11170 9380 11182
rect 9324 11118 9326 11170
rect 9378 11118 9380 11170
rect 8540 9828 8596 9838
rect 8876 9828 8932 10556
rect 8988 10388 9044 10398
rect 9324 10388 9380 11118
rect 8988 10386 9380 10388
rect 8988 10334 8990 10386
rect 9042 10334 9380 10386
rect 8988 10332 9380 10334
rect 9884 10610 9940 11230
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 8988 10052 9044 10332
rect 9192 10220 9456 10230
rect 9192 10154 9456 10164
rect 8988 9986 9044 9996
rect 9884 9940 9940 10558
rect 9996 11172 10052 11182
rect 10444 11172 10500 11452
rect 10668 11442 10724 11452
rect 10556 11284 10612 11294
rect 12124 11284 12180 11294
rect 12236 11284 12292 11294
rect 10556 11282 10724 11284
rect 10556 11230 10558 11282
rect 10610 11230 10724 11282
rect 10556 11228 10724 11230
rect 10556 11218 10612 11228
rect 9996 11170 10500 11172
rect 9996 11118 9998 11170
rect 10050 11118 10500 11170
rect 9996 11116 10500 11118
rect 9996 10386 10052 11116
rect 9996 10334 9998 10386
rect 10050 10334 10052 10386
rect 9996 10164 10052 10334
rect 9996 10098 10052 10108
rect 10556 10610 10612 10622
rect 10556 10558 10558 10610
rect 10610 10558 10612 10610
rect 9212 9884 10052 9940
rect 9212 9828 9268 9884
rect 8316 9826 9268 9828
rect 8316 9774 8542 9826
rect 8594 9774 9214 9826
rect 9266 9774 9268 9826
rect 8316 9772 9268 9774
rect 8540 9762 8596 9772
rect 7252 9714 7364 9716
rect 7252 9662 7310 9714
rect 7362 9662 7364 9714
rect 7252 9660 7364 9662
rect 7196 9622 7252 9660
rect 5964 9602 6244 9604
rect 5964 9550 5966 9602
rect 6018 9550 6244 9602
rect 5964 9548 6244 9550
rect 5964 9492 6020 9548
rect 5404 9042 5796 9044
rect 5404 8990 5406 9042
rect 5458 8990 5796 9042
rect 5404 8988 5796 8990
rect 5852 9436 6020 9492
rect 6532 9436 6796 9446
rect 4956 8484 5012 8522
rect 4956 8418 5012 8428
rect 5404 8484 5460 8988
rect 5404 8418 5460 8428
rect 5516 8818 5572 8830
rect 5516 8766 5518 8818
rect 5570 8766 5572 8818
rect 4844 8094 4846 8146
rect 4898 8094 4900 8146
rect 4844 8036 4900 8094
rect 4844 7476 4900 7980
rect 5516 8148 5572 8766
rect 5852 8148 5908 9436
rect 6532 9370 6796 9380
rect 7308 9156 7364 9660
rect 7980 9604 8036 9614
rect 8652 9604 8708 9614
rect 7980 9602 8260 9604
rect 7980 9550 7982 9602
rect 8034 9550 8260 9602
rect 7980 9548 8260 9550
rect 7420 9156 7476 9166
rect 7532 9156 7588 9166
rect 7308 9154 7588 9156
rect 7308 9102 7422 9154
rect 7474 9102 7534 9154
rect 7586 9102 7588 9154
rect 7308 9100 7588 9102
rect 6076 9044 6132 9054
rect 6188 9044 6244 9054
rect 6748 9044 6804 9054
rect 6860 9044 6916 9054
rect 6076 9042 6244 9044
rect 6076 8990 6078 9042
rect 6130 8990 6190 9042
rect 6242 8990 6244 9042
rect 6076 8988 6244 8990
rect 5964 8484 6020 8522
rect 6076 8428 6132 8988
rect 6188 8978 6244 8988
rect 6636 9042 6916 9044
rect 6636 8990 6750 9042
rect 6802 8990 6862 9042
rect 6914 8990 6916 9042
rect 6636 8988 6916 8990
rect 5964 8372 6132 8428
rect 5516 8146 5908 8148
rect 5516 8094 5854 8146
rect 5906 8094 5908 8146
rect 5516 8092 5908 8094
rect 4844 7382 4900 7420
rect 5404 7476 5460 7486
rect 5516 7476 5572 8092
rect 5852 8082 5908 8092
rect 6076 7700 6132 8372
rect 6524 8484 6580 8494
rect 6636 8484 6692 8988
rect 6748 8978 6804 8988
rect 6580 8482 6692 8484
rect 6580 8430 6638 8482
rect 6690 8430 6692 8482
rect 6580 8428 6692 8430
rect 6524 8258 6580 8428
rect 6636 8418 6692 8428
rect 6524 8206 6526 8258
rect 6578 8206 6580 8258
rect 6524 8194 6580 8206
rect 6532 7868 6796 7878
rect 6532 7802 6796 7812
rect 6188 7700 6244 7710
rect 6076 7698 6244 7700
rect 6076 7646 6190 7698
rect 6242 7646 6244 7698
rect 6076 7644 6244 7646
rect 5460 7420 5572 7476
rect 5404 7344 5460 7420
rect 5516 7250 5572 7420
rect 6076 7476 6132 7486
rect 6076 7382 6132 7420
rect 5516 7198 5518 7250
rect 5570 7198 5572 7250
rect 4956 6916 5012 6926
rect 4732 6914 5012 6916
rect 4732 6862 4958 6914
rect 5010 6862 5012 6914
rect 4732 6860 5012 6862
rect 4956 6850 5012 6860
rect 3724 6738 3780 6748
rect 4620 6804 4676 6814
rect 5516 6804 5572 7198
rect 4676 6748 4788 6804
rect 4620 6738 4676 6748
rect 3612 6414 3614 6466
rect 3666 6414 3668 6466
rect 3388 5058 3444 5068
rect 3500 5684 3556 5694
rect 3612 5684 3668 6414
rect 4172 6578 4228 6590
rect 4172 6526 4174 6578
rect 4226 6526 4228 6578
rect 4060 5908 4116 5918
rect 4060 5796 4116 5852
rect 3500 5682 3668 5684
rect 3500 5630 3502 5682
rect 3554 5630 3668 5682
rect 3500 5628 3668 5630
rect 3724 5740 4116 5796
rect 2828 5012 2884 5022
rect 2828 5010 2996 5012
rect 2828 4958 2830 5010
rect 2882 4958 2996 5010
rect 2828 4956 2996 4958
rect 2828 4946 2884 4956
rect 2268 4846 2270 4898
rect 2322 4846 2324 4898
rect 2268 4788 2324 4846
rect 2940 4900 2996 4956
rect 3500 5010 3556 5628
rect 3500 4958 3502 5010
rect 3554 4958 3556 5010
rect 2940 4898 3108 4900
rect 2940 4846 2942 4898
rect 2994 4846 3108 4898
rect 2940 4844 3108 4846
rect 2940 4834 2996 4844
rect 2268 4732 2548 4788
rect 2380 4452 2436 4462
rect 2156 4396 2380 4452
rect 2380 4358 2436 4396
rect 2492 4340 2548 4732
rect 3052 4452 3108 4844
rect 2492 4246 2548 4284
rect 2828 4340 2884 4350
rect 2156 3556 2212 3566
rect 2156 800 2212 3500
rect 2828 3556 2884 4284
rect 3052 4338 3108 4396
rect 3052 4286 3054 4338
rect 3106 4286 3108 4338
rect 2940 3780 2996 3790
rect 3052 3780 3108 4286
rect 3164 4340 3220 4350
rect 3164 4246 3220 4284
rect 3500 4340 3556 4958
rect 3612 5012 3668 5022
rect 3724 5012 3780 5740
rect 4172 5684 4228 6526
rect 4732 5908 4788 6748
rect 5516 6738 5572 6748
rect 5740 6804 5796 6814
rect 5740 6692 5796 6748
rect 5852 6692 5908 6702
rect 5740 6690 5908 6692
rect 5740 6638 5742 6690
rect 5794 6638 5854 6690
rect 5906 6638 5908 6690
rect 5740 6636 5908 6638
rect 5740 6626 5796 6636
rect 5852 6626 5908 6636
rect 4732 5814 4788 5852
rect 4844 6578 4900 6590
rect 4844 6526 4846 6578
rect 4898 6526 4900 6578
rect 4844 5684 4900 6526
rect 5516 6132 5572 6142
rect 6188 6132 6244 7644
rect 6860 7698 6916 8988
rect 7196 8484 7252 8494
rect 7196 8258 7252 8428
rect 7420 8428 7476 9100
rect 7532 9090 7588 9100
rect 7980 8484 8036 9548
rect 8204 9154 8260 9548
rect 8204 9102 8206 9154
rect 8258 9102 8260 9154
rect 8204 9090 8260 9102
rect 8540 9548 8652 9604
rect 7420 8372 7588 8428
rect 7196 8206 7198 8258
rect 7250 8206 7252 8258
rect 7196 8194 7252 8206
rect 6860 7646 6862 7698
rect 6914 7646 6916 7698
rect 6860 7634 6916 7646
rect 7308 8036 7364 8046
rect 6748 7476 6804 7486
rect 6412 6804 6468 6814
rect 6412 6692 6468 6748
rect 6524 6692 6580 6702
rect 6748 6692 6804 7420
rect 7308 7476 7364 7980
rect 7308 7410 7364 7420
rect 7420 7474 7476 7486
rect 7420 7422 7422 7474
rect 7474 7422 7476 7474
rect 7420 7252 7476 7422
rect 7532 7252 7588 8372
rect 7868 8372 8036 8428
rect 8316 8818 8372 8830
rect 8316 8766 8318 8818
rect 8370 8766 8372 8818
rect 7868 8258 7924 8372
rect 7868 8206 7870 8258
rect 7922 8206 7924 8258
rect 7868 8194 7924 8206
rect 7980 8036 8036 8046
rect 7980 7942 8036 7980
rect 8316 8036 8372 8766
rect 8540 8484 8596 9548
rect 8652 9472 8708 9548
rect 8988 9266 9044 9772
rect 9212 9762 9268 9772
rect 9884 9714 9940 9726
rect 9884 9662 9886 9714
rect 9938 9662 9940 9714
rect 9324 9604 9380 9614
rect 9324 9510 9380 9548
rect 8988 9214 8990 9266
rect 9042 9214 9044 9266
rect 8988 9202 9044 9214
rect 8540 8148 8596 8428
rect 8876 9042 8932 9054
rect 8876 8990 8878 9042
rect 8930 8990 8932 9042
rect 8876 8428 8932 8990
rect 9192 8652 9456 8662
rect 9192 8586 9456 8596
rect 9324 8484 9380 8522
rect 8876 8372 9044 8428
rect 9324 8418 9380 8428
rect 8316 7970 8372 7980
rect 8428 8146 8596 8148
rect 8428 8094 8542 8146
rect 8594 8094 8596 8146
rect 8428 8092 8596 8094
rect 8204 7476 8260 7486
rect 8428 7476 8484 8092
rect 8540 8082 8596 8092
rect 8652 8036 8708 8046
rect 8652 8034 8820 8036
rect 8652 7982 8654 8034
rect 8706 7982 8820 8034
rect 8652 7980 8820 7982
rect 8652 7970 8708 7980
rect 8204 7474 8484 7476
rect 8204 7422 8206 7474
rect 8258 7422 8484 7474
rect 8204 7420 8484 7422
rect 8204 7410 8260 7420
rect 7420 7250 7588 7252
rect 7420 7198 7534 7250
rect 7586 7198 7588 7250
rect 7420 7196 7588 7198
rect 7532 6916 7588 7196
rect 6412 6690 6916 6692
rect 6412 6638 6414 6690
rect 6466 6638 6526 6690
rect 6578 6638 6916 6690
rect 6412 6636 6916 6638
rect 6412 6626 6468 6636
rect 6524 6626 6580 6636
rect 6860 6580 6916 6636
rect 7084 6580 7140 6590
rect 6860 6578 7140 6580
rect 6860 6526 7086 6578
rect 7138 6526 7140 6578
rect 6860 6524 7140 6526
rect 6532 6300 6796 6310
rect 6532 6234 6796 6244
rect 5516 6130 6580 6132
rect 5516 6078 5518 6130
rect 5570 6078 6190 6130
rect 6242 6078 6580 6130
rect 5516 6076 6580 6078
rect 5516 6066 5572 6076
rect 4172 5682 4900 5684
rect 4172 5630 4174 5682
rect 4226 5630 4846 5682
rect 4898 5630 4900 5682
rect 4172 5628 4900 5630
rect 4172 5618 4228 5628
rect 3872 5516 4136 5526
rect 3872 5450 4136 5460
rect 4172 5124 4228 5134
rect 4172 5030 4228 5068
rect 3668 4956 3780 5012
rect 3612 4564 3668 4956
rect 4284 4900 4340 4910
rect 4732 4900 4788 5628
rect 4844 5618 4900 5628
rect 5404 5906 5460 5918
rect 5404 5854 5406 5906
rect 5458 5854 5460 5906
rect 4284 4898 4452 4900
rect 4284 4846 4286 4898
rect 4338 4846 4452 4898
rect 4284 4844 4452 4846
rect 4284 4834 4340 4844
rect 3836 4564 3892 4574
rect 3612 4508 3836 4564
rect 3836 4432 3892 4508
rect 3500 4274 3556 4284
rect 3724 4340 3780 4350
rect 2940 3778 3108 3780
rect 2940 3726 2942 3778
rect 2994 3726 3108 3778
rect 2940 3724 3108 3726
rect 2940 3714 2996 3724
rect 2828 3424 2884 3500
rect 3052 3556 3108 3724
rect 3612 3780 3668 3790
rect 3724 3780 3780 4284
rect 4396 4340 4452 4844
rect 4732 4834 4788 4844
rect 4844 5122 4900 5134
rect 4844 5070 4846 5122
rect 4898 5070 4900 5122
rect 4508 4564 4564 4574
rect 4508 4470 4564 4508
rect 4844 4564 4900 5070
rect 4956 5124 5012 5134
rect 5012 5068 5124 5124
rect 4956 5058 5012 5068
rect 4956 4900 5012 4910
rect 4956 4806 5012 4844
rect 4284 4116 4340 4126
rect 3872 3948 4136 3958
rect 3872 3882 4136 3892
rect 3612 3778 3780 3780
rect 3612 3726 3614 3778
rect 3666 3726 3780 3778
rect 3612 3724 3780 3726
rect 4284 3778 4340 4060
rect 4284 3726 4286 3778
rect 4338 3726 4340 3778
rect 3612 3714 3668 3724
rect 3052 3490 3108 3500
rect 3500 3556 3556 3566
rect 3500 3462 3556 3500
rect 4172 3556 4228 3566
rect 4284 3556 4340 3726
rect 4228 3500 4340 3556
rect 4172 3424 4228 3500
rect 4396 3444 4452 4284
rect 4844 3780 4900 4508
rect 5068 4450 5124 5068
rect 5404 4900 5460 5854
rect 5852 5348 5908 6076
rect 6188 6066 6244 6076
rect 6076 5906 6132 5918
rect 6076 5854 6078 5906
rect 6130 5854 6132 5906
rect 5852 5346 6020 5348
rect 5852 5294 5854 5346
rect 5906 5294 6020 5346
rect 5852 5292 6020 5294
rect 5852 5282 5908 5292
rect 5740 5012 5796 5022
rect 5740 5010 5908 5012
rect 5740 4958 5742 5010
rect 5794 4958 5908 5010
rect 5740 4956 5908 4958
rect 5740 4946 5796 4956
rect 5404 4834 5460 4844
rect 5852 4900 5908 4956
rect 5068 4398 5070 4450
rect 5122 4398 5124 4450
rect 5068 4386 5124 4398
rect 5740 4564 5796 4574
rect 5740 4450 5796 4508
rect 5740 4398 5742 4450
rect 5794 4398 5796 4450
rect 5740 4386 5796 4398
rect 5180 4114 5236 4126
rect 5180 4062 5182 4114
rect 5234 4062 5236 4114
rect 4956 3780 5012 3790
rect 4844 3778 5012 3780
rect 4844 3726 4958 3778
rect 5010 3726 5012 3778
rect 4844 3724 5012 3726
rect 4956 3714 5012 3724
rect 4396 3378 4452 3388
rect 4844 3444 4900 3454
rect 4844 3350 4900 3388
rect 5180 3444 5236 4062
rect 5852 4116 5908 4844
rect 5852 4022 5908 4060
rect 5964 4340 6020 5292
rect 6076 4900 6132 5854
rect 6524 5348 6580 6076
rect 6748 6020 6804 6030
rect 6860 6020 6916 6524
rect 6748 6018 6916 6020
rect 6748 5966 6750 6018
rect 6802 5966 6862 6018
rect 6914 5966 6916 6018
rect 6748 5964 6916 5966
rect 6748 5954 6804 5964
rect 6860 5954 6916 5964
rect 7084 6020 7140 6524
rect 7084 5572 7140 5964
rect 7196 6466 7252 6478
rect 7196 6414 7198 6466
rect 7250 6414 7252 6466
rect 7196 5684 7252 6414
rect 7420 6020 7476 6030
rect 7420 5926 7476 5964
rect 7532 5684 7588 6860
rect 8316 7250 8372 7262
rect 8316 7198 8318 7250
rect 8370 7198 8372 7250
rect 7756 6578 7812 6590
rect 7756 6526 7758 6578
rect 7810 6526 7812 6578
rect 7756 6020 7812 6526
rect 7756 5954 7812 5964
rect 7868 6466 7924 6478
rect 7868 6414 7870 6466
rect 7922 6414 7924 6466
rect 7868 5684 7924 6414
rect 8092 6020 8148 6030
rect 8316 6020 8372 7198
rect 8428 6580 8484 7420
rect 8764 7476 8820 7980
rect 8988 7698 9044 8316
rect 9884 8372 9940 9662
rect 9212 8260 9268 8270
rect 9212 8166 9268 8204
rect 9884 8258 9940 8316
rect 9884 8206 9886 8258
rect 9938 8206 9940 8258
rect 8988 7646 8990 7698
rect 9042 7646 9044 7698
rect 8988 7634 9044 7646
rect 9884 7700 9940 8206
rect 9996 9602 10052 9884
rect 10556 9828 10612 10558
rect 9996 9550 9998 9602
rect 10050 9550 10052 9602
rect 9996 8596 10052 9550
rect 10332 9826 10612 9828
rect 10332 9774 10558 9826
rect 10610 9774 10612 9826
rect 10332 9772 10612 9774
rect 10332 9156 10388 9772
rect 10556 9762 10612 9772
rect 10668 10388 10724 11228
rect 12124 11282 12292 11284
rect 12124 11230 12126 11282
rect 12178 11230 12238 11282
rect 12290 11230 12292 11282
rect 12124 11228 12292 11230
rect 12124 11218 12180 11228
rect 11852 11004 12116 11014
rect 11852 10938 12116 10948
rect 11228 10610 11284 10622
rect 11228 10558 11230 10610
rect 11282 10558 11284 10610
rect 11228 10388 11284 10558
rect 12012 10610 12068 10622
rect 12012 10558 12014 10610
rect 12066 10558 12068 10610
rect 10668 10386 11284 10388
rect 10668 10334 10670 10386
rect 10722 10334 11284 10386
rect 10668 10332 11284 10334
rect 11340 10386 11396 10398
rect 11340 10334 11342 10386
rect 11394 10334 11396 10386
rect 10668 9604 10724 10332
rect 11340 10052 11396 10334
rect 12012 10388 12068 10558
rect 12236 10612 12292 11228
rect 12796 11282 12852 11294
rect 12796 11230 12798 11282
rect 12850 11230 12852 11282
rect 12796 11172 12852 11230
rect 13692 11282 13748 11294
rect 13692 11230 13694 11282
rect 13746 11230 13748 11282
rect 12908 11172 12964 11182
rect 12796 11170 12964 11172
rect 12796 11118 12910 11170
rect 12962 11118 12964 11170
rect 12796 11116 12964 11118
rect 12684 10612 12740 10622
rect 12796 10612 12852 11116
rect 12908 11106 12964 11116
rect 13692 11172 13748 11230
rect 13804 11172 13860 11182
rect 13692 11170 13860 11172
rect 13692 11118 13806 11170
rect 13858 11118 13860 11170
rect 13692 11116 13860 11118
rect 13356 10612 13412 10622
rect 13468 10612 13524 10622
rect 13692 10612 13748 11116
rect 13804 11106 13860 11116
rect 14028 10612 14084 10622
rect 14140 10612 14196 12126
rect 14812 12180 14868 12190
rect 14812 12086 14868 12124
rect 14252 11956 14308 11966
rect 14252 11862 14308 11900
rect 14924 11956 14980 11966
rect 14512 11788 14776 11798
rect 14512 11722 14776 11732
rect 14924 11396 14980 11900
rect 14924 11302 14980 11340
rect 14812 11282 14868 11294
rect 14812 11230 14814 11282
rect 14866 11230 14868 11282
rect 14700 10612 14756 10622
rect 14812 10612 14868 11230
rect 12236 10610 14868 10612
rect 12236 10558 12686 10610
rect 12738 10558 12798 10610
rect 12850 10558 13358 10610
rect 13410 10558 13470 10610
rect 13522 10558 14030 10610
rect 14082 10558 14142 10610
rect 14194 10558 14702 10610
rect 14754 10558 14814 10610
rect 14866 10558 14868 10610
rect 12236 10556 14868 10558
rect 12124 10388 12180 10398
rect 12236 10388 12292 10556
rect 12684 10546 12740 10556
rect 12796 10546 12852 10556
rect 13356 10546 13412 10556
rect 13468 10546 13524 10556
rect 14028 10546 14084 10556
rect 14140 10546 14196 10556
rect 14700 10546 14756 10556
rect 14812 10546 14868 10556
rect 12012 10386 12292 10388
rect 12012 10334 12126 10386
rect 12178 10334 12292 10386
rect 12012 10332 12292 10334
rect 11564 10052 11620 10062
rect 11396 10050 11620 10052
rect 11396 9998 11566 10050
rect 11618 9998 11620 10050
rect 11396 9996 11620 9998
rect 11340 9986 11396 9996
rect 11564 9986 11620 9996
rect 12012 10052 12068 10332
rect 12124 10322 12180 10332
rect 14512 10220 14776 10230
rect 14512 10154 14776 10164
rect 12012 9828 12068 9996
rect 12124 9828 12180 9838
rect 12236 9828 12292 9838
rect 14476 9828 14532 9838
rect 15036 9828 15092 12796
rect 15484 12850 15540 12862
rect 15484 12798 15486 12850
rect 15538 12798 15540 12850
rect 15484 12180 15540 12798
rect 16156 12850 16212 12862
rect 16156 12798 16158 12850
rect 16210 12798 16212 12850
rect 15484 11282 15540 12124
rect 15596 12738 15652 12750
rect 15596 12686 15598 12738
rect 15650 12686 15652 12738
rect 15596 11954 15652 12686
rect 15596 11902 15598 11954
rect 15650 11902 15652 11954
rect 15596 11396 15652 11902
rect 15596 11302 15652 11340
rect 16156 12180 16212 12798
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15372 10612 15428 10622
rect 15484 10612 15540 11230
rect 16156 11282 16212 12124
rect 16268 12738 16324 13020
rect 16828 12852 16884 13694
rect 16940 13524 16996 14366
rect 16940 13430 16996 13468
rect 17052 14308 17108 14588
rect 17612 14418 17668 14430
rect 17612 14366 17614 14418
rect 17666 14366 17668 14418
rect 17500 14308 17556 14318
rect 17052 14306 17556 14308
rect 17052 14254 17502 14306
rect 17554 14254 17556 14306
rect 17052 14252 17556 14254
rect 17052 13188 17108 14252
rect 17500 14242 17556 14252
rect 17172 14140 17436 14150
rect 17172 14074 17436 14084
rect 17052 13122 17108 13132
rect 17388 13524 17444 13534
rect 16828 12850 16996 12852
rect 16828 12798 16830 12850
rect 16882 12798 16996 12850
rect 16828 12796 16996 12798
rect 16828 12786 16884 12796
rect 16268 12686 16270 12738
rect 16322 12686 16324 12738
rect 16268 11954 16324 12686
rect 16940 12738 16996 12796
rect 16940 12686 16942 12738
rect 16994 12686 16996 12738
rect 16828 12180 16884 12190
rect 16828 12086 16884 12124
rect 16268 11902 16270 11954
rect 16322 11902 16324 11954
rect 16268 11396 16324 11902
rect 16940 11954 16996 12686
rect 17388 12740 17444 13468
rect 17612 13524 17668 14366
rect 17612 13458 17668 13468
rect 17724 13746 17780 13758
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13188 17780 13694
rect 18396 13746 18452 13758
rect 18396 13694 18398 13746
rect 18450 13694 18452 13746
rect 17724 13122 17780 13132
rect 17836 13522 17892 13534
rect 17836 13470 17838 13522
rect 17890 13470 17892 13522
rect 17500 12964 17556 12974
rect 17836 12964 17892 13470
rect 18396 13524 18452 13694
rect 18396 13458 18452 13468
rect 18508 13522 18564 13534
rect 18508 13470 18510 13522
rect 18562 13470 18564 13522
rect 18508 13300 18564 13470
rect 18508 13234 18564 13244
rect 18956 13524 19012 13534
rect 18284 13188 18340 13198
rect 18284 13094 18340 13132
rect 18844 13188 18900 13198
rect 17500 12962 17892 12964
rect 17500 12910 17502 12962
rect 17554 12910 17892 12962
rect 17500 12908 17892 12910
rect 17500 12898 17556 12908
rect 17612 12740 17668 12750
rect 17388 12738 17668 12740
rect 17388 12686 17614 12738
rect 17666 12686 17668 12738
rect 17388 12684 17668 12686
rect 17172 12572 17436 12582
rect 17172 12506 17436 12516
rect 16940 11902 16942 11954
rect 16994 11902 16996 11954
rect 16268 11302 16324 11340
rect 16828 11396 16884 11406
rect 16940 11396 16996 11902
rect 17612 11844 17668 12684
rect 17612 11778 17668 11788
rect 17724 12292 17780 12302
rect 17836 12292 17892 12908
rect 18844 12962 18900 13132
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 12898 18900 12910
rect 18956 13186 19012 13468
rect 19628 13524 19684 14700
rect 22492 14140 22756 14150
rect 22492 14074 22756 14084
rect 18956 13134 18958 13186
rect 19010 13134 19012 13186
rect 18172 12850 18228 12862
rect 18172 12798 18174 12850
rect 18226 12798 18228 12850
rect 18172 12292 18228 12798
rect 18396 12292 18452 12302
rect 17724 12290 18396 12292
rect 17724 12238 17726 12290
rect 17778 12238 17838 12290
rect 17890 12238 18396 12290
rect 17724 12236 18396 12238
rect 17612 11620 17668 11630
rect 17724 11620 17780 12236
rect 17836 12226 17892 12236
rect 17612 11618 17780 11620
rect 17612 11566 17614 11618
rect 17666 11566 17780 11618
rect 17612 11564 17780 11566
rect 16828 11394 16940 11396
rect 16828 11342 16830 11394
rect 16882 11342 16940 11394
rect 16828 11340 16940 11342
rect 16156 11230 16158 11282
rect 16210 11230 16212 11282
rect 16044 10612 16100 10622
rect 12012 9826 12404 9828
rect 12012 9774 12126 9826
rect 12178 9774 12238 9826
rect 12290 9774 12404 9826
rect 12012 9772 12404 9774
rect 12124 9762 12180 9772
rect 12236 9762 12292 9772
rect 11452 9716 11508 9726
rect 9996 8482 10052 8540
rect 9996 8430 9998 8482
rect 10050 8430 10052 8482
rect 9996 8260 10052 8430
rect 10108 9154 10388 9156
rect 10108 9102 10334 9154
rect 10386 9102 10388 9154
rect 10108 9100 10388 9102
rect 10108 8428 10164 9100
rect 10332 9090 10388 9100
rect 10556 9602 10724 9604
rect 10556 9550 10670 9602
rect 10722 9550 10724 9602
rect 10556 9548 10724 9550
rect 10444 8932 10500 8942
rect 10556 8932 10612 9548
rect 10668 9538 10724 9548
rect 11340 9714 11508 9716
rect 11340 9662 11454 9714
rect 11506 9662 11508 9714
rect 11340 9660 11508 9662
rect 11004 9044 11060 9054
rect 11004 9042 11172 9044
rect 11004 8990 11006 9042
rect 11058 8990 11172 9042
rect 11004 8988 11172 8990
rect 11004 8978 11060 8988
rect 10444 8930 10612 8932
rect 10444 8878 10446 8930
rect 10498 8878 10612 8930
rect 10444 8876 10612 8878
rect 10444 8866 10500 8876
rect 10556 8596 10612 8876
rect 11116 8820 11172 8988
rect 11340 8820 11396 9660
rect 11452 9650 11508 9660
rect 11852 9436 12116 9446
rect 11852 9370 12116 9380
rect 12348 9156 12404 9772
rect 14476 9826 15092 9828
rect 14476 9774 14478 9826
rect 14530 9774 15038 9826
rect 15090 9774 15092 9826
rect 14476 9772 15092 9774
rect 12796 9716 12852 9726
rect 12908 9716 12964 9726
rect 12796 9714 12964 9716
rect 12796 9662 12798 9714
rect 12850 9662 12910 9714
rect 12962 9662 12964 9714
rect 12796 9660 12964 9662
rect 12796 9156 12852 9660
rect 12908 9650 12964 9660
rect 13692 9716 13748 9726
rect 13804 9716 13860 9726
rect 13692 9714 13860 9716
rect 13692 9662 13694 9714
rect 13746 9662 13806 9714
rect 13858 9662 13860 9714
rect 13692 9660 13860 9662
rect 13020 9156 13076 9166
rect 12348 9154 13076 9156
rect 12348 9102 12350 9154
rect 12402 9102 13022 9154
rect 13074 9102 13076 9154
rect 12348 9100 13076 9102
rect 12348 9090 12404 9100
rect 11116 8818 11396 8820
rect 11116 8766 11118 8818
rect 11170 8766 11396 8818
rect 11116 8764 11396 8766
rect 11676 9042 11732 9054
rect 11676 8990 11678 9042
rect 11730 8990 11732 9042
rect 11676 8820 11732 8990
rect 11788 8820 11844 8830
rect 11676 8818 11844 8820
rect 11676 8766 11790 8818
rect 11842 8766 11844 8818
rect 11676 8764 11844 8766
rect 11116 8754 11172 8764
rect 10556 8484 10612 8540
rect 10668 8484 10724 8494
rect 10556 8482 10836 8484
rect 10556 8430 10670 8482
rect 10722 8430 10836 8482
rect 10556 8428 10836 8430
rect 11340 8428 11396 8764
rect 11788 8428 11844 8764
rect 12460 8818 12516 8830
rect 12460 8766 12462 8818
rect 12514 8766 12516 8818
rect 10108 8372 10388 8428
rect 10668 8418 10724 8428
rect 10780 8372 11284 8428
rect 10388 8316 10612 8372
rect 10332 8306 10388 8316
rect 9996 8194 10052 8204
rect 10556 8258 10612 8316
rect 10556 8206 10558 8258
rect 10610 8206 10612 8258
rect 9996 7700 10052 7710
rect 9884 7698 10052 7700
rect 9884 7646 9998 7698
rect 10050 7646 10052 7698
rect 9884 7644 10052 7646
rect 9996 7634 10052 7644
rect 10556 7586 10612 8206
rect 10668 7700 10724 7710
rect 10780 7700 10836 8372
rect 10668 7698 10836 7700
rect 10668 7646 10670 7698
rect 10722 7646 10836 7698
rect 10668 7644 10836 7646
rect 11228 8370 11284 8372
rect 11228 8318 11230 8370
rect 11282 8318 11284 8370
rect 11228 7698 11284 8318
rect 11228 7646 11230 7698
rect 11282 7646 11284 7698
rect 10668 7634 10724 7644
rect 11228 7634 11284 7646
rect 11340 8372 12180 8428
rect 11340 8146 11396 8372
rect 12124 8260 12180 8372
rect 12236 8260 12292 8270
rect 12460 8260 12516 8766
rect 12124 8258 12460 8260
rect 12124 8206 12126 8258
rect 12178 8206 12238 8258
rect 12290 8206 12460 8258
rect 12124 8204 12460 8206
rect 12124 8194 12180 8204
rect 12236 8194 12292 8204
rect 11340 8094 11342 8146
rect 11394 8094 11396 8146
rect 12460 8128 12516 8204
rect 12796 8484 12852 9100
rect 13020 9090 13076 9100
rect 13692 9042 13748 9660
rect 13804 9650 13860 9660
rect 14364 9714 14420 9726
rect 14364 9662 14366 9714
rect 14418 9662 14420 9714
rect 13692 8990 13694 9042
rect 13746 8990 13748 9042
rect 12796 8146 12852 8428
rect 13132 8818 13188 8830
rect 13132 8766 13134 8818
rect 13186 8766 13188 8818
rect 13132 8428 13188 8766
rect 13692 8484 13748 8990
rect 14364 9044 14420 9662
rect 14476 9266 14532 9772
rect 14476 9214 14478 9266
rect 14530 9214 14532 9266
rect 14476 9202 14532 9214
rect 15036 9268 15092 9772
rect 15260 10610 15540 10612
rect 15260 10558 15374 10610
rect 15426 10558 15486 10610
rect 15538 10558 15540 10610
rect 15260 10556 15540 10558
rect 15148 9604 15204 9614
rect 15260 9604 15316 10556
rect 15372 10546 15428 10556
rect 15484 10546 15540 10556
rect 15708 10610 16100 10612
rect 15708 10558 16046 10610
rect 16098 10558 16100 10610
rect 15708 10556 16100 10558
rect 15148 9602 15316 9604
rect 15148 9550 15150 9602
rect 15202 9550 15316 9602
rect 15148 9548 15316 9550
rect 15148 9538 15204 9548
rect 15148 9268 15204 9278
rect 15036 9266 15204 9268
rect 15036 9214 15150 9266
rect 15202 9214 15204 9266
rect 15036 9212 15204 9214
rect 13132 8372 13412 8428
rect 12908 8260 12964 8270
rect 12908 8166 12964 8204
rect 13356 8260 13412 8372
rect 10556 7534 10558 7586
rect 10610 7534 10612 7586
rect 8876 7476 8932 7486
rect 8764 7474 8932 7476
rect 8764 7422 8878 7474
rect 8930 7422 8932 7474
rect 8764 7420 8932 7422
rect 8428 6486 8484 6524
rect 8540 6692 8596 6702
rect 8148 5964 8372 6020
rect 8092 5926 8148 5964
rect 8204 5684 8260 5694
rect 7196 5682 8260 5684
rect 7196 5630 7534 5682
rect 7586 5630 8206 5682
rect 8258 5630 8260 5682
rect 7196 5628 8260 5630
rect 7084 5516 7252 5572
rect 7196 5348 7252 5516
rect 6524 5346 7140 5348
rect 6524 5294 6526 5346
rect 6578 5294 7140 5346
rect 6524 5292 7140 5294
rect 6524 5282 6580 5292
rect 7084 5124 7140 5292
rect 7196 5346 7364 5348
rect 7196 5294 7198 5346
rect 7250 5294 7364 5346
rect 7196 5292 7364 5294
rect 7196 5282 7252 5292
rect 7308 5124 7364 5292
rect 7084 5122 7252 5124
rect 7084 5070 7086 5122
rect 7138 5070 7252 5122
rect 7084 5068 7252 5070
rect 7084 5058 7140 5068
rect 6076 4834 6132 4844
rect 6412 5010 6468 5022
rect 6412 4958 6414 5010
rect 6466 4958 6468 5010
rect 6300 4564 6356 4574
rect 6412 4564 6468 4958
rect 6532 4732 6796 4742
rect 6532 4666 6796 4676
rect 6412 4508 6580 4564
rect 6300 4340 6356 4508
rect 6412 4340 6468 4350
rect 5964 4284 6244 4340
rect 6300 4338 6468 4340
rect 6300 4286 6414 4338
rect 6466 4286 6468 4338
rect 6300 4284 6468 4286
rect 5964 3892 6020 4284
rect 5852 3836 6020 3892
rect 6076 4116 6132 4126
rect 5852 3554 5908 3836
rect 5852 3502 5854 3554
rect 5906 3502 5908 3554
rect 5852 3490 5908 3502
rect 5180 3378 5236 3388
rect 5740 3444 5796 3454
rect 5740 3350 5796 3388
rect 6076 800 6132 4060
rect 6188 3668 6244 4284
rect 6412 4274 6468 4284
rect 6524 4116 6580 4508
rect 7196 4562 7252 5068
rect 7196 4510 7198 4562
rect 7250 4510 7252 4562
rect 7196 4498 7252 4510
rect 6524 4022 6580 4060
rect 7084 4340 7140 4350
rect 7084 4116 7140 4284
rect 6412 3780 6468 3790
rect 6412 3778 6692 3780
rect 6412 3726 6414 3778
rect 6466 3726 6692 3778
rect 6412 3724 6692 3726
rect 6412 3714 6468 3724
rect 6188 3612 6356 3668
rect 6300 3556 6356 3612
rect 6524 3556 6580 3566
rect 6300 3554 6580 3556
rect 6300 3502 6526 3554
rect 6578 3502 6580 3554
rect 6300 3500 6580 3502
rect 6524 3490 6580 3500
rect 6636 3444 6692 3724
rect 7084 3778 7140 4060
rect 7084 3726 7086 3778
rect 7138 3726 7140 3778
rect 7084 3556 7140 3726
rect 7084 3490 7140 3500
rect 7196 3556 7252 3566
rect 7308 3556 7364 5068
rect 7532 4116 7588 5628
rect 8204 5618 8260 5628
rect 8540 5346 8596 6636
rect 8764 6692 8820 7420
rect 8876 7410 8932 7420
rect 9884 7474 9940 7486
rect 9884 7422 9886 7474
rect 9938 7422 9940 7474
rect 9192 7084 9456 7094
rect 9192 7018 9456 7028
rect 8764 6018 8820 6636
rect 8876 6916 8932 6926
rect 8876 6130 8932 6860
rect 9212 6692 9268 6702
rect 9212 6598 9268 6636
rect 9772 6692 9828 6702
rect 9884 6692 9940 7422
rect 9772 6690 9884 6692
rect 9772 6638 9774 6690
rect 9826 6638 9884 6690
rect 9772 6636 9884 6638
rect 8876 6078 8878 6130
rect 8930 6078 8932 6130
rect 8876 6066 8932 6078
rect 9100 6580 9156 6590
rect 8764 5966 8766 6018
rect 8818 5966 8820 6018
rect 8764 5954 8820 5966
rect 9100 5908 9156 6524
rect 9772 6132 9828 6636
rect 9884 6626 9940 6636
rect 9996 6916 10052 6926
rect 9884 6468 9940 6478
rect 9884 6374 9940 6412
rect 9884 6132 9940 6142
rect 9772 6130 9940 6132
rect 9772 6078 9886 6130
rect 9938 6078 9940 6130
rect 9772 6076 9940 6078
rect 9884 6066 9940 6076
rect 9100 5842 9156 5852
rect 9772 5908 9828 5918
rect 9772 5814 9828 5852
rect 9192 5516 9456 5526
rect 9192 5450 9456 5460
rect 8540 5294 8542 5346
rect 8594 5294 8596 5346
rect 7756 5124 7812 5134
rect 7868 5124 7924 5134
rect 7812 5122 7924 5124
rect 7812 5070 7870 5122
rect 7922 5070 7924 5122
rect 7812 5068 7924 5070
rect 7756 5030 7812 5068
rect 7868 5058 7924 5068
rect 8428 5124 8484 5134
rect 8540 5124 8596 5294
rect 9884 5348 9940 5358
rect 9996 5348 10052 6860
rect 10556 6916 10612 7534
rect 11340 7476 11396 8094
rect 12796 8094 12798 8146
rect 12850 8094 12852 8146
rect 11852 7868 12116 7878
rect 11852 7802 12116 7812
rect 10444 6692 10500 6702
rect 10444 6132 10500 6636
rect 10556 6468 10612 6860
rect 11228 7474 11396 7476
rect 11228 7422 11342 7474
rect 11394 7422 11396 7474
rect 11228 7420 11396 7422
rect 11228 6916 11284 7420
rect 11340 7410 11396 7420
rect 11900 7474 11956 7486
rect 11900 7422 11902 7474
rect 11954 7422 11956 7474
rect 10556 6402 10612 6412
rect 11116 6692 11172 6702
rect 10556 6132 10612 6142
rect 10444 6130 10612 6132
rect 10444 6078 10558 6130
rect 10610 6078 10612 6130
rect 10444 6076 10612 6078
rect 9884 5346 10052 5348
rect 9884 5294 9886 5346
rect 9938 5294 10052 5346
rect 9884 5292 10052 5294
rect 10444 5908 10500 5918
rect 9884 5282 9940 5292
rect 8428 5122 8540 5124
rect 8428 5070 8430 5122
rect 8482 5070 8540 5122
rect 8428 5068 8540 5070
rect 8428 5058 8484 5068
rect 8540 4564 8596 5068
rect 9100 5124 9156 5134
rect 9212 5124 9268 5134
rect 9156 5122 9268 5124
rect 9156 5070 9214 5122
rect 9266 5070 9268 5122
rect 9156 5068 9268 5070
rect 9100 5030 9156 5068
rect 9212 5058 9268 5068
rect 9660 5124 9716 5134
rect 10444 5124 10500 5852
rect 8428 4562 8596 4564
rect 8428 4510 8542 4562
rect 8594 4510 8596 4562
rect 8428 4508 8596 4510
rect 8428 4450 8484 4508
rect 8428 4398 8430 4450
rect 8482 4398 8484 4450
rect 8428 4386 8484 4398
rect 7756 4340 7812 4350
rect 7756 4246 7812 4284
rect 7868 4116 7924 4126
rect 7532 4114 7924 4116
rect 7532 4062 7870 4114
rect 7922 4062 7924 4114
rect 7532 4060 7924 4062
rect 7868 3778 7924 4060
rect 7868 3726 7870 3778
rect 7922 3726 7924 3778
rect 7868 3714 7924 3726
rect 7196 3554 7364 3556
rect 7196 3502 7198 3554
rect 7250 3502 7364 3554
rect 7196 3500 7364 3502
rect 7756 3556 7812 3566
rect 7196 3490 7252 3500
rect 7756 3462 7812 3500
rect 8428 3556 8484 3566
rect 8428 3462 8484 3500
rect 8540 3554 8596 4508
rect 9660 4452 9716 5068
rect 9996 5122 10500 5124
rect 9996 5070 10446 5122
rect 10498 5070 10500 5122
rect 9996 5068 10500 5070
rect 9772 5012 9828 5022
rect 9772 5010 9940 5012
rect 9772 4958 9774 5010
rect 9826 4958 9940 5010
rect 9772 4956 9940 4958
rect 9772 4946 9828 4956
rect 9772 4452 9828 4462
rect 9660 4450 9828 4452
rect 9660 4398 9774 4450
rect 9826 4398 9828 4450
rect 9660 4396 9828 4398
rect 9192 3948 9456 3958
rect 9192 3882 9456 3892
rect 8540 3502 8542 3554
rect 8594 3502 8596 3554
rect 8540 3490 8596 3502
rect 9660 3556 9716 3566
rect 9660 3462 9716 3500
rect 9772 3554 9828 4396
rect 9772 3502 9774 3554
rect 9826 3502 9828 3554
rect 9772 3490 9828 3502
rect 9884 4114 9940 4956
rect 9884 4062 9886 4114
rect 9938 4062 9940 4114
rect 9884 3556 9940 4062
rect 9884 3490 9940 3500
rect 6636 3378 6692 3388
rect 6532 3164 6796 3174
rect 6532 3098 6796 3108
rect 9996 800 10052 5068
rect 10444 5058 10500 5068
rect 10556 5346 10612 6076
rect 11116 6018 11172 6636
rect 11228 6130 11284 6860
rect 11788 6692 11844 6702
rect 11900 6692 11956 7422
rect 12572 7474 12628 7486
rect 12572 7422 12574 7474
rect 12626 7422 12628 7474
rect 11228 6078 11230 6130
rect 11282 6078 11284 6130
rect 11228 6066 11284 6078
rect 11676 6690 11900 6692
rect 11676 6638 11790 6690
rect 11842 6638 11900 6690
rect 11676 6636 11900 6638
rect 11116 5966 11118 6018
rect 11170 5966 11172 6018
rect 11116 5954 11172 5966
rect 11676 6020 11732 6636
rect 11788 6626 11844 6636
rect 11900 6626 11956 6636
rect 12012 7250 12068 7262
rect 12012 7198 12014 7250
rect 12066 7198 12068 7250
rect 12012 6916 12068 7198
rect 11900 6468 11956 6478
rect 12012 6468 12068 6860
rect 12572 7252 12628 7422
rect 12796 7476 12852 8094
rect 13356 7698 13412 8204
rect 13692 8258 13748 8428
rect 13692 8206 13694 8258
rect 13746 8206 13748 8258
rect 13692 8194 13748 8206
rect 13804 8818 13860 8830
rect 13804 8766 13806 8818
rect 13858 8766 13860 8818
rect 13804 8260 13860 8766
rect 13356 7646 13358 7698
rect 13410 7646 13412 7698
rect 13356 7634 13412 7646
rect 13244 7476 13300 7486
rect 12796 7474 13300 7476
rect 12796 7422 13246 7474
rect 13298 7422 13300 7474
rect 12796 7420 13300 7422
rect 12684 7252 12740 7262
rect 12572 7250 12740 7252
rect 12572 7198 12686 7250
rect 12738 7198 12740 7250
rect 12572 7196 12740 7198
rect 12460 6692 12516 6702
rect 12460 6598 12516 6636
rect 12572 6468 12628 7196
rect 12684 7186 12740 7196
rect 11900 6466 12628 6468
rect 11900 6414 11902 6466
rect 11954 6414 12574 6466
rect 12626 6414 12628 6466
rect 11900 6412 12628 6414
rect 11900 6402 11956 6412
rect 11852 6300 12116 6310
rect 11852 6234 12116 6244
rect 11900 6132 11956 6142
rect 12236 6132 12292 6412
rect 11900 6130 12292 6132
rect 11900 6078 11902 6130
rect 11954 6078 12292 6130
rect 11900 6076 12292 6078
rect 11900 6066 11956 6076
rect 11788 6020 11844 6030
rect 11676 6018 11844 6020
rect 11676 5966 11790 6018
rect 11842 5966 11844 6018
rect 11676 5964 11844 5966
rect 11788 5954 11844 5964
rect 12572 6018 12628 6412
rect 13244 6132 13300 7420
rect 13804 7364 13860 8204
rect 13916 8484 13972 8494
rect 13916 7588 13972 8428
rect 14364 8484 14420 8988
rect 15036 9044 15092 9054
rect 15036 8950 15092 8988
rect 15148 8820 15204 9212
rect 15260 9044 15316 9548
rect 15708 9826 15764 10556
rect 16044 10546 16100 10556
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9156 15764 9774
rect 16156 10386 16212 11230
rect 16716 10724 16772 10734
rect 16828 10724 16884 11340
rect 16940 11302 16996 11340
rect 17500 11396 17556 11406
rect 17612 11396 17668 11564
rect 17556 11340 17668 11396
rect 17500 11264 17556 11340
rect 17172 11004 17436 11014
rect 17172 10938 17436 10948
rect 16716 10722 16884 10724
rect 16716 10670 16718 10722
rect 16770 10670 16884 10722
rect 16716 10668 16884 10670
rect 17724 10722 17780 11564
rect 18172 11396 18228 12236
rect 18396 12198 18452 12236
rect 18956 12292 19012 13134
rect 19180 13188 19236 13198
rect 19180 12852 19236 13132
rect 19628 12964 19684 13468
rect 19832 13356 20096 13366
rect 19832 13290 20096 13300
rect 19628 12908 19908 12964
rect 19516 12852 19572 12862
rect 19180 12850 19684 12852
rect 19180 12798 19518 12850
rect 19570 12798 19684 12850
rect 19180 12796 19684 12798
rect 19180 12402 19236 12796
rect 19516 12786 19572 12796
rect 19180 12350 19182 12402
rect 19234 12350 19236 12402
rect 19068 12292 19124 12302
rect 19012 12290 19124 12292
rect 19012 12238 19070 12290
rect 19122 12238 19124 12290
rect 19012 12236 19124 12238
rect 18508 11954 18564 11966
rect 18508 11902 18510 11954
rect 18562 11902 18564 11954
rect 18508 11732 18564 11902
rect 18172 11394 18452 11396
rect 18172 11342 18174 11394
rect 18226 11342 18452 11394
rect 18172 11340 18452 11342
rect 18172 11330 18228 11340
rect 17724 10670 17726 10722
rect 17778 10670 17780 10722
rect 16716 10658 16772 10668
rect 16156 10334 16158 10386
rect 16210 10334 16212 10386
rect 15260 8978 15316 8988
rect 15596 9154 15764 9156
rect 15596 9102 15710 9154
rect 15762 9102 15764 9154
rect 15596 9100 15764 9102
rect 15036 8764 15204 8820
rect 14512 8652 14776 8662
rect 14512 8586 14776 8596
rect 14364 8258 14420 8428
rect 14364 8206 14366 8258
rect 14418 8206 14420 8258
rect 14364 7700 14420 8206
rect 14476 8260 14532 8270
rect 14476 8166 14532 8204
rect 15036 8260 15092 8764
rect 15148 8484 15204 8522
rect 15148 8372 15316 8428
rect 15036 8166 15092 8204
rect 14700 7700 14756 7710
rect 14364 7698 14980 7700
rect 14364 7646 14702 7698
rect 14754 7646 14980 7698
rect 14364 7644 14980 7646
rect 14700 7634 14756 7644
rect 13916 7586 14196 7588
rect 13916 7534 13918 7586
rect 13970 7534 14196 7586
rect 13916 7532 14196 7534
rect 13916 7522 13972 7532
rect 14028 7364 14084 7374
rect 13804 7362 14084 7364
rect 13804 7310 14030 7362
rect 14082 7310 14084 7362
rect 13804 7308 14084 7310
rect 14028 6916 14084 7308
rect 14028 6850 14084 6860
rect 14140 6690 14196 7532
rect 14588 7476 14644 7486
rect 14364 7474 14644 7476
rect 14364 7422 14590 7474
rect 14642 7422 14644 7474
rect 14364 7420 14644 7422
rect 14252 6916 14308 6926
rect 14364 6916 14420 7420
rect 14588 7410 14644 7420
rect 14512 7084 14776 7094
rect 14512 7018 14776 7028
rect 14308 6860 14420 6916
rect 14588 6916 14644 6926
rect 14252 6822 14308 6860
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 13356 6132 13412 6142
rect 13244 6130 13412 6132
rect 13244 6078 13358 6130
rect 13410 6078 13412 6130
rect 13244 6076 13412 6078
rect 13356 6066 13412 6076
rect 14028 6132 14084 6142
rect 14140 6132 14196 6638
rect 14028 6130 14196 6132
rect 14028 6078 14030 6130
rect 14082 6078 14196 6130
rect 14028 6076 14196 6078
rect 14028 6066 14084 6076
rect 12572 5966 12574 6018
rect 12626 5966 12628 6018
rect 10556 5294 10558 5346
rect 10610 5294 10612 5346
rect 10444 4452 10500 4462
rect 10556 4452 10612 5294
rect 11452 5124 11508 5134
rect 11564 5124 11620 5134
rect 11452 5122 11564 5124
rect 11452 5070 11454 5122
rect 11506 5070 11564 5122
rect 11452 5068 11564 5070
rect 11452 5058 11508 5068
rect 11564 5030 11620 5068
rect 12124 5124 12180 5134
rect 12124 5010 12180 5068
rect 12124 4958 12126 5010
rect 12178 4958 12180 5010
rect 12124 4900 12180 4958
rect 12572 5012 12628 5966
rect 13244 5906 13300 5918
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 12684 5682 12740 5694
rect 12684 5630 12686 5682
rect 12738 5630 12740 5682
rect 12684 5236 12740 5630
rect 13244 5236 13300 5854
rect 12684 5180 13300 5236
rect 13916 5906 13972 5918
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 12796 5012 12852 5022
rect 12572 5010 12852 5012
rect 12572 4958 12798 5010
rect 12850 4958 12852 5010
rect 12572 4956 12852 4958
rect 12236 4900 12292 4910
rect 12348 4900 12404 4910
rect 12124 4898 12348 4900
rect 12124 4846 12238 4898
rect 12290 4846 12348 4898
rect 12124 4844 12348 4846
rect 12236 4834 12292 4844
rect 11852 4732 12116 4742
rect 11852 4666 12116 4676
rect 10444 4450 10612 4452
rect 10444 4398 10446 4450
rect 10498 4398 10612 4450
rect 10444 4396 10612 4398
rect 10444 4386 10500 4396
rect 11116 4340 11172 4350
rect 12348 4340 12404 4844
rect 12684 4340 12740 4956
rect 12796 4946 12852 4956
rect 12908 4900 12964 5180
rect 12908 4806 12964 4844
rect 13916 5012 13972 5854
rect 14140 5346 14196 6076
rect 14588 6692 14644 6860
rect 14924 6914 14980 7644
rect 15260 7586 15316 8372
rect 15596 8260 15652 9100
rect 15708 9090 15764 9100
rect 15820 9604 15876 9614
rect 16156 9604 16212 10334
rect 16828 10388 16884 10398
rect 15820 9602 16212 9604
rect 15820 9550 15822 9602
rect 15874 9550 16212 9602
rect 15820 9548 16212 9550
rect 16380 9714 16436 9726
rect 16380 9662 16382 9714
rect 16434 9662 16436 9714
rect 15820 8820 15876 9548
rect 16380 9044 16436 9662
rect 16828 9716 16884 10332
rect 17724 9828 17780 10670
rect 18284 11172 18340 11182
rect 17836 10388 17892 10398
rect 17836 10294 17892 10332
rect 18284 10388 18340 11116
rect 18284 10322 18340 10332
rect 18396 10722 18452 11340
rect 18508 11172 18564 11676
rect 18844 11396 18900 11406
rect 18956 11396 19012 12236
rect 19068 12226 19124 12236
rect 18844 11394 18956 11396
rect 18844 11342 18846 11394
rect 18898 11342 18956 11394
rect 18844 11340 18956 11342
rect 19012 11340 19124 11396
rect 18844 11330 18900 11340
rect 18956 11330 19012 11340
rect 18508 11106 18564 11116
rect 18956 11172 19012 11182
rect 18956 11078 19012 11116
rect 18396 10670 18398 10722
rect 18450 10670 18452 10722
rect 18396 10052 18452 10670
rect 19068 10722 19124 11340
rect 19068 10670 19070 10722
rect 19122 10670 19124 10722
rect 19068 10658 19124 10670
rect 19180 10834 19236 12350
rect 19628 12738 19684 12796
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19628 12292 19684 12686
rect 19852 12402 19908 12908
rect 22492 12572 22756 12582
rect 22492 12506 22756 12516
rect 19852 12350 19854 12402
rect 19906 12350 19908 12402
rect 19852 12338 19908 12350
rect 19740 12292 19796 12302
rect 19628 12236 19740 12292
rect 19628 11618 19684 12236
rect 19740 12160 19796 12236
rect 20412 12292 20468 12302
rect 20524 12292 20580 12302
rect 20468 12290 20580 12292
rect 20468 12238 20526 12290
rect 20578 12238 20580 12290
rect 20468 12236 20580 12238
rect 20412 12198 20468 12236
rect 20524 12226 20580 12236
rect 21084 12292 21140 12302
rect 19832 11788 20096 11798
rect 19832 11722 20096 11732
rect 19628 11566 19630 11618
rect 19682 11566 19684 11618
rect 19516 11396 19572 11406
rect 19516 11302 19572 11340
rect 19180 10782 19182 10834
rect 19234 10782 19236 10834
rect 18508 10388 18564 10398
rect 18508 10294 18564 10332
rect 18508 10052 18564 10062
rect 18396 10050 18564 10052
rect 18396 9998 18510 10050
rect 18562 9998 18564 10050
rect 18396 9996 18564 9998
rect 18508 9986 18564 9996
rect 17836 9828 17892 9838
rect 17724 9826 17892 9828
rect 17724 9774 17838 9826
rect 17890 9774 17892 9826
rect 17724 9772 17892 9774
rect 17836 9762 17892 9772
rect 19068 9828 19124 9838
rect 19180 9828 19236 10782
rect 19068 9826 19236 9828
rect 19068 9774 19070 9826
rect 19122 9774 19236 9826
rect 19068 9772 19236 9774
rect 19628 10724 19684 11566
rect 19852 11396 19908 11406
rect 19852 10834 19908 11340
rect 19852 10782 19854 10834
rect 19906 10782 19908 10834
rect 19740 10724 19796 10734
rect 19628 10722 19796 10724
rect 19628 10670 19742 10722
rect 19794 10670 19796 10722
rect 19628 10668 19796 10670
rect 19628 9828 19684 10668
rect 19740 10658 19796 10668
rect 19852 10724 19908 10782
rect 19852 10658 19908 10668
rect 20188 11282 20244 11294
rect 20188 11230 20190 11282
rect 20242 11230 20244 11282
rect 20188 10724 20244 11230
rect 20300 11170 20356 11182
rect 20300 11118 20302 11170
rect 20354 11118 20356 11170
rect 20300 10724 20356 11118
rect 20412 10724 20468 10734
rect 20300 10722 20468 10724
rect 20300 10670 20414 10722
rect 20466 10670 20468 10722
rect 20300 10668 20468 10670
rect 20188 10658 20244 10668
rect 19832 10220 20096 10230
rect 19832 10154 20096 10164
rect 19852 10052 19908 10062
rect 19740 9828 19796 9838
rect 19628 9826 19796 9828
rect 19628 9774 19742 9826
rect 19794 9774 19796 9826
rect 19628 9772 19796 9774
rect 17052 9716 17108 9726
rect 16828 9714 17108 9716
rect 16828 9662 17054 9714
rect 17106 9662 17108 9714
rect 16828 9660 17108 9662
rect 15596 8194 15652 8204
rect 15708 8818 15876 8820
rect 15708 8766 15822 8818
rect 15874 8766 15876 8818
rect 15708 8764 15876 8766
rect 15708 8484 15764 8764
rect 15820 8754 15876 8764
rect 16268 9042 16436 9044
rect 16268 8990 16382 9042
rect 16434 8990 16436 9042
rect 16268 8988 16436 8990
rect 15260 7534 15262 7586
rect 15314 7534 15316 7586
rect 15260 7522 15316 7534
rect 15708 8146 15764 8428
rect 15708 8094 15710 8146
rect 15762 8094 15764 8146
rect 15372 7252 15428 7262
rect 14924 6862 14926 6914
rect 14978 6862 14980 6914
rect 14812 6692 14868 6702
rect 14588 6690 14868 6692
rect 14588 6638 14814 6690
rect 14866 6638 14868 6690
rect 14588 6636 14868 6638
rect 14588 6132 14644 6636
rect 14812 6626 14868 6636
rect 14700 6132 14756 6142
rect 14588 6130 14756 6132
rect 14588 6078 14702 6130
rect 14754 6078 14756 6130
rect 14588 6076 14756 6078
rect 14588 6020 14644 6076
rect 14700 6066 14756 6076
rect 14140 5294 14142 5346
rect 14194 5294 14196 5346
rect 14140 5282 14196 5294
rect 14364 6018 14644 6020
rect 14364 5966 14590 6018
rect 14642 5966 14644 6018
rect 14364 5964 14644 5966
rect 14028 5012 14084 5022
rect 13916 5010 14084 5012
rect 13916 4958 14030 5010
rect 14082 4958 14084 5010
rect 13916 4956 14084 4958
rect 13020 4340 13076 4350
rect 13692 4340 13748 4350
rect 11116 4338 11284 4340
rect 11116 4286 11118 4338
rect 11170 4286 11284 4338
rect 11116 4284 11284 4286
rect 11116 4274 11172 4284
rect 10556 4116 10612 4126
rect 10444 4114 10612 4116
rect 10444 4062 10558 4114
rect 10610 4062 10612 4114
rect 10444 4060 10612 4062
rect 10332 3556 10388 3566
rect 10444 3556 10500 4060
rect 10556 4050 10612 4060
rect 11228 4114 11284 4284
rect 12348 4338 12516 4340
rect 12348 4286 12350 4338
rect 12402 4286 12516 4338
rect 12348 4284 12516 4286
rect 12684 4338 13748 4340
rect 12684 4286 13022 4338
rect 13074 4286 13694 4338
rect 13746 4286 13748 4338
rect 12684 4284 13748 4286
rect 12348 4274 12404 4284
rect 11228 4062 11230 4114
rect 11282 4062 11284 4114
rect 10388 3554 10500 3556
rect 10388 3502 10446 3554
rect 10498 3502 10500 3554
rect 10388 3500 10500 3502
rect 10332 3462 10388 3500
rect 10444 3490 10500 3500
rect 11116 3556 11172 3566
rect 11228 3556 11284 4062
rect 12460 4116 12516 4284
rect 13020 4274 13076 4284
rect 12460 4022 12516 4060
rect 13132 4116 13188 4126
rect 13132 4022 13188 4060
rect 11172 3500 11284 3556
rect 11676 3556 11732 3566
rect 11116 3462 11172 3500
rect 11676 3462 11732 3500
rect 11004 3444 11060 3454
rect 11004 3350 11060 3388
rect 11788 3444 11844 3454
rect 11788 3350 11844 3388
rect 11852 3164 12116 3174
rect 11852 3098 12116 3108
rect 13692 2996 13748 4284
rect 13804 4116 13860 4126
rect 13916 4116 13972 4956
rect 14028 4946 14084 4956
rect 13860 4060 13972 4116
rect 13804 3984 13860 4060
rect 13916 3444 13972 4060
rect 14364 4450 14420 5964
rect 14588 5954 14644 5964
rect 14512 5516 14776 5526
rect 14512 5450 14776 5460
rect 14812 5348 14868 5358
rect 14924 5348 14980 6862
rect 15260 7250 15428 7252
rect 15260 7198 15374 7250
rect 15426 7198 15428 7250
rect 15260 7196 15428 7198
rect 15260 6916 15316 7196
rect 15372 7186 15428 7196
rect 15260 6692 15316 6860
rect 15596 6916 15652 6926
rect 15708 6916 15764 8094
rect 15820 8260 15876 8270
rect 15820 7588 15876 8204
rect 16268 8260 16324 8988
rect 16380 8978 16436 8988
rect 16492 9604 16548 9614
rect 16492 8820 16548 9548
rect 16268 8194 16324 8204
rect 16380 8818 16548 8820
rect 16380 8766 16494 8818
rect 16546 8766 16548 8818
rect 16380 8764 16548 8766
rect 16380 8484 16436 8764
rect 16492 8754 16548 8764
rect 16380 8146 16436 8428
rect 16492 8260 16548 8270
rect 16492 8166 16548 8204
rect 17052 8260 17108 9660
rect 18396 9714 18452 9726
rect 18396 9662 18398 9714
rect 18450 9662 18452 9714
rect 17164 9604 17220 9642
rect 17164 9538 17220 9548
rect 17724 9602 17780 9614
rect 17724 9550 17726 9602
rect 17778 9550 17780 9602
rect 17172 9436 17436 9446
rect 17172 9370 17436 9380
rect 17724 9154 17780 9550
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17164 8484 17220 8522
rect 17724 8428 17780 9102
rect 18396 9042 18452 9662
rect 18396 8990 18398 9042
rect 18450 8990 18452 9042
rect 17164 8418 17220 8428
rect 17052 8166 17108 8204
rect 17612 8372 17780 8428
rect 17836 8818 17892 8830
rect 17836 8766 17838 8818
rect 17890 8766 17892 8818
rect 17836 8484 17892 8766
rect 17836 8418 17892 8428
rect 18396 8372 18452 8990
rect 19068 9154 19124 9772
rect 19068 9102 19070 9154
rect 19122 9102 19124 9154
rect 18508 8818 18564 8830
rect 18508 8766 18510 8818
rect 18562 8766 18564 8818
rect 18508 8484 18564 8766
rect 18508 8418 18564 8428
rect 18956 8820 19012 8830
rect 18956 8484 19012 8764
rect 19068 8484 19124 9102
rect 19180 9604 19236 9614
rect 19180 8820 19236 9548
rect 19740 9268 19796 9772
rect 19852 9604 19908 9996
rect 19852 9510 19908 9548
rect 20412 9826 20468 10668
rect 21084 10724 21140 12236
rect 21084 10592 21140 10668
rect 21756 11172 21812 11182
rect 21756 10722 21812 11116
rect 22492 11004 22756 11014
rect 22492 10938 22756 10948
rect 21756 10670 21758 10722
rect 21810 10670 21812 10722
rect 21756 10658 21812 10670
rect 21868 10724 21924 10734
rect 20524 10388 20580 10398
rect 21196 10388 21252 10398
rect 20524 10386 21252 10388
rect 20524 10334 20526 10386
rect 20578 10334 21198 10386
rect 21250 10334 21252 10386
rect 20524 10332 21252 10334
rect 20524 10052 20580 10332
rect 21196 10322 21252 10332
rect 21868 10276 21924 10668
rect 20524 9920 20580 9996
rect 21756 10220 21924 10276
rect 21756 10050 21812 10220
rect 21756 9998 21758 10050
rect 21810 9998 21812 10050
rect 20412 9774 20414 9826
rect 20466 9774 20468 9826
rect 19852 9268 19908 9278
rect 20412 9268 20468 9774
rect 21644 9828 21700 9838
rect 21756 9828 21812 9998
rect 21644 9826 21812 9828
rect 21644 9774 21646 9826
rect 21698 9774 21812 9826
rect 21644 9772 21812 9774
rect 21644 9762 21700 9772
rect 20524 9268 20580 9278
rect 19740 9266 20580 9268
rect 19740 9214 19854 9266
rect 19906 9214 20526 9266
rect 20578 9214 20580 9266
rect 19740 9212 20580 9214
rect 19852 9202 19908 9212
rect 20412 9154 20468 9212
rect 20524 9202 20580 9212
rect 20412 9102 20414 9154
rect 20466 9102 20468 9154
rect 20412 9090 20468 9102
rect 19740 9044 19796 9054
rect 19180 8726 19236 8764
rect 19628 9042 19796 9044
rect 19628 8990 19742 9042
rect 19794 8990 19796 9042
rect 19628 8988 19796 8990
rect 19180 8484 19236 8494
rect 19068 8482 19236 8484
rect 19068 8430 19182 8482
rect 19234 8430 19236 8482
rect 19068 8428 19236 8430
rect 17612 8260 17668 8372
rect 17612 8194 17668 8204
rect 18396 8258 18452 8316
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 16380 8094 16382 8146
rect 16434 8094 16436 8146
rect 16380 7700 16436 8094
rect 17724 8148 17780 8158
rect 17724 8146 17892 8148
rect 17724 8094 17726 8146
rect 17778 8094 17892 8146
rect 17724 8092 17892 8094
rect 17724 8082 17780 8092
rect 17172 7868 17436 7878
rect 17172 7802 17436 7812
rect 16716 7700 16772 7710
rect 17836 7700 17892 8092
rect 16380 7698 16772 7700
rect 16380 7646 16718 7698
rect 16770 7646 16772 7698
rect 16380 7644 16772 7646
rect 16716 7634 16772 7644
rect 17612 7644 17836 7700
rect 15932 7588 15988 7598
rect 15820 7586 15988 7588
rect 15820 7534 15934 7586
rect 15986 7534 15988 7586
rect 15820 7532 15988 7534
rect 15932 7522 15988 7532
rect 16604 7476 16660 7486
rect 16604 7382 16660 7420
rect 17612 7476 17668 7644
rect 17836 7606 17892 7644
rect 18396 7700 18452 8206
rect 18508 7700 18564 7710
rect 18452 7698 18564 7700
rect 18452 7646 18510 7698
rect 18562 7646 18564 7698
rect 18452 7644 18564 7646
rect 18396 7634 18452 7644
rect 18508 7634 18564 7644
rect 16044 7250 16100 7262
rect 16044 7198 16046 7250
rect 16098 7198 16100 7250
rect 16044 6916 16100 7198
rect 15596 6914 16100 6916
rect 15596 6862 15598 6914
rect 15650 6862 16100 6914
rect 15596 6860 16100 6862
rect 17612 6914 17668 7420
rect 17612 6862 17614 6914
rect 17666 6862 17668 6914
rect 15596 6850 15652 6860
rect 17612 6850 17668 6862
rect 17724 7474 17780 7486
rect 17724 7422 17726 7474
rect 17778 7422 17780 7474
rect 17724 7364 17780 7422
rect 15484 6692 15540 6702
rect 15260 6690 15540 6692
rect 15260 6638 15486 6690
rect 15538 6638 15540 6690
rect 15260 6636 15540 6638
rect 15260 6132 15316 6636
rect 15484 6626 15540 6636
rect 16156 6580 16212 6590
rect 16268 6580 16324 6590
rect 16828 6580 16884 6590
rect 16940 6580 16996 6590
rect 16044 6578 16940 6580
rect 16044 6526 16158 6578
rect 16210 6526 16270 6578
rect 16322 6526 16830 6578
rect 16882 6526 16940 6578
rect 16044 6524 16940 6526
rect 15372 6132 15428 6142
rect 16044 6132 16100 6524
rect 16156 6514 16212 6524
rect 16268 6514 16324 6524
rect 15260 6130 16100 6132
rect 15260 6078 15374 6130
rect 15426 6078 16046 6130
rect 16098 6078 16100 6130
rect 15260 6076 16100 6078
rect 15260 6018 15316 6076
rect 15372 6066 15428 6076
rect 15260 5966 15262 6018
rect 15314 5966 15316 6018
rect 15260 5954 15316 5966
rect 14812 5346 15204 5348
rect 14812 5294 14814 5346
rect 14866 5294 15204 5346
rect 14812 5292 15204 5294
rect 14812 5282 14868 5292
rect 14364 4398 14366 4450
rect 14418 4398 14420 4450
rect 14364 3780 14420 4398
rect 14700 5012 14756 5022
rect 14476 4340 14532 4350
rect 14476 4246 14532 4284
rect 14700 4340 14756 4956
rect 15148 4564 15204 5292
rect 15484 5346 15540 6076
rect 15932 6018 15988 6076
rect 16044 6066 16100 6076
rect 16604 6132 16660 6524
rect 16828 6514 16884 6524
rect 16940 6448 16996 6524
rect 17500 6580 17556 6590
rect 17724 6580 17780 7308
rect 18396 7474 18452 7486
rect 18396 7422 18398 7474
rect 18450 7422 18452 7474
rect 18396 7364 18452 7422
rect 18956 7476 19012 8428
rect 19180 8372 19236 8428
rect 19180 8306 19236 8316
rect 19068 8260 19124 8270
rect 19068 8166 19124 8204
rect 19628 8260 19684 8988
rect 19740 8978 19796 8988
rect 19832 8652 20096 8662
rect 19832 8586 20096 8596
rect 21756 8428 21812 9772
rect 22492 9436 22756 9446
rect 22492 9370 22756 9380
rect 21756 8372 22036 8428
rect 19740 8260 19796 8270
rect 19852 8260 19908 8270
rect 19684 8258 19908 8260
rect 19684 8206 19742 8258
rect 19794 8206 19854 8258
rect 19906 8206 19908 8258
rect 19684 8204 19908 8206
rect 19628 8194 19684 8204
rect 19740 8194 19796 8204
rect 19852 8194 19908 8204
rect 20524 8146 20580 8158
rect 20524 8094 20526 8146
rect 20578 8094 20580 8146
rect 20412 8036 20468 8046
rect 20524 8036 20580 8094
rect 20412 8034 20580 8036
rect 20412 7982 20414 8034
rect 20466 7982 20580 8034
rect 20412 7980 20580 7982
rect 20412 7970 20468 7980
rect 19068 7476 19124 7486
rect 19740 7476 19796 7486
rect 20412 7476 20468 7486
rect 18956 7474 19124 7476
rect 18956 7422 19070 7474
rect 19122 7422 19124 7474
rect 18956 7420 19124 7422
rect 18396 7298 18452 7308
rect 18956 6692 19012 6702
rect 18956 6598 19012 6636
rect 17556 6524 17780 6580
rect 18172 6578 18228 6590
rect 18172 6526 18174 6578
rect 18226 6526 18228 6578
rect 17500 6486 17556 6524
rect 17172 6300 17436 6310
rect 17172 6234 17436 6244
rect 16716 6132 16772 6142
rect 16604 6130 16772 6132
rect 16604 6078 16718 6130
rect 16770 6078 16772 6130
rect 16604 6076 16772 6078
rect 15932 5966 15934 6018
rect 15986 5966 15988 6018
rect 15932 5954 15988 5966
rect 16604 6018 16660 6076
rect 16716 6066 16772 6076
rect 16604 5966 16606 6018
rect 16658 5966 16660 6018
rect 16604 5954 16660 5966
rect 15484 5294 15486 5346
rect 15538 5294 15540 5346
rect 15372 5124 15428 5134
rect 15484 5124 15540 5294
rect 15372 5122 15540 5124
rect 15372 5070 15374 5122
rect 15426 5070 15540 5122
rect 15372 5068 15540 5070
rect 16156 5124 16212 5134
rect 15372 5058 15428 5068
rect 16044 5012 16100 5022
rect 16044 4918 16100 4956
rect 16156 4898 16212 5068
rect 16828 5124 16884 5134
rect 16828 5030 16884 5068
rect 17388 5124 17444 5134
rect 17388 5030 17444 5068
rect 17612 5124 17668 6524
rect 18172 6132 18228 6526
rect 18844 6578 18900 6590
rect 18844 6526 18846 6578
rect 18898 6526 18900 6578
rect 18284 6468 18340 6478
rect 18844 6468 18900 6526
rect 18284 6466 18900 6468
rect 18284 6414 18286 6466
rect 18338 6414 18900 6466
rect 18284 6412 18900 6414
rect 18284 6402 18340 6412
rect 16716 5012 16772 5022
rect 16716 4918 16772 4956
rect 16156 4846 16158 4898
rect 16210 4846 16212 4898
rect 15820 4564 15876 4574
rect 16156 4564 16212 4846
rect 17500 4898 17556 4910
rect 17500 4846 17502 4898
rect 17554 4846 17556 4898
rect 17172 4732 17436 4742
rect 17172 4666 17436 4676
rect 15148 4562 16436 4564
rect 15148 4510 15150 4562
rect 15202 4510 15822 4562
rect 15874 4510 16436 4562
rect 15148 4508 16436 4510
rect 15148 4498 15204 4508
rect 15820 4498 15876 4508
rect 16380 4450 16436 4508
rect 16380 4398 16382 4450
rect 16434 4398 16436 4450
rect 16380 4386 16436 4398
rect 16492 4452 16548 4462
rect 16492 4358 16548 4396
rect 17500 4452 17556 4846
rect 17612 4788 17668 5068
rect 17724 6076 18228 6132
rect 17724 5906 17780 6076
rect 17724 5854 17726 5906
rect 17778 5854 17780 5906
rect 17724 5012 17780 5854
rect 17836 5908 17892 5918
rect 17836 5682 17892 5852
rect 18396 5908 18452 6412
rect 18844 6020 18900 6412
rect 19068 6020 19124 7420
rect 19516 7474 20468 7476
rect 19516 7422 19742 7474
rect 19794 7422 20414 7474
rect 20466 7422 20468 7474
rect 19516 7420 20468 7422
rect 19180 7250 19236 7262
rect 19180 7198 19182 7250
rect 19234 7198 19236 7250
rect 19180 6692 19236 7198
rect 19180 6626 19236 6636
rect 19516 6578 19572 7420
rect 19740 7410 19796 7420
rect 20412 7410 20468 7420
rect 19852 7252 19908 7262
rect 19516 6526 19518 6578
rect 19570 6526 19572 6578
rect 19516 6020 19572 6526
rect 18844 6018 19572 6020
rect 18844 5966 19070 6018
rect 19122 5966 19572 6018
rect 18844 5964 19572 5966
rect 19628 7250 19908 7252
rect 19628 7198 19854 7250
rect 19906 7198 19908 7250
rect 19628 7196 19908 7198
rect 19628 6914 19684 7196
rect 19852 7186 19908 7196
rect 20524 7250 20580 7980
rect 20524 7198 20526 7250
rect 20578 7198 20580 7250
rect 19832 7084 20096 7094
rect 19832 7018 20096 7028
rect 19628 6862 19630 6914
rect 19682 6862 19684 6914
rect 19628 6692 19684 6862
rect 19628 6020 19684 6636
rect 20300 6578 20356 6590
rect 20300 6526 20302 6578
rect 20354 6526 20356 6578
rect 20188 6466 20244 6478
rect 20188 6414 20190 6466
rect 20242 6414 20244 6466
rect 19740 6020 19796 6030
rect 19628 6018 19796 6020
rect 19628 5966 19742 6018
rect 19794 5966 19796 6018
rect 19628 5964 19796 5966
rect 19068 5954 19124 5964
rect 19628 5908 19684 5964
rect 19740 5954 19796 5964
rect 18396 5814 18452 5852
rect 19180 5852 19684 5908
rect 17836 5630 17838 5682
rect 17890 5630 17892 5682
rect 17836 5124 17892 5630
rect 18172 5796 18228 5806
rect 18172 5348 18228 5740
rect 18508 5796 18564 5806
rect 18508 5702 18564 5740
rect 18732 5796 18788 5806
rect 18172 5346 18452 5348
rect 18172 5294 18174 5346
rect 18226 5294 18452 5346
rect 18172 5292 18452 5294
rect 18172 5282 18228 5292
rect 18060 5124 18116 5134
rect 17836 5122 18116 5124
rect 17836 5070 18062 5122
rect 18114 5070 18116 5122
rect 17836 5068 18116 5070
rect 18060 5058 18116 5068
rect 17724 4946 17780 4956
rect 17612 4732 17892 4788
rect 17836 4562 17892 4732
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17724 4452 17780 4462
rect 17500 4396 17724 4452
rect 14700 4274 14756 4284
rect 15036 4340 15092 4350
rect 15036 4246 15092 4284
rect 15708 4340 15764 4350
rect 14512 3948 14776 3958
rect 14512 3882 14776 3892
rect 14364 3724 14644 3780
rect 14588 3668 14644 3724
rect 14588 3612 15652 3668
rect 14588 3554 14644 3612
rect 14588 3502 14590 3554
rect 14642 3502 14644 3554
rect 14588 3490 14644 3502
rect 15260 3554 15316 3612
rect 15260 3502 15262 3554
rect 15314 3502 15316 3554
rect 15260 3490 15316 3502
rect 15596 3554 15652 3612
rect 15596 3502 15598 3554
rect 15650 3502 15652 3554
rect 15596 3490 15652 3502
rect 14028 3444 14084 3454
rect 13916 3442 14028 3444
rect 13916 3390 13918 3442
rect 13970 3390 14028 3442
rect 13916 3388 14028 3390
rect 13916 3378 13972 3388
rect 14028 3350 14084 3388
rect 14700 3444 14756 3454
rect 14700 3350 14756 3388
rect 15372 3444 15428 3454
rect 15372 3350 15428 3388
rect 15708 3444 15764 4284
rect 15932 3612 16660 3668
rect 15820 3556 15876 3566
rect 15932 3556 15988 3612
rect 15820 3554 15988 3556
rect 15820 3502 15822 3554
rect 15874 3502 15988 3554
rect 15820 3500 15988 3502
rect 15820 3490 15876 3500
rect 15708 3378 15764 3388
rect 15932 3442 15988 3500
rect 16604 3554 16660 3612
rect 16604 3502 16606 3554
rect 16658 3502 16660 3554
rect 16604 3490 16660 3502
rect 17500 3554 17556 4396
rect 17724 4358 17780 4396
rect 17836 4228 17892 4510
rect 17612 4172 17892 4228
rect 18172 4452 18228 4462
rect 17612 3778 17668 4172
rect 17612 3726 17614 3778
rect 17666 3726 17668 3778
rect 17612 3714 17668 3726
rect 17500 3502 17502 3554
rect 17554 3502 17556 3554
rect 17500 3490 17556 3502
rect 18172 3554 18228 4396
rect 18396 4452 18452 5292
rect 18508 5124 18564 5134
rect 18508 4562 18564 5068
rect 18732 5122 18788 5740
rect 19180 5796 19236 5852
rect 19180 5664 19236 5740
rect 18732 5070 18734 5122
rect 18786 5070 18788 5122
rect 18732 5058 18788 5070
rect 18844 5124 18900 5134
rect 18844 5030 18900 5068
rect 19068 5124 19124 5134
rect 18508 4510 18510 4562
rect 18562 4510 18564 4562
rect 18508 4498 18564 4510
rect 19068 4452 19124 5068
rect 19404 5124 19460 5852
rect 19852 5684 19908 5760
rect 19628 5628 19852 5684
rect 19516 5236 19572 5246
rect 19628 5236 19684 5628
rect 19852 5618 19908 5628
rect 19832 5516 20096 5526
rect 19832 5450 20096 5460
rect 19572 5180 19684 5236
rect 20188 5346 20244 6414
rect 20300 5684 20356 6526
rect 20300 5618 20356 5628
rect 20412 5908 20468 5918
rect 20524 5908 20580 7198
rect 20412 5906 20580 5908
rect 20412 5854 20414 5906
rect 20466 5854 20580 5906
rect 20412 5852 20580 5854
rect 21084 7474 21140 7486
rect 21084 7422 21086 7474
rect 21138 7422 21140 7474
rect 21084 5906 21140 7422
rect 21084 5854 21086 5906
rect 21138 5854 21140 5906
rect 20188 5294 20190 5346
rect 20242 5294 20244 5346
rect 19516 5142 19572 5180
rect 19404 4992 19460 5068
rect 19852 5124 19908 5134
rect 19852 4564 19908 5068
rect 18396 4320 18452 4396
rect 18844 4450 19124 4452
rect 18844 4398 19070 4450
rect 19122 4398 19124 4450
rect 18844 4396 19124 4398
rect 18172 3502 18174 3554
rect 18226 3502 18228 3554
rect 18172 3490 18228 3502
rect 18844 3554 18900 4396
rect 19068 4386 19124 4396
rect 19628 4562 19908 4564
rect 19628 4510 19854 4562
rect 19906 4510 19908 4562
rect 19628 4508 19908 4510
rect 20076 5124 20132 5134
rect 20076 4564 20132 5068
rect 20188 5012 20244 5294
rect 20412 5348 20468 5852
rect 20524 5684 20580 5694
rect 20524 5590 20580 5628
rect 20412 5292 20580 5348
rect 20188 4946 20244 4956
rect 20412 5012 20468 5022
rect 20076 4508 20356 4564
rect 18844 3502 18846 3554
rect 18898 3502 18900 3554
rect 18844 3490 18900 3502
rect 19180 4340 19236 4350
rect 19180 4114 19236 4284
rect 19180 4062 19182 4114
rect 19234 4062 19236 4114
rect 15932 3390 15934 3442
rect 15986 3390 15988 3442
rect 15932 3378 15988 3390
rect 16044 3444 16100 3454
rect 16044 3350 16100 3388
rect 16716 3444 16772 3454
rect 16716 3350 16772 3388
rect 17836 3444 17892 3454
rect 17172 3164 17436 3174
rect 17172 3098 17436 3108
rect 13692 2940 13972 2996
rect 13916 800 13972 2940
rect 17836 800 17892 3388
rect 18284 3444 18340 3454
rect 18284 3350 18340 3388
rect 18956 3444 19012 3454
rect 18956 3350 19012 3388
rect 19180 3444 19236 4062
rect 19628 3778 19684 4508
rect 19852 4498 19908 4508
rect 19740 4340 19796 4350
rect 19740 4246 19796 4284
rect 20300 4116 20356 4508
rect 20412 4450 20468 4956
rect 20412 4398 20414 4450
rect 20466 4398 20468 4450
rect 20412 4340 20468 4398
rect 20412 4274 20468 4284
rect 20524 4564 20580 5292
rect 20748 5012 20804 5022
rect 20748 4918 20804 4956
rect 20860 4898 20916 4910
rect 20860 4846 20862 4898
rect 20914 4846 20916 4898
rect 20860 4564 20916 4846
rect 20524 4562 20916 4564
rect 20524 4510 20526 4562
rect 20578 4510 20916 4562
rect 20524 4508 20916 4510
rect 20524 4116 20580 4508
rect 20860 4452 20916 4508
rect 21084 4452 21140 5854
rect 21196 7250 21252 7262
rect 21196 7198 21198 7250
rect 21250 7198 21252 7250
rect 21196 5684 21252 7198
rect 21644 6692 21700 6702
rect 21644 6690 21924 6692
rect 21644 6638 21646 6690
rect 21698 6638 21924 6690
rect 21644 6636 21924 6638
rect 21644 6626 21700 6636
rect 21756 6466 21812 6478
rect 21756 6414 21758 6466
rect 21810 6414 21812 6466
rect 21756 6244 21812 6414
rect 21196 5590 21252 5628
rect 21644 6188 21812 6244
rect 21644 5684 21700 6188
rect 21868 5906 21924 6636
rect 21868 5854 21870 5906
rect 21922 5854 21924 5906
rect 21644 5618 21700 5628
rect 21756 5682 21812 5694
rect 21756 5630 21758 5682
rect 21810 5630 21812 5682
rect 21756 5124 21812 5630
rect 21644 5068 21812 5124
rect 21644 5012 21700 5068
rect 21644 4918 21700 4956
rect 21756 4900 21812 4910
rect 21868 4900 21924 5854
rect 21980 5012 22036 8372
rect 22492 7868 22756 7878
rect 22492 7802 22756 7812
rect 22492 6300 22756 6310
rect 22492 6234 22756 6244
rect 21980 4946 22036 4956
rect 21756 4898 21924 4900
rect 21756 4846 21758 4898
rect 21810 4846 21924 4898
rect 21756 4844 21924 4846
rect 21196 4564 21252 4574
rect 21756 4564 21812 4844
rect 22492 4732 22756 4742
rect 22492 4666 22756 4676
rect 21196 4562 21812 4564
rect 21196 4510 21198 4562
rect 21250 4510 21812 4562
rect 21196 4508 21812 4510
rect 21196 4452 21252 4508
rect 20860 4450 21252 4452
rect 20860 4398 21086 4450
rect 21138 4398 21252 4450
rect 20860 4396 21252 4398
rect 21084 4386 21140 4396
rect 20300 4060 20580 4116
rect 21756 4340 21812 4508
rect 21868 4340 21924 4350
rect 21756 4338 21924 4340
rect 21756 4286 21870 4338
rect 21922 4286 21924 4338
rect 21756 4284 21924 4286
rect 21756 4114 21812 4284
rect 21868 4274 21924 4284
rect 21756 4062 21758 4114
rect 21810 4062 21812 4114
rect 19832 3948 20096 3958
rect 19832 3882 20096 3892
rect 19628 3726 19630 3778
rect 19682 3726 19684 3778
rect 19628 3714 19684 3726
rect 20300 3778 20356 4060
rect 20300 3726 20302 3778
rect 20354 3726 20356 3778
rect 20188 3556 20244 3566
rect 20300 3556 20356 3726
rect 20188 3554 20356 3556
rect 20188 3502 20190 3554
rect 20242 3502 20356 3554
rect 20188 3500 20356 3502
rect 20188 3490 20244 3500
rect 19180 3378 19236 3388
rect 19516 3444 19572 3454
rect 19516 3350 19572 3388
rect 21756 800 21812 4062
rect 22492 3164 22756 3174
rect 22492 3098 22756 3108
rect 2128 0 2240 800
rect 6048 0 6160 800
rect 9968 0 10080 800
rect 13888 0 14000 800
rect 17808 0 17920 800
rect 21728 0 21840 800
<< via2 >>
rect 3872 16490 4136 16492
rect 3872 16438 3874 16490
rect 3874 16438 4134 16490
rect 4134 16438 4136 16490
rect 3872 16436 4136 16438
rect 9192 16490 9456 16492
rect 9192 16438 9194 16490
rect 9194 16438 9454 16490
rect 9454 16438 9456 16490
rect 9192 16436 9456 16438
rect 14512 16490 14776 16492
rect 14512 16438 14514 16490
rect 14514 16438 14774 16490
rect 14774 16438 14776 16490
rect 14512 16436 14776 16438
rect 19832 16490 20096 16492
rect 19832 16438 19834 16490
rect 19834 16438 20094 16490
rect 20094 16438 20096 16490
rect 19832 16436 20096 16438
rect 6532 15706 6796 15708
rect 6532 15654 6534 15706
rect 6534 15654 6794 15706
rect 6794 15654 6796 15706
rect 6532 15652 6796 15654
rect 11852 15706 12116 15708
rect 11852 15654 11854 15706
rect 11854 15654 12114 15706
rect 12114 15654 12116 15706
rect 11852 15652 12116 15654
rect 17172 15706 17436 15708
rect 17172 15654 17174 15706
rect 17174 15654 17434 15706
rect 17434 15654 17436 15706
rect 17172 15652 17436 15654
rect 22492 15706 22756 15708
rect 22492 15654 22494 15706
rect 22494 15654 22754 15706
rect 22754 15654 22756 15706
rect 22492 15652 22756 15654
rect 3612 14924 3668 14980
rect 3500 9154 3556 9156
rect 3500 9102 3502 9154
rect 3502 9102 3554 9154
rect 3554 9102 3556 9154
rect 3500 9100 3556 9102
rect 3872 14922 4136 14924
rect 3872 14870 3874 14922
rect 3874 14870 4134 14922
rect 4134 14870 4136 14922
rect 3872 14868 4136 14870
rect 9192 14922 9456 14924
rect 9192 14870 9194 14922
rect 9194 14870 9454 14922
rect 9454 14870 9456 14922
rect 9192 14868 9456 14870
rect 14512 14922 14776 14924
rect 14512 14870 14514 14922
rect 14514 14870 14774 14922
rect 14774 14870 14776 14922
rect 14512 14868 14776 14870
rect 19832 14922 20096 14924
rect 19832 14870 19834 14922
rect 19834 14870 20094 14922
rect 20094 14870 20096 14922
rect 19832 14868 20096 14870
rect 19628 14700 19684 14756
rect 6532 14138 6796 14140
rect 6532 14086 6534 14138
rect 6534 14086 6794 14138
rect 6794 14086 6796 14138
rect 6532 14084 6796 14086
rect 11852 14138 12116 14140
rect 11852 14086 11854 14138
rect 11854 14086 12114 14138
rect 12114 14086 12116 14138
rect 11852 14084 12116 14086
rect 3872 13354 4136 13356
rect 3872 13302 3874 13354
rect 3874 13302 4134 13354
rect 4134 13302 4136 13354
rect 3872 13300 4136 13302
rect 9192 13354 9456 13356
rect 9192 13302 9194 13354
rect 9194 13302 9454 13354
rect 9454 13302 9456 13354
rect 9192 13300 9456 13302
rect 14512 13354 14776 13356
rect 14512 13302 14514 13354
rect 14514 13302 14774 13354
rect 14774 13302 14776 13354
rect 14512 13300 14776 13302
rect 14924 13186 14980 13188
rect 14924 13134 14926 13186
rect 14926 13134 14978 13186
rect 14978 13134 14980 13186
rect 14924 13132 14980 13134
rect 16268 13522 16324 13524
rect 16268 13470 16270 13522
rect 16270 13470 16322 13522
rect 16322 13470 16324 13522
rect 16268 13468 16324 13470
rect 6532 12570 6796 12572
rect 6532 12518 6534 12570
rect 6534 12518 6794 12570
rect 6794 12518 6796 12570
rect 6532 12516 6796 12518
rect 11852 12570 12116 12572
rect 11852 12518 11854 12570
rect 11854 12518 12114 12570
rect 12114 12518 12116 12570
rect 11852 12516 12116 12518
rect 3872 11786 4136 11788
rect 3872 11734 3874 11786
rect 3874 11734 4134 11786
rect 4134 11734 4136 11786
rect 3872 11732 4136 11734
rect 9192 11786 9456 11788
rect 9192 11734 9194 11786
rect 9194 11734 9454 11786
rect 9454 11734 9456 11786
rect 9192 11732 9456 11734
rect 6188 11282 6244 11284
rect 6188 11230 6190 11282
rect 6190 11230 6242 11282
rect 6242 11230 6244 11282
rect 6188 11228 6244 11230
rect 5516 10722 5572 10724
rect 5516 10670 5518 10722
rect 5518 10670 5570 10722
rect 5570 10670 5572 10722
rect 5516 10668 5572 10670
rect 3872 10218 4136 10220
rect 3872 10166 3874 10218
rect 3874 10166 4134 10218
rect 4134 10166 4136 10218
rect 3872 10164 4136 10166
rect 4284 9826 4340 9828
rect 4284 9774 4286 9826
rect 4286 9774 4338 9826
rect 4338 9774 4340 9826
rect 4284 9772 4340 9774
rect 4844 9826 4900 9828
rect 4844 9774 4846 9826
rect 4846 9774 4898 9826
rect 4898 9774 4900 9826
rect 4844 9772 4900 9774
rect 6972 11282 7028 11284
rect 6972 11230 6974 11282
rect 6974 11230 7026 11282
rect 7026 11230 7028 11282
rect 6972 11228 7028 11230
rect 6532 11002 6796 11004
rect 6532 10950 6534 11002
rect 6534 10950 6794 11002
rect 6794 10950 6796 11002
rect 6532 10948 6796 10950
rect 6076 10722 6132 10724
rect 6076 10670 6078 10722
rect 6078 10670 6130 10722
rect 6130 10670 6132 10722
rect 6076 10668 6132 10670
rect 5404 9772 5460 9828
rect 5852 9714 5908 9716
rect 5852 9662 5854 9714
rect 5854 9662 5906 9714
rect 5906 9662 5908 9714
rect 5852 9660 5908 9662
rect 4060 9154 4116 9156
rect 4060 9102 4062 9154
rect 4062 9102 4114 9154
rect 4114 9102 4116 9154
rect 4060 9100 4116 9102
rect 3872 8650 4136 8652
rect 3872 8598 3874 8650
rect 3874 8598 4134 8650
rect 4134 8598 4136 8650
rect 3872 8596 4136 8598
rect 3612 8428 3668 8484
rect 4172 8428 4228 8484
rect 2156 7474 2212 7476
rect 2156 7422 2158 7474
rect 2158 7422 2210 7474
rect 2210 7422 2212 7474
rect 2156 7420 2212 7422
rect 2716 7474 2772 7476
rect 2716 7422 2718 7474
rect 2718 7422 2770 7474
rect 2770 7422 2772 7474
rect 2716 7420 2772 7422
rect 2156 6578 2212 6580
rect 2156 6526 2158 6578
rect 2158 6526 2210 6578
rect 2210 6526 2212 6578
rect 2156 6524 2212 6526
rect 2828 6748 2884 6804
rect 2828 6578 2884 6580
rect 2828 6526 2830 6578
rect 2830 6526 2882 6578
rect 2882 6526 2884 6578
rect 2828 6524 2884 6526
rect 3612 7196 3668 7252
rect 3388 6524 3444 6580
rect 2716 5068 2772 5124
rect 4284 8034 4340 8036
rect 4284 7982 4286 8034
rect 4286 7982 4338 8034
rect 4338 7982 4340 8034
rect 4284 7980 4340 7982
rect 4732 8428 4788 8484
rect 4172 7250 4228 7252
rect 4172 7198 4174 7250
rect 4174 7198 4226 7250
rect 4226 7198 4228 7250
rect 4172 7196 4228 7198
rect 3872 7082 4136 7084
rect 3872 7030 3874 7082
rect 3874 7030 4134 7082
rect 4134 7030 4136 7082
rect 3872 7028 4136 7030
rect 6524 9714 6580 9716
rect 6524 9662 6526 9714
rect 6526 9662 6578 9714
rect 6578 9662 6580 9714
rect 6524 9660 6580 9662
rect 9192 10218 9456 10220
rect 9192 10166 9194 10218
rect 9194 10166 9454 10218
rect 9454 10166 9456 10218
rect 9192 10164 9456 10166
rect 8988 9996 9044 10052
rect 9996 10108 10052 10164
rect 7196 9714 7252 9716
rect 7196 9662 7198 9714
rect 7198 9662 7250 9714
rect 7250 9662 7252 9714
rect 7196 9660 7252 9662
rect 4956 8482 5012 8484
rect 4956 8430 4958 8482
rect 4958 8430 5010 8482
rect 5010 8430 5012 8482
rect 4956 8428 5012 8430
rect 5404 8428 5460 8484
rect 4844 7980 4900 8036
rect 6532 9434 6796 9436
rect 6532 9382 6534 9434
rect 6534 9382 6794 9434
rect 6794 9382 6796 9434
rect 6532 9380 6796 9382
rect 5964 8482 6020 8484
rect 5964 8430 5966 8482
rect 5966 8430 6018 8482
rect 6018 8430 6020 8482
rect 5964 8428 6020 8430
rect 4844 7474 4900 7476
rect 4844 7422 4846 7474
rect 4846 7422 4898 7474
rect 4898 7422 4900 7474
rect 4844 7420 4900 7422
rect 6524 8428 6580 8484
rect 6532 7866 6796 7868
rect 6532 7814 6534 7866
rect 6534 7814 6794 7866
rect 6794 7814 6796 7866
rect 6532 7812 6796 7814
rect 5404 7474 5460 7476
rect 5404 7422 5406 7474
rect 5406 7422 5458 7474
rect 5458 7422 5460 7474
rect 5404 7420 5460 7422
rect 6076 7474 6132 7476
rect 6076 7422 6078 7474
rect 6078 7422 6130 7474
rect 6130 7422 6132 7474
rect 6076 7420 6132 7422
rect 3724 6748 3780 6804
rect 4620 6748 4676 6804
rect 3388 5068 3444 5124
rect 4060 5906 4116 5908
rect 4060 5854 4062 5906
rect 4062 5854 4114 5906
rect 4114 5854 4116 5906
rect 4060 5852 4116 5854
rect 2380 4450 2436 4452
rect 2380 4398 2382 4450
rect 2382 4398 2434 4450
rect 2434 4398 2436 4450
rect 2380 4396 2436 4398
rect 3052 4396 3108 4452
rect 2492 4338 2548 4340
rect 2492 4286 2494 4338
rect 2494 4286 2546 4338
rect 2546 4286 2548 4338
rect 2492 4284 2548 4286
rect 2828 4284 2884 4340
rect 2156 3500 2212 3556
rect 3164 4338 3220 4340
rect 3164 4286 3166 4338
rect 3166 4286 3218 4338
rect 3218 4286 3220 4338
rect 3164 4284 3220 4286
rect 5516 6748 5572 6804
rect 5740 6748 5796 6804
rect 4732 5906 4788 5908
rect 4732 5854 4734 5906
rect 4734 5854 4786 5906
rect 4786 5854 4788 5906
rect 4732 5852 4788 5854
rect 7196 8428 7252 8484
rect 8652 9602 8708 9604
rect 8652 9550 8654 9602
rect 8654 9550 8706 9602
rect 8706 9550 8708 9602
rect 8652 9548 8708 9550
rect 7980 8428 8036 8484
rect 7308 8034 7364 8036
rect 7308 7982 7310 8034
rect 7310 7982 7362 8034
rect 7362 7982 7364 8034
rect 7308 7980 7364 7982
rect 6748 7474 6804 7476
rect 6748 7422 6750 7474
rect 6750 7422 6802 7474
rect 6802 7422 6804 7474
rect 6748 7420 6804 7422
rect 6412 6748 6468 6804
rect 7308 7420 7364 7476
rect 7980 8034 8036 8036
rect 7980 7982 7982 8034
rect 7982 7982 8034 8034
rect 8034 7982 8036 8034
rect 7980 7980 8036 7982
rect 9324 9602 9380 9604
rect 9324 9550 9326 9602
rect 9326 9550 9378 9602
rect 9378 9550 9380 9602
rect 9324 9548 9380 9550
rect 8540 8428 8596 8484
rect 9192 8650 9456 8652
rect 9192 8598 9194 8650
rect 9194 8598 9454 8650
rect 9454 8598 9456 8650
rect 9192 8596 9456 8598
rect 9324 8482 9380 8484
rect 9324 8430 9326 8482
rect 9326 8430 9378 8482
rect 9378 8430 9380 8482
rect 9324 8428 9380 8430
rect 8316 7980 8372 8036
rect 8988 8316 9044 8372
rect 7532 6860 7588 6916
rect 6532 6298 6796 6300
rect 6532 6246 6534 6298
rect 6534 6246 6794 6298
rect 6794 6246 6796 6298
rect 6532 6244 6796 6246
rect 3872 5514 4136 5516
rect 3872 5462 3874 5514
rect 3874 5462 4134 5514
rect 4134 5462 4136 5514
rect 3872 5460 4136 5462
rect 4172 5122 4228 5124
rect 4172 5070 4174 5122
rect 4174 5070 4226 5122
rect 4226 5070 4228 5122
rect 4172 5068 4228 5070
rect 3612 5010 3668 5012
rect 3612 4958 3614 5010
rect 3614 4958 3666 5010
rect 3666 4958 3668 5010
rect 3612 4956 3668 4958
rect 3836 4562 3892 4564
rect 3836 4510 3838 4562
rect 3838 4510 3890 4562
rect 3890 4510 3892 4562
rect 3836 4508 3892 4510
rect 3500 4284 3556 4340
rect 3724 4338 3780 4340
rect 3724 4286 3726 4338
rect 3726 4286 3778 4338
rect 3778 4286 3780 4338
rect 3724 4284 3780 4286
rect 2828 3554 2884 3556
rect 2828 3502 2830 3554
rect 2830 3502 2882 3554
rect 2882 3502 2884 3554
rect 2828 3500 2884 3502
rect 4732 4844 4788 4900
rect 4508 4562 4564 4564
rect 4508 4510 4510 4562
rect 4510 4510 4562 4562
rect 4562 4510 4564 4562
rect 4508 4508 4564 4510
rect 4956 5068 5012 5124
rect 4956 4898 5012 4900
rect 4956 4846 4958 4898
rect 4958 4846 5010 4898
rect 5010 4846 5012 4898
rect 4956 4844 5012 4846
rect 4844 4508 4900 4564
rect 4396 4338 4452 4340
rect 4396 4286 4398 4338
rect 4398 4286 4450 4338
rect 4450 4286 4452 4338
rect 4396 4284 4452 4286
rect 4284 4060 4340 4116
rect 3872 3946 4136 3948
rect 3872 3894 3874 3946
rect 3874 3894 4134 3946
rect 4134 3894 4136 3946
rect 3872 3892 4136 3894
rect 3052 3500 3108 3556
rect 3500 3554 3556 3556
rect 3500 3502 3502 3554
rect 3502 3502 3554 3554
rect 3554 3502 3556 3554
rect 3500 3500 3556 3502
rect 4172 3554 4228 3556
rect 4172 3502 4174 3554
rect 4174 3502 4226 3554
rect 4226 3502 4228 3554
rect 4172 3500 4228 3502
rect 5404 4844 5460 4900
rect 5852 4844 5908 4900
rect 5740 4508 5796 4564
rect 4396 3388 4452 3444
rect 4844 3442 4900 3444
rect 4844 3390 4846 3442
rect 4846 3390 4898 3442
rect 4898 3390 4900 3442
rect 4844 3388 4900 3390
rect 5852 4114 5908 4116
rect 5852 4062 5854 4114
rect 5854 4062 5906 4114
rect 5906 4062 5908 4114
rect 5852 4060 5908 4062
rect 7084 5964 7140 6020
rect 7420 6018 7476 6020
rect 7420 5966 7422 6018
rect 7422 5966 7474 6018
rect 7474 5966 7476 6018
rect 7420 5964 7476 5966
rect 7756 5964 7812 6020
rect 9884 8316 9940 8372
rect 9212 8258 9268 8260
rect 9212 8206 9214 8258
rect 9214 8206 9266 8258
rect 9266 8206 9268 8258
rect 9212 8204 9268 8206
rect 11852 11002 12116 11004
rect 11852 10950 11854 11002
rect 11854 10950 12114 11002
rect 12114 10950 12116 11002
rect 11852 10948 12116 10950
rect 14812 12178 14868 12180
rect 14812 12126 14814 12178
rect 14814 12126 14866 12178
rect 14866 12126 14868 12178
rect 14812 12124 14868 12126
rect 14252 11954 14308 11956
rect 14252 11902 14254 11954
rect 14254 11902 14306 11954
rect 14306 11902 14308 11954
rect 14252 11900 14308 11902
rect 14924 11954 14980 11956
rect 14924 11902 14926 11954
rect 14926 11902 14978 11954
rect 14978 11902 14980 11954
rect 14924 11900 14980 11902
rect 14512 11786 14776 11788
rect 14512 11734 14514 11786
rect 14514 11734 14774 11786
rect 14774 11734 14776 11786
rect 14512 11732 14776 11734
rect 14924 11394 14980 11396
rect 14924 11342 14926 11394
rect 14926 11342 14978 11394
rect 14978 11342 14980 11394
rect 14924 11340 14980 11342
rect 11340 9996 11396 10052
rect 14512 10218 14776 10220
rect 14512 10166 14514 10218
rect 14514 10166 14774 10218
rect 14774 10166 14776 10218
rect 14512 10164 14776 10166
rect 12012 9996 12068 10052
rect 15484 12178 15540 12180
rect 15484 12126 15486 12178
rect 15486 12126 15538 12178
rect 15538 12126 15540 12178
rect 15484 12124 15540 12126
rect 15596 11394 15652 11396
rect 15596 11342 15598 11394
rect 15598 11342 15650 11394
rect 15650 11342 15652 11394
rect 15596 11340 15652 11342
rect 16156 12178 16212 12180
rect 16156 12126 16158 12178
rect 16158 12126 16210 12178
rect 16210 12126 16212 12178
rect 16156 12124 16212 12126
rect 16940 13522 16996 13524
rect 16940 13470 16942 13522
rect 16942 13470 16994 13522
rect 16994 13470 16996 13522
rect 16940 13468 16996 13470
rect 17172 14138 17436 14140
rect 17172 14086 17174 14138
rect 17174 14086 17434 14138
rect 17434 14086 17436 14138
rect 17172 14084 17436 14086
rect 17052 13132 17108 13188
rect 17388 13468 17444 13524
rect 16828 12178 16884 12180
rect 16828 12126 16830 12178
rect 16830 12126 16882 12178
rect 16882 12126 16884 12178
rect 16828 12124 16884 12126
rect 17612 13468 17668 13524
rect 17724 13132 17780 13188
rect 18396 13468 18452 13524
rect 18508 13244 18564 13300
rect 18956 13468 19012 13524
rect 18284 13186 18340 13188
rect 18284 13134 18286 13186
rect 18286 13134 18338 13186
rect 18338 13134 18340 13186
rect 18284 13132 18340 13134
rect 18844 13132 18900 13188
rect 17172 12570 17436 12572
rect 17172 12518 17174 12570
rect 17174 12518 17434 12570
rect 17434 12518 17436 12570
rect 17172 12516 17436 12518
rect 16268 11394 16324 11396
rect 16268 11342 16270 11394
rect 16270 11342 16322 11394
rect 16322 11342 16324 11394
rect 16268 11340 16324 11342
rect 17612 11788 17668 11844
rect 22492 14138 22756 14140
rect 22492 14086 22494 14138
rect 22494 14086 22754 14138
rect 22754 14086 22756 14138
rect 22492 14084 22756 14086
rect 19628 13468 19684 13524
rect 18396 12290 18452 12292
rect 18396 12238 18398 12290
rect 18398 12238 18450 12290
rect 18450 12238 18452 12290
rect 18396 12236 18452 12238
rect 16940 11394 16996 11396
rect 16940 11342 16942 11394
rect 16942 11342 16994 11394
rect 16994 11342 16996 11394
rect 16940 11340 16996 11342
rect 9996 8540 10052 8596
rect 11852 9434 12116 9436
rect 11852 9382 11854 9434
rect 11854 9382 12114 9434
rect 12114 9382 12116 9434
rect 11852 9380 12116 9382
rect 10556 8540 10612 8596
rect 10332 8316 10388 8372
rect 9996 8204 10052 8260
rect 12460 8204 12516 8260
rect 12796 8428 12852 8484
rect 14364 9042 14420 9044
rect 14364 8990 14366 9042
rect 14366 8990 14418 9042
rect 14418 8990 14420 9042
rect 14364 8988 14420 8990
rect 13692 8428 13748 8484
rect 12908 8258 12964 8260
rect 12908 8206 12910 8258
rect 12910 8206 12962 8258
rect 12962 8206 12964 8258
rect 12908 8204 12964 8206
rect 13356 8204 13412 8260
rect 8428 6578 8484 6580
rect 8428 6526 8430 6578
rect 8430 6526 8482 6578
rect 8482 6526 8484 6578
rect 8428 6524 8484 6526
rect 8540 6690 8596 6692
rect 8540 6638 8542 6690
rect 8542 6638 8594 6690
rect 8594 6638 8596 6690
rect 8540 6636 8596 6638
rect 8092 6018 8148 6020
rect 8092 5966 8094 6018
rect 8094 5966 8146 6018
rect 8146 5966 8148 6018
rect 8092 5964 8148 5966
rect 6076 4844 6132 4900
rect 6300 4508 6356 4564
rect 6532 4730 6796 4732
rect 6532 4678 6534 4730
rect 6534 4678 6794 4730
rect 6794 4678 6796 4730
rect 6532 4676 6796 4678
rect 6076 4060 6132 4116
rect 5180 3388 5236 3444
rect 5740 3442 5796 3444
rect 5740 3390 5742 3442
rect 5742 3390 5794 3442
rect 5794 3390 5796 3442
rect 5740 3388 5796 3390
rect 7308 5068 7364 5124
rect 6524 4114 6580 4116
rect 6524 4062 6526 4114
rect 6526 4062 6578 4114
rect 6578 4062 6580 4114
rect 6524 4060 6580 4062
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 7084 4060 7140 4116
rect 7084 3500 7140 3556
rect 9192 7082 9456 7084
rect 9192 7030 9194 7082
rect 9194 7030 9454 7082
rect 9454 7030 9456 7082
rect 9192 7028 9456 7030
rect 8764 6636 8820 6692
rect 8876 6860 8932 6916
rect 9212 6690 9268 6692
rect 9212 6638 9214 6690
rect 9214 6638 9266 6690
rect 9266 6638 9268 6690
rect 9212 6636 9268 6638
rect 9884 6636 9940 6692
rect 9100 6578 9156 6580
rect 9100 6526 9102 6578
rect 9102 6526 9154 6578
rect 9154 6526 9156 6578
rect 9100 6524 9156 6526
rect 9996 6860 10052 6916
rect 9884 6466 9940 6468
rect 9884 6414 9886 6466
rect 9886 6414 9938 6466
rect 9938 6414 9940 6466
rect 9884 6412 9940 6414
rect 9100 5852 9156 5908
rect 9772 5906 9828 5908
rect 9772 5854 9774 5906
rect 9774 5854 9826 5906
rect 9826 5854 9828 5906
rect 9772 5852 9828 5854
rect 9192 5514 9456 5516
rect 9192 5462 9194 5514
rect 9194 5462 9454 5514
rect 9454 5462 9456 5514
rect 9192 5460 9456 5462
rect 7756 5122 7812 5124
rect 7756 5070 7758 5122
rect 7758 5070 7810 5122
rect 7810 5070 7812 5122
rect 7756 5068 7812 5070
rect 11852 7866 12116 7868
rect 11852 7814 11854 7866
rect 11854 7814 12114 7866
rect 12114 7814 12116 7866
rect 11852 7812 12116 7814
rect 10556 6914 10612 6916
rect 10556 6862 10558 6914
rect 10558 6862 10610 6914
rect 10610 6862 10612 6914
rect 10556 6860 10612 6862
rect 10444 6690 10500 6692
rect 10444 6638 10446 6690
rect 10446 6638 10498 6690
rect 10498 6638 10500 6690
rect 10444 6636 10500 6638
rect 11228 6914 11284 6916
rect 11228 6862 11230 6914
rect 11230 6862 11282 6914
rect 11282 6862 11284 6914
rect 11228 6860 11284 6862
rect 10556 6412 10612 6468
rect 11116 6690 11172 6692
rect 11116 6638 11118 6690
rect 11118 6638 11170 6690
rect 11170 6638 11172 6690
rect 11116 6636 11172 6638
rect 10444 5906 10500 5908
rect 10444 5854 10446 5906
rect 10446 5854 10498 5906
rect 10498 5854 10500 5906
rect 10444 5852 10500 5854
rect 8540 5068 8596 5124
rect 9100 5122 9156 5124
rect 9100 5070 9102 5122
rect 9102 5070 9154 5122
rect 9154 5070 9156 5122
rect 9100 5068 9156 5070
rect 9660 5068 9716 5124
rect 7756 4338 7812 4340
rect 7756 4286 7758 4338
rect 7758 4286 7810 4338
rect 7810 4286 7812 4338
rect 7756 4284 7812 4286
rect 7756 3554 7812 3556
rect 7756 3502 7758 3554
rect 7758 3502 7810 3554
rect 7810 3502 7812 3554
rect 7756 3500 7812 3502
rect 8428 3554 8484 3556
rect 8428 3502 8430 3554
rect 8430 3502 8482 3554
rect 8482 3502 8484 3554
rect 8428 3500 8484 3502
rect 9192 3946 9456 3948
rect 9192 3894 9194 3946
rect 9194 3894 9454 3946
rect 9454 3894 9456 3946
rect 9192 3892 9456 3894
rect 9660 3554 9716 3556
rect 9660 3502 9662 3554
rect 9662 3502 9714 3554
rect 9714 3502 9716 3554
rect 9660 3500 9716 3502
rect 9884 3500 9940 3556
rect 6636 3388 6692 3444
rect 6532 3162 6796 3164
rect 6532 3110 6534 3162
rect 6534 3110 6794 3162
rect 6794 3110 6796 3162
rect 6532 3108 6796 3110
rect 11900 6636 11956 6692
rect 12012 6860 12068 6916
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 12460 6690 12516 6692
rect 12460 6638 12462 6690
rect 12462 6638 12514 6690
rect 12514 6638 12516 6690
rect 12460 6636 12516 6638
rect 11852 6298 12116 6300
rect 11852 6246 11854 6298
rect 11854 6246 12114 6298
rect 12114 6246 12116 6298
rect 11852 6244 12116 6246
rect 13916 8428 13972 8484
rect 15036 9042 15092 9044
rect 15036 8990 15038 9042
rect 15038 8990 15090 9042
rect 15090 8990 15092 9042
rect 15036 8988 15092 8990
rect 17500 11394 17556 11396
rect 17500 11342 17502 11394
rect 17502 11342 17554 11394
rect 17554 11342 17556 11394
rect 17500 11340 17556 11342
rect 17172 11002 17436 11004
rect 17172 10950 17174 11002
rect 17174 10950 17434 11002
rect 17434 10950 17436 11002
rect 17172 10948 17436 10950
rect 19180 13132 19236 13188
rect 19832 13354 20096 13356
rect 19832 13302 19834 13354
rect 19834 13302 20094 13354
rect 20094 13302 20096 13354
rect 19832 13300 20096 13302
rect 18956 12236 19012 12292
rect 18508 11676 18564 11732
rect 15260 8988 15316 9044
rect 14512 8650 14776 8652
rect 14512 8598 14514 8650
rect 14514 8598 14774 8650
rect 14774 8598 14776 8650
rect 14512 8596 14776 8598
rect 14364 8428 14420 8484
rect 14476 8258 14532 8260
rect 14476 8206 14478 8258
rect 14478 8206 14530 8258
rect 14530 8206 14532 8258
rect 14476 8204 14532 8206
rect 15148 8482 15204 8484
rect 15148 8430 15150 8482
rect 15150 8430 15202 8482
rect 15202 8430 15204 8482
rect 15148 8428 15204 8430
rect 15036 8258 15092 8260
rect 15036 8206 15038 8258
rect 15038 8206 15090 8258
rect 15090 8206 15092 8258
rect 15036 8204 15092 8206
rect 14028 6860 14084 6916
rect 14512 7082 14776 7084
rect 14512 7030 14514 7082
rect 14514 7030 14774 7082
rect 14774 7030 14776 7082
rect 14512 7028 14776 7030
rect 14252 6914 14308 6916
rect 14252 6862 14254 6914
rect 14254 6862 14306 6914
rect 14306 6862 14308 6914
rect 14252 6860 14308 6862
rect 14588 6860 14644 6916
rect 11564 5122 11620 5124
rect 11564 5070 11566 5122
rect 11566 5070 11618 5122
rect 11618 5070 11620 5122
rect 11564 5068 11620 5070
rect 12124 5068 12180 5124
rect 12348 4844 12404 4900
rect 11852 4730 12116 4732
rect 11852 4678 11854 4730
rect 11854 4678 12114 4730
rect 12114 4678 12116 4730
rect 11852 4676 12116 4678
rect 12908 4898 12964 4900
rect 12908 4846 12910 4898
rect 12910 4846 12962 4898
rect 12962 4846 12964 4898
rect 12908 4844 12964 4846
rect 16828 10386 16884 10388
rect 16828 10334 16830 10386
rect 16830 10334 16882 10386
rect 16882 10334 16884 10386
rect 16828 10332 16884 10334
rect 18284 11170 18340 11172
rect 18284 11118 18286 11170
rect 18286 11118 18338 11170
rect 18338 11118 18340 11170
rect 18284 11116 18340 11118
rect 17836 10386 17892 10388
rect 17836 10334 17838 10386
rect 17838 10334 17890 10386
rect 17890 10334 17892 10386
rect 17836 10332 17892 10334
rect 18284 10332 18340 10388
rect 18956 11340 19012 11396
rect 18508 11116 18564 11172
rect 18956 11170 19012 11172
rect 18956 11118 18958 11170
rect 18958 11118 19010 11170
rect 19010 11118 19012 11170
rect 18956 11116 19012 11118
rect 22492 12570 22756 12572
rect 22492 12518 22494 12570
rect 22494 12518 22754 12570
rect 22754 12518 22756 12570
rect 22492 12516 22756 12518
rect 19740 12290 19796 12292
rect 19740 12238 19742 12290
rect 19742 12238 19794 12290
rect 19794 12238 19796 12290
rect 19740 12236 19796 12238
rect 20412 12290 20468 12292
rect 20412 12238 20414 12290
rect 20414 12238 20466 12290
rect 20466 12238 20468 12290
rect 20412 12236 20468 12238
rect 21084 12236 21140 12292
rect 19832 11786 20096 11788
rect 19832 11734 19834 11786
rect 19834 11734 20094 11786
rect 20094 11734 20096 11786
rect 19832 11732 20096 11734
rect 19516 11394 19572 11396
rect 19516 11342 19518 11394
rect 19518 11342 19570 11394
rect 19570 11342 19572 11394
rect 19516 11340 19572 11342
rect 18508 10386 18564 10388
rect 18508 10334 18510 10386
rect 18510 10334 18562 10386
rect 18562 10334 18564 10386
rect 18508 10332 18564 10334
rect 19852 11340 19908 11396
rect 19852 10668 19908 10724
rect 20188 10668 20244 10724
rect 19832 10218 20096 10220
rect 19832 10166 19834 10218
rect 19834 10166 20094 10218
rect 20094 10166 20096 10218
rect 19832 10164 20096 10166
rect 19852 9996 19908 10052
rect 15596 8204 15652 8260
rect 15708 8428 15764 8484
rect 10332 3554 10388 3556
rect 10332 3502 10334 3554
rect 10334 3502 10386 3554
rect 10386 3502 10388 3554
rect 10332 3500 10388 3502
rect 12460 4114 12516 4116
rect 12460 4062 12462 4114
rect 12462 4062 12514 4114
rect 12514 4062 12516 4114
rect 12460 4060 12516 4062
rect 13132 4114 13188 4116
rect 13132 4062 13134 4114
rect 13134 4062 13186 4114
rect 13186 4062 13188 4114
rect 13132 4060 13188 4062
rect 11116 3554 11172 3556
rect 11116 3502 11118 3554
rect 11118 3502 11170 3554
rect 11170 3502 11172 3554
rect 11116 3500 11172 3502
rect 11676 3554 11732 3556
rect 11676 3502 11678 3554
rect 11678 3502 11730 3554
rect 11730 3502 11732 3554
rect 11676 3500 11732 3502
rect 11004 3442 11060 3444
rect 11004 3390 11006 3442
rect 11006 3390 11058 3442
rect 11058 3390 11060 3442
rect 11004 3388 11060 3390
rect 11788 3442 11844 3444
rect 11788 3390 11790 3442
rect 11790 3390 11842 3442
rect 11842 3390 11844 3442
rect 11788 3388 11844 3390
rect 11852 3162 12116 3164
rect 11852 3110 11854 3162
rect 11854 3110 12114 3162
rect 12114 3110 12116 3162
rect 11852 3108 12116 3110
rect 13804 4114 13860 4116
rect 13804 4062 13806 4114
rect 13806 4062 13858 4114
rect 13858 4062 13860 4114
rect 13804 4060 13860 4062
rect 14512 5514 14776 5516
rect 14512 5462 14514 5514
rect 14514 5462 14774 5514
rect 14774 5462 14776 5514
rect 14512 5460 14776 5462
rect 15260 6860 15316 6916
rect 15820 8258 15876 8260
rect 15820 8206 15822 8258
rect 15822 8206 15874 8258
rect 15874 8206 15876 8258
rect 15820 8204 15876 8206
rect 16492 9602 16548 9604
rect 16492 9550 16494 9602
rect 16494 9550 16546 9602
rect 16546 9550 16548 9602
rect 16492 9548 16548 9550
rect 16268 8204 16324 8260
rect 16380 8428 16436 8484
rect 16492 8258 16548 8260
rect 16492 8206 16494 8258
rect 16494 8206 16546 8258
rect 16546 8206 16548 8258
rect 16492 8204 16548 8206
rect 17164 9602 17220 9604
rect 17164 9550 17166 9602
rect 17166 9550 17218 9602
rect 17218 9550 17220 9602
rect 17164 9548 17220 9550
rect 17172 9434 17436 9436
rect 17172 9382 17174 9434
rect 17174 9382 17434 9434
rect 17434 9382 17436 9434
rect 17172 9380 17436 9382
rect 17164 8482 17220 8484
rect 17164 8430 17166 8482
rect 17166 8430 17218 8482
rect 17218 8430 17220 8482
rect 17164 8428 17220 8430
rect 17052 8258 17108 8260
rect 17052 8206 17054 8258
rect 17054 8206 17106 8258
rect 17106 8206 17108 8258
rect 17052 8204 17108 8206
rect 17836 8482 17892 8484
rect 17836 8430 17838 8482
rect 17838 8430 17890 8482
rect 17890 8430 17892 8482
rect 17836 8428 17892 8430
rect 18508 8482 18564 8484
rect 18508 8430 18510 8482
rect 18510 8430 18562 8482
rect 18562 8430 18564 8482
rect 18508 8428 18564 8430
rect 18956 8764 19012 8820
rect 18956 8428 19012 8484
rect 19180 9602 19236 9604
rect 19180 9550 19182 9602
rect 19182 9550 19234 9602
rect 19234 9550 19236 9602
rect 19180 9548 19236 9550
rect 19852 9602 19908 9604
rect 19852 9550 19854 9602
rect 19854 9550 19906 9602
rect 19906 9550 19908 9602
rect 19852 9548 19908 9550
rect 21084 10722 21140 10724
rect 21084 10670 21086 10722
rect 21086 10670 21138 10722
rect 21138 10670 21140 10722
rect 21084 10668 21140 10670
rect 21756 11116 21812 11172
rect 22492 11002 22756 11004
rect 22492 10950 22494 11002
rect 22494 10950 22754 11002
rect 22754 10950 22756 11002
rect 22492 10948 22756 10950
rect 21868 10722 21924 10724
rect 21868 10670 21870 10722
rect 21870 10670 21922 10722
rect 21922 10670 21924 10722
rect 21868 10668 21924 10670
rect 20524 10050 20580 10052
rect 20524 9998 20526 10050
rect 20526 9998 20578 10050
rect 20578 9998 20580 10050
rect 20524 9996 20580 9998
rect 19180 8818 19236 8820
rect 19180 8766 19182 8818
rect 19182 8766 19234 8818
rect 19234 8766 19236 8818
rect 19180 8764 19236 8766
rect 17612 8204 17668 8260
rect 18396 8316 18452 8372
rect 17172 7866 17436 7868
rect 17172 7814 17174 7866
rect 17174 7814 17434 7866
rect 17434 7814 17436 7866
rect 17172 7812 17436 7814
rect 17836 7698 17892 7700
rect 17836 7646 17838 7698
rect 17838 7646 17890 7698
rect 17890 7646 17892 7698
rect 17836 7644 17892 7646
rect 16604 7474 16660 7476
rect 16604 7422 16606 7474
rect 16606 7422 16658 7474
rect 16658 7422 16660 7474
rect 16604 7420 16660 7422
rect 18396 7644 18452 7700
rect 17612 7420 17668 7476
rect 17724 7308 17780 7364
rect 16940 6578 16996 6580
rect 16940 6526 16942 6578
rect 16942 6526 16994 6578
rect 16994 6526 16996 6578
rect 16940 6524 16996 6526
rect 14700 5010 14756 5012
rect 14700 4958 14702 5010
rect 14702 4958 14754 5010
rect 14754 4958 14756 5010
rect 14700 4956 14756 4958
rect 14476 4338 14532 4340
rect 14476 4286 14478 4338
rect 14478 4286 14530 4338
rect 14530 4286 14532 4338
rect 14476 4284 14532 4286
rect 19180 8316 19236 8372
rect 19068 8258 19124 8260
rect 19068 8206 19070 8258
rect 19070 8206 19122 8258
rect 19122 8206 19124 8258
rect 19068 8204 19124 8206
rect 19832 8650 20096 8652
rect 19832 8598 19834 8650
rect 19834 8598 20094 8650
rect 20094 8598 20096 8650
rect 19832 8596 20096 8598
rect 22492 9434 22756 9436
rect 22492 9382 22494 9434
rect 22494 9382 22754 9434
rect 22754 9382 22756 9434
rect 22492 9380 22756 9382
rect 19628 8204 19684 8260
rect 18396 7308 18452 7364
rect 18956 6690 19012 6692
rect 18956 6638 18958 6690
rect 18958 6638 19010 6690
rect 19010 6638 19012 6690
rect 18956 6636 19012 6638
rect 17500 6578 17556 6580
rect 17500 6526 17502 6578
rect 17502 6526 17554 6578
rect 17554 6526 17556 6578
rect 17500 6524 17556 6526
rect 17172 6298 17436 6300
rect 17172 6246 17174 6298
rect 17174 6246 17434 6298
rect 17434 6246 17436 6298
rect 17172 6244 17436 6246
rect 16156 5068 16212 5124
rect 16044 5010 16100 5012
rect 16044 4958 16046 5010
rect 16046 4958 16098 5010
rect 16098 4958 16100 5010
rect 16044 4956 16100 4958
rect 16828 5122 16884 5124
rect 16828 5070 16830 5122
rect 16830 5070 16882 5122
rect 16882 5070 16884 5122
rect 16828 5068 16884 5070
rect 17388 5122 17444 5124
rect 17388 5070 17390 5122
rect 17390 5070 17442 5122
rect 17442 5070 17444 5122
rect 17388 5068 17444 5070
rect 17612 5068 17668 5124
rect 16716 5010 16772 5012
rect 16716 4958 16718 5010
rect 16718 4958 16770 5010
rect 16770 4958 16772 5010
rect 16716 4956 16772 4958
rect 17172 4730 17436 4732
rect 17172 4678 17174 4730
rect 17174 4678 17434 4730
rect 17434 4678 17436 4730
rect 17172 4676 17436 4678
rect 16492 4450 16548 4452
rect 16492 4398 16494 4450
rect 16494 4398 16546 4450
rect 16546 4398 16548 4450
rect 16492 4396 16548 4398
rect 17836 5852 17892 5908
rect 19180 6636 19236 6692
rect 19832 7082 20096 7084
rect 19832 7030 19834 7082
rect 19834 7030 20094 7082
rect 20094 7030 20096 7082
rect 19832 7028 20096 7030
rect 19628 6636 19684 6692
rect 18396 5906 18452 5908
rect 18396 5854 18398 5906
rect 18398 5854 18450 5906
rect 18450 5854 18452 5906
rect 18396 5852 18452 5854
rect 18172 5740 18228 5796
rect 18508 5794 18564 5796
rect 18508 5742 18510 5794
rect 18510 5742 18562 5794
rect 18562 5742 18564 5794
rect 18508 5740 18564 5742
rect 18732 5740 18788 5796
rect 17724 4956 17780 5012
rect 17724 4450 17780 4452
rect 17724 4398 17726 4450
rect 17726 4398 17778 4450
rect 17778 4398 17780 4450
rect 17724 4396 17780 4398
rect 14700 4284 14756 4340
rect 15036 4338 15092 4340
rect 15036 4286 15038 4338
rect 15038 4286 15090 4338
rect 15090 4286 15092 4338
rect 15036 4284 15092 4286
rect 15708 4338 15764 4340
rect 15708 4286 15710 4338
rect 15710 4286 15762 4338
rect 15762 4286 15764 4338
rect 15708 4284 15764 4286
rect 14512 3946 14776 3948
rect 14512 3894 14514 3946
rect 14514 3894 14774 3946
rect 14774 3894 14776 3946
rect 14512 3892 14776 3894
rect 14028 3442 14084 3444
rect 14028 3390 14030 3442
rect 14030 3390 14082 3442
rect 14082 3390 14084 3442
rect 14028 3388 14084 3390
rect 14700 3442 14756 3444
rect 14700 3390 14702 3442
rect 14702 3390 14754 3442
rect 14754 3390 14756 3442
rect 14700 3388 14756 3390
rect 15372 3442 15428 3444
rect 15372 3390 15374 3442
rect 15374 3390 15426 3442
rect 15426 3390 15428 3442
rect 15372 3388 15428 3390
rect 15708 3388 15764 3444
rect 18172 4396 18228 4452
rect 18508 5068 18564 5124
rect 19180 5794 19236 5796
rect 19180 5742 19182 5794
rect 19182 5742 19234 5794
rect 19234 5742 19236 5794
rect 19180 5740 19236 5742
rect 18844 5122 18900 5124
rect 18844 5070 18846 5122
rect 18846 5070 18898 5122
rect 18898 5070 18900 5122
rect 18844 5068 18900 5070
rect 19068 5068 19124 5124
rect 19852 5682 19908 5684
rect 19852 5630 19854 5682
rect 19854 5630 19906 5682
rect 19906 5630 19908 5682
rect 19852 5628 19908 5630
rect 19832 5514 20096 5516
rect 19832 5462 19834 5514
rect 19834 5462 20094 5514
rect 20094 5462 20096 5514
rect 19832 5460 20096 5462
rect 19516 5234 19572 5236
rect 19516 5182 19518 5234
rect 19518 5182 19570 5234
rect 19570 5182 19572 5234
rect 19516 5180 19572 5182
rect 20300 5628 20356 5684
rect 19404 5122 19460 5124
rect 19404 5070 19406 5122
rect 19406 5070 19458 5122
rect 19458 5070 19460 5122
rect 19404 5068 19460 5070
rect 19852 5068 19908 5124
rect 18396 4450 18452 4452
rect 18396 4398 18398 4450
rect 18398 4398 18450 4450
rect 18450 4398 18452 4450
rect 18396 4396 18452 4398
rect 20076 5122 20132 5124
rect 20076 5070 20078 5122
rect 20078 5070 20130 5122
rect 20130 5070 20132 5122
rect 20076 5068 20132 5070
rect 20524 5682 20580 5684
rect 20524 5630 20526 5682
rect 20526 5630 20578 5682
rect 20578 5630 20580 5682
rect 20524 5628 20580 5630
rect 20188 4956 20244 5012
rect 20412 4956 20468 5012
rect 19180 4284 19236 4340
rect 16044 3442 16100 3444
rect 16044 3390 16046 3442
rect 16046 3390 16098 3442
rect 16098 3390 16100 3442
rect 16044 3388 16100 3390
rect 16716 3442 16772 3444
rect 16716 3390 16718 3442
rect 16718 3390 16770 3442
rect 16770 3390 16772 3442
rect 16716 3388 16772 3390
rect 17836 3388 17892 3444
rect 17172 3162 17436 3164
rect 17172 3110 17174 3162
rect 17174 3110 17434 3162
rect 17434 3110 17436 3162
rect 17172 3108 17436 3110
rect 18284 3442 18340 3444
rect 18284 3390 18286 3442
rect 18286 3390 18338 3442
rect 18338 3390 18340 3442
rect 18284 3388 18340 3390
rect 18956 3442 19012 3444
rect 18956 3390 18958 3442
rect 18958 3390 19010 3442
rect 19010 3390 19012 3442
rect 18956 3388 19012 3390
rect 19740 4338 19796 4340
rect 19740 4286 19742 4338
rect 19742 4286 19794 4338
rect 19794 4286 19796 4338
rect 19740 4284 19796 4286
rect 20412 4284 20468 4340
rect 20748 5010 20804 5012
rect 20748 4958 20750 5010
rect 20750 4958 20802 5010
rect 20802 4958 20804 5010
rect 20748 4956 20804 4958
rect 21196 5682 21252 5684
rect 21196 5630 21198 5682
rect 21198 5630 21250 5682
rect 21250 5630 21252 5682
rect 21196 5628 21252 5630
rect 21644 5628 21700 5684
rect 21644 5010 21700 5012
rect 21644 4958 21646 5010
rect 21646 4958 21698 5010
rect 21698 4958 21700 5010
rect 21644 4956 21700 4958
rect 22492 7866 22756 7868
rect 22492 7814 22494 7866
rect 22494 7814 22754 7866
rect 22754 7814 22756 7866
rect 22492 7812 22756 7814
rect 22492 6298 22756 6300
rect 22492 6246 22494 6298
rect 22494 6246 22754 6298
rect 22754 6246 22756 6298
rect 22492 6244 22756 6246
rect 21980 4956 22036 5012
rect 22492 4730 22756 4732
rect 22492 4678 22494 4730
rect 22494 4678 22754 4730
rect 22754 4678 22756 4730
rect 22492 4676 22756 4678
rect 19832 3946 20096 3948
rect 19832 3894 19834 3946
rect 19834 3894 20094 3946
rect 20094 3894 20096 3946
rect 19832 3892 20096 3894
rect 19180 3388 19236 3444
rect 19516 3442 19572 3444
rect 19516 3390 19518 3442
rect 19518 3390 19570 3442
rect 19570 3390 19572 3442
rect 19516 3388 19572 3390
rect 22492 3162 22756 3164
rect 22492 3110 22494 3162
rect 22494 3110 22754 3162
rect 22754 3110 22756 3162
rect 22492 3108 22756 3110
<< metal3 >>
rect 3862 16436 3872 16492
rect 4136 16436 4146 16492
rect 9182 16436 9192 16492
rect 9456 16436 9466 16492
rect 14502 16436 14512 16492
rect 14776 16436 14786 16492
rect 19822 16436 19832 16492
rect 20096 16436 20106 16492
rect 6522 15652 6532 15708
rect 6796 15652 6806 15708
rect 11842 15652 11852 15708
rect 12116 15652 12126 15708
rect 17162 15652 17172 15708
rect 17436 15652 17446 15708
rect 22482 15652 22492 15708
rect 22756 15652 22766 15708
rect 0 14980 800 15008
rect 23200 14980 24000 15008
rect 0 14924 3612 14980
rect 3668 14924 3678 14980
rect 21644 14924 24000 14980
rect 0 14896 800 14924
rect 3862 14868 3872 14924
rect 4136 14868 4146 14924
rect 9182 14868 9192 14924
rect 9456 14868 9466 14924
rect 14502 14868 14512 14924
rect 14776 14868 14786 14924
rect 19822 14868 19832 14924
rect 20096 14868 20106 14924
rect 21644 14756 21700 14924
rect 23200 14896 24000 14924
rect 19618 14700 19628 14756
rect 19684 14700 21700 14756
rect 6522 14084 6532 14140
rect 6796 14084 6806 14140
rect 11842 14084 11852 14140
rect 12116 14084 12126 14140
rect 17162 14084 17172 14140
rect 17436 14084 17446 14140
rect 22482 14084 22492 14140
rect 22756 14084 22766 14140
rect 16258 13468 16268 13524
rect 16324 13468 16940 13524
rect 16996 13468 17388 13524
rect 17444 13468 17612 13524
rect 17668 13468 18396 13524
rect 18452 13468 18462 13524
rect 18946 13468 18956 13524
rect 19012 13468 19628 13524
rect 19684 13468 19694 13524
rect 3862 13300 3872 13356
rect 4136 13300 4146 13356
rect 9182 13300 9192 13356
rect 9456 13300 9466 13356
rect 14502 13300 14512 13356
rect 14776 13300 14786 13356
rect 19822 13300 19832 13356
rect 20096 13300 20106 13356
rect 18498 13244 18508 13300
rect 18564 13244 18574 13300
rect 18508 13188 18564 13244
rect 14914 13132 14924 13188
rect 14980 13132 17052 13188
rect 17108 13132 17724 13188
rect 17780 13132 18284 13188
rect 18340 13132 18844 13188
rect 18900 13132 19180 13188
rect 19236 13132 19246 13188
rect 6522 12516 6532 12572
rect 6796 12516 6806 12572
rect 11842 12516 11852 12572
rect 12116 12516 12126 12572
rect 17162 12516 17172 12572
rect 17436 12516 17446 12572
rect 22482 12516 22492 12572
rect 22756 12516 22766 12572
rect 18386 12236 18396 12292
rect 18452 12236 18956 12292
rect 19012 12236 19022 12292
rect 19730 12236 19740 12292
rect 19796 12236 20412 12292
rect 20468 12236 21084 12292
rect 21140 12236 21150 12292
rect 14802 12124 14812 12180
rect 14868 12124 15484 12180
rect 15540 12124 15550 12180
rect 16146 12124 16156 12180
rect 16212 12124 16828 12180
rect 16884 12124 16894 12180
rect 14242 11900 14252 11956
rect 14308 11900 14924 11956
rect 14980 11900 14990 11956
rect 17602 11788 17612 11844
rect 17668 11788 17678 11844
rect 3862 11732 3872 11788
rect 4136 11732 4146 11788
rect 9182 11732 9192 11788
rect 9456 11732 9466 11788
rect 14502 11732 14512 11788
rect 14776 11732 14786 11788
rect 17612 11732 17668 11788
rect 19822 11732 19832 11788
rect 20096 11732 20106 11788
rect 17612 11676 18508 11732
rect 18564 11676 18574 11732
rect 14914 11340 14924 11396
rect 14980 11340 15596 11396
rect 15652 11340 16268 11396
rect 16324 11340 16940 11396
rect 16996 11340 17500 11396
rect 17556 11340 17566 11396
rect 18946 11340 18956 11396
rect 19012 11340 19516 11396
rect 19572 11340 19852 11396
rect 19908 11340 19918 11396
rect 6178 11228 6188 11284
rect 6244 11228 6972 11284
rect 7028 11228 7038 11284
rect 18274 11116 18284 11172
rect 18340 11116 18508 11172
rect 18564 11116 18956 11172
rect 19012 11116 21756 11172
rect 21812 11116 21822 11172
rect 6522 10948 6532 11004
rect 6796 10948 6806 11004
rect 11842 10948 11852 11004
rect 12116 10948 12126 11004
rect 17162 10948 17172 11004
rect 17436 10948 17446 11004
rect 22482 10948 22492 11004
rect 22756 10948 22766 11004
rect 5506 10668 5516 10724
rect 5572 10668 6076 10724
rect 6132 10668 6142 10724
rect 19842 10668 19852 10724
rect 19908 10668 20188 10724
rect 20244 10668 20254 10724
rect 21074 10668 21084 10724
rect 21140 10668 21868 10724
rect 21924 10668 21934 10724
rect 16818 10332 16828 10388
rect 16884 10332 17836 10388
rect 17892 10332 18284 10388
rect 18340 10332 18508 10388
rect 18564 10332 18574 10388
rect 3862 10164 3872 10220
rect 4136 10164 4146 10220
rect 9182 10164 9192 10220
rect 9456 10164 9466 10220
rect 14502 10164 14512 10220
rect 14776 10164 14786 10220
rect 19822 10164 19832 10220
rect 20096 10164 20106 10220
rect 9986 10108 9996 10164
rect 10052 10108 10062 10164
rect 9996 10052 10052 10108
rect 8978 9996 8988 10052
rect 9044 9996 11340 10052
rect 11396 9996 12012 10052
rect 12068 9996 12078 10052
rect 19842 9996 19852 10052
rect 19908 9996 20524 10052
rect 20580 9996 20590 10052
rect 4274 9772 4284 9828
rect 4340 9772 4844 9828
rect 4900 9772 5404 9828
rect 5460 9772 5470 9828
rect 5842 9660 5852 9716
rect 5908 9660 6524 9716
rect 6580 9660 7196 9716
rect 7252 9660 7262 9716
rect 8988 9604 9044 9996
rect 8642 9548 8652 9604
rect 8708 9548 9324 9604
rect 9380 9548 9390 9604
rect 16482 9548 16492 9604
rect 16548 9548 17164 9604
rect 17220 9548 17230 9604
rect 19170 9548 19180 9604
rect 19236 9548 19852 9604
rect 19908 9548 19918 9604
rect 6522 9380 6532 9436
rect 6796 9380 6806 9436
rect 11842 9380 11852 9436
rect 12116 9380 12126 9436
rect 17162 9380 17172 9436
rect 17436 9380 17446 9436
rect 22482 9380 22492 9436
rect 22756 9380 22766 9436
rect 3490 9100 3500 9156
rect 3556 9100 4060 9156
rect 4116 9100 4126 9156
rect 14354 8988 14364 9044
rect 14420 8988 15036 9044
rect 15092 8988 15260 9044
rect 15316 8988 15326 9044
rect 18946 8764 18956 8820
rect 19012 8764 19180 8820
rect 19236 8764 19246 8820
rect 3862 8596 3872 8652
rect 4136 8596 4146 8652
rect 9182 8596 9192 8652
rect 9456 8596 9466 8652
rect 14502 8596 14512 8652
rect 14776 8596 14786 8652
rect 19822 8596 19832 8652
rect 20096 8596 20106 8652
rect 9986 8540 9996 8596
rect 10052 8540 10556 8596
rect 10612 8540 10622 8596
rect 3602 8428 3612 8484
rect 3668 8428 4172 8484
rect 4228 8428 4732 8484
rect 4788 8428 4956 8484
rect 5012 8428 5404 8484
rect 5460 8428 5964 8484
rect 6020 8428 6524 8484
rect 6580 8428 6590 8484
rect 7186 8428 7196 8484
rect 7252 8428 7980 8484
rect 8036 8428 8540 8484
rect 8596 8428 9324 8484
rect 9380 8428 9390 8484
rect 12786 8428 12796 8484
rect 12852 8428 13692 8484
rect 13748 8428 13916 8484
rect 13972 8428 14364 8484
rect 14420 8428 15148 8484
rect 15204 8428 15708 8484
rect 15764 8428 16380 8484
rect 16436 8428 17164 8484
rect 17220 8428 17836 8484
rect 17892 8428 18508 8484
rect 18564 8428 18956 8484
rect 19012 8428 19022 8484
rect 8978 8316 8988 8372
rect 9044 8316 9884 8372
rect 9940 8316 10332 8372
rect 10388 8316 10398 8372
rect 18386 8316 18396 8372
rect 18452 8316 19180 8372
rect 19236 8316 19246 8372
rect 9202 8204 9212 8260
rect 9268 8204 9996 8260
rect 10052 8204 10062 8260
rect 12450 8204 12460 8260
rect 12516 8204 12908 8260
rect 12964 8204 13356 8260
rect 13412 8204 13804 8260
rect 13860 8204 14476 8260
rect 14532 8204 15036 8260
rect 15092 8204 15596 8260
rect 15652 8204 15820 8260
rect 15876 8204 16268 8260
rect 16324 8204 16492 8260
rect 16548 8204 17052 8260
rect 17108 8204 17612 8260
rect 17668 8204 19068 8260
rect 19124 8204 19628 8260
rect 19684 8204 19694 8260
rect 4274 7980 4284 8036
rect 4340 7980 4844 8036
rect 4900 7980 4910 8036
rect 7298 7980 7308 8036
rect 7364 7980 7980 8036
rect 8036 7980 8316 8036
rect 8372 7980 8382 8036
rect 6522 7812 6532 7868
rect 6796 7812 6806 7868
rect 11842 7812 11852 7868
rect 12116 7812 12126 7868
rect 17162 7812 17172 7868
rect 17436 7812 17446 7868
rect 22482 7812 22492 7868
rect 22756 7812 22766 7868
rect 17826 7644 17836 7700
rect 17892 7644 18396 7700
rect 18452 7644 18462 7700
rect 2146 7420 2156 7476
rect 2212 7420 2716 7476
rect 2772 7420 2782 7476
rect 4834 7420 4844 7476
rect 4900 7420 5404 7476
rect 5460 7420 6076 7476
rect 6132 7420 6142 7476
rect 6738 7420 6748 7476
rect 6804 7420 7308 7476
rect 7364 7420 7374 7476
rect 16594 7420 16604 7476
rect 16660 7420 17612 7476
rect 17668 7420 17678 7476
rect 17714 7308 17724 7364
rect 17780 7308 18396 7364
rect 18452 7308 18462 7364
rect 3602 7196 3612 7252
rect 3668 7196 4172 7252
rect 4228 7196 4238 7252
rect 3862 7028 3872 7084
rect 4136 7028 4146 7084
rect 9182 7028 9192 7084
rect 9456 7028 9466 7084
rect 14502 7028 14512 7084
rect 14776 7028 14786 7084
rect 19822 7028 19832 7084
rect 20096 7028 20106 7084
rect 7522 6860 7532 6916
rect 7588 6860 8876 6916
rect 8932 6860 9996 6916
rect 10052 6860 10062 6916
rect 10546 6860 10556 6916
rect 10612 6860 11228 6916
rect 11284 6860 12012 6916
rect 12068 6860 12078 6916
rect 14018 6860 14028 6916
rect 14084 6860 14252 6916
rect 14308 6860 14588 6916
rect 14644 6860 15260 6916
rect 15316 6860 15326 6916
rect 2818 6748 2828 6804
rect 2884 6748 3724 6804
rect 3780 6748 4620 6804
rect 4676 6748 5516 6804
rect 5572 6748 5740 6804
rect 5796 6748 6412 6804
rect 6468 6748 6478 6804
rect 8530 6636 8540 6692
rect 8596 6636 8764 6692
rect 8820 6636 9212 6692
rect 9268 6636 9884 6692
rect 9940 6636 10444 6692
rect 10500 6636 11116 6692
rect 11172 6636 11900 6692
rect 11956 6636 12460 6692
rect 12516 6636 12526 6692
rect 18946 6636 18956 6692
rect 19012 6636 19180 6692
rect 19236 6636 19628 6692
rect 19684 6636 19694 6692
rect 2146 6524 2156 6580
rect 2212 6524 2828 6580
rect 2884 6524 3388 6580
rect 3444 6524 3454 6580
rect 8418 6524 8428 6580
rect 8484 6524 9100 6580
rect 9156 6524 9166 6580
rect 16930 6524 16940 6580
rect 16996 6524 17500 6580
rect 17556 6524 17566 6580
rect 9874 6412 9884 6468
rect 9940 6412 10556 6468
rect 10612 6412 10622 6468
rect 6522 6244 6532 6300
rect 6796 6244 6806 6300
rect 11842 6244 11852 6300
rect 12116 6244 12126 6300
rect 17162 6244 17172 6300
rect 17436 6244 17446 6300
rect 22482 6244 22492 6300
rect 22756 6244 22766 6300
rect 7074 5964 7084 6020
rect 7140 5964 7420 6020
rect 7476 5964 7756 6020
rect 7812 5964 8092 6020
rect 8148 5964 8158 6020
rect 4050 5852 4060 5908
rect 4116 5852 4732 5908
rect 4788 5852 4798 5908
rect 9090 5852 9100 5908
rect 9156 5852 9772 5908
rect 9828 5852 10444 5908
rect 10500 5852 10510 5908
rect 17826 5852 17836 5908
rect 17892 5852 18396 5908
rect 18452 5852 18462 5908
rect 18162 5740 18172 5796
rect 18228 5740 18508 5796
rect 18564 5740 18732 5796
rect 18788 5740 19180 5796
rect 19236 5740 19246 5796
rect 19842 5628 19852 5684
rect 19908 5628 20300 5684
rect 20356 5628 20524 5684
rect 20580 5628 21196 5684
rect 21252 5628 21644 5684
rect 21700 5628 21710 5684
rect 3862 5460 3872 5516
rect 4136 5460 4146 5516
rect 9182 5460 9192 5516
rect 9456 5460 9466 5516
rect 14502 5460 14512 5516
rect 14776 5460 14786 5516
rect 19822 5460 19832 5516
rect 20096 5460 20106 5516
rect 18844 5180 19516 5236
rect 19572 5180 19582 5236
rect 18844 5124 18900 5180
rect 2706 5068 2716 5124
rect 2772 5068 2782 5124
rect 3378 5068 3388 5124
rect 3444 5068 4172 5124
rect 4228 5068 4956 5124
rect 5012 5068 5022 5124
rect 7298 5068 7308 5124
rect 7364 5068 7756 5124
rect 7812 5068 8540 5124
rect 8596 5068 9100 5124
rect 9156 5068 9660 5124
rect 9716 5068 9726 5124
rect 11554 5068 11564 5124
rect 11620 5068 12124 5124
rect 12180 5068 12190 5124
rect 16146 5068 16156 5124
rect 16212 5068 16828 5124
rect 16884 5068 17388 5124
rect 17444 5068 17454 5124
rect 17602 5068 17612 5124
rect 17668 5068 18508 5124
rect 18564 5068 18844 5124
rect 18900 5068 18910 5124
rect 19058 5068 19068 5124
rect 19124 5068 19404 5124
rect 19460 5068 19852 5124
rect 19908 5068 20076 5124
rect 20132 5068 20142 5124
rect 0 5012 800 5040
rect 2716 5012 2772 5068
rect 23200 5012 24000 5040
rect 0 4956 3612 5012
rect 3668 4956 3678 5012
rect 14690 4956 14700 5012
rect 14756 4956 16044 5012
rect 16100 4956 16716 5012
rect 16772 4956 17724 5012
rect 17780 4956 17790 5012
rect 20178 4956 20188 5012
rect 20244 4956 20412 5012
rect 20468 4956 20748 5012
rect 20804 4956 21644 5012
rect 21700 4956 21710 5012
rect 21970 4956 21980 5012
rect 22036 4956 24000 5012
rect 0 4928 800 4956
rect 23200 4928 24000 4956
rect 4722 4844 4732 4900
rect 4788 4844 4956 4900
rect 5012 4844 5404 4900
rect 5460 4844 5852 4900
rect 5908 4844 6076 4900
rect 6132 4844 6142 4900
rect 12338 4844 12348 4900
rect 12404 4844 12908 4900
rect 12964 4844 12974 4900
rect 6522 4676 6532 4732
rect 6796 4676 6806 4732
rect 11842 4676 11852 4732
rect 12116 4676 12126 4732
rect 17162 4676 17172 4732
rect 17436 4676 17446 4732
rect 22482 4676 22492 4732
rect 22756 4676 22766 4732
rect 3826 4508 3836 4564
rect 3892 4508 4508 4564
rect 4564 4508 4844 4564
rect 4900 4508 5740 4564
rect 5796 4508 6300 4564
rect 6356 4508 6366 4564
rect 2370 4396 2380 4452
rect 2436 4396 3052 4452
rect 3108 4396 3118 4452
rect 16482 4396 16492 4452
rect 16548 4396 17724 4452
rect 17780 4396 18172 4452
rect 18228 4396 18396 4452
rect 18452 4396 18462 4452
rect 2482 4284 2492 4340
rect 2548 4284 2828 4340
rect 2884 4284 3164 4340
rect 3220 4284 3500 4340
rect 3556 4284 3724 4340
rect 3780 4284 4396 4340
rect 4452 4284 4462 4340
rect 7074 4284 7084 4340
rect 7140 4284 7756 4340
rect 7812 4284 7822 4340
rect 14466 4284 14476 4340
rect 14532 4284 14700 4340
rect 14756 4284 15036 4340
rect 15092 4284 15708 4340
rect 15764 4284 15774 4340
rect 19170 4284 19180 4340
rect 19236 4284 19740 4340
rect 19796 4284 20412 4340
rect 20468 4284 20478 4340
rect 4274 4060 4284 4116
rect 4340 4060 5852 4116
rect 5908 4060 6076 4116
rect 6132 4060 6524 4116
rect 6580 4060 7084 4116
rect 7140 4060 7150 4116
rect 12450 4060 12460 4116
rect 12516 4060 13132 4116
rect 13188 4060 13804 4116
rect 13860 4060 13870 4116
rect 3862 3892 3872 3948
rect 4136 3892 4146 3948
rect 9182 3892 9192 3948
rect 9456 3892 9466 3948
rect 14502 3892 14512 3948
rect 14776 3892 14786 3948
rect 19822 3892 19832 3948
rect 20096 3892 20106 3948
rect 2146 3500 2156 3556
rect 2212 3500 2828 3556
rect 2884 3500 2894 3556
rect 3042 3500 3052 3556
rect 3108 3500 3500 3556
rect 3556 3500 4172 3556
rect 4228 3500 4238 3556
rect 7074 3500 7084 3556
rect 7140 3500 7756 3556
rect 7812 3500 8428 3556
rect 8484 3500 9660 3556
rect 9716 3500 9884 3556
rect 9940 3500 10332 3556
rect 10388 3500 11116 3556
rect 11172 3500 11676 3556
rect 11732 3500 11742 3556
rect 4386 3388 4396 3444
rect 4452 3388 4844 3444
rect 4900 3388 5180 3444
rect 5236 3388 5740 3444
rect 5796 3388 6636 3444
rect 6692 3388 11004 3444
rect 11060 3388 11788 3444
rect 11844 3388 11854 3444
rect 14018 3388 14028 3444
rect 14084 3388 14700 3444
rect 14756 3388 15372 3444
rect 15428 3388 15708 3444
rect 15764 3388 16044 3444
rect 16100 3388 16716 3444
rect 16772 3388 17836 3444
rect 17892 3388 18284 3444
rect 18340 3388 18956 3444
rect 19012 3388 19180 3444
rect 19236 3388 19516 3444
rect 19572 3388 19582 3444
rect 6522 3108 6532 3164
rect 6796 3108 6806 3164
rect 11842 3108 11852 3164
rect 12116 3108 12126 3164
rect 17162 3108 17172 3164
rect 17436 3108 17446 3164
rect 22482 3108 22492 3164
rect 22756 3108 22766 3164
<< via3 >>
rect 3872 16436 4136 16492
rect 9192 16436 9456 16492
rect 14512 16436 14776 16492
rect 19832 16436 20096 16492
rect 6532 15652 6796 15708
rect 11852 15652 12116 15708
rect 17172 15652 17436 15708
rect 22492 15652 22756 15708
rect 3872 14868 4136 14924
rect 9192 14868 9456 14924
rect 14512 14868 14776 14924
rect 19832 14868 20096 14924
rect 6532 14084 6796 14140
rect 11852 14084 12116 14140
rect 17172 14084 17436 14140
rect 22492 14084 22756 14140
rect 3872 13300 4136 13356
rect 9192 13300 9456 13356
rect 14512 13300 14776 13356
rect 19832 13300 20096 13356
rect 6532 12516 6796 12572
rect 11852 12516 12116 12572
rect 17172 12516 17436 12572
rect 22492 12516 22756 12572
rect 3872 11732 4136 11788
rect 9192 11732 9456 11788
rect 14512 11732 14776 11788
rect 19832 11732 20096 11788
rect 6532 10948 6796 11004
rect 11852 10948 12116 11004
rect 17172 10948 17436 11004
rect 22492 10948 22756 11004
rect 3872 10164 4136 10220
rect 9192 10164 9456 10220
rect 14512 10164 14776 10220
rect 19832 10164 20096 10220
rect 6532 9380 6796 9436
rect 11852 9380 12116 9436
rect 17172 9380 17436 9436
rect 22492 9380 22756 9436
rect 3872 8596 4136 8652
rect 9192 8596 9456 8652
rect 14512 8596 14776 8652
rect 19832 8596 20096 8652
rect 6532 7812 6796 7868
rect 11852 7812 12116 7868
rect 17172 7812 17436 7868
rect 22492 7812 22756 7868
rect 3872 7028 4136 7084
rect 9192 7028 9456 7084
rect 14512 7028 14776 7084
rect 19832 7028 20096 7084
rect 6532 6244 6796 6300
rect 11852 6244 12116 6300
rect 17172 6244 17436 6300
rect 22492 6244 22756 6300
rect 3872 5460 4136 5516
rect 9192 5460 9456 5516
rect 14512 5460 14776 5516
rect 19832 5460 20096 5516
rect 6532 4676 6796 4732
rect 11852 4676 12116 4732
rect 17172 4676 17436 4732
rect 22492 4676 22756 4732
rect 3872 3892 4136 3948
rect 9192 3892 9456 3948
rect 14512 3892 14776 3948
rect 19832 3892 20096 3948
rect 6532 3108 6796 3164
rect 11852 3108 12116 3164
rect 17172 3108 17436 3164
rect 22492 3108 22756 3164
<< metal4 >>
rect 3844 16492 4164 16524
rect 3844 16436 3872 16492
rect 4136 16436 4164 16492
rect 3844 14924 4164 16436
rect 3844 14868 3872 14924
rect 4136 14868 4164 14924
rect 3844 13356 4164 14868
rect 3844 13300 3872 13356
rect 4136 13300 4164 13356
rect 3844 11788 4164 13300
rect 3844 11732 3872 11788
rect 4136 11732 4164 11788
rect 3844 10220 4164 11732
rect 3844 10164 3872 10220
rect 4136 10164 4164 10220
rect 3844 8652 4164 10164
rect 3844 8596 3872 8652
rect 4136 8596 4164 8652
rect 3844 7084 4164 8596
rect 3844 7028 3872 7084
rect 4136 7028 4164 7084
rect 3844 5516 4164 7028
rect 3844 5460 3872 5516
rect 4136 5460 4164 5516
rect 3844 3948 4164 5460
rect 3844 3892 3872 3948
rect 4136 3892 4164 3948
rect 3844 3076 4164 3892
rect 6504 15708 6824 16524
rect 6504 15652 6532 15708
rect 6796 15652 6824 15708
rect 6504 14140 6824 15652
rect 6504 14084 6532 14140
rect 6796 14084 6824 14140
rect 6504 12572 6824 14084
rect 6504 12516 6532 12572
rect 6796 12516 6824 12572
rect 6504 11004 6824 12516
rect 6504 10948 6532 11004
rect 6796 10948 6824 11004
rect 6504 9436 6824 10948
rect 6504 9380 6532 9436
rect 6796 9380 6824 9436
rect 6504 7868 6824 9380
rect 6504 7812 6532 7868
rect 6796 7812 6824 7868
rect 6504 6300 6824 7812
rect 6504 6244 6532 6300
rect 6796 6244 6824 6300
rect 6504 4732 6824 6244
rect 6504 4676 6532 4732
rect 6796 4676 6824 4732
rect 6504 3164 6824 4676
rect 6504 3108 6532 3164
rect 6796 3108 6824 3164
rect 6504 3076 6824 3108
rect 9164 16492 9484 16524
rect 9164 16436 9192 16492
rect 9456 16436 9484 16492
rect 9164 14924 9484 16436
rect 9164 14868 9192 14924
rect 9456 14868 9484 14924
rect 9164 13356 9484 14868
rect 9164 13300 9192 13356
rect 9456 13300 9484 13356
rect 9164 11788 9484 13300
rect 9164 11732 9192 11788
rect 9456 11732 9484 11788
rect 9164 10220 9484 11732
rect 9164 10164 9192 10220
rect 9456 10164 9484 10220
rect 9164 8652 9484 10164
rect 9164 8596 9192 8652
rect 9456 8596 9484 8652
rect 9164 7084 9484 8596
rect 9164 7028 9192 7084
rect 9456 7028 9484 7084
rect 9164 5516 9484 7028
rect 9164 5460 9192 5516
rect 9456 5460 9484 5516
rect 9164 3948 9484 5460
rect 9164 3892 9192 3948
rect 9456 3892 9484 3948
rect 9164 3076 9484 3892
rect 11824 15708 12144 16524
rect 11824 15652 11852 15708
rect 12116 15652 12144 15708
rect 11824 14140 12144 15652
rect 11824 14084 11852 14140
rect 12116 14084 12144 14140
rect 11824 12572 12144 14084
rect 11824 12516 11852 12572
rect 12116 12516 12144 12572
rect 11824 11004 12144 12516
rect 11824 10948 11852 11004
rect 12116 10948 12144 11004
rect 11824 9436 12144 10948
rect 11824 9380 11852 9436
rect 12116 9380 12144 9436
rect 11824 7868 12144 9380
rect 11824 7812 11852 7868
rect 12116 7812 12144 7868
rect 11824 6300 12144 7812
rect 11824 6244 11852 6300
rect 12116 6244 12144 6300
rect 11824 4732 12144 6244
rect 11824 4676 11852 4732
rect 12116 4676 12144 4732
rect 11824 3164 12144 4676
rect 11824 3108 11852 3164
rect 12116 3108 12144 3164
rect 11824 3076 12144 3108
rect 14484 16492 14804 16524
rect 14484 16436 14512 16492
rect 14776 16436 14804 16492
rect 14484 14924 14804 16436
rect 14484 14868 14512 14924
rect 14776 14868 14804 14924
rect 14484 13356 14804 14868
rect 14484 13300 14512 13356
rect 14776 13300 14804 13356
rect 14484 11788 14804 13300
rect 14484 11732 14512 11788
rect 14776 11732 14804 11788
rect 14484 10220 14804 11732
rect 14484 10164 14512 10220
rect 14776 10164 14804 10220
rect 14484 8652 14804 10164
rect 14484 8596 14512 8652
rect 14776 8596 14804 8652
rect 14484 7084 14804 8596
rect 14484 7028 14512 7084
rect 14776 7028 14804 7084
rect 14484 5516 14804 7028
rect 14484 5460 14512 5516
rect 14776 5460 14804 5516
rect 14484 3948 14804 5460
rect 14484 3892 14512 3948
rect 14776 3892 14804 3948
rect 14484 3076 14804 3892
rect 17144 15708 17464 16524
rect 17144 15652 17172 15708
rect 17436 15652 17464 15708
rect 17144 14140 17464 15652
rect 17144 14084 17172 14140
rect 17436 14084 17464 14140
rect 17144 12572 17464 14084
rect 17144 12516 17172 12572
rect 17436 12516 17464 12572
rect 17144 11004 17464 12516
rect 17144 10948 17172 11004
rect 17436 10948 17464 11004
rect 17144 9436 17464 10948
rect 17144 9380 17172 9436
rect 17436 9380 17464 9436
rect 17144 7868 17464 9380
rect 17144 7812 17172 7868
rect 17436 7812 17464 7868
rect 17144 6300 17464 7812
rect 17144 6244 17172 6300
rect 17436 6244 17464 6300
rect 17144 4732 17464 6244
rect 17144 4676 17172 4732
rect 17436 4676 17464 4732
rect 17144 3164 17464 4676
rect 17144 3108 17172 3164
rect 17436 3108 17464 3164
rect 17144 3076 17464 3108
rect 19804 16492 20124 16524
rect 19804 16436 19832 16492
rect 20096 16436 20124 16492
rect 19804 14924 20124 16436
rect 19804 14868 19832 14924
rect 20096 14868 20124 14924
rect 19804 13356 20124 14868
rect 19804 13300 19832 13356
rect 20096 13300 20124 13356
rect 19804 11788 20124 13300
rect 19804 11732 19832 11788
rect 20096 11732 20124 11788
rect 19804 10220 20124 11732
rect 19804 10164 19832 10220
rect 20096 10164 20124 10220
rect 19804 8652 20124 10164
rect 19804 8596 19832 8652
rect 20096 8596 20124 8652
rect 19804 7084 20124 8596
rect 19804 7028 19832 7084
rect 20096 7028 20124 7084
rect 19804 5516 20124 7028
rect 19804 5460 19832 5516
rect 20096 5460 20124 5516
rect 19804 3948 20124 5460
rect 19804 3892 19832 3948
rect 20096 3892 20124 3948
rect 19804 3076 20124 3892
rect 22464 15708 22784 16524
rect 22464 15652 22492 15708
rect 22756 15652 22784 15708
rect 22464 14140 22784 15652
rect 22464 14084 22492 14140
rect 22756 14084 22784 14140
rect 22464 12572 22784 14084
rect 22464 12516 22492 12572
rect 22756 12516 22784 12572
rect 22464 11004 22784 12516
rect 22464 10948 22492 11004
rect 22756 10948 22784 11004
rect 22464 9436 22784 10948
rect 22464 9380 22492 9436
rect 22756 9380 22784 9436
rect 22464 7868 22784 9380
rect 22464 7812 22492 7868
rect 22756 7812 22784 7868
rect 22464 6300 22784 7812
rect 22464 6244 22492 6300
rect 22756 6244 22784 6300
rect 22464 4732 22784 6244
rect 22464 4676 22492 4732
rect 22756 4676 22784 4732
rect 22464 3164 22784 4676
rect 22464 3108 22492 3164
rect 22756 3108 22784 3164
rect 22464 3076 22784 3108
<< labels >>
rlabel metal1 s 11984 16464 11984 16464 4 vdd
rlabel metal2 s 12064 15680 12064 15680 4 vss
rlabel metal3 s 4592 5096 4592 5096 4 nbusin_nshunt
rlabel metal2 s 20216 10976 20216 10976 4 nbusout
rlabel metal3 s 20888 5656 20888 5656 4 nseries_gy
rlabel metal2 s 21784 2422 21784 2422 4 nseries_gygy
rlabel metal3 s 5992 4088 5992 4088 4 nshunt_gy
rlabel metal2 s 2856 5600 2856 5600 4 pbusin_pshunt
rlabel metal3 s 22610 4984 22610 4984 4 pbusout
rlabel metal2 s 7896 8316 7896 8316 4 pseries_gy
rlabel metal2 s 20216 5880 20216 5880 4 pseries_gygy
rlabel metal2 s 6552 3752 6552 3752 4 pshunt_gy
flabel metal3 s 0 14896 800 15008 0 FreeSans 560 0 0 0 nbusin_nshunt
port 1 nsew
flabel metal3 s 23200 14896 24000 15008 0 FreeSans 560 0 0 0 nbusout
port 2 nsew
flabel metal2 s 13888 0 14000 800 0 FreeSans 560 90 0 0 nseries_gy
port 3 nsew
flabel metal2 s 21728 0 21840 800 0 FreeSans 560 90 0 0 nseries_gygy
port 4 nsew
flabel metal2 s 6048 0 6160 800 0 FreeSans 560 90 0 0 nshunt_gy
port 5 nsew
flabel metal3 s 0 4928 800 5040 0 FreeSans 560 0 0 0 pbusin_pshunt
port 6 nsew
flabel metal3 s 23200 4928 24000 5040 0 FreeSans 560 0 0 0 pbusout
port 7 nsew
flabel metal2 s 9968 0 10080 800 0 FreeSans 560 90 0 0 pseries_gy
port 8 nsew
flabel metal2 s 17808 0 17920 800 0 FreeSans 560 90 0 0 pseries_gygy
port 9 nsew
flabel metal2 s 2128 0 2240 800 0 FreeSans 560 90 0 0 pshunt_gy
port 10 nsew
flabel metal4 s 3844 3076 4164 16524 0 FreeSans 1600 90 0 0 vdd
port 11 nsew
flabel metal4 s 9164 3076 9484 16524 0 FreeSans 1600 90 0 0 vdd
port 11 nsew
flabel metal4 s 14484 3076 14804 16524 0 FreeSans 1600 90 0 0 vdd
port 11 nsew
flabel metal4 s 19804 3076 20124 16524 0 FreeSans 1600 90 0 0 vdd
port 11 nsew
flabel metal4 s 6504 3076 6824 16524 0 FreeSans 1600 90 0 0 vss
port 12 nsew
flabel metal4 s 11824 3076 12144 16524 0 FreeSans 1600 90 0 0 vss
port 12 nsew
flabel metal4 s 17144 3076 17464 16524 0 FreeSans 1600 90 0 0 vss
port 12 nsew
flabel metal4 s 22464 3076 22784 16524 0 FreeSans 1600 90 0 0 vss
port 12 nsew
<< end >>
