magic
tech gf180mcuC
magscale 1 5
timestamp 1669922097
<< metal1 >>
rect 672 28237 19320 28254
rect 672 28211 9919 28237
rect 9945 28211 9971 28237
rect 9997 28211 10023 28237
rect 10049 28211 19320 28237
rect 672 28194 19320 28211
rect 672 27845 19320 27862
rect 672 27819 2239 27845
rect 2265 27819 2291 27845
rect 2317 27819 2343 27845
rect 2369 27819 17599 27845
rect 17625 27819 17651 27845
rect 17677 27819 17703 27845
rect 17729 27819 19320 27845
rect 672 27802 19320 27819
rect 672 27453 19320 27470
rect 672 27427 9919 27453
rect 9945 27427 9971 27453
rect 9997 27427 10023 27453
rect 10049 27427 19320 27453
rect 672 27410 19320 27427
rect 672 27061 19320 27078
rect 672 27035 2239 27061
rect 2265 27035 2291 27061
rect 2317 27035 2343 27061
rect 2369 27035 17599 27061
rect 17625 27035 17651 27061
rect 17677 27035 17703 27061
rect 17729 27035 19320 27061
rect 672 27018 19320 27035
rect 3369 26839 3375 26865
rect 3401 26839 3407 26865
rect 3817 26839 3823 26865
rect 3849 26839 3855 26865
rect 4489 26839 4495 26865
rect 4521 26839 4527 26865
rect 672 26669 19320 26686
rect 672 26643 9919 26669
rect 9945 26643 9971 26669
rect 9997 26643 10023 26669
rect 10049 26643 19320 26669
rect 672 26626 19320 26643
rect 4489 26503 4495 26529
rect 4521 26503 4527 26529
rect 5833 26503 5839 26529
rect 5865 26503 5871 26529
rect 3313 26447 3319 26473
rect 3345 26447 3351 26473
rect 4489 26447 4495 26473
rect 4521 26447 4527 26473
rect 5161 26447 5167 26473
rect 5193 26447 5199 26473
rect 5721 26447 5727 26473
rect 5753 26447 5759 26473
rect 672 26277 19320 26294
rect 672 26251 2239 26277
rect 2265 26251 2291 26277
rect 2317 26251 2343 26277
rect 2369 26251 17599 26277
rect 17625 26251 17651 26277
rect 17677 26251 17703 26277
rect 17729 26251 19320 26277
rect 672 26234 19320 26251
rect 3089 26055 3095 26081
rect 3121 26055 3127 26081
rect 3537 26055 3543 26081
rect 3569 26055 3575 26081
rect 3761 26055 3767 26081
rect 3793 26055 3799 26081
rect 4825 26055 4831 26081
rect 4857 26055 4863 26081
rect 5721 26055 5727 26081
rect 5753 26055 5759 26081
rect 5721 25999 5727 26025
rect 5753 25999 5759 26025
rect 672 25885 19320 25902
rect 672 25859 9919 25885
rect 9945 25859 9971 25885
rect 9997 25859 10023 25885
rect 10049 25859 19320 25885
rect 672 25842 19320 25859
rect 2809 25719 2815 25745
rect 2841 25719 2847 25745
rect 5833 25719 5839 25745
rect 5865 25719 5871 25745
rect 18551 25689 18577 25695
rect 1633 25663 1639 25689
rect 1665 25663 1671 25689
rect 2809 25663 2815 25689
rect 2841 25663 2847 25689
rect 3089 25663 3095 25689
rect 3121 25663 3127 25689
rect 3537 25663 3543 25689
rect 3569 25663 3575 25689
rect 3761 25663 3767 25689
rect 3793 25663 3799 25689
rect 5161 25663 5167 25689
rect 5193 25663 5199 25689
rect 5721 25663 5727 25689
rect 5753 25663 5759 25689
rect 18551 25657 18577 25663
rect 18663 25689 18689 25695
rect 18663 25657 18689 25663
rect 18831 25689 18857 25695
rect 18831 25657 18857 25663
rect 672 25493 19320 25510
rect 672 25467 2239 25493
rect 2265 25467 2291 25493
rect 2317 25467 2343 25493
rect 2369 25467 17599 25493
rect 17625 25467 17651 25493
rect 17677 25467 17703 25493
rect 17729 25467 19320 25493
rect 672 25450 19320 25467
rect 18775 25297 18801 25303
rect 1577 25271 1583 25297
rect 1609 25271 1615 25297
rect 2473 25271 2479 25297
rect 2505 25271 2511 25297
rect 3089 25271 3095 25297
rect 3121 25271 3127 25297
rect 3537 25271 3543 25297
rect 3569 25271 3575 25297
rect 3761 25271 3767 25297
rect 3793 25271 3799 25297
rect 4881 25271 4887 25297
rect 4913 25271 4919 25297
rect 5777 25271 5783 25297
rect 5809 25271 5815 25297
rect 7121 25271 7127 25297
rect 7153 25271 7159 25297
rect 8017 25271 8023 25297
rect 8049 25271 8055 25297
rect 18775 25265 18801 25271
rect 18887 25297 18913 25303
rect 18887 25265 18913 25271
rect 19055 25297 19081 25303
rect 19055 25265 19081 25271
rect 18103 25241 18129 25247
rect 2473 25215 2479 25241
rect 2505 25215 2511 25241
rect 5777 25215 5783 25241
rect 5809 25215 5815 25241
rect 8017 25215 8023 25241
rect 8049 25215 8055 25241
rect 18103 25209 18129 25215
rect 18215 25241 18241 25247
rect 18215 25209 18241 25215
rect 18383 25241 18409 25247
rect 18383 25209 18409 25215
rect 672 25101 19320 25118
rect 672 25075 9919 25101
rect 9945 25075 9971 25101
rect 9997 25075 10023 25101
rect 10049 25075 19320 25101
rect 672 25058 19320 25075
rect 17823 24961 17849 24967
rect 5833 24935 5839 24961
rect 5865 24935 5871 24961
rect 7513 24935 7519 24961
rect 7545 24935 7551 24961
rect 17823 24929 17849 24935
rect 17991 24961 18017 24967
rect 17991 24929 18017 24935
rect 18383 24961 18409 24967
rect 18383 24929 18409 24935
rect 18551 24961 18577 24967
rect 18551 24929 18577 24935
rect 17711 24905 17737 24911
rect 1633 24879 1639 24905
rect 1665 24879 1671 24905
rect 2081 24879 2087 24905
rect 2113 24879 2119 24905
rect 2305 24879 2311 24905
rect 2337 24879 2343 24905
rect 3089 24879 3095 24905
rect 3121 24879 3127 24905
rect 3537 24879 3543 24905
rect 3569 24879 3575 24905
rect 3761 24879 3767 24905
rect 3793 24879 3799 24905
rect 4881 24879 4887 24905
rect 4913 24879 4919 24905
rect 5833 24879 5839 24905
rect 5865 24879 5871 24905
rect 6617 24879 6623 24905
rect 6649 24879 6655 24905
rect 7513 24879 7519 24905
rect 7545 24879 7551 24905
rect 17711 24873 17737 24879
rect 18327 24905 18353 24911
rect 18327 24873 18353 24879
rect 672 24709 19320 24726
rect 672 24683 2239 24709
rect 2265 24683 2291 24709
rect 2317 24683 2343 24709
rect 2369 24683 17599 24709
rect 17625 24683 17651 24709
rect 17677 24683 17703 24709
rect 17729 24683 19320 24709
rect 672 24666 19320 24683
rect 17151 24513 17177 24519
rect 1577 24487 1583 24513
rect 1609 24487 1615 24513
rect 2137 24487 2143 24513
rect 2169 24487 2175 24513
rect 3089 24487 3095 24513
rect 3121 24487 3127 24513
rect 3537 24487 3543 24513
rect 3569 24487 3575 24513
rect 3761 24487 3767 24513
rect 3793 24487 3799 24513
rect 4881 24487 4887 24513
rect 4913 24487 4919 24513
rect 5777 24487 5783 24513
rect 5809 24487 5815 24513
rect 7065 24487 7071 24513
rect 7097 24487 7103 24513
rect 7961 24487 7967 24513
rect 7993 24487 7999 24513
rect 8577 24487 8583 24513
rect 8609 24487 8615 24513
rect 9473 24487 9479 24513
rect 9505 24487 9511 24513
rect 17151 24481 17177 24487
rect 17319 24513 17345 24519
rect 17319 24481 17345 24487
rect 17543 24513 17569 24519
rect 17543 24481 17569 24487
rect 17711 24513 17737 24519
rect 17711 24481 17737 24487
rect 17879 24513 17905 24519
rect 17879 24481 17905 24487
rect 18271 24513 18297 24519
rect 18271 24481 18297 24487
rect 18439 24513 18465 24519
rect 18439 24481 18465 24487
rect 18775 24513 18801 24519
rect 18775 24481 18801 24487
rect 18887 24513 18913 24519
rect 18887 24481 18913 24487
rect 18999 24513 19025 24519
rect 18999 24481 19025 24487
rect 16983 24457 17009 24463
rect 2249 24431 2255 24457
rect 2281 24431 2287 24457
rect 5777 24431 5783 24457
rect 5809 24431 5815 24457
rect 7961 24431 7967 24457
rect 7993 24431 7999 24457
rect 9473 24431 9479 24457
rect 9505 24431 9511 24457
rect 16983 24425 17009 24431
rect 18103 24457 18129 24463
rect 18103 24425 18129 24431
rect 672 24317 19320 24334
rect 672 24291 9919 24317
rect 9945 24291 9971 24317
rect 9997 24291 10023 24317
rect 10049 24291 19320 24317
rect 672 24274 19320 24291
rect 17263 24177 17289 24183
rect 5833 24151 5839 24177
rect 5865 24151 5871 24177
rect 7513 24151 7519 24177
rect 7545 24151 7551 24177
rect 9809 24151 9815 24177
rect 9841 24151 9847 24177
rect 17263 24145 17289 24151
rect 17431 24177 17457 24183
rect 17431 24145 17457 24151
rect 17711 24177 17737 24183
rect 17711 24145 17737 24151
rect 17823 24177 17849 24183
rect 17823 24145 17849 24151
rect 17991 24177 18017 24183
rect 17991 24145 18017 24151
rect 18383 24177 18409 24183
rect 18383 24145 18409 24151
rect 18551 24177 18577 24183
rect 18551 24145 18577 24151
rect 17207 24121 17233 24127
rect 1857 24095 1863 24121
rect 1889 24095 1895 24121
rect 2305 24095 2311 24121
rect 2337 24095 2343 24121
rect 2529 24095 2535 24121
rect 2561 24095 2567 24121
rect 3313 24095 3319 24121
rect 3345 24095 3351 24121
rect 3761 24095 3767 24121
rect 3793 24095 3799 24121
rect 3985 24095 3991 24121
rect 4017 24095 4023 24121
rect 5161 24095 5167 24121
rect 5193 24095 5199 24121
rect 5833 24095 5839 24121
rect 5865 24095 5871 24121
rect 6337 24095 6343 24121
rect 6369 24095 6375 24121
rect 7513 24095 7519 24121
rect 7545 24095 7551 24121
rect 9137 24095 9143 24121
rect 9169 24095 9175 24121
rect 9809 24095 9815 24121
rect 9841 24095 9847 24121
rect 17207 24089 17233 24095
rect 18327 24121 18353 24127
rect 18327 24089 18353 24095
rect 672 23925 19320 23942
rect 672 23899 2239 23925
rect 2265 23899 2291 23925
rect 2317 23899 2343 23925
rect 2369 23899 17599 23925
rect 17625 23899 17651 23925
rect 17677 23899 17703 23925
rect 17729 23899 19320 23925
rect 672 23882 19320 23899
rect 16479 23729 16505 23735
rect 1577 23703 1583 23729
rect 1609 23703 1615 23729
rect 2473 23703 2479 23729
rect 2505 23703 2511 23729
rect 3145 23703 3151 23729
rect 3177 23703 3183 23729
rect 3593 23703 3599 23729
rect 3625 23703 3631 23729
rect 3817 23703 3823 23729
rect 3849 23703 3855 23729
rect 4881 23703 4887 23729
rect 4913 23703 4919 23729
rect 5777 23703 5783 23729
rect 5809 23703 5815 23729
rect 7121 23703 7127 23729
rect 7153 23703 7159 23729
rect 8017 23703 8023 23729
rect 8049 23703 8055 23729
rect 8577 23703 8583 23729
rect 8609 23703 8615 23729
rect 9417 23703 9423 23729
rect 9449 23703 9455 23729
rect 16479 23697 16505 23703
rect 16591 23729 16617 23735
rect 16591 23697 16617 23703
rect 16759 23729 16785 23735
rect 16759 23697 16785 23703
rect 17039 23729 17065 23735
rect 17039 23697 17065 23703
rect 17151 23729 17177 23735
rect 17151 23697 17177 23703
rect 17263 23729 17289 23735
rect 17263 23697 17289 23703
rect 17599 23729 17625 23735
rect 17599 23697 17625 23703
rect 17711 23729 17737 23735
rect 17711 23697 17737 23703
rect 17879 23729 17905 23735
rect 17879 23697 17905 23703
rect 18159 23729 18185 23735
rect 18159 23697 18185 23703
rect 18383 23729 18409 23735
rect 18383 23697 18409 23703
rect 18719 23729 18745 23735
rect 18719 23697 18745 23703
rect 18999 23729 19025 23735
rect 18999 23697 19025 23703
rect 18215 23673 18241 23679
rect 2473 23647 2479 23673
rect 2505 23647 2511 23673
rect 5777 23647 5783 23673
rect 5809 23647 5815 23673
rect 8017 23647 8023 23673
rect 8049 23647 8055 23673
rect 9417 23647 9423 23673
rect 9449 23647 9455 23673
rect 18215 23641 18241 23647
rect 18943 23673 18969 23679
rect 18943 23641 18969 23647
rect 672 23533 19320 23550
rect 672 23507 9919 23533
rect 9945 23507 9971 23533
rect 9997 23507 10023 23533
rect 10049 23507 19320 23533
rect 672 23490 19320 23507
rect 17431 23393 17457 23399
rect 4433 23367 4439 23393
rect 4465 23367 4471 23393
rect 8185 23367 8191 23393
rect 8217 23367 8223 23393
rect 11489 23367 11495 23393
rect 11521 23367 11527 23393
rect 17431 23361 17457 23367
rect 17711 23393 17737 23399
rect 17711 23361 17737 23367
rect 17991 23393 18017 23399
rect 17991 23361 18017 23367
rect 18383 23393 18409 23399
rect 18383 23361 18409 23367
rect 18551 23393 18577 23399
rect 18551 23361 18577 23367
rect 16199 23337 16225 23343
rect 1913 23311 1919 23337
rect 1945 23311 1951 23337
rect 2417 23311 2423 23337
rect 2449 23311 2455 23337
rect 2529 23311 2535 23337
rect 2561 23311 2567 23337
rect 3593 23311 3599 23337
rect 3625 23311 3631 23337
rect 4433 23311 4439 23337
rect 4465 23311 4471 23337
rect 6057 23311 6063 23337
rect 6089 23311 6095 23337
rect 6337 23311 6343 23337
rect 6369 23311 6375 23337
rect 6449 23311 6455 23337
rect 6481 23311 6487 23337
rect 7233 23311 7239 23337
rect 7265 23311 7271 23337
rect 8017 23311 8023 23337
rect 8049 23311 8055 23337
rect 9081 23311 9087 23337
rect 9113 23311 9119 23337
rect 9417 23311 9423 23337
rect 9449 23311 9455 23337
rect 9529 23311 9535 23337
rect 9561 23311 9567 23337
rect 10593 23311 10599 23337
rect 10625 23311 10631 23337
rect 11489 23311 11495 23337
rect 11521 23311 11527 23337
rect 16199 23305 16225 23311
rect 16311 23337 16337 23343
rect 16311 23305 16337 23311
rect 16479 23337 16505 23343
rect 16479 23305 16505 23311
rect 17207 23337 17233 23343
rect 17207 23305 17233 23311
rect 17319 23337 17345 23343
rect 17319 23305 17345 23311
rect 17879 23337 17905 23343
rect 17879 23305 17905 23311
rect 18327 23337 18353 23343
rect 18327 23305 18353 23311
rect 672 23141 19320 23158
rect 672 23115 2239 23141
rect 2265 23115 2291 23141
rect 2317 23115 2343 23141
rect 2369 23115 17599 23141
rect 17625 23115 17651 23141
rect 17677 23115 17703 23141
rect 17729 23115 19320 23141
rect 672 23098 19320 23115
rect 16199 22945 16225 22951
rect 1409 22919 1415 22945
rect 1441 22919 1447 22945
rect 2473 22919 2479 22945
rect 2505 22919 2511 22945
rect 3929 22919 3935 22945
rect 3961 22919 3967 22945
rect 4377 22919 4383 22945
rect 4409 22919 4415 22945
rect 4489 22919 4495 22945
rect 4521 22919 4527 22945
rect 5273 22919 5279 22945
rect 5305 22919 5311 22945
rect 6337 22919 6343 22945
rect 6369 22919 6375 22945
rect 7121 22919 7127 22945
rect 7153 22919 7159 22945
rect 8017 22919 8023 22945
rect 8049 22919 8055 22945
rect 8409 22919 8415 22945
rect 8441 22919 8447 22945
rect 9473 22919 9479 22945
rect 9505 22919 9511 22945
rect 11097 22919 11103 22945
rect 11129 22919 11135 22945
rect 11377 22919 11383 22945
rect 11409 22919 11415 22945
rect 11489 22919 11495 22945
rect 11521 22919 11527 22945
rect 16199 22913 16225 22919
rect 16423 22945 16449 22951
rect 16423 22913 16449 22919
rect 16535 22945 16561 22951
rect 16535 22913 16561 22919
rect 16703 22945 16729 22951
rect 16703 22913 16729 22919
rect 17039 22945 17065 22951
rect 17039 22913 17065 22919
rect 17151 22945 17177 22951
rect 17151 22913 17177 22919
rect 17319 22945 17345 22951
rect 17319 22913 17345 22919
rect 17543 22945 17569 22951
rect 17543 22913 17569 22919
rect 17711 22945 17737 22951
rect 17711 22913 17737 22919
rect 17879 22945 17905 22951
rect 17879 22913 17905 22919
rect 18159 22945 18185 22951
rect 18159 22913 18185 22919
rect 18271 22945 18297 22951
rect 18271 22913 18297 22919
rect 18383 22945 18409 22951
rect 18383 22913 18409 22919
rect 18775 22945 18801 22951
rect 18775 22913 18801 22919
rect 18887 22945 18913 22951
rect 18887 22913 18913 22919
rect 15303 22889 15329 22895
rect 2473 22863 2479 22889
rect 2505 22863 2511 22889
rect 6337 22863 6343 22889
rect 6369 22863 6375 22889
rect 8017 22863 8023 22889
rect 8049 22863 8055 22889
rect 9473 22863 9479 22889
rect 9505 22863 9511 22889
rect 15303 22857 15329 22863
rect 15471 22889 15497 22895
rect 15471 22857 15497 22863
rect 15583 22889 15609 22895
rect 15583 22857 15609 22863
rect 15863 22889 15889 22895
rect 15863 22857 15889 22863
rect 15975 22889 16001 22895
rect 15975 22857 16001 22863
rect 19055 22889 19081 22895
rect 19055 22857 19081 22863
rect 672 22749 19320 22766
rect 672 22723 9919 22749
rect 9945 22723 9971 22749
rect 9997 22723 10023 22749
rect 10049 22723 19320 22749
rect 672 22706 19320 22723
rect 15583 22609 15609 22615
rect 4433 22583 4439 22609
rect 4465 22583 4471 22609
rect 8353 22583 8359 22609
rect 8385 22583 8391 22609
rect 9809 22583 9815 22609
rect 9841 22583 9847 22609
rect 11265 22583 11271 22609
rect 11297 22583 11303 22609
rect 15583 22577 15609 22583
rect 15751 22609 15777 22615
rect 15751 22577 15777 22583
rect 16143 22609 16169 22615
rect 16143 22577 16169 22583
rect 16871 22609 16897 22615
rect 16871 22577 16897 22583
rect 17151 22609 17177 22615
rect 17151 22577 17177 22583
rect 17711 22609 17737 22615
rect 17711 22577 17737 22583
rect 18103 22609 18129 22615
rect 18103 22577 18129 22583
rect 18271 22609 18297 22615
rect 18271 22577 18297 22583
rect 15863 22553 15889 22559
rect 1913 22527 1919 22553
rect 1945 22527 1951 22553
rect 2417 22527 2423 22553
rect 2449 22527 2455 22553
rect 2529 22527 2535 22553
rect 2561 22527 2567 22553
rect 3593 22527 3599 22553
rect 3625 22527 3631 22553
rect 4433 22527 4439 22553
rect 4465 22527 4471 22553
rect 6057 22527 6063 22553
rect 6089 22527 6095 22553
rect 6337 22527 6343 22553
rect 6369 22527 6375 22553
rect 6449 22527 6455 22553
rect 6481 22527 6487 22553
rect 7457 22527 7463 22553
rect 7489 22527 7495 22553
rect 8353 22527 8359 22553
rect 8385 22527 8391 22553
rect 9137 22527 9143 22553
rect 9169 22527 9175 22553
rect 9809 22527 9815 22553
rect 9841 22527 9847 22553
rect 10369 22527 10375 22553
rect 10401 22527 10407 22553
rect 11265 22527 11271 22553
rect 11297 22527 11303 22553
rect 15863 22521 15889 22527
rect 16311 22553 16337 22559
rect 16311 22521 16337 22527
rect 16479 22553 16505 22559
rect 16479 22521 16505 22527
rect 17039 22553 17065 22559
rect 17039 22521 17065 22527
rect 17487 22553 17513 22559
rect 17487 22521 17513 22527
rect 17543 22553 17569 22559
rect 17543 22521 17569 22527
rect 18047 22553 18073 22559
rect 18047 22521 18073 22527
rect 18551 22553 18577 22559
rect 18551 22521 18577 22527
rect 18719 22553 18745 22559
rect 18719 22521 18745 22527
rect 18831 22553 18857 22559
rect 18831 22521 18857 22527
rect 672 22357 19320 22374
rect 672 22331 2239 22357
rect 2265 22331 2291 22357
rect 2317 22331 2343 22357
rect 2369 22331 17599 22357
rect 17625 22331 17651 22357
rect 17677 22331 17703 22357
rect 17729 22331 19320 22357
rect 672 22314 19320 22331
rect 16423 22161 16449 22167
rect 1409 22135 1415 22161
rect 1441 22135 1447 22161
rect 2249 22135 2255 22161
rect 2281 22135 2287 22161
rect 3929 22135 3935 22161
rect 3961 22135 3967 22161
rect 4769 22135 4775 22161
rect 4801 22135 4807 22161
rect 5273 22135 5279 22161
rect 5305 22135 5311 22161
rect 6337 22135 6343 22161
rect 6369 22135 6375 22161
rect 7121 22135 7127 22161
rect 7153 22135 7159 22161
rect 7793 22135 7799 22161
rect 7825 22135 7831 22161
rect 8409 22135 8415 22161
rect 8441 22135 8447 22161
rect 9473 22135 9479 22161
rect 9505 22135 9511 22161
rect 11097 22135 11103 22161
rect 11129 22135 11135 22161
rect 11265 22135 11271 22161
rect 11297 22135 11303 22161
rect 11489 22135 11495 22161
rect 11521 22135 11527 22161
rect 12553 22135 12559 22161
rect 12585 22135 12591 22161
rect 12833 22135 12839 22161
rect 12865 22135 12871 22161
rect 12945 22135 12951 22161
rect 12977 22135 12983 22161
rect 16423 22129 16449 22135
rect 16535 22161 16561 22167
rect 16535 22129 16561 22135
rect 16703 22161 16729 22167
rect 16703 22129 16729 22135
rect 16983 22161 17009 22167
rect 16983 22129 17009 22135
rect 17151 22161 17177 22167
rect 17151 22129 17177 22135
rect 17319 22161 17345 22167
rect 17319 22129 17345 22135
rect 17487 22161 17513 22167
rect 17487 22129 17513 22135
rect 18159 22161 18185 22167
rect 18159 22129 18185 22135
rect 18271 22161 18297 22167
rect 18271 22129 18297 22135
rect 18383 22161 18409 22167
rect 18383 22129 18409 22135
rect 18887 22161 18913 22167
rect 18887 22129 18913 22135
rect 17711 22105 17737 22111
rect 2249 22079 2255 22105
rect 2281 22079 2287 22105
rect 4769 22079 4775 22105
rect 4801 22079 4807 22105
rect 6337 22079 6343 22105
rect 6369 22079 6375 22105
rect 7793 22079 7799 22105
rect 7825 22079 7831 22105
rect 9473 22079 9479 22105
rect 9505 22079 9511 22105
rect 17711 22073 17737 22079
rect 17823 22105 17849 22111
rect 17823 22073 17849 22079
rect 18775 22105 18801 22111
rect 18775 22073 18801 22079
rect 19055 22105 19081 22111
rect 19055 22073 19081 22079
rect 672 21965 19320 21982
rect 672 21939 9919 21965
rect 9945 21939 9971 21965
rect 9997 21939 10023 21965
rect 10049 21939 19320 21965
rect 672 21922 19320 21939
rect 18551 21825 18577 21831
rect 3033 21799 3039 21825
rect 3065 21799 3071 21825
rect 4265 21799 4271 21825
rect 4297 21799 4303 21825
rect 9977 21799 9983 21825
rect 10009 21799 10015 21825
rect 11489 21799 11495 21825
rect 11521 21799 11527 21825
rect 18551 21793 18577 21799
rect 16871 21769 16897 21775
rect 1857 21743 1863 21769
rect 1889 21743 1895 21769
rect 3033 21743 3039 21769
rect 3065 21743 3071 21769
rect 3369 21743 3375 21769
rect 3401 21743 3407 21769
rect 4209 21743 4215 21769
rect 4241 21743 4247 21769
rect 6057 21743 6063 21769
rect 6089 21743 6095 21769
rect 6337 21743 6343 21769
rect 6369 21743 6375 21769
rect 6449 21743 6455 21769
rect 6481 21743 6487 21769
rect 7457 21743 7463 21769
rect 7489 21743 7495 21769
rect 7681 21743 7687 21769
rect 7713 21743 7719 21769
rect 7905 21743 7911 21769
rect 7937 21743 7943 21769
rect 9137 21743 9143 21769
rect 9169 21743 9175 21769
rect 9977 21743 9983 21769
rect 10009 21743 10015 21769
rect 10593 21743 10599 21769
rect 10625 21743 10631 21769
rect 11489 21743 11495 21769
rect 11521 21743 11527 21769
rect 12833 21743 12839 21769
rect 12865 21743 12871 21769
rect 13393 21743 13399 21769
rect 13425 21743 13431 21769
rect 13561 21743 13567 21769
rect 13593 21743 13599 21769
rect 16871 21737 16897 21743
rect 17039 21769 17065 21775
rect 17039 21737 17065 21743
rect 17151 21769 17177 21775
rect 17151 21737 17177 21743
rect 17487 21769 17513 21775
rect 17487 21737 17513 21743
rect 17599 21769 17625 21775
rect 17599 21737 17625 21743
rect 17711 21769 17737 21775
rect 17711 21737 17737 21743
rect 18047 21769 18073 21775
rect 18047 21737 18073 21743
rect 18159 21769 18185 21775
rect 18159 21737 18185 21743
rect 18327 21769 18353 21775
rect 18327 21737 18353 21743
rect 18719 21769 18745 21775
rect 18719 21737 18745 21743
rect 18831 21769 18857 21775
rect 18831 21737 18857 21743
rect 672 21573 19320 21590
rect 672 21547 2239 21573
rect 2265 21547 2291 21573
rect 2317 21547 2343 21573
rect 2369 21547 17599 21573
rect 17625 21547 17651 21573
rect 17677 21547 17703 21573
rect 17729 21547 19320 21573
rect 672 21530 19320 21547
rect 16983 21377 17009 21383
rect 1577 21351 1583 21377
rect 1609 21351 1615 21377
rect 2473 21351 2479 21377
rect 2505 21351 2511 21377
rect 3817 21351 3823 21377
rect 3849 21351 3855 21377
rect 4769 21351 4775 21377
rect 4801 21351 4807 21377
rect 5273 21351 5279 21377
rect 5305 21351 5311 21377
rect 6449 21351 6455 21377
rect 6481 21351 6487 21377
rect 7121 21351 7127 21377
rect 7153 21351 7159 21377
rect 7569 21351 7575 21377
rect 7601 21351 7607 21377
rect 8577 21351 8583 21377
rect 8609 21351 8615 21377
rect 8745 21351 8751 21377
rect 8777 21351 8783 21377
rect 8969 21351 8975 21377
rect 9001 21351 9007 21377
rect 11097 21351 11103 21377
rect 11129 21351 11135 21377
rect 11377 21351 11383 21377
rect 11409 21351 11415 21377
rect 11545 21351 11551 21377
rect 11577 21351 11583 21377
rect 12553 21351 12559 21377
rect 12585 21351 12591 21377
rect 12721 21351 12727 21377
rect 12753 21351 12759 21377
rect 12945 21351 12951 21377
rect 12977 21351 12983 21377
rect 16983 21345 17009 21351
rect 17151 21377 17177 21383
rect 17151 21345 17177 21351
rect 17263 21377 17289 21383
rect 17263 21345 17289 21351
rect 17543 21377 17569 21383
rect 17543 21345 17569 21351
rect 17711 21377 17737 21383
rect 17711 21345 17737 21351
rect 17879 21377 17905 21383
rect 17879 21345 17905 21351
rect 18103 21377 18129 21383
rect 18103 21345 18129 21351
rect 18887 21377 18913 21383
rect 18887 21345 18913 21351
rect 18999 21377 19025 21383
rect 18999 21345 19025 21351
rect 18215 21321 18241 21327
rect 2473 21295 2479 21321
rect 2505 21295 2511 21321
rect 4769 21295 4775 21321
rect 4801 21295 4807 21321
rect 6449 21295 6455 21321
rect 6481 21295 6487 21321
rect 7793 21295 7799 21321
rect 7825 21295 7831 21321
rect 18215 21289 18241 21295
rect 18383 21321 18409 21327
rect 18383 21289 18409 21295
rect 18775 21321 18801 21327
rect 18775 21289 18801 21295
rect 672 21181 19320 21198
rect 672 21155 9919 21181
rect 9945 21155 9971 21181
rect 9997 21155 10023 21181
rect 10049 21155 19320 21181
rect 672 21138 19320 21155
rect 17655 21041 17681 21047
rect 3033 21015 3039 21041
rect 3065 21015 3071 21041
rect 4489 21015 4495 21041
rect 4521 21015 4527 21041
rect 11321 21015 11327 21041
rect 11353 21015 11359 21041
rect 17655 21009 17681 21015
rect 17767 21041 17793 21047
rect 17767 21009 17793 21015
rect 17935 21041 17961 21047
rect 17935 21009 17961 21015
rect 18215 21041 18241 21047
rect 18215 21009 18241 21015
rect 18383 21041 18409 21047
rect 18383 21009 18409 21015
rect 18495 20985 18521 20991
rect 1857 20959 1863 20985
rect 1889 20959 1895 20985
rect 3033 20959 3039 20985
rect 3065 20959 3071 20985
rect 3369 20959 3375 20985
rect 3401 20959 3407 20985
rect 4489 20959 4495 20985
rect 4521 20959 4527 20985
rect 6057 20959 6063 20985
rect 6089 20959 6095 20985
rect 6337 20959 6343 20985
rect 6369 20959 6375 20985
rect 6449 20959 6455 20985
rect 6481 20959 6487 20985
rect 7513 20959 7519 20985
rect 7545 20959 7551 20985
rect 7681 20959 7687 20985
rect 7713 20959 7719 20985
rect 7905 20959 7911 20985
rect 7937 20959 7943 20985
rect 9137 20959 9143 20985
rect 9169 20959 9175 20985
rect 9305 20959 9311 20985
rect 9337 20959 9343 20985
rect 9529 20959 9535 20985
rect 9561 20959 9567 20985
rect 10593 20959 10599 20985
rect 10625 20959 10631 20985
rect 11321 20959 11327 20985
rect 11353 20959 11359 20985
rect 13113 20959 13119 20985
rect 13145 20959 13151 20985
rect 13281 20959 13287 20985
rect 13313 20959 13319 20985
rect 13505 20959 13511 20985
rect 13537 20959 13543 20985
rect 18495 20953 18521 20959
rect 18775 20985 18801 20991
rect 18775 20953 18801 20959
rect 18887 20985 18913 20991
rect 18887 20953 18913 20959
rect 18999 20985 19025 20991
rect 18999 20953 19025 20959
rect 672 20789 19320 20806
rect 672 20763 2239 20789
rect 2265 20763 2291 20789
rect 2317 20763 2343 20789
rect 2369 20763 17599 20789
rect 17625 20763 17651 20789
rect 17677 20763 17703 20789
rect 17729 20763 19320 20789
rect 672 20746 19320 20763
rect 18103 20593 18129 20599
rect 1577 20567 1583 20593
rect 1609 20567 1615 20593
rect 2473 20567 2479 20593
rect 2505 20567 2511 20593
rect 3817 20567 3823 20593
rect 3849 20567 3855 20593
rect 4377 20567 4383 20593
rect 4409 20567 4415 20593
rect 4489 20567 4495 20593
rect 4521 20567 4527 20593
rect 5273 20567 5279 20593
rect 5305 20567 5311 20593
rect 6449 20567 6455 20593
rect 6481 20567 6487 20593
rect 7121 20567 7127 20593
rect 7153 20567 7159 20593
rect 7569 20567 7575 20593
rect 7601 20567 7607 20593
rect 8577 20567 8583 20593
rect 8609 20567 8615 20593
rect 8745 20567 8751 20593
rect 8777 20567 8783 20593
rect 8969 20567 8975 20593
rect 9001 20567 9007 20593
rect 11097 20567 11103 20593
rect 11129 20567 11135 20593
rect 11321 20567 11327 20593
rect 11353 20567 11359 20593
rect 11489 20567 11495 20593
rect 11521 20567 11527 20593
rect 12553 20567 12559 20593
rect 12585 20567 12591 20593
rect 12721 20567 12727 20593
rect 12753 20567 12759 20593
rect 12945 20567 12951 20593
rect 12977 20567 12983 20593
rect 18103 20561 18129 20567
rect 18271 20593 18297 20599
rect 18271 20561 18297 20567
rect 18439 20593 18465 20599
rect 18439 20561 18465 20567
rect 18999 20593 19025 20599
rect 18999 20561 19025 20567
rect 18775 20537 18801 20543
rect 2473 20511 2479 20537
rect 2505 20511 2511 20537
rect 6449 20511 6455 20537
rect 6481 20511 6487 20537
rect 7793 20511 7799 20537
rect 7825 20511 7831 20537
rect 18775 20505 18801 20511
rect 18943 20537 18969 20543
rect 18943 20505 18969 20511
rect 672 20397 19320 20414
rect 672 20371 9919 20397
rect 9945 20371 9971 20397
rect 9997 20371 10023 20397
rect 10049 20371 19320 20397
rect 672 20354 19320 20371
rect 4433 20231 4439 20257
rect 4465 20231 4471 20257
rect 11489 20231 11495 20257
rect 11521 20231 11527 20257
rect 15241 20231 15247 20257
rect 15273 20231 15279 20257
rect 18719 20201 18745 20207
rect 1857 20175 1863 20201
rect 1889 20175 1895 20201
rect 2417 20175 2423 20201
rect 2449 20175 2455 20201
rect 2529 20175 2535 20201
rect 2561 20175 2567 20201
rect 3369 20175 3375 20201
rect 3401 20175 3407 20201
rect 4433 20175 4439 20201
rect 4465 20175 4471 20201
rect 6057 20175 6063 20201
rect 6089 20175 6095 20201
rect 6337 20175 6343 20201
rect 6369 20175 6375 20201
rect 6449 20175 6455 20201
rect 6481 20175 6487 20201
rect 7457 20175 7463 20201
rect 7489 20175 7495 20201
rect 7681 20175 7687 20201
rect 7713 20175 7719 20201
rect 7905 20175 7911 20201
rect 7937 20175 7943 20201
rect 9137 20175 9143 20201
rect 9169 20175 9175 20201
rect 9305 20175 9311 20201
rect 9337 20175 9343 20201
rect 9529 20175 9535 20201
rect 9561 20175 9567 20201
rect 10593 20175 10599 20201
rect 10625 20175 10631 20201
rect 11489 20175 11495 20201
rect 11521 20175 11527 20201
rect 13057 20175 13063 20201
rect 13089 20175 13095 20201
rect 13281 20175 13287 20201
rect 13313 20175 13319 20201
rect 13505 20175 13511 20201
rect 13537 20175 13543 20201
rect 14569 20175 14575 20201
rect 14601 20175 14607 20201
rect 15241 20175 15247 20201
rect 15273 20175 15279 20201
rect 18719 20169 18745 20175
rect 18887 20201 18913 20207
rect 18887 20169 18913 20175
rect 19055 20201 19081 20207
rect 19055 20169 19081 20175
rect 672 20005 19320 20022
rect 672 19979 2239 20005
rect 2265 19979 2291 20005
rect 2317 19979 2343 20005
rect 2369 19979 17599 20005
rect 17625 19979 17651 20005
rect 17677 19979 17703 20005
rect 17729 19979 19320 20005
rect 672 19962 19320 19979
rect 18103 19809 18129 19815
rect 1577 19783 1583 19809
rect 1609 19783 1615 19809
rect 2417 19783 2423 19809
rect 2449 19783 2455 19809
rect 3817 19783 3823 19809
rect 3849 19783 3855 19809
rect 4377 19783 4383 19809
rect 4409 19783 4415 19809
rect 4489 19783 4495 19809
rect 4521 19783 4527 19809
rect 5273 19783 5279 19809
rect 5305 19783 5311 19809
rect 6393 19783 6399 19809
rect 6425 19783 6431 19809
rect 6953 19783 6959 19809
rect 6985 19783 6991 19809
rect 7345 19783 7351 19809
rect 7377 19783 7383 19809
rect 7569 19783 7575 19809
rect 7601 19783 7607 19809
rect 8577 19783 8583 19809
rect 8609 19783 8615 19809
rect 8745 19783 8751 19809
rect 8777 19783 8783 19809
rect 8969 19783 8975 19809
rect 9001 19783 9007 19809
rect 11097 19783 11103 19809
rect 11129 19783 11135 19809
rect 11377 19783 11383 19809
rect 11409 19783 11415 19809
rect 11489 19783 11495 19809
rect 11521 19783 11527 19809
rect 12553 19783 12559 19809
rect 12585 19783 12591 19809
rect 12721 19783 12727 19809
rect 12753 19783 12759 19809
rect 12945 19783 12951 19809
rect 12977 19783 12983 19809
rect 15073 19783 15079 19809
rect 15105 19783 15111 19809
rect 15241 19783 15247 19809
rect 15273 19783 15279 19809
rect 15465 19783 15471 19809
rect 15497 19783 15503 19809
rect 18103 19777 18129 19783
rect 18271 19809 18297 19815
rect 18271 19777 18297 19783
rect 18383 19753 18409 19759
rect 2417 19727 2423 19753
rect 2449 19727 2455 19753
rect 6393 19727 6399 19753
rect 6425 19727 6431 19753
rect 18383 19721 18409 19727
rect 18775 19753 18801 19759
rect 18775 19721 18801 19727
rect 18943 19753 18969 19759
rect 18943 19721 18969 19727
rect 19055 19753 19081 19759
rect 19055 19721 19081 19727
rect 672 19613 19320 19630
rect 672 19587 9919 19613
rect 9945 19587 9971 19613
rect 9997 19587 10023 19613
rect 10049 19587 19320 19613
rect 672 19570 19320 19587
rect 18775 19473 18801 19479
rect 4433 19447 4439 19473
rect 4465 19447 4471 19473
rect 6393 19447 6399 19473
rect 6425 19447 6431 19473
rect 11489 19447 11495 19473
rect 11521 19447 11527 19473
rect 15465 19447 15471 19473
rect 15497 19447 15503 19473
rect 18775 19441 18801 19447
rect 18943 19417 18969 19423
rect 1857 19391 1863 19417
rect 1889 19391 1895 19417
rect 2417 19391 2423 19417
rect 2449 19391 2455 19417
rect 2529 19391 2535 19417
rect 2561 19391 2567 19417
rect 3369 19391 3375 19417
rect 3401 19391 3407 19417
rect 4433 19391 4439 19417
rect 4465 19391 4471 19417
rect 5273 19391 5279 19417
rect 5305 19391 5311 19417
rect 6393 19391 6399 19417
rect 6425 19391 6431 19417
rect 6953 19391 6959 19417
rect 6985 19391 6991 19417
rect 7233 19391 7239 19417
rect 7265 19391 7271 19417
rect 7345 19391 7351 19417
rect 7377 19391 7383 19417
rect 9137 19391 9143 19417
rect 9169 19391 9175 19417
rect 9305 19391 9311 19417
rect 9337 19391 9343 19417
rect 9529 19391 9535 19417
rect 9561 19391 9567 19417
rect 10593 19391 10599 19417
rect 10625 19391 10631 19417
rect 11489 19391 11495 19417
rect 11521 19391 11527 19417
rect 13113 19391 13119 19417
rect 13145 19391 13151 19417
rect 13393 19391 13399 19417
rect 13425 19391 13431 19417
rect 13561 19391 13567 19417
rect 13593 19391 13599 19417
rect 14569 19391 14575 19417
rect 14601 19391 14607 19417
rect 15465 19391 15471 19417
rect 15497 19391 15503 19417
rect 18943 19385 18969 19391
rect 19055 19417 19081 19423
rect 19055 19385 19081 19391
rect 672 19221 19320 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 19320 19221
rect 672 19178 19320 19195
rect 1577 18999 1583 19025
rect 1609 18999 1615 19025
rect 2473 18999 2479 19025
rect 2505 18999 2511 19025
rect 3817 18999 3823 19025
rect 3849 18999 3855 19025
rect 4377 18999 4383 19025
rect 4409 18999 4415 19025
rect 4489 18999 4495 19025
rect 4521 18999 4527 19025
rect 5273 18999 5279 19025
rect 5305 18999 5311 19025
rect 6393 18999 6399 19025
rect 6425 18999 6431 19025
rect 7121 18999 7127 19025
rect 7153 18999 7159 19025
rect 7345 18999 7351 19025
rect 7377 18999 7383 19025
rect 7569 18999 7575 19025
rect 7601 18999 7607 19025
rect 8409 18999 8415 19025
rect 8441 18999 8447 19025
rect 8745 18999 8751 19025
rect 8777 18999 8783 19025
rect 8969 18999 8975 19025
rect 9001 18999 9007 19025
rect 11097 18999 11103 19025
rect 11129 18999 11135 19025
rect 11377 18999 11383 19025
rect 11409 18999 11415 19025
rect 11489 18999 11495 19025
rect 11521 18999 11527 19025
rect 12553 18999 12559 19025
rect 12585 18999 12591 19025
rect 13393 18999 13399 19025
rect 13425 18999 13431 19025
rect 14849 18999 14855 19025
rect 14881 18999 14887 19025
rect 15913 18999 15919 19025
rect 15945 18999 15951 19025
rect 16249 18999 16255 19025
rect 16281 18999 16287 19025
rect 16809 18999 16815 19025
rect 16841 18999 16847 19025
rect 16921 18999 16927 19025
rect 16953 18999 16959 19025
rect 2473 18943 2479 18969
rect 2505 18943 2511 18969
rect 6393 18943 6399 18969
rect 6425 18943 6431 18969
rect 13393 18943 13399 18969
rect 13425 18943 13431 18969
rect 15913 18943 15919 18969
rect 15945 18943 15951 18969
rect 672 18829 19320 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 19320 18829
rect 672 18786 19320 18803
rect 3033 18663 3039 18689
rect 3065 18663 3071 18689
rect 4433 18663 4439 18689
rect 4465 18663 4471 18689
rect 6393 18663 6399 18689
rect 6425 18663 6431 18689
rect 11489 18663 11495 18689
rect 11521 18663 11527 18689
rect 15241 18663 15247 18689
rect 15273 18663 15279 18689
rect 17985 18663 17991 18689
rect 18017 18663 18023 18689
rect 1857 18607 1863 18633
rect 1889 18607 1895 18633
rect 3033 18607 3039 18633
rect 3065 18607 3071 18633
rect 3369 18607 3375 18633
rect 3401 18607 3407 18633
rect 4433 18607 4439 18633
rect 4465 18607 4471 18633
rect 5273 18607 5279 18633
rect 5305 18607 5311 18633
rect 6393 18607 6399 18633
rect 6425 18607 6431 18633
rect 6953 18607 6959 18633
rect 6985 18607 6991 18633
rect 7233 18607 7239 18633
rect 7265 18607 7271 18633
rect 7345 18607 7351 18633
rect 7377 18607 7383 18633
rect 8857 18607 8863 18633
rect 8889 18607 8895 18633
rect 9305 18607 9311 18633
rect 9337 18607 9343 18633
rect 9529 18607 9535 18633
rect 9561 18607 9567 18633
rect 10593 18607 10599 18633
rect 10625 18607 10631 18633
rect 11489 18607 11495 18633
rect 11521 18607 11527 18633
rect 13113 18607 13119 18633
rect 13145 18607 13151 18633
rect 13393 18607 13399 18633
rect 13425 18607 13431 18633
rect 13505 18607 13511 18633
rect 13537 18607 13543 18633
rect 14569 18607 14575 18633
rect 14601 18607 14607 18633
rect 15241 18607 15247 18633
rect 15273 18607 15279 18633
rect 17985 18607 17991 18633
rect 18017 18607 18023 18633
rect 18769 18607 18775 18633
rect 18801 18607 18807 18633
rect 672 18437 19320 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 19320 18437
rect 672 18394 19320 18411
rect 1577 18215 1583 18241
rect 1609 18215 1615 18241
rect 2473 18215 2479 18241
rect 2505 18215 2511 18241
rect 3817 18215 3823 18241
rect 3849 18215 3855 18241
rect 4377 18215 4383 18241
rect 4409 18215 4415 18241
rect 4489 18215 4495 18241
rect 4521 18215 4527 18241
rect 5273 18215 5279 18241
rect 5305 18215 5311 18241
rect 6393 18215 6399 18241
rect 6425 18215 6431 18241
rect 7121 18215 7127 18241
rect 7153 18215 7159 18241
rect 7345 18215 7351 18241
rect 7377 18215 7383 18241
rect 7569 18215 7575 18241
rect 7601 18215 7607 18241
rect 8409 18215 8415 18241
rect 8441 18215 8447 18241
rect 8745 18215 8751 18241
rect 8777 18215 8783 18241
rect 8969 18215 8975 18241
rect 9001 18215 9007 18241
rect 11097 18215 11103 18241
rect 11129 18215 11135 18241
rect 11377 18215 11383 18241
rect 11409 18215 11415 18241
rect 11489 18215 11495 18241
rect 11521 18215 11527 18241
rect 12553 18215 12559 18241
rect 12585 18215 12591 18241
rect 13393 18215 13399 18241
rect 13425 18215 13431 18241
rect 14849 18215 14855 18241
rect 14881 18215 14887 18241
rect 15913 18215 15919 18241
rect 15945 18215 15951 18241
rect 16249 18215 16255 18241
rect 16281 18215 16287 18241
rect 16753 18215 16759 18241
rect 16785 18215 16791 18241
rect 16921 18215 16927 18241
rect 16953 18215 16959 18241
rect 2473 18159 2479 18185
rect 2505 18159 2511 18185
rect 6393 18159 6399 18185
rect 6425 18159 6431 18185
rect 13393 18159 13399 18185
rect 13425 18159 13431 18185
rect 15913 18159 15919 18185
rect 15945 18159 15951 18185
rect 672 18045 19320 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 19320 18045
rect 672 18002 19320 18019
rect 3033 17879 3039 17905
rect 3065 17879 3071 17905
rect 4433 17879 4439 17905
rect 4465 17879 4471 17905
rect 6393 17879 6399 17905
rect 6425 17879 6431 17905
rect 11489 17879 11495 17905
rect 11521 17879 11527 17905
rect 15241 17879 15247 17905
rect 15273 17879 15279 17905
rect 1857 17823 1863 17849
rect 1889 17823 1895 17849
rect 3033 17823 3039 17849
rect 3065 17823 3071 17849
rect 3369 17823 3375 17849
rect 3401 17823 3407 17849
rect 4433 17823 4439 17849
rect 4465 17823 4471 17849
rect 5273 17823 5279 17849
rect 5305 17823 5311 17849
rect 6393 17823 6399 17849
rect 6425 17823 6431 17849
rect 6953 17823 6959 17849
rect 6985 17823 6991 17849
rect 7177 17823 7183 17849
rect 7209 17823 7215 17849
rect 7345 17823 7351 17849
rect 7377 17823 7383 17849
rect 8857 17823 8863 17849
rect 8889 17823 8895 17849
rect 9305 17823 9311 17849
rect 9337 17823 9343 17849
rect 9529 17823 9535 17849
rect 9561 17823 9567 17849
rect 10593 17823 10599 17849
rect 10625 17823 10631 17849
rect 11489 17823 11495 17849
rect 11521 17823 11527 17849
rect 13113 17823 13119 17849
rect 13145 17823 13151 17849
rect 13393 17823 13399 17849
rect 13425 17823 13431 17849
rect 13505 17823 13511 17849
rect 13537 17823 13543 17849
rect 14569 17823 14575 17849
rect 14601 17823 14607 17849
rect 15241 17823 15247 17849
rect 15273 17823 15279 17849
rect 16809 17823 16815 17849
rect 16841 17823 16847 17849
rect 17257 17823 17263 17849
rect 17289 17823 17295 17849
rect 17481 17823 17487 17849
rect 17513 17823 17519 17849
rect 672 17653 19320 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 19320 17653
rect 672 17610 19320 17627
rect 1577 17431 1583 17457
rect 1609 17431 1615 17457
rect 2417 17431 2423 17457
rect 2449 17431 2455 17457
rect 3873 17431 3879 17457
rect 3905 17431 3911 17457
rect 4377 17431 4383 17457
rect 4409 17431 4415 17457
rect 4489 17431 4495 17457
rect 4521 17431 4527 17457
rect 5273 17431 5279 17457
rect 5305 17431 5311 17457
rect 6393 17431 6399 17457
rect 6425 17431 6431 17457
rect 7121 17431 7127 17457
rect 7153 17431 7159 17457
rect 7793 17431 7799 17457
rect 7825 17431 7831 17457
rect 8409 17431 8415 17457
rect 8441 17431 8447 17457
rect 9305 17431 9311 17457
rect 9337 17431 9343 17457
rect 11097 17431 11103 17457
rect 11129 17431 11135 17457
rect 11377 17431 11383 17457
rect 11409 17431 11415 17457
rect 11489 17431 11495 17457
rect 11521 17431 11527 17457
rect 12553 17431 12559 17457
rect 12585 17431 12591 17457
rect 13393 17431 13399 17457
rect 13425 17431 13431 17457
rect 14793 17431 14799 17457
rect 14825 17431 14831 17457
rect 15241 17431 15247 17457
rect 15273 17431 15279 17457
rect 15465 17431 15471 17457
rect 15497 17431 15503 17457
rect 16249 17431 16255 17457
rect 16281 17431 16287 17457
rect 17257 17431 17263 17457
rect 17289 17431 17295 17457
rect 2417 17375 2423 17401
rect 2449 17375 2455 17401
rect 6393 17375 6399 17401
rect 6425 17375 6431 17401
rect 7793 17375 7799 17401
rect 7825 17375 7831 17401
rect 9305 17375 9311 17401
rect 9337 17375 9343 17401
rect 13393 17375 13399 17401
rect 13425 17375 13431 17401
rect 17257 17375 17263 17401
rect 17289 17375 17295 17401
rect 672 17261 19320 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 19320 17261
rect 672 17218 19320 17235
rect 4433 17095 4439 17121
rect 4465 17095 4471 17121
rect 6393 17095 6399 17121
rect 6425 17095 6431 17121
rect 7793 17095 7799 17121
rect 7825 17095 7831 17121
rect 11265 17095 11271 17121
rect 11297 17095 11303 17121
rect 15241 17095 15247 17121
rect 15273 17095 15279 17121
rect 18775 17065 18801 17071
rect 1857 17039 1863 17065
rect 1889 17039 1895 17065
rect 2417 17039 2423 17065
rect 2449 17039 2455 17065
rect 2585 17039 2591 17065
rect 2617 17039 2623 17065
rect 3425 17039 3431 17065
rect 3457 17039 3463 17065
rect 4433 17039 4439 17065
rect 4465 17039 4471 17065
rect 5273 17039 5279 17065
rect 5305 17039 5311 17065
rect 6393 17039 6399 17065
rect 6425 17039 6431 17065
rect 6953 17039 6959 17065
rect 6985 17039 6991 17065
rect 7793 17039 7799 17065
rect 7825 17039 7831 17065
rect 8857 17039 8863 17065
rect 8889 17039 8895 17065
rect 9305 17039 9311 17065
rect 9337 17039 9343 17065
rect 9529 17039 9535 17065
rect 9561 17039 9567 17065
rect 10593 17039 10599 17065
rect 10625 17039 10631 17065
rect 11265 17039 11271 17065
rect 11297 17039 11303 17065
rect 13113 17039 13119 17065
rect 13145 17039 13151 17065
rect 13393 17039 13399 17065
rect 13425 17039 13431 17065
rect 13505 17039 13511 17065
rect 13537 17039 13543 17065
rect 14569 17039 14575 17065
rect 14601 17039 14607 17065
rect 15241 17039 15247 17065
rect 15273 17039 15279 17065
rect 16809 17039 16815 17065
rect 16841 17039 16847 17065
rect 17257 17039 17263 17065
rect 17289 17039 17295 17065
rect 17481 17039 17487 17065
rect 17513 17039 17519 17065
rect 18775 17033 18801 17039
rect 18887 17065 18913 17071
rect 18887 17033 18913 17039
rect 19055 17065 19081 17071
rect 19055 17033 19081 17039
rect 672 16869 19320 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 19320 16869
rect 672 16826 19320 16843
rect 18775 16673 18801 16679
rect 1577 16647 1583 16673
rect 1609 16647 1615 16673
rect 2305 16647 2311 16673
rect 2337 16647 2343 16673
rect 3873 16647 3879 16673
rect 3905 16647 3911 16673
rect 4377 16647 4383 16673
rect 4409 16647 4415 16673
rect 4489 16647 4495 16673
rect 4521 16647 4527 16673
rect 5273 16647 5279 16673
rect 5305 16647 5311 16673
rect 6393 16647 6399 16673
rect 6425 16647 6431 16673
rect 7121 16647 7127 16673
rect 7153 16647 7159 16673
rect 7793 16647 7799 16673
rect 7825 16647 7831 16673
rect 8409 16647 8415 16673
rect 8441 16647 8447 16673
rect 9305 16647 9311 16673
rect 9337 16647 9343 16673
rect 10817 16647 10823 16673
rect 10849 16647 10855 16673
rect 11265 16647 11271 16673
rect 11297 16647 11303 16673
rect 11489 16647 11495 16673
rect 11521 16647 11527 16673
rect 12553 16647 12559 16673
rect 12585 16647 12591 16673
rect 13393 16647 13399 16673
rect 13425 16647 13431 16673
rect 14793 16647 14799 16673
rect 14825 16647 14831 16673
rect 15241 16647 15247 16673
rect 15273 16647 15279 16673
rect 15465 16647 15471 16673
rect 15497 16647 15503 16673
rect 16249 16647 16255 16673
rect 16281 16647 16287 16673
rect 17257 16647 17263 16673
rect 17289 16647 17295 16673
rect 18775 16641 18801 16647
rect 18887 16673 18913 16679
rect 18887 16641 18913 16647
rect 19055 16617 19081 16623
rect 2305 16591 2311 16617
rect 2337 16591 2343 16617
rect 6393 16591 6399 16617
rect 6425 16591 6431 16617
rect 7793 16591 7799 16617
rect 7825 16591 7831 16617
rect 9305 16591 9311 16617
rect 9337 16591 9343 16617
rect 13393 16591 13399 16617
rect 13425 16591 13431 16617
rect 17257 16591 17263 16617
rect 17289 16591 17295 16617
rect 19055 16585 19081 16591
rect 672 16477 19320 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 19320 16477
rect 672 16434 19320 16451
rect 4433 16311 4439 16337
rect 4465 16311 4471 16337
rect 6393 16311 6399 16337
rect 6425 16311 6431 16337
rect 7793 16311 7799 16337
rect 7825 16311 7831 16337
rect 11265 16311 11271 16337
rect 11297 16311 11303 16337
rect 15241 16311 15247 16337
rect 15273 16311 15279 16337
rect 1857 16255 1863 16281
rect 1889 16255 1895 16281
rect 2305 16255 2311 16281
rect 2337 16255 2343 16281
rect 2529 16255 2535 16281
rect 2561 16255 2567 16281
rect 3425 16255 3431 16281
rect 3457 16255 3463 16281
rect 4433 16255 4439 16281
rect 4465 16255 4471 16281
rect 5273 16255 5279 16281
rect 5305 16255 5311 16281
rect 6393 16255 6399 16281
rect 6425 16255 6431 16281
rect 6953 16255 6959 16281
rect 6985 16255 6991 16281
rect 7793 16255 7799 16281
rect 7825 16255 7831 16281
rect 8857 16255 8863 16281
rect 8889 16255 8895 16281
rect 9305 16255 9311 16281
rect 9337 16255 9343 16281
rect 9529 16255 9535 16281
rect 9561 16255 9567 16281
rect 10593 16255 10599 16281
rect 10625 16255 10631 16281
rect 11265 16255 11271 16281
rect 11297 16255 11303 16281
rect 13113 16255 13119 16281
rect 13145 16255 13151 16281
rect 13393 16255 13399 16281
rect 13425 16255 13431 16281
rect 13505 16255 13511 16281
rect 13537 16255 13543 16281
rect 14289 16255 14295 16281
rect 14321 16255 14327 16281
rect 15241 16255 15247 16281
rect 15273 16255 15279 16281
rect 16809 16255 16815 16281
rect 16841 16255 16847 16281
rect 17257 16255 17263 16281
rect 17289 16255 17295 16281
rect 17481 16255 17487 16281
rect 17513 16255 17519 16281
rect 672 16085 19320 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 19320 16085
rect 672 16042 19320 16059
rect 1353 15863 1359 15889
rect 1385 15863 1391 15889
rect 2473 15863 2479 15889
rect 2505 15863 2511 15889
rect 4041 15863 4047 15889
rect 4073 15863 4079 15889
rect 4265 15863 4271 15889
rect 4297 15863 4303 15889
rect 4489 15863 4495 15889
rect 4521 15863 4527 15889
rect 5273 15863 5279 15889
rect 5305 15863 5311 15889
rect 6169 15863 6175 15889
rect 6201 15863 6207 15889
rect 7121 15863 7127 15889
rect 7153 15863 7159 15889
rect 7625 15863 7631 15889
rect 7657 15863 7663 15889
rect 8409 15863 8415 15889
rect 8441 15863 8447 15889
rect 8801 15863 8807 15889
rect 8833 15863 8839 15889
rect 8969 15863 8975 15889
rect 9001 15863 9007 15889
rect 10817 15863 10823 15889
rect 10849 15863 10855 15889
rect 11489 15863 11495 15889
rect 11521 15863 11527 15889
rect 12273 15863 12279 15889
rect 12305 15863 12311 15889
rect 12721 15863 12727 15889
rect 12753 15863 12759 15889
rect 12945 15863 12951 15889
rect 12977 15863 12983 15889
rect 14793 15863 14799 15889
rect 14825 15863 14831 15889
rect 15241 15863 15247 15889
rect 15273 15863 15279 15889
rect 15465 15863 15471 15889
rect 15497 15863 15503 15889
rect 16249 15863 16255 15889
rect 16281 15863 16287 15889
rect 16809 15863 16815 15889
rect 16841 15863 16847 15889
rect 16921 15863 16927 15889
rect 16953 15863 16959 15889
rect 2473 15807 2479 15833
rect 2505 15807 2511 15833
rect 6225 15807 6231 15833
rect 6257 15807 6263 15833
rect 7793 15807 7799 15833
rect 7825 15807 7831 15833
rect 11769 15807 11775 15833
rect 11801 15807 11807 15833
rect 672 15693 19320 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 19320 15693
rect 672 15650 19320 15667
rect 4489 15527 4495 15553
rect 4521 15527 4527 15553
rect 6169 15527 6175 15553
rect 6201 15527 6207 15553
rect 7625 15527 7631 15553
rect 7657 15527 7663 15553
rect 11433 15527 11439 15553
rect 11465 15527 11471 15553
rect 15297 15527 15303 15553
rect 15329 15527 15335 15553
rect 1857 15471 1863 15497
rect 1889 15471 1895 15497
rect 2417 15471 2423 15497
rect 2449 15471 2455 15497
rect 2529 15471 2535 15497
rect 2561 15471 2567 15497
rect 3593 15471 3599 15497
rect 3625 15471 3631 15497
rect 4489 15471 4495 15497
rect 4521 15471 4527 15497
rect 5273 15471 5279 15497
rect 5305 15471 5311 15497
rect 6169 15471 6175 15497
rect 6201 15471 6207 15497
rect 6953 15471 6959 15497
rect 6985 15471 6991 15497
rect 7625 15471 7631 15497
rect 7657 15471 7663 15497
rect 8857 15471 8863 15497
rect 8889 15471 8895 15497
rect 9305 15471 9311 15497
rect 9337 15471 9343 15497
rect 9529 15471 9535 15497
rect 9561 15471 9567 15497
rect 10369 15471 10375 15497
rect 10401 15471 10407 15497
rect 11433 15471 11439 15497
rect 11465 15471 11471 15497
rect 12833 15471 12839 15497
rect 12865 15471 12871 15497
rect 13393 15471 13399 15497
rect 13425 15471 13431 15497
rect 13505 15471 13511 15497
rect 13537 15471 13543 15497
rect 14289 15471 14295 15497
rect 14321 15471 14327 15497
rect 15185 15471 15191 15497
rect 15217 15471 15223 15497
rect 16809 15471 16815 15497
rect 16841 15471 16847 15497
rect 17257 15471 17263 15497
rect 17289 15471 17295 15497
rect 17481 15471 17487 15497
rect 17513 15471 17519 15497
rect 672 15301 19320 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 19320 15301
rect 672 15258 19320 15275
rect 1353 15079 1359 15105
rect 1385 15079 1391 15105
rect 2473 15079 2479 15105
rect 2505 15079 2511 15105
rect 4041 15079 4047 15105
rect 4073 15079 4079 15105
rect 4377 15079 4383 15105
rect 4409 15079 4415 15105
rect 4489 15079 4495 15105
rect 4521 15079 4527 15105
rect 5273 15079 5279 15105
rect 5305 15079 5311 15105
rect 6169 15079 6175 15105
rect 6201 15079 6207 15105
rect 6953 15079 6959 15105
rect 6985 15079 6991 15105
rect 7625 15079 7631 15105
rect 7657 15079 7663 15105
rect 8409 15079 8415 15105
rect 8441 15079 8447 15105
rect 8801 15079 8807 15105
rect 8833 15079 8839 15105
rect 8969 15079 8975 15105
rect 9001 15079 9007 15105
rect 10817 15079 10823 15105
rect 10849 15079 10855 15105
rect 11489 15079 11495 15105
rect 11521 15079 11527 15105
rect 12273 15079 12279 15105
rect 12305 15079 12311 15105
rect 13337 15079 13343 15105
rect 13369 15079 13375 15105
rect 14793 15079 14799 15105
rect 14825 15079 14831 15105
rect 15241 15079 15247 15105
rect 15273 15079 15279 15105
rect 15465 15079 15471 15105
rect 15497 15079 15503 15105
rect 16529 15079 16535 15105
rect 16561 15079 16567 15105
rect 17257 15079 17263 15105
rect 17289 15079 17295 15105
rect 2473 15023 2479 15049
rect 2505 15023 2511 15049
rect 6225 15023 6231 15049
rect 6257 15023 6263 15049
rect 7793 15023 7799 15049
rect 7825 15023 7831 15049
rect 11769 15023 11775 15049
rect 11801 15023 11807 15049
rect 13337 15023 13343 15049
rect 13369 15023 13375 15049
rect 17257 15023 17263 15049
rect 17289 15023 17295 15049
rect 672 14909 19320 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 19320 14909
rect 672 14866 19320 14883
rect 4489 14743 4495 14769
rect 4521 14743 4527 14769
rect 6169 14743 6175 14769
rect 6201 14743 6207 14769
rect 7625 14743 7631 14769
rect 7657 14743 7663 14769
rect 11433 14743 11439 14769
rect 11465 14743 11471 14769
rect 15241 14743 15247 14769
rect 15273 14743 15279 14769
rect 1857 14687 1863 14713
rect 1889 14687 1895 14713
rect 2417 14687 2423 14713
rect 2449 14687 2455 14713
rect 2529 14687 2535 14713
rect 2561 14687 2567 14713
rect 3593 14687 3599 14713
rect 3625 14687 3631 14713
rect 4489 14687 4495 14713
rect 4521 14687 4527 14713
rect 5217 14687 5223 14713
rect 5249 14687 5255 14713
rect 5945 14687 5951 14713
rect 5977 14687 5983 14713
rect 6953 14687 6959 14713
rect 6985 14687 6991 14713
rect 7625 14687 7631 14713
rect 7657 14687 7663 14713
rect 8857 14687 8863 14713
rect 8889 14687 8895 14713
rect 9305 14687 9311 14713
rect 9337 14687 9343 14713
rect 9529 14687 9535 14713
rect 9561 14687 9567 14713
rect 10369 14687 10375 14713
rect 10401 14687 10407 14713
rect 11433 14687 11439 14713
rect 11465 14687 11471 14713
rect 12833 14687 12839 14713
rect 12865 14687 12871 14713
rect 13393 14687 13399 14713
rect 13425 14687 13431 14713
rect 13505 14687 13511 14713
rect 13537 14687 13543 14713
rect 14289 14687 14295 14713
rect 14321 14687 14327 14713
rect 15241 14687 15247 14713
rect 15273 14687 15279 14713
rect 16809 14687 16815 14713
rect 16841 14687 16847 14713
rect 17257 14687 17263 14713
rect 17289 14687 17295 14713
rect 17481 14687 17487 14713
rect 17513 14687 17519 14713
rect 672 14517 19320 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 19320 14517
rect 672 14474 19320 14491
rect 1353 14295 1359 14321
rect 1385 14295 1391 14321
rect 2473 14295 2479 14321
rect 2505 14295 2511 14321
rect 4041 14295 4047 14321
rect 4073 14295 4079 14321
rect 4377 14295 4383 14321
rect 4409 14295 4415 14321
rect 4489 14295 4495 14321
rect 4521 14295 4527 14321
rect 5273 14295 5279 14321
rect 5305 14295 5311 14321
rect 5833 14295 5839 14321
rect 5865 14295 5871 14321
rect 5945 14295 5951 14321
rect 5977 14295 5983 14321
rect 6953 14295 6959 14321
rect 6985 14295 6991 14321
rect 7625 14295 7631 14321
rect 7657 14295 7663 14321
rect 8409 14295 8415 14321
rect 8441 14295 8447 14321
rect 8801 14295 8807 14321
rect 8833 14295 8839 14321
rect 8969 14295 8975 14321
rect 9001 14295 9007 14321
rect 10817 14295 10823 14321
rect 10849 14295 10855 14321
rect 11489 14295 11495 14321
rect 11521 14295 11527 14321
rect 12273 14295 12279 14321
rect 12305 14295 12311 14321
rect 13393 14295 13399 14321
rect 13425 14295 13431 14321
rect 14793 14295 14799 14321
rect 14825 14295 14831 14321
rect 15241 14295 15247 14321
rect 15273 14295 15279 14321
rect 15465 14295 15471 14321
rect 15497 14295 15503 14321
rect 16529 14295 16535 14321
rect 16561 14295 16567 14321
rect 17257 14295 17263 14321
rect 17289 14295 17295 14321
rect 2473 14239 2479 14265
rect 2505 14239 2511 14265
rect 7793 14239 7799 14265
rect 7825 14239 7831 14265
rect 11769 14239 11775 14265
rect 11801 14239 11807 14265
rect 13393 14239 13399 14265
rect 13425 14239 13431 14265
rect 17257 14239 17263 14265
rect 17289 14239 17295 14265
rect 672 14125 19320 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 19320 14125
rect 672 14082 19320 14099
rect 4489 13959 4495 13985
rect 4521 13959 4527 13985
rect 7625 13959 7631 13985
rect 7657 13959 7663 13985
rect 11489 13959 11495 13985
rect 11521 13959 11527 13985
rect 15241 13959 15247 13985
rect 15273 13959 15279 13985
rect 1857 13903 1863 13929
rect 1889 13903 1895 13929
rect 2417 13903 2423 13929
rect 2449 13903 2455 13929
rect 2585 13903 2591 13929
rect 2617 13903 2623 13929
rect 3593 13903 3599 13929
rect 3625 13903 3631 13929
rect 4489 13903 4495 13929
rect 4521 13903 4527 13929
rect 5217 13903 5223 13929
rect 5249 13903 5255 13929
rect 5777 13903 5783 13929
rect 5809 13903 5815 13929
rect 5889 13903 5895 13929
rect 5921 13903 5927 13929
rect 6953 13903 6959 13929
rect 6985 13903 6991 13929
rect 7625 13903 7631 13929
rect 7657 13903 7663 13929
rect 8857 13903 8863 13929
rect 8889 13903 8895 13929
rect 9305 13903 9311 13929
rect 9337 13903 9343 13929
rect 9529 13903 9535 13929
rect 9561 13903 9567 13929
rect 10369 13903 10375 13929
rect 10401 13903 10407 13929
rect 11489 13903 11495 13929
rect 11521 13903 11527 13929
rect 12833 13903 12839 13929
rect 12865 13903 12871 13929
rect 13393 13903 13399 13929
rect 13425 13903 13431 13929
rect 13505 13903 13511 13929
rect 13537 13903 13543 13929
rect 14289 13903 14295 13929
rect 14321 13903 14327 13929
rect 15241 13903 15247 13929
rect 15273 13903 15279 13929
rect 16809 13903 16815 13929
rect 16841 13903 16847 13929
rect 17257 13903 17263 13929
rect 17289 13903 17295 13929
rect 17481 13903 17487 13929
rect 17513 13903 17519 13929
rect 672 13733 19320 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 19320 13733
rect 672 13690 19320 13707
rect 1353 13511 1359 13537
rect 1385 13511 1391 13537
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 4041 13511 4047 13537
rect 4073 13511 4079 13537
rect 4377 13511 4383 13537
rect 4409 13511 4415 13537
rect 4489 13511 4495 13537
rect 4521 13511 4527 13537
rect 5273 13511 5279 13537
rect 5305 13511 5311 13537
rect 5833 13511 5839 13537
rect 5865 13511 5871 13537
rect 5945 13511 5951 13537
rect 5977 13511 5983 13537
rect 6953 13511 6959 13537
rect 6985 13511 6991 13537
rect 7625 13511 7631 13537
rect 7657 13511 7663 13537
rect 8409 13511 8415 13537
rect 8441 13511 8447 13537
rect 8801 13511 8807 13537
rect 8833 13511 8839 13537
rect 8969 13511 8975 13537
rect 9001 13511 9007 13537
rect 10817 13511 10823 13537
rect 10849 13511 10855 13537
rect 11713 13511 11719 13537
rect 11745 13511 11751 13537
rect 12273 13511 12279 13537
rect 12305 13511 12311 13537
rect 13449 13511 13455 13537
rect 13481 13511 13487 13537
rect 14793 13511 14799 13537
rect 14825 13511 14831 13537
rect 15241 13511 15247 13537
rect 15273 13511 15279 13537
rect 15465 13511 15471 13537
rect 15497 13511 15503 13537
rect 16529 13511 16535 13537
rect 16561 13511 16567 13537
rect 16809 13511 16815 13537
rect 16841 13511 16847 13537
rect 16921 13511 16927 13537
rect 16953 13511 16959 13537
rect 2249 13455 2255 13481
rect 2281 13455 2287 13481
rect 7793 13455 7799 13481
rect 7825 13455 7831 13481
rect 11769 13455 11775 13481
rect 11801 13455 11807 13481
rect 13449 13455 13455 13481
rect 13481 13455 13487 13481
rect 672 13341 19320 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 19320 13341
rect 672 13298 19320 13315
rect 4489 13175 4495 13201
rect 4521 13175 4527 13201
rect 7625 13175 7631 13201
rect 7657 13175 7663 13201
rect 11489 13175 11495 13201
rect 11521 13175 11527 13201
rect 15241 13175 15247 13201
rect 15273 13175 15279 13201
rect 17873 13175 17879 13201
rect 17905 13175 17911 13201
rect 1857 13119 1863 13145
rect 1889 13119 1895 13145
rect 2305 13119 2311 13145
rect 2337 13119 2343 13145
rect 2529 13119 2535 13145
rect 2561 13119 2567 13145
rect 3593 13119 3599 13145
rect 3625 13119 3631 13145
rect 4489 13119 4495 13145
rect 4521 13119 4527 13145
rect 5217 13119 5223 13145
rect 5249 13119 5255 13145
rect 5777 13119 5783 13145
rect 5809 13119 5815 13145
rect 5889 13119 5895 13145
rect 5921 13119 5927 13145
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 7625 13119 7631 13145
rect 7657 13119 7663 13145
rect 8857 13119 8863 13145
rect 8889 13119 8895 13145
rect 9305 13119 9311 13145
rect 9337 13119 9343 13145
rect 9529 13119 9535 13145
rect 9561 13119 9567 13145
rect 10369 13119 10375 13145
rect 10401 13119 10407 13145
rect 11489 13119 11495 13145
rect 11521 13119 11527 13145
rect 12833 13119 12839 13145
rect 12865 13119 12871 13145
rect 13393 13119 13399 13145
rect 13425 13119 13431 13145
rect 13505 13119 13511 13145
rect 13537 13119 13543 13145
rect 14289 13119 14295 13145
rect 14321 13119 14327 13145
rect 15241 13119 15247 13145
rect 15273 13119 15279 13145
rect 17873 13119 17879 13145
rect 17905 13119 17911 13145
rect 19049 13119 19055 13145
rect 19081 13119 19087 13145
rect 672 12949 19320 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 19320 12949
rect 672 12906 19320 12923
rect 1353 12727 1359 12753
rect 1385 12727 1391 12753
rect 2473 12727 2479 12753
rect 2505 12727 2511 12753
rect 4041 12727 4047 12753
rect 4073 12727 4079 12753
rect 4377 12727 4383 12753
rect 4409 12727 4415 12753
rect 4489 12727 4495 12753
rect 4521 12727 4527 12753
rect 5273 12727 5279 12753
rect 5305 12727 5311 12753
rect 5833 12727 5839 12753
rect 5865 12727 5871 12753
rect 5945 12727 5951 12753
rect 5977 12727 5983 12753
rect 6953 12727 6959 12753
rect 6985 12727 6991 12753
rect 7625 12727 7631 12753
rect 7657 12727 7663 12753
rect 8409 12727 8415 12753
rect 8441 12727 8447 12753
rect 8801 12727 8807 12753
rect 8833 12727 8839 12753
rect 8969 12727 8975 12753
rect 9001 12727 9007 12753
rect 10929 12727 10935 12753
rect 10961 12727 10967 12753
rect 11713 12727 11719 12753
rect 11745 12727 11751 12753
rect 12273 12727 12279 12753
rect 12305 12727 12311 12753
rect 13449 12727 13455 12753
rect 13481 12727 13487 12753
rect 14793 12727 14799 12753
rect 14825 12727 14831 12753
rect 15241 12727 15247 12753
rect 15273 12727 15279 12753
rect 15465 12727 15471 12753
rect 15497 12727 15503 12753
rect 16249 12727 16255 12753
rect 16281 12727 16287 12753
rect 16809 12727 16815 12753
rect 16841 12727 16847 12753
rect 16921 12727 16927 12753
rect 16953 12727 16959 12753
rect 2473 12671 2479 12697
rect 2505 12671 2511 12697
rect 7793 12671 7799 12697
rect 7825 12671 7831 12697
rect 11769 12671 11775 12697
rect 11801 12671 11807 12697
rect 13449 12671 13455 12697
rect 13481 12671 13487 12697
rect 672 12557 19320 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 19320 12557
rect 672 12514 19320 12531
rect 6169 12391 6175 12417
rect 6201 12391 6207 12417
rect 7625 12391 7631 12417
rect 7657 12391 7663 12417
rect 11489 12391 11495 12417
rect 11521 12391 11527 12417
rect 15241 12391 15247 12417
rect 15273 12391 15279 12417
rect 17873 12391 17879 12417
rect 17905 12391 17911 12417
rect 1857 12335 1863 12361
rect 1889 12335 1895 12361
rect 2417 12335 2423 12361
rect 2449 12335 2455 12361
rect 2529 12335 2535 12361
rect 2561 12335 2567 12361
rect 3593 12335 3599 12361
rect 3625 12335 3631 12361
rect 3761 12335 3767 12361
rect 3793 12335 3799 12361
rect 3985 12335 3991 12361
rect 4017 12335 4023 12361
rect 5217 12335 5223 12361
rect 5249 12335 5255 12361
rect 5945 12335 5951 12361
rect 5977 12335 5983 12361
rect 6953 12335 6959 12361
rect 6985 12335 6991 12361
rect 7569 12335 7575 12361
rect 7601 12335 7607 12361
rect 8857 12335 8863 12361
rect 8889 12335 8895 12361
rect 9305 12335 9311 12361
rect 9337 12335 9343 12361
rect 9529 12335 9535 12361
rect 9561 12335 9567 12361
rect 10313 12335 10319 12361
rect 10345 12335 10351 12361
rect 11489 12335 11495 12361
rect 11521 12335 11527 12361
rect 12833 12335 12839 12361
rect 12865 12335 12871 12361
rect 13393 12335 13399 12361
rect 13425 12335 13431 12361
rect 13505 12335 13511 12361
rect 13537 12335 13543 12361
rect 14289 12335 14295 12361
rect 14321 12335 14327 12361
rect 15241 12335 15247 12361
rect 15273 12335 15279 12361
rect 17873 12335 17879 12361
rect 17905 12335 17911 12361
rect 19049 12335 19055 12361
rect 19081 12335 19087 12361
rect 672 12165 19320 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 19320 12165
rect 672 12122 19320 12139
rect 1353 11943 1359 11969
rect 1385 11943 1391 11969
rect 2473 11943 2479 11969
rect 2505 11943 2511 11969
rect 4097 11943 4103 11969
rect 4129 11943 4135 11969
rect 4769 11943 4775 11969
rect 4801 11943 4807 11969
rect 5273 11943 5279 11969
rect 5305 11943 5311 11969
rect 5833 11943 5839 11969
rect 5865 11943 5871 11969
rect 5945 11943 5951 11969
rect 5977 11943 5983 11969
rect 6953 11943 6959 11969
rect 6985 11943 6991 11969
rect 7569 11943 7575 11969
rect 7601 11943 7607 11969
rect 8409 11943 8415 11969
rect 8441 11943 8447 11969
rect 8745 11943 8751 11969
rect 8777 11943 8783 11969
rect 8969 11943 8975 11969
rect 9001 11943 9007 11969
rect 10929 11943 10935 11969
rect 10961 11943 10967 11969
rect 11377 11943 11383 11969
rect 11409 11943 11415 11969
rect 11489 11943 11495 11969
rect 11521 11943 11527 11969
rect 12273 11943 12279 11969
rect 12305 11943 12311 11969
rect 13393 11943 13399 11969
rect 13425 11943 13431 11969
rect 15073 11943 15079 11969
rect 15105 11943 15111 11969
rect 15241 11943 15247 11969
rect 15273 11943 15279 11969
rect 15465 11943 15471 11969
rect 15497 11943 15503 11969
rect 17481 11943 17487 11969
rect 17513 11943 17519 11969
rect 17761 11943 17767 11969
rect 17793 11943 17799 11969
rect 17873 11943 17879 11969
rect 17905 11943 17911 11969
rect 2473 11887 2479 11913
rect 2505 11887 2511 11913
rect 4769 11887 4775 11913
rect 4801 11887 4807 11913
rect 7793 11887 7799 11913
rect 7825 11887 7831 11913
rect 13393 11887 13399 11913
rect 13425 11887 13431 11913
rect 672 11773 19320 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 19320 11773
rect 672 11730 19320 11747
rect 6169 11607 6175 11633
rect 6201 11607 6207 11633
rect 7625 11607 7631 11633
rect 7657 11607 7663 11633
rect 11489 11607 11495 11633
rect 11521 11607 11527 11633
rect 15241 11607 15247 11633
rect 15273 11607 15279 11633
rect 17873 11607 17879 11633
rect 17905 11607 17911 11633
rect 1857 11551 1863 11577
rect 1889 11551 1895 11577
rect 2417 11551 2423 11577
rect 2449 11551 2455 11577
rect 2529 11551 2535 11577
rect 2561 11551 2567 11577
rect 3313 11551 3319 11577
rect 3345 11551 3351 11577
rect 3873 11551 3879 11577
rect 3905 11551 3911 11577
rect 3985 11551 3991 11577
rect 4017 11551 4023 11577
rect 5217 11551 5223 11577
rect 5249 11551 5255 11577
rect 5945 11551 5951 11577
rect 5977 11551 5983 11577
rect 6953 11551 6959 11577
rect 6985 11551 6991 11577
rect 7569 11551 7575 11577
rect 7601 11551 7607 11577
rect 9025 11551 9031 11577
rect 9057 11551 9063 11577
rect 9305 11551 9311 11577
rect 9337 11551 9343 11577
rect 9529 11551 9535 11577
rect 9561 11551 9567 11577
rect 10313 11551 10319 11577
rect 10345 11551 10351 11577
rect 11489 11551 11495 11577
rect 11521 11551 11527 11577
rect 12833 11551 12839 11577
rect 12865 11551 12871 11577
rect 13393 11551 13399 11577
rect 13425 11551 13431 11577
rect 13505 11551 13511 11577
rect 13537 11551 13543 11577
rect 14569 11551 14575 11577
rect 14601 11551 14607 11577
rect 15129 11551 15135 11577
rect 15161 11551 15167 11577
rect 17873 11551 17879 11577
rect 17905 11551 17911 11577
rect 19049 11551 19055 11577
rect 19081 11551 19087 11577
rect 672 11381 19320 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 19320 11381
rect 672 11338 19320 11355
rect 1409 11159 1415 11185
rect 1441 11159 1447 11185
rect 2473 11159 2479 11185
rect 2505 11159 2511 11185
rect 3313 11159 3319 11185
rect 3345 11159 3351 11185
rect 3985 11159 3991 11185
rect 4017 11159 4023 11185
rect 4657 11159 4663 11185
rect 4689 11159 4695 11185
rect 5049 11159 5055 11185
rect 5081 11159 5087 11185
rect 5273 11159 5279 11185
rect 5305 11159 5311 11185
rect 6953 11159 6959 11185
rect 6985 11159 6991 11185
rect 7569 11159 7575 11185
rect 7601 11159 7607 11185
rect 8409 11159 8415 11185
rect 8441 11159 8447 11185
rect 8745 11159 8751 11185
rect 8777 11159 8783 11185
rect 8969 11159 8975 11185
rect 9001 11159 9007 11185
rect 10817 11159 10823 11185
rect 10849 11159 10855 11185
rect 11377 11159 11383 11185
rect 11409 11159 11415 11185
rect 11489 11159 11495 11185
rect 11521 11159 11527 11185
rect 12273 11159 12279 11185
rect 12305 11159 12311 11185
rect 13449 11159 13455 11185
rect 13481 11159 13487 11185
rect 15969 11159 15975 11185
rect 16001 11159 16007 11185
rect 16921 11159 16927 11185
rect 16953 11159 16959 11185
rect 17481 11159 17487 11185
rect 17513 11159 17519 11185
rect 17761 11159 17767 11185
rect 17793 11159 17799 11185
rect 17873 11159 17879 11185
rect 17905 11159 17911 11185
rect 2473 11103 2479 11129
rect 2505 11103 2511 11129
rect 4097 11103 4103 11129
rect 4129 11103 4135 11129
rect 7793 11103 7799 11129
rect 7825 11103 7831 11129
rect 13449 11103 13455 11129
rect 13481 11103 13487 11129
rect 15969 11103 15975 11129
rect 16001 11103 16007 11129
rect 672 10989 19320 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 19320 10989
rect 672 10946 19320 10963
rect 5833 10823 5839 10849
rect 5865 10823 5871 10849
rect 7793 10823 7799 10849
rect 7825 10823 7831 10849
rect 9809 10823 9815 10849
rect 9841 10823 9847 10849
rect 11489 10823 11495 10849
rect 11521 10823 11527 10849
rect 15465 10823 15471 10849
rect 15497 10823 15503 10849
rect 17873 10823 17879 10849
rect 17905 10823 17911 10849
rect 1913 10767 1919 10793
rect 1945 10767 1951 10793
rect 2417 10767 2423 10793
rect 2449 10767 2455 10793
rect 2529 10767 2535 10793
rect 2561 10767 2567 10793
rect 3369 10767 3375 10793
rect 3401 10767 3407 10793
rect 3873 10767 3879 10793
rect 3905 10767 3911 10793
rect 3985 10767 3991 10793
rect 4017 10767 4023 10793
rect 4881 10767 4887 10793
rect 4913 10767 4919 10793
rect 5833 10767 5839 10793
rect 5865 10767 5871 10793
rect 6953 10767 6959 10793
rect 6985 10767 6991 10793
rect 7793 10767 7799 10793
rect 7825 10767 7831 10793
rect 9025 10767 9031 10793
rect 9057 10767 9063 10793
rect 9753 10767 9759 10793
rect 9785 10767 9791 10793
rect 10313 10767 10319 10793
rect 10345 10767 10351 10793
rect 11489 10767 11495 10793
rect 11521 10767 11527 10793
rect 12833 10767 12839 10793
rect 12865 10767 12871 10793
rect 13393 10767 13399 10793
rect 13425 10767 13431 10793
rect 13505 10767 13511 10793
rect 13537 10767 13543 10793
rect 15465 10767 15471 10793
rect 15497 10767 15503 10793
rect 16417 10767 16423 10793
rect 16449 10767 16455 10793
rect 17873 10767 17879 10793
rect 17905 10767 17911 10793
rect 19049 10767 19055 10793
rect 19081 10767 19087 10793
rect 672 10597 19320 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 19320 10597
rect 672 10554 19320 10571
rect 1409 10375 1415 10401
rect 1441 10375 1447 10401
rect 2473 10375 2479 10401
rect 2505 10375 2511 10401
rect 3369 10375 3375 10401
rect 3401 10375 3407 10401
rect 3761 10375 3767 10401
rect 3793 10375 3799 10401
rect 3985 10375 3991 10401
rect 4017 10375 4023 10401
rect 4657 10375 4663 10401
rect 4689 10375 4695 10401
rect 5105 10375 5111 10401
rect 5137 10375 5143 10401
rect 5833 10375 5839 10401
rect 5865 10375 5871 10401
rect 6953 10375 6959 10401
rect 6985 10375 6991 10401
rect 7793 10375 7799 10401
rect 7825 10375 7831 10401
rect 8409 10375 8415 10401
rect 8441 10375 8447 10401
rect 9249 10375 9255 10401
rect 9281 10375 9287 10401
rect 10817 10375 10823 10401
rect 10849 10375 10855 10401
rect 11377 10375 11383 10401
rect 11409 10375 11415 10401
rect 11489 10375 11495 10401
rect 11521 10375 11527 10401
rect 12273 10375 12279 10401
rect 12305 10375 12311 10401
rect 13449 10375 13455 10401
rect 13481 10375 13487 10401
rect 15745 10375 15751 10401
rect 15777 10375 15783 10401
rect 16921 10375 16927 10401
rect 16953 10375 16959 10401
rect 17481 10375 17487 10401
rect 17513 10375 17519 10401
rect 17761 10375 17767 10401
rect 17793 10375 17799 10401
rect 17873 10375 17879 10401
rect 17905 10375 17911 10401
rect 2473 10319 2479 10345
rect 2505 10319 2511 10345
rect 7793 10319 7799 10345
rect 7825 10319 7831 10345
rect 9249 10319 9255 10345
rect 9281 10319 9287 10345
rect 13449 10319 13455 10345
rect 13481 10319 13487 10345
rect 15745 10319 15751 10345
rect 15777 10319 15783 10345
rect 672 10205 19320 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 19320 10205
rect 672 10162 19320 10179
rect 3033 10039 3039 10065
rect 3065 10039 3071 10065
rect 11265 10039 11271 10065
rect 11297 10039 11303 10065
rect 17873 10039 17879 10065
rect 17905 10039 17911 10065
rect 1913 9983 1919 10009
rect 1945 9983 1951 10009
rect 3033 9983 3039 10009
rect 3065 9983 3071 10009
rect 3369 9983 3375 10009
rect 3401 9983 3407 10009
rect 3761 9983 3767 10009
rect 3793 9983 3799 10009
rect 3985 9983 3991 10009
rect 4017 9983 4023 10009
rect 4993 9983 4999 10009
rect 5025 9983 5031 10009
rect 5441 9983 5447 10009
rect 5473 9983 5479 10009
rect 5553 9983 5559 10009
rect 5585 9983 5591 10009
rect 6337 9983 6343 10009
rect 6369 9983 6375 10009
rect 6897 9983 6903 10009
rect 6929 9983 6935 10009
rect 7009 9983 7015 10009
rect 7041 9983 7047 10009
rect 9081 9983 9087 10009
rect 9113 9983 9119 10009
rect 9305 9983 9311 10009
rect 9337 9983 9343 10009
rect 9529 9983 9535 10009
rect 9561 9983 9567 10009
rect 10313 9983 10319 10009
rect 10345 9983 10351 10009
rect 11265 9983 11271 10009
rect 11297 9983 11303 10009
rect 12833 9983 12839 10009
rect 12865 9983 12871 10009
rect 13393 9983 13399 10009
rect 13425 9983 13431 10009
rect 13505 9983 13511 10009
rect 13537 9983 13543 10009
rect 15745 9983 15751 10009
rect 15777 9983 15783 10009
rect 15969 9983 15975 10009
rect 16001 9983 16007 10009
rect 16417 9983 16423 10009
rect 16449 9983 16455 10009
rect 17873 9983 17879 10009
rect 17905 9983 17911 10009
rect 18769 9983 18775 10009
rect 18801 9983 18807 10009
rect 672 9813 19320 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 19320 9813
rect 672 9770 19320 9787
rect 1577 9591 1583 9617
rect 1609 9591 1615 9617
rect 2473 9591 2479 9617
rect 2505 9591 2511 9617
rect 3313 9591 3319 9617
rect 3345 9591 3351 9617
rect 3649 9591 3655 9617
rect 3681 9591 3687 9617
rect 3761 9591 3767 9617
rect 3793 9591 3799 9617
rect 4937 9591 4943 9617
rect 4969 9591 4975 9617
rect 5105 9591 5111 9617
rect 5137 9591 5143 9617
rect 5553 9591 5559 9617
rect 5585 9591 5591 9617
rect 6841 9591 6847 9617
rect 6873 9591 6879 9617
rect 7289 9591 7295 9617
rect 7321 9591 7327 9617
rect 7513 9591 7519 9617
rect 7545 9591 7551 9617
rect 8409 9591 8415 9617
rect 8441 9591 8447 9617
rect 8745 9591 8751 9617
rect 8777 9591 8783 9617
rect 8969 9591 8975 9617
rect 9001 9591 9007 9617
rect 10817 9591 10823 9617
rect 10849 9591 10855 9617
rect 11265 9591 11271 9617
rect 11297 9591 11303 9617
rect 11489 9591 11495 9617
rect 11521 9591 11527 9617
rect 12553 9591 12559 9617
rect 12585 9591 12591 9617
rect 13337 9591 13343 9617
rect 13369 9591 13375 9617
rect 16249 9591 16255 9617
rect 16281 9591 16287 9617
rect 16473 9591 16479 9617
rect 16505 9591 16511 9617
rect 16753 9591 16759 9617
rect 16785 9591 16791 9617
rect 17201 9591 17207 9617
rect 17233 9591 17239 9617
rect 17761 9591 17767 9617
rect 17793 9591 17799 9617
rect 17873 9591 17879 9617
rect 17905 9591 17911 9617
rect 2473 9535 2479 9561
rect 2505 9535 2511 9561
rect 13337 9535 13343 9561
rect 13369 9535 13375 9561
rect 672 9421 19320 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 19320 9421
rect 672 9378 19320 9395
rect 2809 9255 2815 9281
rect 2841 9255 2847 9281
rect 11265 9255 11271 9281
rect 11297 9255 11303 9281
rect 17873 9255 17879 9281
rect 17905 9255 17911 9281
rect 1913 9199 1919 9225
rect 1945 9199 1951 9225
rect 2809 9199 2815 9225
rect 2841 9199 2847 9225
rect 3313 9199 3319 9225
rect 3345 9199 3351 9225
rect 3649 9199 3655 9225
rect 3681 9199 3687 9225
rect 3761 9199 3767 9225
rect 3793 9199 3799 9225
rect 4993 9199 4999 9225
rect 5025 9199 5031 9225
rect 5441 9199 5447 9225
rect 5473 9199 5479 9225
rect 5553 9199 5559 9225
rect 5585 9199 5591 9225
rect 6337 9199 6343 9225
rect 6369 9199 6375 9225
rect 6897 9199 6903 9225
rect 6929 9199 6935 9225
rect 7009 9199 7015 9225
rect 7041 9199 7047 9225
rect 9081 9199 9087 9225
rect 9113 9199 9119 9225
rect 9305 9199 9311 9225
rect 9337 9199 9343 9225
rect 9529 9199 9535 9225
rect 9561 9199 9567 9225
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 10985 9199 10991 9225
rect 11017 9199 11023 9225
rect 12833 9199 12839 9225
rect 12865 9199 12871 9225
rect 13337 9199 13343 9225
rect 13369 9199 13375 9225
rect 13505 9199 13511 9225
rect 13537 9199 13543 9225
rect 14289 9199 14295 9225
rect 14321 9199 14327 9225
rect 14737 9199 14743 9225
rect 14769 9199 14775 9225
rect 14961 9199 14967 9225
rect 14993 9199 14999 9225
rect 17873 9199 17879 9225
rect 17905 9199 17911 9225
rect 18769 9199 18775 9225
rect 18801 9199 18807 9225
rect 672 9029 19320 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 19320 9029
rect 672 8986 19320 9003
rect 1577 8807 1583 8833
rect 1609 8807 1615 8833
rect 2473 8807 2479 8833
rect 2505 8807 2511 8833
rect 3313 8807 3319 8833
rect 3345 8807 3351 8833
rect 3649 8807 3655 8833
rect 3681 8807 3687 8833
rect 3761 8807 3767 8833
rect 3793 8807 3799 8833
rect 4937 8807 4943 8833
rect 4969 8807 4975 8833
rect 5105 8807 5111 8833
rect 5137 8807 5143 8833
rect 5553 8807 5559 8833
rect 5585 8807 5591 8833
rect 6841 8807 6847 8833
rect 6873 8807 6879 8833
rect 7289 8807 7295 8833
rect 7321 8807 7327 8833
rect 7513 8807 7519 8833
rect 7545 8807 7551 8833
rect 8409 8807 8415 8833
rect 8441 8807 8447 8833
rect 8745 8807 8751 8833
rect 8777 8807 8783 8833
rect 8969 8807 8975 8833
rect 9001 8807 9007 8833
rect 11097 8807 11103 8833
rect 11129 8807 11135 8833
rect 11265 8807 11271 8833
rect 11297 8807 11303 8833
rect 11489 8807 11495 8833
rect 11521 8807 11527 8833
rect 12273 8807 12279 8833
rect 12305 8807 12311 8833
rect 13393 8807 13399 8833
rect 13425 8807 13431 8833
rect 14793 8807 14799 8833
rect 14825 8807 14831 8833
rect 15241 8807 15247 8833
rect 15273 8807 15279 8833
rect 15465 8807 15471 8833
rect 15497 8807 15503 8833
rect 17201 8807 17207 8833
rect 17233 8807 17239 8833
rect 17761 8807 17767 8833
rect 17793 8807 17799 8833
rect 17873 8807 17879 8833
rect 17905 8807 17911 8833
rect 2473 8751 2479 8777
rect 2505 8751 2511 8777
rect 13393 8751 13399 8777
rect 13425 8751 13431 8777
rect 672 8637 19320 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 19320 8637
rect 672 8594 19320 8611
rect 2809 8471 2815 8497
rect 2841 8471 2847 8497
rect 11265 8471 11271 8497
rect 11297 8471 11303 8497
rect 15353 8471 15359 8497
rect 15385 8471 15391 8497
rect 17873 8471 17879 8497
rect 17905 8471 17911 8497
rect 1913 8415 1919 8441
rect 1945 8415 1951 8441
rect 2809 8415 2815 8441
rect 2841 8415 2847 8441
rect 3313 8415 3319 8441
rect 3345 8415 3351 8441
rect 3649 8415 3655 8441
rect 3681 8415 3687 8441
rect 3761 8415 3767 8441
rect 3793 8415 3799 8441
rect 4993 8415 4999 8441
rect 5025 8415 5031 8441
rect 5441 8415 5447 8441
rect 5473 8415 5479 8441
rect 5553 8415 5559 8441
rect 5585 8415 5591 8441
rect 6337 8415 6343 8441
rect 6369 8415 6375 8441
rect 6897 8415 6903 8441
rect 6929 8415 6935 8441
rect 7009 8415 7015 8441
rect 7041 8415 7047 8441
rect 9081 8415 9087 8441
rect 9113 8415 9119 8441
rect 9305 8415 9311 8441
rect 9337 8415 9343 8441
rect 9529 8415 9535 8441
rect 9561 8415 9567 8441
rect 10593 8415 10599 8441
rect 10625 8415 10631 8441
rect 11265 8415 11271 8441
rect 11297 8415 11303 8441
rect 12833 8415 12839 8441
rect 12865 8415 12871 8441
rect 13393 8415 13399 8441
rect 13425 8415 13431 8441
rect 13505 8415 13511 8441
rect 13537 8415 13543 8441
rect 14289 8415 14295 8441
rect 14321 8415 14327 8441
rect 15353 8415 15359 8441
rect 15385 8415 15391 8441
rect 17873 8415 17879 8441
rect 17905 8415 17911 8441
rect 18769 8415 18775 8441
rect 18801 8415 18807 8441
rect 672 8245 19320 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 19320 8245
rect 672 8202 19320 8219
rect 1577 8023 1583 8049
rect 1609 8023 1615 8049
rect 2473 8023 2479 8049
rect 2505 8023 2511 8049
rect 3313 8023 3319 8049
rect 3345 8023 3351 8049
rect 3649 8023 3655 8049
rect 3681 8023 3687 8049
rect 3817 8023 3823 8049
rect 3849 8023 3855 8049
rect 4993 8023 4999 8049
rect 5025 8023 5031 8049
rect 5553 8023 5559 8049
rect 5585 8023 5591 8049
rect 6841 8023 6847 8049
rect 6873 8023 6879 8049
rect 7289 8023 7295 8049
rect 7321 8023 7327 8049
rect 7513 8023 7519 8049
rect 7545 8023 7551 8049
rect 8409 8023 8415 8049
rect 8441 8023 8447 8049
rect 8745 8023 8751 8049
rect 8777 8023 8783 8049
rect 8969 8023 8975 8049
rect 9001 8023 9007 8049
rect 11097 8023 11103 8049
rect 11129 8023 11135 8049
rect 11993 8023 11999 8049
rect 12025 8023 12031 8049
rect 12273 8023 12279 8049
rect 12305 8023 12311 8049
rect 13337 8023 13343 8049
rect 13369 8023 13375 8049
rect 15185 8023 15191 8049
rect 15217 8023 15223 8049
rect 15409 8023 15415 8049
rect 15441 8023 15447 8049
rect 15689 8023 15695 8049
rect 15721 8023 15727 8049
rect 17201 8023 17207 8049
rect 17233 8023 17239 8049
rect 17761 8023 17767 8049
rect 17793 8023 17799 8049
rect 17873 8023 17879 8049
rect 17905 8023 17911 8049
rect 2473 7967 2479 7993
rect 2505 7967 2511 7993
rect 5665 7967 5671 7993
rect 5697 7967 5703 7993
rect 11993 7967 11999 7993
rect 12025 7967 12031 7993
rect 13337 7967 13343 7993
rect 13369 7967 13375 7993
rect 672 7853 19320 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 19320 7853
rect 672 7810 19320 7827
rect 3033 7687 3039 7713
rect 3065 7687 3071 7713
rect 11489 7687 11495 7713
rect 11521 7687 11527 7713
rect 15353 7687 15359 7713
rect 15385 7687 15391 7713
rect 17873 7687 17879 7713
rect 17905 7687 17911 7713
rect 2137 7631 2143 7657
rect 2169 7631 2175 7657
rect 3033 7631 3039 7657
rect 3065 7631 3071 7657
rect 3593 7631 3599 7657
rect 3625 7631 3631 7657
rect 3817 7631 3823 7657
rect 3849 7631 3855 7657
rect 3985 7631 3991 7657
rect 4017 7631 4023 7657
rect 4993 7631 4999 7657
rect 5025 7631 5031 7657
rect 5441 7631 5447 7657
rect 5473 7631 5479 7657
rect 5553 7631 5559 7657
rect 5585 7631 5591 7657
rect 6337 7631 6343 7657
rect 6369 7631 6375 7657
rect 6897 7631 6903 7657
rect 6929 7631 6935 7657
rect 7009 7631 7015 7657
rect 7041 7631 7047 7657
rect 9081 7631 9087 7657
rect 9113 7631 9119 7657
rect 9305 7631 9311 7657
rect 9337 7631 9343 7657
rect 9529 7631 9535 7657
rect 9561 7631 9567 7657
rect 10593 7631 10599 7657
rect 10625 7631 10631 7657
rect 11489 7631 11495 7657
rect 11521 7631 11527 7657
rect 12833 7631 12839 7657
rect 12865 7631 12871 7657
rect 13393 7631 13399 7657
rect 13425 7631 13431 7657
rect 13505 7631 13511 7657
rect 13537 7631 13543 7657
rect 14289 7631 14295 7657
rect 14321 7631 14327 7657
rect 15353 7631 15359 7657
rect 15385 7631 15391 7657
rect 17873 7631 17879 7657
rect 17905 7631 17911 7657
rect 18769 7631 18775 7657
rect 18801 7631 18807 7657
rect 672 7461 19320 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 19320 7461
rect 672 7418 19320 7435
rect 1577 7239 1583 7265
rect 1609 7239 1615 7265
rect 2473 7239 2479 7265
rect 2505 7239 2511 7265
rect 3537 7239 3543 7265
rect 3569 7239 3575 7265
rect 3817 7239 3823 7265
rect 3849 7239 3855 7265
rect 3929 7239 3935 7265
rect 3961 7239 3967 7265
rect 4993 7239 4999 7265
rect 5025 7239 5031 7265
rect 5553 7239 5559 7265
rect 5585 7239 5591 7265
rect 6841 7239 6847 7265
rect 6873 7239 6879 7265
rect 7289 7239 7295 7265
rect 7321 7239 7327 7265
rect 7513 7239 7519 7265
rect 7545 7239 7551 7265
rect 8409 7239 8415 7265
rect 8441 7239 8447 7265
rect 8745 7239 8751 7265
rect 8777 7239 8783 7265
rect 8969 7239 8975 7265
rect 9001 7239 9007 7265
rect 11097 7239 11103 7265
rect 11129 7239 11135 7265
rect 11993 7239 11999 7265
rect 12025 7239 12031 7265
rect 12273 7239 12279 7265
rect 12305 7239 12311 7265
rect 13393 7239 13399 7265
rect 13425 7239 13431 7265
rect 14793 7239 14799 7265
rect 14825 7239 14831 7265
rect 15241 7239 15247 7265
rect 15273 7239 15279 7265
rect 15465 7239 15471 7265
rect 15497 7239 15503 7265
rect 16249 7239 16255 7265
rect 16281 7239 16287 7265
rect 17145 7239 17151 7265
rect 17177 7239 17183 7265
rect 2473 7183 2479 7209
rect 2505 7183 2511 7209
rect 5665 7183 5671 7209
rect 5697 7183 5703 7209
rect 11993 7183 11999 7209
rect 12025 7183 12031 7209
rect 13393 7183 13399 7209
rect 13425 7183 13431 7209
rect 16249 7183 16255 7209
rect 16281 7183 16287 7209
rect 672 7069 19320 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 19320 7069
rect 672 7026 19320 7043
rect 10985 6903 10991 6929
rect 11017 6903 11023 6929
rect 12441 6903 12447 6929
rect 12473 6903 12479 6929
rect 14009 6903 14015 6929
rect 14041 6903 14047 6929
rect 15241 6903 15247 6929
rect 15273 6903 15279 6929
rect 17873 6903 17879 6929
rect 17905 6903 17911 6929
rect 2081 6847 2087 6873
rect 2113 6847 2119 6873
rect 2417 6847 2423 6873
rect 2449 6847 2455 6873
rect 2529 6847 2535 6873
rect 2561 6847 2567 6873
rect 3537 6847 3543 6873
rect 3569 6847 3575 6873
rect 3817 6847 3823 6873
rect 3849 6847 3855 6873
rect 3985 6847 3991 6873
rect 4017 6847 4023 6873
rect 4993 6847 4999 6873
rect 5025 6847 5031 6873
rect 5441 6847 5447 6873
rect 5473 6847 5479 6873
rect 5553 6847 5559 6873
rect 5585 6847 5591 6873
rect 6337 6847 6343 6873
rect 6369 6847 6375 6873
rect 6897 6847 6903 6873
rect 6929 6847 6935 6873
rect 7009 6847 7015 6873
rect 7041 6847 7047 6873
rect 9809 6847 9815 6873
rect 9841 6847 9847 6873
rect 10985 6847 10991 6873
rect 11017 6847 11023 6873
rect 11265 6847 11271 6873
rect 11297 6847 11303 6873
rect 12441 6847 12447 6873
rect 12473 6847 12479 6873
rect 12833 6847 12839 6873
rect 12865 6847 12871 6873
rect 14009 6847 14015 6873
rect 14041 6847 14047 6873
rect 14289 6847 14295 6873
rect 14321 6847 14327 6873
rect 15241 6847 15247 6873
rect 15273 6847 15279 6873
rect 17873 6847 17879 6873
rect 17905 6847 17911 6873
rect 18769 6847 18775 6873
rect 18801 6847 18807 6873
rect 672 6677 19320 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 19320 6677
rect 672 6634 19320 6651
rect 1577 6455 1583 6481
rect 1609 6455 1615 6481
rect 2417 6455 2423 6481
rect 2449 6455 2455 6481
rect 3537 6455 3543 6481
rect 3569 6455 3575 6481
rect 3817 6455 3823 6481
rect 3849 6455 3855 6481
rect 3929 6455 3935 6481
rect 3961 6455 3967 6481
rect 4993 6455 4999 6481
rect 5025 6455 5031 6481
rect 5553 6455 5559 6481
rect 5585 6455 5591 6481
rect 6841 6455 6847 6481
rect 6873 6455 6879 6481
rect 7289 6455 7295 6481
rect 7321 6455 7327 6481
rect 7513 6455 7519 6481
rect 7545 6455 7551 6481
rect 9529 6455 9535 6481
rect 9561 6455 9567 6481
rect 10425 6455 10431 6481
rect 10457 6455 10463 6481
rect 11097 6455 11103 6481
rect 11129 6455 11135 6481
rect 11993 6455 11999 6481
rect 12025 6455 12031 6481
rect 12273 6455 12279 6481
rect 12305 6455 12311 6481
rect 13393 6455 13399 6481
rect 13425 6455 13431 6481
rect 15241 6455 15247 6481
rect 15273 6455 15279 6481
rect 15409 6455 15415 6481
rect 15441 6455 15447 6481
rect 15689 6455 15695 6481
rect 15721 6455 15727 6481
rect 17201 6455 17207 6481
rect 17233 6455 17239 6481
rect 17985 6455 17991 6481
rect 18017 6455 18023 6481
rect 2417 6399 2423 6425
rect 2449 6399 2455 6425
rect 5665 6399 5671 6425
rect 5697 6399 5703 6425
rect 10425 6399 10431 6425
rect 10457 6399 10463 6425
rect 11993 6399 11999 6425
rect 12025 6399 12031 6425
rect 13393 6399 13399 6425
rect 13425 6399 13431 6425
rect 18153 6399 18159 6425
rect 18185 6399 18191 6425
rect 672 6285 19320 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 19320 6285
rect 672 6242 19320 6259
rect 2417 6119 2423 6145
rect 2449 6119 2455 6145
rect 10985 6119 10991 6145
rect 11017 6119 11023 6145
rect 12441 6119 12447 6145
rect 12473 6119 12479 6145
rect 15241 6119 15247 6145
rect 15273 6119 15279 6145
rect 18097 6119 18103 6145
rect 18129 6119 18135 6145
rect 1633 6063 1639 6089
rect 1665 6063 1671 6089
rect 2417 6063 2423 6089
rect 2449 6063 2455 6089
rect 3537 6063 3543 6089
rect 3569 6063 3575 6089
rect 3873 6063 3879 6089
rect 3905 6063 3911 6089
rect 3985 6063 3991 6089
rect 4017 6063 4023 6089
rect 4993 6063 4999 6089
rect 5025 6063 5031 6089
rect 5441 6063 5447 6089
rect 5473 6063 5479 6089
rect 5553 6063 5559 6089
rect 5585 6063 5591 6089
rect 6337 6063 6343 6089
rect 6369 6063 6375 6089
rect 6785 6063 6791 6089
rect 6817 6063 6823 6089
rect 7009 6063 7015 6089
rect 7041 6063 7047 6089
rect 9809 6063 9815 6089
rect 9841 6063 9847 6089
rect 10985 6063 10991 6089
rect 11017 6063 11023 6089
rect 11265 6063 11271 6089
rect 11297 6063 11303 6089
rect 12441 6063 12447 6089
rect 12473 6063 12479 6089
rect 12833 6063 12839 6089
rect 12865 6063 12871 6089
rect 13393 6063 13399 6089
rect 13425 6063 13431 6089
rect 13505 6063 13511 6089
rect 13537 6063 13543 6089
rect 14569 6063 14575 6089
rect 14601 6063 14607 6089
rect 15241 6063 15247 6089
rect 15273 6063 15279 6089
rect 18097 6063 18103 6089
rect 18129 6063 18135 6089
rect 18769 6063 18775 6089
rect 18801 6063 18807 6089
rect 672 5893 19320 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 19320 5893
rect 672 5850 19320 5867
rect 1577 5671 1583 5697
rect 1609 5671 1615 5697
rect 2417 5671 2423 5697
rect 2449 5671 2455 5697
rect 2865 5671 2871 5697
rect 2897 5671 2903 5697
rect 3369 5671 3375 5697
rect 3401 5671 3407 5697
rect 3537 5671 3543 5697
rect 3569 5671 3575 5697
rect 4993 5671 4999 5697
rect 5025 5671 5031 5697
rect 5553 5671 5559 5697
rect 5585 5671 5591 5697
rect 8297 5671 8303 5697
rect 8329 5671 8335 5697
rect 8409 5671 8415 5697
rect 8441 5671 8447 5697
rect 8969 5671 8975 5697
rect 9001 5671 9007 5697
rect 9529 5671 9535 5697
rect 9561 5671 9567 5697
rect 10425 5671 10431 5697
rect 10457 5671 10463 5697
rect 11097 5671 11103 5697
rect 11129 5671 11135 5697
rect 11993 5671 11999 5697
rect 12025 5671 12031 5697
rect 12273 5671 12279 5697
rect 12305 5671 12311 5697
rect 13393 5671 13399 5697
rect 13425 5671 13431 5697
rect 14905 5671 14911 5697
rect 14937 5671 14943 5697
rect 15969 5671 15975 5697
rect 16001 5671 16007 5697
rect 16249 5671 16255 5697
rect 16281 5671 16287 5697
rect 17145 5671 17151 5697
rect 17177 5671 17183 5697
rect 2417 5615 2423 5641
rect 2449 5615 2455 5641
rect 5665 5615 5671 5641
rect 5697 5615 5703 5641
rect 10425 5615 10431 5641
rect 10457 5615 10463 5641
rect 11993 5615 11999 5641
rect 12025 5615 12031 5641
rect 13393 5615 13399 5641
rect 13425 5615 13431 5641
rect 15969 5615 15975 5641
rect 16001 5615 16007 5641
rect 16249 5615 16255 5641
rect 16281 5615 16287 5641
rect 672 5501 19320 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 19320 5501
rect 672 5458 19320 5475
rect 2417 5335 2423 5361
rect 2449 5335 2455 5361
rect 8353 5335 8359 5361
rect 8385 5335 8391 5361
rect 10985 5335 10991 5361
rect 11017 5335 11023 5361
rect 12273 5335 12279 5361
rect 12305 5335 12311 5361
rect 14009 5335 14015 5361
rect 14041 5335 14047 5361
rect 15465 5335 15471 5361
rect 15497 5335 15503 5361
rect 18097 5335 18103 5361
rect 18129 5335 18135 5361
rect 1633 5279 1639 5305
rect 1665 5279 1671 5305
rect 2417 5279 2423 5305
rect 2449 5279 2455 5305
rect 2865 5279 2871 5305
rect 2897 5279 2903 5305
rect 3425 5279 3431 5305
rect 3457 5279 3463 5305
rect 3537 5279 3543 5305
rect 3569 5279 3575 5305
rect 4993 5279 4999 5305
rect 5025 5279 5031 5305
rect 5385 5279 5391 5305
rect 5417 5279 5423 5305
rect 5553 5279 5559 5305
rect 5585 5279 5591 5305
rect 7513 5279 7519 5305
rect 7545 5279 7551 5305
rect 8353 5279 8359 5305
rect 8385 5279 8391 5305
rect 10033 5279 10039 5305
rect 10065 5279 10071 5305
rect 10985 5279 10991 5305
rect 11017 5279 11023 5305
rect 11377 5279 11383 5305
rect 11409 5279 11415 5305
rect 12273 5279 12279 5305
rect 12305 5279 12311 5305
rect 13113 5279 13119 5305
rect 13145 5279 13151 5305
rect 14009 5279 14015 5305
rect 14041 5279 14047 5305
rect 14569 5279 14575 5305
rect 14601 5279 14607 5305
rect 15465 5279 15471 5305
rect 15497 5279 15503 5305
rect 18097 5279 18103 5305
rect 18129 5279 18135 5305
rect 18769 5279 18775 5305
rect 18801 5279 18807 5305
rect 672 5109 19320 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 19320 5109
rect 672 5066 19320 5083
rect 1577 4887 1583 4913
rect 1609 4887 1615 4913
rect 2417 4887 2423 4913
rect 2449 4887 2455 4913
rect 2865 4887 2871 4913
rect 2897 4887 2903 4913
rect 3425 4887 3431 4913
rect 3457 4887 3463 4913
rect 3537 4887 3543 4913
rect 3569 4887 3575 4913
rect 4993 4887 4999 4913
rect 5025 4887 5031 4913
rect 5161 4887 5167 4913
rect 5193 4887 5199 4913
rect 5385 4887 5391 4913
rect 5417 4887 5423 4913
rect 7793 4887 7799 4913
rect 7825 4887 7831 4913
rect 8353 4887 8359 4913
rect 8385 4887 8391 4913
rect 8465 4887 8471 4913
rect 8497 4887 8503 4913
rect 9529 4887 9535 4913
rect 9561 4887 9567 4913
rect 10425 4887 10431 4913
rect 10457 4887 10463 4913
rect 11097 4887 11103 4913
rect 11129 4887 11135 4913
rect 11993 4887 11999 4913
rect 12025 4887 12031 4913
rect 12553 4887 12559 4913
rect 12585 4887 12591 4913
rect 13393 4887 13399 4913
rect 13425 4887 13431 4913
rect 14849 4887 14855 4913
rect 14881 4887 14887 4913
rect 15913 4887 15919 4913
rect 15945 4887 15951 4913
rect 17705 4887 17711 4913
rect 17737 4887 17743 4913
rect 17929 4887 17935 4913
rect 17961 4887 17967 4913
rect 18377 4887 18383 4913
rect 18409 4887 18415 4913
rect 2417 4831 2423 4857
rect 2449 4831 2455 4857
rect 10425 4831 10431 4857
rect 10457 4831 10463 4857
rect 11993 4831 11999 4857
rect 12025 4831 12031 4857
rect 13393 4831 13399 4857
rect 13425 4831 13431 4857
rect 14849 4831 14855 4857
rect 14881 4831 14887 4857
rect 672 4717 19320 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 19320 4717
rect 672 4674 19320 4691
rect 2417 4551 2423 4577
rect 2449 4551 2455 4577
rect 6057 4551 6063 4577
rect 6089 4551 6095 4577
rect 8465 4551 8471 4577
rect 8497 4551 8503 4577
rect 10761 4551 10767 4577
rect 10793 4551 10799 4577
rect 12273 4551 12279 4577
rect 12305 4551 12311 4577
rect 14009 4551 14015 4577
rect 14041 4551 14047 4577
rect 17985 4551 17991 4577
rect 18017 4551 18023 4577
rect 1577 4495 1583 4521
rect 1609 4495 1615 4521
rect 2417 4495 2423 4521
rect 2449 4495 2455 4521
rect 2865 4495 2871 4521
rect 2897 4495 2903 4521
rect 3369 4495 3375 4521
rect 3401 4495 3407 4521
rect 3537 4495 3543 4521
rect 3569 4495 3575 4521
rect 6057 4495 6063 4521
rect 6089 4495 6095 4521
rect 7009 4495 7015 4521
rect 7041 4495 7047 4521
rect 7569 4495 7575 4521
rect 7601 4495 7607 4521
rect 8465 4495 8471 4521
rect 8497 4495 8503 4521
rect 10033 4495 10039 4521
rect 10065 4495 10071 4521
rect 10761 4495 10767 4521
rect 10793 4495 10799 4521
rect 11377 4495 11383 4521
rect 11409 4495 11415 4521
rect 11993 4495 11999 4521
rect 12025 4495 12031 4521
rect 13113 4495 13119 4521
rect 13145 4495 13151 4521
rect 14009 4495 14015 4521
rect 14041 4495 14047 4521
rect 14569 4495 14575 4521
rect 14601 4495 14607 4521
rect 14849 4495 14855 4521
rect 14881 4495 14887 4521
rect 14961 4495 14967 4521
rect 14993 4495 14999 4521
rect 17985 4495 17991 4521
rect 18017 4495 18023 4521
rect 18769 4495 18775 4521
rect 18801 4495 18807 4521
rect 672 4325 19320 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 19320 4325
rect 672 4282 19320 4299
rect 905 4103 911 4129
rect 937 4103 943 4129
rect 2081 4103 2087 4129
rect 2113 4103 2119 4129
rect 3873 4103 3879 4129
rect 3905 4103 3911 4129
rect 4993 4103 4999 4129
rect 5025 4103 5031 4129
rect 5777 4103 5783 4129
rect 5809 4103 5815 4129
rect 6001 4103 6007 4129
rect 6033 4103 6039 4129
rect 6449 4103 6455 4129
rect 6481 4103 6487 4129
rect 7793 4103 7799 4129
rect 7825 4103 7831 4129
rect 8465 4103 8471 4129
rect 8497 4103 8503 4129
rect 9529 4103 9535 4129
rect 9561 4103 9567 4129
rect 10425 4103 10431 4129
rect 10457 4103 10463 4129
rect 11097 4103 11103 4129
rect 11129 4103 11135 4129
rect 11769 4103 11775 4129
rect 11801 4103 11807 4129
rect 12553 4103 12559 4129
rect 12585 4103 12591 4129
rect 13225 4103 13231 4129
rect 13257 4103 13263 4129
rect 16249 4103 16255 4129
rect 16281 4103 16287 4129
rect 16473 4103 16479 4129
rect 16505 4103 16511 4129
rect 16753 4103 16759 4129
rect 16785 4103 16791 4129
rect 17705 4103 17711 4129
rect 17737 4103 17743 4129
rect 17873 4103 17879 4129
rect 17905 4103 17911 4129
rect 18377 4103 18383 4129
rect 18409 4103 18415 4129
rect 2081 4047 2087 4073
rect 2113 4047 2119 4073
rect 3873 4047 3879 4073
rect 3905 4047 3911 4073
rect 8745 4047 8751 4073
rect 8777 4047 8783 4073
rect 10425 4047 10431 4073
rect 10457 4047 10463 4073
rect 11769 4047 11775 4073
rect 11801 4047 11807 4073
rect 13225 4047 13231 4073
rect 13257 4047 13263 4073
rect 672 3933 19320 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 19320 3933
rect 672 3890 19320 3907
rect 2081 3767 2087 3793
rect 2113 3767 2119 3793
rect 8353 3767 8359 3793
rect 8385 3767 8391 3793
rect 12441 3767 12447 3793
rect 12473 3767 12479 3793
rect 15409 3767 15415 3793
rect 15441 3767 15447 3793
rect 17873 3767 17879 3793
rect 17905 3767 17911 3793
rect 905 3711 911 3737
rect 937 3711 943 3737
rect 2081 3711 2087 3737
rect 2113 3711 2119 3737
rect 3817 3711 3823 3737
rect 3849 3711 3855 3737
rect 4041 3711 4047 3737
rect 4073 3711 4079 3737
rect 4489 3711 4495 3737
rect 4521 3711 4527 3737
rect 6337 3711 6343 3737
rect 6369 3711 6375 3737
rect 6561 3711 6567 3737
rect 6593 3711 6599 3737
rect 7009 3711 7015 3737
rect 7041 3711 7047 3737
rect 7513 3711 7519 3737
rect 7545 3711 7551 3737
rect 8353 3711 8359 3737
rect 8385 3711 8391 3737
rect 9809 3711 9815 3737
rect 9841 3711 9847 3737
rect 10369 3711 10375 3737
rect 10401 3711 10407 3737
rect 10481 3711 10487 3737
rect 10513 3711 10519 3737
rect 11545 3711 11551 3737
rect 11577 3711 11583 3737
rect 12441 3711 12447 3737
rect 12473 3711 12479 3737
rect 13113 3711 13119 3737
rect 13145 3711 13151 3737
rect 13281 3711 13287 3737
rect 13313 3711 13319 3737
rect 13561 3711 13567 3737
rect 13593 3711 13599 3737
rect 14513 3711 14519 3737
rect 14545 3711 14551 3737
rect 15353 3711 15359 3737
rect 15385 3711 15391 3737
rect 17873 3711 17879 3737
rect 17905 3711 17911 3737
rect 18825 3711 18831 3737
rect 18857 3711 18863 3737
rect 672 3541 19320 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 19320 3541
rect 672 3498 19320 3515
rect 905 3319 911 3345
rect 937 3319 943 3345
rect 2081 3319 2087 3345
rect 2113 3319 2119 3345
rect 3817 3319 3823 3345
rect 3849 3319 3855 3345
rect 4993 3319 4999 3345
rect 5025 3319 5031 3345
rect 5553 3319 5559 3345
rect 5585 3319 5591 3345
rect 5833 3319 5839 3345
rect 5865 3319 5871 3345
rect 5945 3319 5951 3345
rect 5977 3319 5983 3345
rect 7793 3319 7799 3345
rect 7825 3319 7831 3345
rect 8801 3319 8807 3345
rect 8833 3319 8839 3345
rect 9249 3319 9255 3345
rect 9281 3319 9287 3345
rect 9753 3319 9759 3345
rect 9785 3319 9791 3345
rect 9921 3319 9927 3345
rect 9953 3319 9959 3345
rect 11097 3319 11103 3345
rect 11129 3319 11135 3345
rect 11377 3319 11383 3345
rect 11409 3319 11415 3345
rect 11489 3319 11495 3345
rect 11521 3319 11527 3345
rect 12553 3319 12559 3345
rect 12585 3319 12591 3345
rect 12721 3319 12727 3345
rect 12753 3319 12759 3345
rect 12945 3319 12951 3345
rect 12977 3319 12983 3345
rect 16249 3319 16255 3345
rect 16281 3319 16287 3345
rect 16361 3319 16367 3345
rect 16393 3319 16399 3345
rect 16921 3319 16927 3345
rect 16953 3319 16959 3345
rect 17705 3319 17711 3345
rect 17737 3319 17743 3345
rect 17817 3319 17823 3345
rect 17849 3319 17855 3345
rect 18377 3319 18383 3345
rect 18409 3319 18415 3345
rect 2081 3263 2087 3289
rect 2113 3263 2119 3289
rect 3817 3263 3823 3289
rect 3849 3263 3855 3289
rect 8801 3263 8807 3289
rect 8833 3263 8839 3289
rect 672 3149 19320 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 19320 3149
rect 672 3106 19320 3123
rect 2025 2983 2031 3009
rect 2057 2983 2063 3009
rect 11713 2983 11719 3009
rect 11745 2983 11751 3009
rect 14009 2983 14015 3009
rect 14041 2983 14047 3009
rect 15241 2983 15247 3009
rect 15273 2983 15279 3009
rect 17985 2983 17991 3009
rect 18017 2983 18023 3009
rect 905 2927 911 2953
rect 937 2927 943 2953
rect 2025 2927 2031 2953
rect 2057 2927 2063 2953
rect 3817 2927 3823 2953
rect 3849 2927 3855 2953
rect 3929 2927 3935 2953
rect 3961 2927 3967 2953
rect 4489 2927 4495 2953
rect 4521 2927 4527 2953
rect 6113 2927 6119 2953
rect 6145 2927 6151 2953
rect 6281 2927 6287 2953
rect 6313 2927 6319 2953
rect 6505 2927 6511 2953
rect 6537 2927 6543 2953
rect 7513 2927 7519 2953
rect 7545 2927 7551 2953
rect 7737 2927 7743 2953
rect 7769 2927 7775 2953
rect 7961 2927 7967 2953
rect 7993 2927 7999 2953
rect 9305 2927 9311 2953
rect 9337 2927 9343 2953
rect 9753 2927 9759 2953
rect 9785 2927 9791 2953
rect 9977 2927 9983 2953
rect 10009 2927 10015 2953
rect 11041 2927 11047 2953
rect 11073 2927 11079 2953
rect 11657 2927 11663 2953
rect 11689 2927 11695 2953
rect 13113 2927 13119 2953
rect 13145 2927 13151 2953
rect 14009 2927 14015 2953
rect 14041 2927 14047 2953
rect 14345 2927 14351 2953
rect 14377 2927 14383 2953
rect 15129 2927 15135 2953
rect 15161 2927 15167 2953
rect 17985 2927 17991 2953
rect 18017 2927 18023 2953
rect 18769 2927 18775 2953
rect 18801 2927 18807 2953
rect 672 2757 19320 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 19320 2757
rect 672 2714 19320 2731
rect 905 2535 911 2561
rect 937 2535 943 2561
rect 2025 2535 2031 2561
rect 2057 2535 2063 2561
rect 3985 2535 3991 2561
rect 4017 2535 4023 2561
rect 4993 2535 4999 2561
rect 5025 2535 5031 2561
rect 5553 2535 5559 2561
rect 5585 2535 5591 2561
rect 6449 2535 6455 2561
rect 6481 2535 6487 2561
rect 8073 2535 8079 2561
rect 8105 2535 8111 2561
rect 8241 2535 8247 2561
rect 8273 2535 8279 2561
rect 8465 2535 8471 2561
rect 8497 2535 8503 2561
rect 9249 2535 9255 2561
rect 9281 2535 9287 2561
rect 10425 2535 10431 2561
rect 10457 2535 10463 2561
rect 11041 2535 11047 2561
rect 11073 2535 11079 2561
rect 11657 2535 11663 2561
rect 11689 2535 11695 2561
rect 12553 2535 12559 2561
rect 12585 2535 12591 2561
rect 13449 2535 13455 2561
rect 13481 2535 13487 2561
rect 14793 2535 14799 2561
rect 14825 2535 14831 2561
rect 15241 2535 15247 2561
rect 15273 2535 15279 2561
rect 15465 2535 15471 2561
rect 15497 2535 15503 2561
rect 17481 2535 17487 2561
rect 17513 2535 17519 2561
rect 17761 2535 17767 2561
rect 17793 2535 17799 2561
rect 17873 2535 17879 2561
rect 17905 2535 17911 2561
rect 2025 2479 2031 2505
rect 2057 2479 2063 2505
rect 3985 2479 3991 2505
rect 4017 2479 4023 2505
rect 6449 2479 6455 2505
rect 6481 2479 6487 2505
rect 10425 2479 10431 2505
rect 10457 2479 10463 2505
rect 11769 2479 11775 2505
rect 11801 2479 11807 2505
rect 13393 2479 13399 2505
rect 13425 2479 13431 2505
rect 672 2365 19320 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 19320 2365
rect 672 2322 19320 2339
rect 2025 2199 2031 2225
rect 2057 2199 2063 2225
rect 7009 2199 7015 2225
rect 7041 2199 7047 2225
rect 8353 2199 8359 2225
rect 8385 2199 8391 2225
rect 10425 2199 10431 2225
rect 10457 2199 10463 2225
rect 13785 2199 13791 2225
rect 13817 2199 13823 2225
rect 15241 2199 15247 2225
rect 15273 2199 15279 2225
rect 17873 2199 17879 2225
rect 17905 2199 17911 2225
rect 905 2143 911 2169
rect 937 2143 943 2169
rect 2025 2143 2031 2169
rect 2057 2143 2063 2169
rect 3817 2143 3823 2169
rect 3849 2143 3855 2169
rect 3929 2143 3935 2169
rect 3961 2143 3967 2169
rect 4489 2143 4495 2169
rect 4521 2143 4527 2169
rect 6113 2143 6119 2169
rect 6145 2143 6151 2169
rect 7009 2143 7015 2169
rect 7041 2143 7047 2169
rect 7513 2143 7519 2169
rect 7545 2143 7551 2169
rect 8353 2143 8359 2169
rect 8385 2143 8391 2169
rect 9249 2143 9255 2169
rect 9281 2143 9287 2169
rect 10425 2143 10431 2169
rect 10457 2143 10463 2169
rect 10873 2143 10879 2169
rect 10905 2143 10911 2169
rect 11153 2143 11159 2169
rect 11185 2143 11191 2169
rect 11377 2143 11383 2169
rect 11409 2143 11415 2169
rect 12833 2143 12839 2169
rect 12865 2143 12871 2169
rect 13617 2143 13623 2169
rect 13649 2143 13655 2169
rect 14289 2143 14295 2169
rect 14321 2143 14327 2169
rect 15241 2143 15247 2169
rect 15273 2143 15279 2169
rect 17873 2143 17879 2169
rect 17905 2143 17911 2169
rect 18769 2143 18775 2169
rect 18801 2143 18807 2169
rect 672 1973 19320 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 19320 1973
rect 672 1930 19320 1947
rect 961 1751 967 1777
rect 993 1751 999 1777
rect 2081 1751 2087 1777
rect 2113 1751 2119 1777
rect 2865 1751 2871 1777
rect 2897 1751 2903 1777
rect 3817 1751 3823 1777
rect 3849 1751 3855 1777
rect 5217 1751 5223 1777
rect 5249 1751 5255 1777
rect 5777 1751 5783 1777
rect 5809 1751 5815 1777
rect 5889 1751 5895 1777
rect 5921 1751 5927 1777
rect 7457 1751 7463 1777
rect 7489 1751 7495 1777
rect 7625 1751 7631 1777
rect 7657 1751 7663 1777
rect 7849 1751 7855 1777
rect 7881 1751 7887 1777
rect 9417 1751 9423 1777
rect 9449 1751 9455 1777
rect 9585 1751 9591 1777
rect 9617 1751 9623 1777
rect 9809 1751 9815 1777
rect 9841 1751 9847 1777
rect 10873 1751 10879 1777
rect 10905 1751 10911 1777
rect 11657 1751 11663 1777
rect 11689 1751 11695 1777
rect 12665 1751 12671 1777
rect 12697 1751 12703 1777
rect 13617 1751 13623 1777
rect 13649 1751 13655 1777
rect 14737 1751 14743 1777
rect 14769 1751 14775 1777
rect 15521 1751 15527 1777
rect 15553 1751 15559 1777
rect 2081 1695 2087 1721
rect 2113 1695 2119 1721
rect 3817 1695 3823 1721
rect 3849 1695 3855 1721
rect 11657 1695 11663 1721
rect 11689 1695 11695 1721
rect 13617 1695 13623 1721
rect 13649 1695 13655 1721
rect 14737 1695 14743 1721
rect 14769 1695 14775 1721
rect 672 1581 19320 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 19320 1581
rect 672 1538 19320 1555
<< via1 >>
rect 9919 28211 9945 28237
rect 9971 28211 9997 28237
rect 10023 28211 10049 28237
rect 2239 27819 2265 27845
rect 2291 27819 2317 27845
rect 2343 27819 2369 27845
rect 17599 27819 17625 27845
rect 17651 27819 17677 27845
rect 17703 27819 17729 27845
rect 9919 27427 9945 27453
rect 9971 27427 9997 27453
rect 10023 27427 10049 27453
rect 2239 27035 2265 27061
rect 2291 27035 2317 27061
rect 2343 27035 2369 27061
rect 17599 27035 17625 27061
rect 17651 27035 17677 27061
rect 17703 27035 17729 27061
rect 3375 26839 3401 26865
rect 3823 26839 3849 26865
rect 4495 26839 4521 26865
rect 9919 26643 9945 26669
rect 9971 26643 9997 26669
rect 10023 26643 10049 26669
rect 4495 26503 4521 26529
rect 5839 26503 5865 26529
rect 3319 26447 3345 26473
rect 4495 26447 4521 26473
rect 5167 26447 5193 26473
rect 5727 26447 5753 26473
rect 2239 26251 2265 26277
rect 2291 26251 2317 26277
rect 2343 26251 2369 26277
rect 17599 26251 17625 26277
rect 17651 26251 17677 26277
rect 17703 26251 17729 26277
rect 3095 26055 3121 26081
rect 3543 26055 3569 26081
rect 3767 26055 3793 26081
rect 4831 26055 4857 26081
rect 5727 26055 5753 26081
rect 5727 25999 5753 26025
rect 9919 25859 9945 25885
rect 9971 25859 9997 25885
rect 10023 25859 10049 25885
rect 2815 25719 2841 25745
rect 5839 25719 5865 25745
rect 1639 25663 1665 25689
rect 2815 25663 2841 25689
rect 3095 25663 3121 25689
rect 3543 25663 3569 25689
rect 3767 25663 3793 25689
rect 5167 25663 5193 25689
rect 5727 25663 5753 25689
rect 18551 25663 18577 25689
rect 18663 25663 18689 25689
rect 18831 25663 18857 25689
rect 2239 25467 2265 25493
rect 2291 25467 2317 25493
rect 2343 25467 2369 25493
rect 17599 25467 17625 25493
rect 17651 25467 17677 25493
rect 17703 25467 17729 25493
rect 1583 25271 1609 25297
rect 2479 25271 2505 25297
rect 3095 25271 3121 25297
rect 3543 25271 3569 25297
rect 3767 25271 3793 25297
rect 4887 25271 4913 25297
rect 5783 25271 5809 25297
rect 7127 25271 7153 25297
rect 8023 25271 8049 25297
rect 18775 25271 18801 25297
rect 18887 25271 18913 25297
rect 19055 25271 19081 25297
rect 2479 25215 2505 25241
rect 5783 25215 5809 25241
rect 8023 25215 8049 25241
rect 18103 25215 18129 25241
rect 18215 25215 18241 25241
rect 18383 25215 18409 25241
rect 9919 25075 9945 25101
rect 9971 25075 9997 25101
rect 10023 25075 10049 25101
rect 5839 24935 5865 24961
rect 7519 24935 7545 24961
rect 17823 24935 17849 24961
rect 17991 24935 18017 24961
rect 18383 24935 18409 24961
rect 18551 24935 18577 24961
rect 1639 24879 1665 24905
rect 2087 24879 2113 24905
rect 2311 24879 2337 24905
rect 3095 24879 3121 24905
rect 3543 24879 3569 24905
rect 3767 24879 3793 24905
rect 4887 24879 4913 24905
rect 5839 24879 5865 24905
rect 6623 24879 6649 24905
rect 7519 24879 7545 24905
rect 17711 24879 17737 24905
rect 18327 24879 18353 24905
rect 2239 24683 2265 24709
rect 2291 24683 2317 24709
rect 2343 24683 2369 24709
rect 17599 24683 17625 24709
rect 17651 24683 17677 24709
rect 17703 24683 17729 24709
rect 1583 24487 1609 24513
rect 2143 24487 2169 24513
rect 3095 24487 3121 24513
rect 3543 24487 3569 24513
rect 3767 24487 3793 24513
rect 4887 24487 4913 24513
rect 5783 24487 5809 24513
rect 7071 24487 7097 24513
rect 7967 24487 7993 24513
rect 8583 24487 8609 24513
rect 9479 24487 9505 24513
rect 17151 24487 17177 24513
rect 17319 24487 17345 24513
rect 17543 24487 17569 24513
rect 17711 24487 17737 24513
rect 17879 24487 17905 24513
rect 18271 24487 18297 24513
rect 18439 24487 18465 24513
rect 18775 24487 18801 24513
rect 18887 24487 18913 24513
rect 18999 24487 19025 24513
rect 2255 24431 2281 24457
rect 5783 24431 5809 24457
rect 7967 24431 7993 24457
rect 9479 24431 9505 24457
rect 16983 24431 17009 24457
rect 18103 24431 18129 24457
rect 9919 24291 9945 24317
rect 9971 24291 9997 24317
rect 10023 24291 10049 24317
rect 5839 24151 5865 24177
rect 7519 24151 7545 24177
rect 9815 24151 9841 24177
rect 17263 24151 17289 24177
rect 17431 24151 17457 24177
rect 17711 24151 17737 24177
rect 17823 24151 17849 24177
rect 17991 24151 18017 24177
rect 18383 24151 18409 24177
rect 18551 24151 18577 24177
rect 1863 24095 1889 24121
rect 2311 24095 2337 24121
rect 2535 24095 2561 24121
rect 3319 24095 3345 24121
rect 3767 24095 3793 24121
rect 3991 24095 4017 24121
rect 5167 24095 5193 24121
rect 5839 24095 5865 24121
rect 6343 24095 6369 24121
rect 7519 24095 7545 24121
rect 9143 24095 9169 24121
rect 9815 24095 9841 24121
rect 17207 24095 17233 24121
rect 18327 24095 18353 24121
rect 2239 23899 2265 23925
rect 2291 23899 2317 23925
rect 2343 23899 2369 23925
rect 17599 23899 17625 23925
rect 17651 23899 17677 23925
rect 17703 23899 17729 23925
rect 1583 23703 1609 23729
rect 2479 23703 2505 23729
rect 3151 23703 3177 23729
rect 3599 23703 3625 23729
rect 3823 23703 3849 23729
rect 4887 23703 4913 23729
rect 5783 23703 5809 23729
rect 7127 23703 7153 23729
rect 8023 23703 8049 23729
rect 8583 23703 8609 23729
rect 9423 23703 9449 23729
rect 16479 23703 16505 23729
rect 16591 23703 16617 23729
rect 16759 23703 16785 23729
rect 17039 23703 17065 23729
rect 17151 23703 17177 23729
rect 17263 23703 17289 23729
rect 17599 23703 17625 23729
rect 17711 23703 17737 23729
rect 17879 23703 17905 23729
rect 18159 23703 18185 23729
rect 18383 23703 18409 23729
rect 18719 23703 18745 23729
rect 18999 23703 19025 23729
rect 2479 23647 2505 23673
rect 5783 23647 5809 23673
rect 8023 23647 8049 23673
rect 9423 23647 9449 23673
rect 18215 23647 18241 23673
rect 18943 23647 18969 23673
rect 9919 23507 9945 23533
rect 9971 23507 9997 23533
rect 10023 23507 10049 23533
rect 4439 23367 4465 23393
rect 8191 23367 8217 23393
rect 11495 23367 11521 23393
rect 17431 23367 17457 23393
rect 17711 23367 17737 23393
rect 17991 23367 18017 23393
rect 18383 23367 18409 23393
rect 18551 23367 18577 23393
rect 1919 23311 1945 23337
rect 2423 23311 2449 23337
rect 2535 23311 2561 23337
rect 3599 23311 3625 23337
rect 4439 23311 4465 23337
rect 6063 23311 6089 23337
rect 6343 23311 6369 23337
rect 6455 23311 6481 23337
rect 7239 23311 7265 23337
rect 8023 23311 8049 23337
rect 9087 23311 9113 23337
rect 9423 23311 9449 23337
rect 9535 23311 9561 23337
rect 10599 23311 10625 23337
rect 11495 23311 11521 23337
rect 16199 23311 16225 23337
rect 16311 23311 16337 23337
rect 16479 23311 16505 23337
rect 17207 23311 17233 23337
rect 17319 23311 17345 23337
rect 17879 23311 17905 23337
rect 18327 23311 18353 23337
rect 2239 23115 2265 23141
rect 2291 23115 2317 23141
rect 2343 23115 2369 23141
rect 17599 23115 17625 23141
rect 17651 23115 17677 23141
rect 17703 23115 17729 23141
rect 1415 22919 1441 22945
rect 2479 22919 2505 22945
rect 3935 22919 3961 22945
rect 4383 22919 4409 22945
rect 4495 22919 4521 22945
rect 5279 22919 5305 22945
rect 6343 22919 6369 22945
rect 7127 22919 7153 22945
rect 8023 22919 8049 22945
rect 8415 22919 8441 22945
rect 9479 22919 9505 22945
rect 11103 22919 11129 22945
rect 11383 22919 11409 22945
rect 11495 22919 11521 22945
rect 16199 22919 16225 22945
rect 16423 22919 16449 22945
rect 16535 22919 16561 22945
rect 16703 22919 16729 22945
rect 17039 22919 17065 22945
rect 17151 22919 17177 22945
rect 17319 22919 17345 22945
rect 17543 22919 17569 22945
rect 17711 22919 17737 22945
rect 17879 22919 17905 22945
rect 18159 22919 18185 22945
rect 18271 22919 18297 22945
rect 18383 22919 18409 22945
rect 18775 22919 18801 22945
rect 18887 22919 18913 22945
rect 2479 22863 2505 22889
rect 6343 22863 6369 22889
rect 8023 22863 8049 22889
rect 9479 22863 9505 22889
rect 15303 22863 15329 22889
rect 15471 22863 15497 22889
rect 15583 22863 15609 22889
rect 15863 22863 15889 22889
rect 15975 22863 16001 22889
rect 19055 22863 19081 22889
rect 9919 22723 9945 22749
rect 9971 22723 9997 22749
rect 10023 22723 10049 22749
rect 4439 22583 4465 22609
rect 8359 22583 8385 22609
rect 9815 22583 9841 22609
rect 11271 22583 11297 22609
rect 15583 22583 15609 22609
rect 15751 22583 15777 22609
rect 16143 22583 16169 22609
rect 16871 22583 16897 22609
rect 17151 22583 17177 22609
rect 17711 22583 17737 22609
rect 18103 22583 18129 22609
rect 18271 22583 18297 22609
rect 1919 22527 1945 22553
rect 2423 22527 2449 22553
rect 2535 22527 2561 22553
rect 3599 22527 3625 22553
rect 4439 22527 4465 22553
rect 6063 22527 6089 22553
rect 6343 22527 6369 22553
rect 6455 22527 6481 22553
rect 7463 22527 7489 22553
rect 8359 22527 8385 22553
rect 9143 22527 9169 22553
rect 9815 22527 9841 22553
rect 10375 22527 10401 22553
rect 11271 22527 11297 22553
rect 15863 22527 15889 22553
rect 16311 22527 16337 22553
rect 16479 22527 16505 22553
rect 17039 22527 17065 22553
rect 17487 22527 17513 22553
rect 17543 22527 17569 22553
rect 18047 22527 18073 22553
rect 18551 22527 18577 22553
rect 18719 22527 18745 22553
rect 18831 22527 18857 22553
rect 2239 22331 2265 22357
rect 2291 22331 2317 22357
rect 2343 22331 2369 22357
rect 17599 22331 17625 22357
rect 17651 22331 17677 22357
rect 17703 22331 17729 22357
rect 1415 22135 1441 22161
rect 2255 22135 2281 22161
rect 3935 22135 3961 22161
rect 4775 22135 4801 22161
rect 5279 22135 5305 22161
rect 6343 22135 6369 22161
rect 7127 22135 7153 22161
rect 7799 22135 7825 22161
rect 8415 22135 8441 22161
rect 9479 22135 9505 22161
rect 11103 22135 11129 22161
rect 11271 22135 11297 22161
rect 11495 22135 11521 22161
rect 12559 22135 12585 22161
rect 12839 22135 12865 22161
rect 12951 22135 12977 22161
rect 16423 22135 16449 22161
rect 16535 22135 16561 22161
rect 16703 22135 16729 22161
rect 16983 22135 17009 22161
rect 17151 22135 17177 22161
rect 17319 22135 17345 22161
rect 17487 22135 17513 22161
rect 18159 22135 18185 22161
rect 18271 22135 18297 22161
rect 18383 22135 18409 22161
rect 18887 22135 18913 22161
rect 2255 22079 2281 22105
rect 4775 22079 4801 22105
rect 6343 22079 6369 22105
rect 7799 22079 7825 22105
rect 9479 22079 9505 22105
rect 17711 22079 17737 22105
rect 17823 22079 17849 22105
rect 18775 22079 18801 22105
rect 19055 22079 19081 22105
rect 9919 21939 9945 21965
rect 9971 21939 9997 21965
rect 10023 21939 10049 21965
rect 3039 21799 3065 21825
rect 4271 21799 4297 21825
rect 9983 21799 10009 21825
rect 11495 21799 11521 21825
rect 18551 21799 18577 21825
rect 1863 21743 1889 21769
rect 3039 21743 3065 21769
rect 3375 21743 3401 21769
rect 4215 21743 4241 21769
rect 6063 21743 6089 21769
rect 6343 21743 6369 21769
rect 6455 21743 6481 21769
rect 7463 21743 7489 21769
rect 7687 21743 7713 21769
rect 7911 21743 7937 21769
rect 9143 21743 9169 21769
rect 9983 21743 10009 21769
rect 10599 21743 10625 21769
rect 11495 21743 11521 21769
rect 12839 21743 12865 21769
rect 13399 21743 13425 21769
rect 13567 21743 13593 21769
rect 16871 21743 16897 21769
rect 17039 21743 17065 21769
rect 17151 21743 17177 21769
rect 17487 21743 17513 21769
rect 17599 21743 17625 21769
rect 17711 21743 17737 21769
rect 18047 21743 18073 21769
rect 18159 21743 18185 21769
rect 18327 21743 18353 21769
rect 18719 21743 18745 21769
rect 18831 21743 18857 21769
rect 2239 21547 2265 21573
rect 2291 21547 2317 21573
rect 2343 21547 2369 21573
rect 17599 21547 17625 21573
rect 17651 21547 17677 21573
rect 17703 21547 17729 21573
rect 1583 21351 1609 21377
rect 2479 21351 2505 21377
rect 3823 21351 3849 21377
rect 4775 21351 4801 21377
rect 5279 21351 5305 21377
rect 6455 21351 6481 21377
rect 7127 21351 7153 21377
rect 7575 21351 7601 21377
rect 8583 21351 8609 21377
rect 8751 21351 8777 21377
rect 8975 21351 9001 21377
rect 11103 21351 11129 21377
rect 11383 21351 11409 21377
rect 11551 21351 11577 21377
rect 12559 21351 12585 21377
rect 12727 21351 12753 21377
rect 12951 21351 12977 21377
rect 16983 21351 17009 21377
rect 17151 21351 17177 21377
rect 17263 21351 17289 21377
rect 17543 21351 17569 21377
rect 17711 21351 17737 21377
rect 17879 21351 17905 21377
rect 18103 21351 18129 21377
rect 18887 21351 18913 21377
rect 18999 21351 19025 21377
rect 2479 21295 2505 21321
rect 4775 21295 4801 21321
rect 6455 21295 6481 21321
rect 7799 21295 7825 21321
rect 18215 21295 18241 21321
rect 18383 21295 18409 21321
rect 18775 21295 18801 21321
rect 9919 21155 9945 21181
rect 9971 21155 9997 21181
rect 10023 21155 10049 21181
rect 3039 21015 3065 21041
rect 4495 21015 4521 21041
rect 11327 21015 11353 21041
rect 17655 21015 17681 21041
rect 17767 21015 17793 21041
rect 17935 21015 17961 21041
rect 18215 21015 18241 21041
rect 18383 21015 18409 21041
rect 1863 20959 1889 20985
rect 3039 20959 3065 20985
rect 3375 20959 3401 20985
rect 4495 20959 4521 20985
rect 6063 20959 6089 20985
rect 6343 20959 6369 20985
rect 6455 20959 6481 20985
rect 7519 20959 7545 20985
rect 7687 20959 7713 20985
rect 7911 20959 7937 20985
rect 9143 20959 9169 20985
rect 9311 20959 9337 20985
rect 9535 20959 9561 20985
rect 10599 20959 10625 20985
rect 11327 20959 11353 20985
rect 13119 20959 13145 20985
rect 13287 20959 13313 20985
rect 13511 20959 13537 20985
rect 18495 20959 18521 20985
rect 18775 20959 18801 20985
rect 18887 20959 18913 20985
rect 18999 20959 19025 20985
rect 2239 20763 2265 20789
rect 2291 20763 2317 20789
rect 2343 20763 2369 20789
rect 17599 20763 17625 20789
rect 17651 20763 17677 20789
rect 17703 20763 17729 20789
rect 1583 20567 1609 20593
rect 2479 20567 2505 20593
rect 3823 20567 3849 20593
rect 4383 20567 4409 20593
rect 4495 20567 4521 20593
rect 5279 20567 5305 20593
rect 6455 20567 6481 20593
rect 7127 20567 7153 20593
rect 7575 20567 7601 20593
rect 8583 20567 8609 20593
rect 8751 20567 8777 20593
rect 8975 20567 9001 20593
rect 11103 20567 11129 20593
rect 11327 20567 11353 20593
rect 11495 20567 11521 20593
rect 12559 20567 12585 20593
rect 12727 20567 12753 20593
rect 12951 20567 12977 20593
rect 18103 20567 18129 20593
rect 18271 20567 18297 20593
rect 18439 20567 18465 20593
rect 18999 20567 19025 20593
rect 2479 20511 2505 20537
rect 6455 20511 6481 20537
rect 7799 20511 7825 20537
rect 18775 20511 18801 20537
rect 18943 20511 18969 20537
rect 9919 20371 9945 20397
rect 9971 20371 9997 20397
rect 10023 20371 10049 20397
rect 4439 20231 4465 20257
rect 11495 20231 11521 20257
rect 15247 20231 15273 20257
rect 1863 20175 1889 20201
rect 2423 20175 2449 20201
rect 2535 20175 2561 20201
rect 3375 20175 3401 20201
rect 4439 20175 4465 20201
rect 6063 20175 6089 20201
rect 6343 20175 6369 20201
rect 6455 20175 6481 20201
rect 7463 20175 7489 20201
rect 7687 20175 7713 20201
rect 7911 20175 7937 20201
rect 9143 20175 9169 20201
rect 9311 20175 9337 20201
rect 9535 20175 9561 20201
rect 10599 20175 10625 20201
rect 11495 20175 11521 20201
rect 13063 20175 13089 20201
rect 13287 20175 13313 20201
rect 13511 20175 13537 20201
rect 14575 20175 14601 20201
rect 15247 20175 15273 20201
rect 18719 20175 18745 20201
rect 18887 20175 18913 20201
rect 19055 20175 19081 20201
rect 2239 19979 2265 20005
rect 2291 19979 2317 20005
rect 2343 19979 2369 20005
rect 17599 19979 17625 20005
rect 17651 19979 17677 20005
rect 17703 19979 17729 20005
rect 1583 19783 1609 19809
rect 2423 19783 2449 19809
rect 3823 19783 3849 19809
rect 4383 19783 4409 19809
rect 4495 19783 4521 19809
rect 5279 19783 5305 19809
rect 6399 19783 6425 19809
rect 6959 19783 6985 19809
rect 7351 19783 7377 19809
rect 7575 19783 7601 19809
rect 8583 19783 8609 19809
rect 8751 19783 8777 19809
rect 8975 19783 9001 19809
rect 11103 19783 11129 19809
rect 11383 19783 11409 19809
rect 11495 19783 11521 19809
rect 12559 19783 12585 19809
rect 12727 19783 12753 19809
rect 12951 19783 12977 19809
rect 15079 19783 15105 19809
rect 15247 19783 15273 19809
rect 15471 19783 15497 19809
rect 18103 19783 18129 19809
rect 18271 19783 18297 19809
rect 2423 19727 2449 19753
rect 6399 19727 6425 19753
rect 18383 19727 18409 19753
rect 18775 19727 18801 19753
rect 18943 19727 18969 19753
rect 19055 19727 19081 19753
rect 9919 19587 9945 19613
rect 9971 19587 9997 19613
rect 10023 19587 10049 19613
rect 4439 19447 4465 19473
rect 6399 19447 6425 19473
rect 11495 19447 11521 19473
rect 15471 19447 15497 19473
rect 18775 19447 18801 19473
rect 1863 19391 1889 19417
rect 2423 19391 2449 19417
rect 2535 19391 2561 19417
rect 3375 19391 3401 19417
rect 4439 19391 4465 19417
rect 5279 19391 5305 19417
rect 6399 19391 6425 19417
rect 6959 19391 6985 19417
rect 7239 19391 7265 19417
rect 7351 19391 7377 19417
rect 9143 19391 9169 19417
rect 9311 19391 9337 19417
rect 9535 19391 9561 19417
rect 10599 19391 10625 19417
rect 11495 19391 11521 19417
rect 13119 19391 13145 19417
rect 13399 19391 13425 19417
rect 13567 19391 13593 19417
rect 14575 19391 14601 19417
rect 15471 19391 15497 19417
rect 18943 19391 18969 19417
rect 19055 19391 19081 19417
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 1583 18999 1609 19025
rect 2479 18999 2505 19025
rect 3823 18999 3849 19025
rect 4383 18999 4409 19025
rect 4495 18999 4521 19025
rect 5279 18999 5305 19025
rect 6399 18999 6425 19025
rect 7127 18999 7153 19025
rect 7351 18999 7377 19025
rect 7575 18999 7601 19025
rect 8415 18999 8441 19025
rect 8751 18999 8777 19025
rect 8975 18999 9001 19025
rect 11103 18999 11129 19025
rect 11383 18999 11409 19025
rect 11495 18999 11521 19025
rect 12559 18999 12585 19025
rect 13399 18999 13425 19025
rect 14855 18999 14881 19025
rect 15919 18999 15945 19025
rect 16255 18999 16281 19025
rect 16815 18999 16841 19025
rect 16927 18999 16953 19025
rect 2479 18943 2505 18969
rect 6399 18943 6425 18969
rect 13399 18943 13425 18969
rect 15919 18943 15945 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 3039 18663 3065 18689
rect 4439 18663 4465 18689
rect 6399 18663 6425 18689
rect 11495 18663 11521 18689
rect 15247 18663 15273 18689
rect 17991 18663 18017 18689
rect 1863 18607 1889 18633
rect 3039 18607 3065 18633
rect 3375 18607 3401 18633
rect 4439 18607 4465 18633
rect 5279 18607 5305 18633
rect 6399 18607 6425 18633
rect 6959 18607 6985 18633
rect 7239 18607 7265 18633
rect 7351 18607 7377 18633
rect 8863 18607 8889 18633
rect 9311 18607 9337 18633
rect 9535 18607 9561 18633
rect 10599 18607 10625 18633
rect 11495 18607 11521 18633
rect 13119 18607 13145 18633
rect 13399 18607 13425 18633
rect 13511 18607 13537 18633
rect 14575 18607 14601 18633
rect 15247 18607 15273 18633
rect 17991 18607 18017 18633
rect 18775 18607 18801 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 1583 18215 1609 18241
rect 2479 18215 2505 18241
rect 3823 18215 3849 18241
rect 4383 18215 4409 18241
rect 4495 18215 4521 18241
rect 5279 18215 5305 18241
rect 6399 18215 6425 18241
rect 7127 18215 7153 18241
rect 7351 18215 7377 18241
rect 7575 18215 7601 18241
rect 8415 18215 8441 18241
rect 8751 18215 8777 18241
rect 8975 18215 9001 18241
rect 11103 18215 11129 18241
rect 11383 18215 11409 18241
rect 11495 18215 11521 18241
rect 12559 18215 12585 18241
rect 13399 18215 13425 18241
rect 14855 18215 14881 18241
rect 15919 18215 15945 18241
rect 16255 18215 16281 18241
rect 16759 18215 16785 18241
rect 16927 18215 16953 18241
rect 2479 18159 2505 18185
rect 6399 18159 6425 18185
rect 13399 18159 13425 18185
rect 15919 18159 15945 18185
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 3039 17879 3065 17905
rect 4439 17879 4465 17905
rect 6399 17879 6425 17905
rect 11495 17879 11521 17905
rect 15247 17879 15273 17905
rect 1863 17823 1889 17849
rect 3039 17823 3065 17849
rect 3375 17823 3401 17849
rect 4439 17823 4465 17849
rect 5279 17823 5305 17849
rect 6399 17823 6425 17849
rect 6959 17823 6985 17849
rect 7183 17823 7209 17849
rect 7351 17823 7377 17849
rect 8863 17823 8889 17849
rect 9311 17823 9337 17849
rect 9535 17823 9561 17849
rect 10599 17823 10625 17849
rect 11495 17823 11521 17849
rect 13119 17823 13145 17849
rect 13399 17823 13425 17849
rect 13511 17823 13537 17849
rect 14575 17823 14601 17849
rect 15247 17823 15273 17849
rect 16815 17823 16841 17849
rect 17263 17823 17289 17849
rect 17487 17823 17513 17849
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 1583 17431 1609 17457
rect 2423 17431 2449 17457
rect 3879 17431 3905 17457
rect 4383 17431 4409 17457
rect 4495 17431 4521 17457
rect 5279 17431 5305 17457
rect 6399 17431 6425 17457
rect 7127 17431 7153 17457
rect 7799 17431 7825 17457
rect 8415 17431 8441 17457
rect 9311 17431 9337 17457
rect 11103 17431 11129 17457
rect 11383 17431 11409 17457
rect 11495 17431 11521 17457
rect 12559 17431 12585 17457
rect 13399 17431 13425 17457
rect 14799 17431 14825 17457
rect 15247 17431 15273 17457
rect 15471 17431 15497 17457
rect 16255 17431 16281 17457
rect 17263 17431 17289 17457
rect 2423 17375 2449 17401
rect 6399 17375 6425 17401
rect 7799 17375 7825 17401
rect 9311 17375 9337 17401
rect 13399 17375 13425 17401
rect 17263 17375 17289 17401
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 4439 17095 4465 17121
rect 6399 17095 6425 17121
rect 7799 17095 7825 17121
rect 11271 17095 11297 17121
rect 15247 17095 15273 17121
rect 1863 17039 1889 17065
rect 2423 17039 2449 17065
rect 2591 17039 2617 17065
rect 3431 17039 3457 17065
rect 4439 17039 4465 17065
rect 5279 17039 5305 17065
rect 6399 17039 6425 17065
rect 6959 17039 6985 17065
rect 7799 17039 7825 17065
rect 8863 17039 8889 17065
rect 9311 17039 9337 17065
rect 9535 17039 9561 17065
rect 10599 17039 10625 17065
rect 11271 17039 11297 17065
rect 13119 17039 13145 17065
rect 13399 17039 13425 17065
rect 13511 17039 13537 17065
rect 14575 17039 14601 17065
rect 15247 17039 15273 17065
rect 16815 17039 16841 17065
rect 17263 17039 17289 17065
rect 17487 17039 17513 17065
rect 18775 17039 18801 17065
rect 18887 17039 18913 17065
rect 19055 17039 19081 17065
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 1583 16647 1609 16673
rect 2311 16647 2337 16673
rect 3879 16647 3905 16673
rect 4383 16647 4409 16673
rect 4495 16647 4521 16673
rect 5279 16647 5305 16673
rect 6399 16647 6425 16673
rect 7127 16647 7153 16673
rect 7799 16647 7825 16673
rect 8415 16647 8441 16673
rect 9311 16647 9337 16673
rect 10823 16647 10849 16673
rect 11271 16647 11297 16673
rect 11495 16647 11521 16673
rect 12559 16647 12585 16673
rect 13399 16647 13425 16673
rect 14799 16647 14825 16673
rect 15247 16647 15273 16673
rect 15471 16647 15497 16673
rect 16255 16647 16281 16673
rect 17263 16647 17289 16673
rect 18775 16647 18801 16673
rect 18887 16647 18913 16673
rect 2311 16591 2337 16617
rect 6399 16591 6425 16617
rect 7799 16591 7825 16617
rect 9311 16591 9337 16617
rect 13399 16591 13425 16617
rect 17263 16591 17289 16617
rect 19055 16591 19081 16617
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 4439 16311 4465 16337
rect 6399 16311 6425 16337
rect 7799 16311 7825 16337
rect 11271 16311 11297 16337
rect 15247 16311 15273 16337
rect 1863 16255 1889 16281
rect 2311 16255 2337 16281
rect 2535 16255 2561 16281
rect 3431 16255 3457 16281
rect 4439 16255 4465 16281
rect 5279 16255 5305 16281
rect 6399 16255 6425 16281
rect 6959 16255 6985 16281
rect 7799 16255 7825 16281
rect 8863 16255 8889 16281
rect 9311 16255 9337 16281
rect 9535 16255 9561 16281
rect 10599 16255 10625 16281
rect 11271 16255 11297 16281
rect 13119 16255 13145 16281
rect 13399 16255 13425 16281
rect 13511 16255 13537 16281
rect 14295 16255 14321 16281
rect 15247 16255 15273 16281
rect 16815 16255 16841 16281
rect 17263 16255 17289 16281
rect 17487 16255 17513 16281
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 1359 15863 1385 15889
rect 2479 15863 2505 15889
rect 4047 15863 4073 15889
rect 4271 15863 4297 15889
rect 4495 15863 4521 15889
rect 5279 15863 5305 15889
rect 6175 15863 6201 15889
rect 7127 15863 7153 15889
rect 7631 15863 7657 15889
rect 8415 15863 8441 15889
rect 8807 15863 8833 15889
rect 8975 15863 9001 15889
rect 10823 15863 10849 15889
rect 11495 15863 11521 15889
rect 12279 15863 12305 15889
rect 12727 15863 12753 15889
rect 12951 15863 12977 15889
rect 14799 15863 14825 15889
rect 15247 15863 15273 15889
rect 15471 15863 15497 15889
rect 16255 15863 16281 15889
rect 16815 15863 16841 15889
rect 16927 15863 16953 15889
rect 2479 15807 2505 15833
rect 6231 15807 6257 15833
rect 7799 15807 7825 15833
rect 11775 15807 11801 15833
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 4495 15527 4521 15553
rect 6175 15527 6201 15553
rect 7631 15527 7657 15553
rect 11439 15527 11465 15553
rect 15303 15527 15329 15553
rect 1863 15471 1889 15497
rect 2423 15471 2449 15497
rect 2535 15471 2561 15497
rect 3599 15471 3625 15497
rect 4495 15471 4521 15497
rect 5279 15471 5305 15497
rect 6175 15471 6201 15497
rect 6959 15471 6985 15497
rect 7631 15471 7657 15497
rect 8863 15471 8889 15497
rect 9311 15471 9337 15497
rect 9535 15471 9561 15497
rect 10375 15471 10401 15497
rect 11439 15471 11465 15497
rect 12839 15471 12865 15497
rect 13399 15471 13425 15497
rect 13511 15471 13537 15497
rect 14295 15471 14321 15497
rect 15191 15471 15217 15497
rect 16815 15471 16841 15497
rect 17263 15471 17289 15497
rect 17487 15471 17513 15497
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 1359 15079 1385 15105
rect 2479 15079 2505 15105
rect 4047 15079 4073 15105
rect 4383 15079 4409 15105
rect 4495 15079 4521 15105
rect 5279 15079 5305 15105
rect 6175 15079 6201 15105
rect 6959 15079 6985 15105
rect 7631 15079 7657 15105
rect 8415 15079 8441 15105
rect 8807 15079 8833 15105
rect 8975 15079 9001 15105
rect 10823 15079 10849 15105
rect 11495 15079 11521 15105
rect 12279 15079 12305 15105
rect 13343 15079 13369 15105
rect 14799 15079 14825 15105
rect 15247 15079 15273 15105
rect 15471 15079 15497 15105
rect 16535 15079 16561 15105
rect 17263 15079 17289 15105
rect 2479 15023 2505 15049
rect 6231 15023 6257 15049
rect 7799 15023 7825 15049
rect 11775 15023 11801 15049
rect 13343 15023 13369 15049
rect 17263 15023 17289 15049
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 4495 14743 4521 14769
rect 6175 14743 6201 14769
rect 7631 14743 7657 14769
rect 11439 14743 11465 14769
rect 15247 14743 15273 14769
rect 1863 14687 1889 14713
rect 2423 14687 2449 14713
rect 2535 14687 2561 14713
rect 3599 14687 3625 14713
rect 4495 14687 4521 14713
rect 5223 14687 5249 14713
rect 5951 14687 5977 14713
rect 6959 14687 6985 14713
rect 7631 14687 7657 14713
rect 8863 14687 8889 14713
rect 9311 14687 9337 14713
rect 9535 14687 9561 14713
rect 10375 14687 10401 14713
rect 11439 14687 11465 14713
rect 12839 14687 12865 14713
rect 13399 14687 13425 14713
rect 13511 14687 13537 14713
rect 14295 14687 14321 14713
rect 15247 14687 15273 14713
rect 16815 14687 16841 14713
rect 17263 14687 17289 14713
rect 17487 14687 17513 14713
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 1359 14295 1385 14321
rect 2479 14295 2505 14321
rect 4047 14295 4073 14321
rect 4383 14295 4409 14321
rect 4495 14295 4521 14321
rect 5279 14295 5305 14321
rect 5839 14295 5865 14321
rect 5951 14295 5977 14321
rect 6959 14295 6985 14321
rect 7631 14295 7657 14321
rect 8415 14295 8441 14321
rect 8807 14295 8833 14321
rect 8975 14295 9001 14321
rect 10823 14295 10849 14321
rect 11495 14295 11521 14321
rect 12279 14295 12305 14321
rect 13399 14295 13425 14321
rect 14799 14295 14825 14321
rect 15247 14295 15273 14321
rect 15471 14295 15497 14321
rect 16535 14295 16561 14321
rect 17263 14295 17289 14321
rect 2479 14239 2505 14265
rect 7799 14239 7825 14265
rect 11775 14239 11801 14265
rect 13399 14239 13425 14265
rect 17263 14239 17289 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 4495 13959 4521 13985
rect 7631 13959 7657 13985
rect 11495 13959 11521 13985
rect 15247 13959 15273 13985
rect 1863 13903 1889 13929
rect 2423 13903 2449 13929
rect 2591 13903 2617 13929
rect 3599 13903 3625 13929
rect 4495 13903 4521 13929
rect 5223 13903 5249 13929
rect 5783 13903 5809 13929
rect 5895 13903 5921 13929
rect 6959 13903 6985 13929
rect 7631 13903 7657 13929
rect 8863 13903 8889 13929
rect 9311 13903 9337 13929
rect 9535 13903 9561 13929
rect 10375 13903 10401 13929
rect 11495 13903 11521 13929
rect 12839 13903 12865 13929
rect 13399 13903 13425 13929
rect 13511 13903 13537 13929
rect 14295 13903 14321 13929
rect 15247 13903 15273 13929
rect 16815 13903 16841 13929
rect 17263 13903 17289 13929
rect 17487 13903 17513 13929
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 1359 13511 1385 13537
rect 2143 13511 2169 13537
rect 4047 13511 4073 13537
rect 4383 13511 4409 13537
rect 4495 13511 4521 13537
rect 5279 13511 5305 13537
rect 5839 13511 5865 13537
rect 5951 13511 5977 13537
rect 6959 13511 6985 13537
rect 7631 13511 7657 13537
rect 8415 13511 8441 13537
rect 8807 13511 8833 13537
rect 8975 13511 9001 13537
rect 10823 13511 10849 13537
rect 11719 13511 11745 13537
rect 12279 13511 12305 13537
rect 13455 13511 13481 13537
rect 14799 13511 14825 13537
rect 15247 13511 15273 13537
rect 15471 13511 15497 13537
rect 16535 13511 16561 13537
rect 16815 13511 16841 13537
rect 16927 13511 16953 13537
rect 2255 13455 2281 13481
rect 7799 13455 7825 13481
rect 11775 13455 11801 13481
rect 13455 13455 13481 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 4495 13175 4521 13201
rect 7631 13175 7657 13201
rect 11495 13175 11521 13201
rect 15247 13175 15273 13201
rect 17879 13175 17905 13201
rect 1863 13119 1889 13145
rect 2311 13119 2337 13145
rect 2535 13119 2561 13145
rect 3599 13119 3625 13145
rect 4495 13119 4521 13145
rect 5223 13119 5249 13145
rect 5783 13119 5809 13145
rect 5895 13119 5921 13145
rect 6959 13119 6985 13145
rect 7631 13119 7657 13145
rect 8863 13119 8889 13145
rect 9311 13119 9337 13145
rect 9535 13119 9561 13145
rect 10375 13119 10401 13145
rect 11495 13119 11521 13145
rect 12839 13119 12865 13145
rect 13399 13119 13425 13145
rect 13511 13119 13537 13145
rect 14295 13119 14321 13145
rect 15247 13119 15273 13145
rect 17879 13119 17905 13145
rect 19055 13119 19081 13145
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 1359 12727 1385 12753
rect 2479 12727 2505 12753
rect 4047 12727 4073 12753
rect 4383 12727 4409 12753
rect 4495 12727 4521 12753
rect 5279 12727 5305 12753
rect 5839 12727 5865 12753
rect 5951 12727 5977 12753
rect 6959 12727 6985 12753
rect 7631 12727 7657 12753
rect 8415 12727 8441 12753
rect 8807 12727 8833 12753
rect 8975 12727 9001 12753
rect 10935 12727 10961 12753
rect 11719 12727 11745 12753
rect 12279 12727 12305 12753
rect 13455 12727 13481 12753
rect 14799 12727 14825 12753
rect 15247 12727 15273 12753
rect 15471 12727 15497 12753
rect 16255 12727 16281 12753
rect 16815 12727 16841 12753
rect 16927 12727 16953 12753
rect 2479 12671 2505 12697
rect 7799 12671 7825 12697
rect 11775 12671 11801 12697
rect 13455 12671 13481 12697
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 6175 12391 6201 12417
rect 7631 12391 7657 12417
rect 11495 12391 11521 12417
rect 15247 12391 15273 12417
rect 17879 12391 17905 12417
rect 1863 12335 1889 12361
rect 2423 12335 2449 12361
rect 2535 12335 2561 12361
rect 3599 12335 3625 12361
rect 3767 12335 3793 12361
rect 3991 12335 4017 12361
rect 5223 12335 5249 12361
rect 5951 12335 5977 12361
rect 6959 12335 6985 12361
rect 7575 12335 7601 12361
rect 8863 12335 8889 12361
rect 9311 12335 9337 12361
rect 9535 12335 9561 12361
rect 10319 12335 10345 12361
rect 11495 12335 11521 12361
rect 12839 12335 12865 12361
rect 13399 12335 13425 12361
rect 13511 12335 13537 12361
rect 14295 12335 14321 12361
rect 15247 12335 15273 12361
rect 17879 12335 17905 12361
rect 19055 12335 19081 12361
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 1359 11943 1385 11969
rect 2479 11943 2505 11969
rect 4103 11943 4129 11969
rect 4775 11943 4801 11969
rect 5279 11943 5305 11969
rect 5839 11943 5865 11969
rect 5951 11943 5977 11969
rect 6959 11943 6985 11969
rect 7575 11943 7601 11969
rect 8415 11943 8441 11969
rect 8751 11943 8777 11969
rect 8975 11943 9001 11969
rect 10935 11943 10961 11969
rect 11383 11943 11409 11969
rect 11495 11943 11521 11969
rect 12279 11943 12305 11969
rect 13399 11943 13425 11969
rect 15079 11943 15105 11969
rect 15247 11943 15273 11969
rect 15471 11943 15497 11969
rect 17487 11943 17513 11969
rect 17767 11943 17793 11969
rect 17879 11943 17905 11969
rect 2479 11887 2505 11913
rect 4775 11887 4801 11913
rect 7799 11887 7825 11913
rect 13399 11887 13425 11913
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 6175 11607 6201 11633
rect 7631 11607 7657 11633
rect 11495 11607 11521 11633
rect 15247 11607 15273 11633
rect 17879 11607 17905 11633
rect 1863 11551 1889 11577
rect 2423 11551 2449 11577
rect 2535 11551 2561 11577
rect 3319 11551 3345 11577
rect 3879 11551 3905 11577
rect 3991 11551 4017 11577
rect 5223 11551 5249 11577
rect 5951 11551 5977 11577
rect 6959 11551 6985 11577
rect 7575 11551 7601 11577
rect 9031 11551 9057 11577
rect 9311 11551 9337 11577
rect 9535 11551 9561 11577
rect 10319 11551 10345 11577
rect 11495 11551 11521 11577
rect 12839 11551 12865 11577
rect 13399 11551 13425 11577
rect 13511 11551 13537 11577
rect 14575 11551 14601 11577
rect 15135 11551 15161 11577
rect 17879 11551 17905 11577
rect 19055 11551 19081 11577
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 1415 11159 1441 11185
rect 2479 11159 2505 11185
rect 3319 11159 3345 11185
rect 3991 11159 4017 11185
rect 4663 11159 4689 11185
rect 5055 11159 5081 11185
rect 5279 11159 5305 11185
rect 6959 11159 6985 11185
rect 7575 11159 7601 11185
rect 8415 11159 8441 11185
rect 8751 11159 8777 11185
rect 8975 11159 9001 11185
rect 10823 11159 10849 11185
rect 11383 11159 11409 11185
rect 11495 11159 11521 11185
rect 12279 11159 12305 11185
rect 13455 11159 13481 11185
rect 15975 11159 16001 11185
rect 16927 11159 16953 11185
rect 17487 11159 17513 11185
rect 17767 11159 17793 11185
rect 17879 11159 17905 11185
rect 2479 11103 2505 11129
rect 4103 11103 4129 11129
rect 7799 11103 7825 11129
rect 13455 11103 13481 11129
rect 15975 11103 16001 11129
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 5839 10823 5865 10849
rect 7799 10823 7825 10849
rect 9815 10823 9841 10849
rect 11495 10823 11521 10849
rect 15471 10823 15497 10849
rect 17879 10823 17905 10849
rect 1919 10767 1945 10793
rect 2423 10767 2449 10793
rect 2535 10767 2561 10793
rect 3375 10767 3401 10793
rect 3879 10767 3905 10793
rect 3991 10767 4017 10793
rect 4887 10767 4913 10793
rect 5839 10767 5865 10793
rect 6959 10767 6985 10793
rect 7799 10767 7825 10793
rect 9031 10767 9057 10793
rect 9759 10767 9785 10793
rect 10319 10767 10345 10793
rect 11495 10767 11521 10793
rect 12839 10767 12865 10793
rect 13399 10767 13425 10793
rect 13511 10767 13537 10793
rect 15471 10767 15497 10793
rect 16423 10767 16449 10793
rect 17879 10767 17905 10793
rect 19055 10767 19081 10793
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 1415 10375 1441 10401
rect 2479 10375 2505 10401
rect 3375 10375 3401 10401
rect 3767 10375 3793 10401
rect 3991 10375 4017 10401
rect 4663 10375 4689 10401
rect 5111 10375 5137 10401
rect 5839 10375 5865 10401
rect 6959 10375 6985 10401
rect 7799 10375 7825 10401
rect 8415 10375 8441 10401
rect 9255 10375 9281 10401
rect 10823 10375 10849 10401
rect 11383 10375 11409 10401
rect 11495 10375 11521 10401
rect 12279 10375 12305 10401
rect 13455 10375 13481 10401
rect 15751 10375 15777 10401
rect 16927 10375 16953 10401
rect 17487 10375 17513 10401
rect 17767 10375 17793 10401
rect 17879 10375 17905 10401
rect 2479 10319 2505 10345
rect 7799 10319 7825 10345
rect 9255 10319 9281 10345
rect 13455 10319 13481 10345
rect 15751 10319 15777 10345
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 3039 10039 3065 10065
rect 11271 10039 11297 10065
rect 17879 10039 17905 10065
rect 1919 9983 1945 10009
rect 3039 9983 3065 10009
rect 3375 9983 3401 10009
rect 3767 9983 3793 10009
rect 3991 9983 4017 10009
rect 4999 9983 5025 10009
rect 5447 9983 5473 10009
rect 5559 9983 5585 10009
rect 6343 9983 6369 10009
rect 6903 9983 6929 10009
rect 7015 9983 7041 10009
rect 9087 9983 9113 10009
rect 9311 9983 9337 10009
rect 9535 9983 9561 10009
rect 10319 9983 10345 10009
rect 11271 9983 11297 10009
rect 12839 9983 12865 10009
rect 13399 9983 13425 10009
rect 13511 9983 13537 10009
rect 15751 9983 15777 10009
rect 15975 9983 16001 10009
rect 16423 9983 16449 10009
rect 17879 9983 17905 10009
rect 18775 9983 18801 10009
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 1583 9591 1609 9617
rect 2479 9591 2505 9617
rect 3319 9591 3345 9617
rect 3655 9591 3681 9617
rect 3767 9591 3793 9617
rect 4943 9591 4969 9617
rect 5111 9591 5137 9617
rect 5559 9591 5585 9617
rect 6847 9591 6873 9617
rect 7295 9591 7321 9617
rect 7519 9591 7545 9617
rect 8415 9591 8441 9617
rect 8751 9591 8777 9617
rect 8975 9591 9001 9617
rect 10823 9591 10849 9617
rect 11271 9591 11297 9617
rect 11495 9591 11521 9617
rect 12559 9591 12585 9617
rect 13343 9591 13369 9617
rect 16255 9591 16281 9617
rect 16479 9591 16505 9617
rect 16759 9591 16785 9617
rect 17207 9591 17233 9617
rect 17767 9591 17793 9617
rect 17879 9591 17905 9617
rect 2479 9535 2505 9561
rect 13343 9535 13369 9561
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 2815 9255 2841 9281
rect 11271 9255 11297 9281
rect 17879 9255 17905 9281
rect 1919 9199 1945 9225
rect 2815 9199 2841 9225
rect 3319 9199 3345 9225
rect 3655 9199 3681 9225
rect 3767 9199 3793 9225
rect 4999 9199 5025 9225
rect 5447 9199 5473 9225
rect 5559 9199 5585 9225
rect 6343 9199 6369 9225
rect 6903 9199 6929 9225
rect 7015 9199 7041 9225
rect 9087 9199 9113 9225
rect 9311 9199 9337 9225
rect 9535 9199 9561 9225
rect 10319 9199 10345 9225
rect 10991 9199 11017 9225
rect 12839 9199 12865 9225
rect 13343 9199 13369 9225
rect 13511 9199 13537 9225
rect 14295 9199 14321 9225
rect 14743 9199 14769 9225
rect 14967 9199 14993 9225
rect 17879 9199 17905 9225
rect 18775 9199 18801 9225
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 1583 8807 1609 8833
rect 2479 8807 2505 8833
rect 3319 8807 3345 8833
rect 3655 8807 3681 8833
rect 3767 8807 3793 8833
rect 4943 8807 4969 8833
rect 5111 8807 5137 8833
rect 5559 8807 5585 8833
rect 6847 8807 6873 8833
rect 7295 8807 7321 8833
rect 7519 8807 7545 8833
rect 8415 8807 8441 8833
rect 8751 8807 8777 8833
rect 8975 8807 9001 8833
rect 11103 8807 11129 8833
rect 11271 8807 11297 8833
rect 11495 8807 11521 8833
rect 12279 8807 12305 8833
rect 13399 8807 13425 8833
rect 14799 8807 14825 8833
rect 15247 8807 15273 8833
rect 15471 8807 15497 8833
rect 17207 8807 17233 8833
rect 17767 8807 17793 8833
rect 17879 8807 17905 8833
rect 2479 8751 2505 8777
rect 13399 8751 13425 8777
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 2815 8471 2841 8497
rect 11271 8471 11297 8497
rect 15359 8471 15385 8497
rect 17879 8471 17905 8497
rect 1919 8415 1945 8441
rect 2815 8415 2841 8441
rect 3319 8415 3345 8441
rect 3655 8415 3681 8441
rect 3767 8415 3793 8441
rect 4999 8415 5025 8441
rect 5447 8415 5473 8441
rect 5559 8415 5585 8441
rect 6343 8415 6369 8441
rect 6903 8415 6929 8441
rect 7015 8415 7041 8441
rect 9087 8415 9113 8441
rect 9311 8415 9337 8441
rect 9535 8415 9561 8441
rect 10599 8415 10625 8441
rect 11271 8415 11297 8441
rect 12839 8415 12865 8441
rect 13399 8415 13425 8441
rect 13511 8415 13537 8441
rect 14295 8415 14321 8441
rect 15359 8415 15385 8441
rect 17879 8415 17905 8441
rect 18775 8415 18801 8441
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 1583 8023 1609 8049
rect 2479 8023 2505 8049
rect 3319 8023 3345 8049
rect 3655 8023 3681 8049
rect 3823 8023 3849 8049
rect 4999 8023 5025 8049
rect 5559 8023 5585 8049
rect 6847 8023 6873 8049
rect 7295 8023 7321 8049
rect 7519 8023 7545 8049
rect 8415 8023 8441 8049
rect 8751 8023 8777 8049
rect 8975 8023 9001 8049
rect 11103 8023 11129 8049
rect 11999 8023 12025 8049
rect 12279 8023 12305 8049
rect 13343 8023 13369 8049
rect 15191 8023 15217 8049
rect 15415 8023 15441 8049
rect 15695 8023 15721 8049
rect 17207 8023 17233 8049
rect 17767 8023 17793 8049
rect 17879 8023 17905 8049
rect 2479 7967 2505 7993
rect 5671 7967 5697 7993
rect 11999 7967 12025 7993
rect 13343 7967 13369 7993
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 3039 7687 3065 7713
rect 11495 7687 11521 7713
rect 15359 7687 15385 7713
rect 17879 7687 17905 7713
rect 2143 7631 2169 7657
rect 3039 7631 3065 7657
rect 3599 7631 3625 7657
rect 3823 7631 3849 7657
rect 3991 7631 4017 7657
rect 4999 7631 5025 7657
rect 5447 7631 5473 7657
rect 5559 7631 5585 7657
rect 6343 7631 6369 7657
rect 6903 7631 6929 7657
rect 7015 7631 7041 7657
rect 9087 7631 9113 7657
rect 9311 7631 9337 7657
rect 9535 7631 9561 7657
rect 10599 7631 10625 7657
rect 11495 7631 11521 7657
rect 12839 7631 12865 7657
rect 13399 7631 13425 7657
rect 13511 7631 13537 7657
rect 14295 7631 14321 7657
rect 15359 7631 15385 7657
rect 17879 7631 17905 7657
rect 18775 7631 18801 7657
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 1583 7239 1609 7265
rect 2479 7239 2505 7265
rect 3543 7239 3569 7265
rect 3823 7239 3849 7265
rect 3935 7239 3961 7265
rect 4999 7239 5025 7265
rect 5559 7239 5585 7265
rect 6847 7239 6873 7265
rect 7295 7239 7321 7265
rect 7519 7239 7545 7265
rect 8415 7239 8441 7265
rect 8751 7239 8777 7265
rect 8975 7239 9001 7265
rect 11103 7239 11129 7265
rect 11999 7239 12025 7265
rect 12279 7239 12305 7265
rect 13399 7239 13425 7265
rect 14799 7239 14825 7265
rect 15247 7239 15273 7265
rect 15471 7239 15497 7265
rect 16255 7239 16281 7265
rect 17151 7239 17177 7265
rect 2479 7183 2505 7209
rect 5671 7183 5697 7209
rect 11999 7183 12025 7209
rect 13399 7183 13425 7209
rect 16255 7183 16281 7209
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 10991 6903 11017 6929
rect 12447 6903 12473 6929
rect 14015 6903 14041 6929
rect 15247 6903 15273 6929
rect 17879 6903 17905 6929
rect 2087 6847 2113 6873
rect 2423 6847 2449 6873
rect 2535 6847 2561 6873
rect 3543 6847 3569 6873
rect 3823 6847 3849 6873
rect 3991 6847 4017 6873
rect 4999 6847 5025 6873
rect 5447 6847 5473 6873
rect 5559 6847 5585 6873
rect 6343 6847 6369 6873
rect 6903 6847 6929 6873
rect 7015 6847 7041 6873
rect 9815 6847 9841 6873
rect 10991 6847 11017 6873
rect 11271 6847 11297 6873
rect 12447 6847 12473 6873
rect 12839 6847 12865 6873
rect 14015 6847 14041 6873
rect 14295 6847 14321 6873
rect 15247 6847 15273 6873
rect 17879 6847 17905 6873
rect 18775 6847 18801 6873
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 1583 6455 1609 6481
rect 2423 6455 2449 6481
rect 3543 6455 3569 6481
rect 3823 6455 3849 6481
rect 3935 6455 3961 6481
rect 4999 6455 5025 6481
rect 5559 6455 5585 6481
rect 6847 6455 6873 6481
rect 7295 6455 7321 6481
rect 7519 6455 7545 6481
rect 9535 6455 9561 6481
rect 10431 6455 10457 6481
rect 11103 6455 11129 6481
rect 11999 6455 12025 6481
rect 12279 6455 12305 6481
rect 13399 6455 13425 6481
rect 15247 6455 15273 6481
rect 15415 6455 15441 6481
rect 15695 6455 15721 6481
rect 17207 6455 17233 6481
rect 17991 6455 18017 6481
rect 2423 6399 2449 6425
rect 5671 6399 5697 6425
rect 10431 6399 10457 6425
rect 11999 6399 12025 6425
rect 13399 6399 13425 6425
rect 18159 6399 18185 6425
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2423 6119 2449 6145
rect 10991 6119 11017 6145
rect 12447 6119 12473 6145
rect 15247 6119 15273 6145
rect 18103 6119 18129 6145
rect 1639 6063 1665 6089
rect 2423 6063 2449 6089
rect 3543 6063 3569 6089
rect 3879 6063 3905 6089
rect 3991 6063 4017 6089
rect 4999 6063 5025 6089
rect 5447 6063 5473 6089
rect 5559 6063 5585 6089
rect 6343 6063 6369 6089
rect 6791 6063 6817 6089
rect 7015 6063 7041 6089
rect 9815 6063 9841 6089
rect 10991 6063 11017 6089
rect 11271 6063 11297 6089
rect 12447 6063 12473 6089
rect 12839 6063 12865 6089
rect 13399 6063 13425 6089
rect 13511 6063 13537 6089
rect 14575 6063 14601 6089
rect 15247 6063 15273 6089
rect 18103 6063 18129 6089
rect 18775 6063 18801 6089
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 1583 5671 1609 5697
rect 2423 5671 2449 5697
rect 2871 5671 2897 5697
rect 3375 5671 3401 5697
rect 3543 5671 3569 5697
rect 4999 5671 5025 5697
rect 5559 5671 5585 5697
rect 8303 5671 8329 5697
rect 8415 5671 8441 5697
rect 8975 5671 9001 5697
rect 9535 5671 9561 5697
rect 10431 5671 10457 5697
rect 11103 5671 11129 5697
rect 11999 5671 12025 5697
rect 12279 5671 12305 5697
rect 13399 5671 13425 5697
rect 14911 5671 14937 5697
rect 15975 5671 16001 5697
rect 16255 5671 16281 5697
rect 17151 5671 17177 5697
rect 2423 5615 2449 5641
rect 5671 5615 5697 5641
rect 10431 5615 10457 5641
rect 11999 5615 12025 5641
rect 13399 5615 13425 5641
rect 15975 5615 16001 5641
rect 16255 5615 16281 5641
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2423 5335 2449 5361
rect 8359 5335 8385 5361
rect 10991 5335 11017 5361
rect 12279 5335 12305 5361
rect 14015 5335 14041 5361
rect 15471 5335 15497 5361
rect 18103 5335 18129 5361
rect 1639 5279 1665 5305
rect 2423 5279 2449 5305
rect 2871 5279 2897 5305
rect 3431 5279 3457 5305
rect 3543 5279 3569 5305
rect 4999 5279 5025 5305
rect 5391 5279 5417 5305
rect 5559 5279 5585 5305
rect 7519 5279 7545 5305
rect 8359 5279 8385 5305
rect 10039 5279 10065 5305
rect 10991 5279 11017 5305
rect 11383 5279 11409 5305
rect 12279 5279 12305 5305
rect 13119 5279 13145 5305
rect 14015 5279 14041 5305
rect 14575 5279 14601 5305
rect 15471 5279 15497 5305
rect 18103 5279 18129 5305
rect 18775 5279 18801 5305
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 1583 4887 1609 4913
rect 2423 4887 2449 4913
rect 2871 4887 2897 4913
rect 3431 4887 3457 4913
rect 3543 4887 3569 4913
rect 4999 4887 5025 4913
rect 5167 4887 5193 4913
rect 5391 4887 5417 4913
rect 7799 4887 7825 4913
rect 8359 4887 8385 4913
rect 8471 4887 8497 4913
rect 9535 4887 9561 4913
rect 10431 4887 10457 4913
rect 11103 4887 11129 4913
rect 11999 4887 12025 4913
rect 12559 4887 12585 4913
rect 13399 4887 13425 4913
rect 14855 4887 14881 4913
rect 15919 4887 15945 4913
rect 17711 4887 17737 4913
rect 17935 4887 17961 4913
rect 18383 4887 18409 4913
rect 2423 4831 2449 4857
rect 10431 4831 10457 4857
rect 11999 4831 12025 4857
rect 13399 4831 13425 4857
rect 14855 4831 14881 4857
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2423 4551 2449 4577
rect 6063 4551 6089 4577
rect 8471 4551 8497 4577
rect 10767 4551 10793 4577
rect 12279 4551 12305 4577
rect 14015 4551 14041 4577
rect 17991 4551 18017 4577
rect 1583 4495 1609 4521
rect 2423 4495 2449 4521
rect 2871 4495 2897 4521
rect 3375 4495 3401 4521
rect 3543 4495 3569 4521
rect 6063 4495 6089 4521
rect 7015 4495 7041 4521
rect 7575 4495 7601 4521
rect 8471 4495 8497 4521
rect 10039 4495 10065 4521
rect 10767 4495 10793 4521
rect 11383 4495 11409 4521
rect 11999 4495 12025 4521
rect 13119 4495 13145 4521
rect 14015 4495 14041 4521
rect 14575 4495 14601 4521
rect 14855 4495 14881 4521
rect 14967 4495 14993 4521
rect 17991 4495 18017 4521
rect 18775 4495 18801 4521
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 911 4103 937 4129
rect 2087 4103 2113 4129
rect 3879 4103 3905 4129
rect 4999 4103 5025 4129
rect 5783 4103 5809 4129
rect 6007 4103 6033 4129
rect 6455 4103 6481 4129
rect 7799 4103 7825 4129
rect 8471 4103 8497 4129
rect 9535 4103 9561 4129
rect 10431 4103 10457 4129
rect 11103 4103 11129 4129
rect 11775 4103 11801 4129
rect 12559 4103 12585 4129
rect 13231 4103 13257 4129
rect 16255 4103 16281 4129
rect 16479 4103 16505 4129
rect 16759 4103 16785 4129
rect 17711 4103 17737 4129
rect 17879 4103 17905 4129
rect 18383 4103 18409 4129
rect 2087 4047 2113 4073
rect 3879 4047 3905 4073
rect 8751 4047 8777 4073
rect 10431 4047 10457 4073
rect 11775 4047 11801 4073
rect 13231 4047 13257 4073
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2087 3767 2113 3793
rect 8359 3767 8385 3793
rect 12447 3767 12473 3793
rect 15415 3767 15441 3793
rect 17879 3767 17905 3793
rect 911 3711 937 3737
rect 2087 3711 2113 3737
rect 3823 3711 3849 3737
rect 4047 3711 4073 3737
rect 4495 3711 4521 3737
rect 6343 3711 6369 3737
rect 6567 3711 6593 3737
rect 7015 3711 7041 3737
rect 7519 3711 7545 3737
rect 8359 3711 8385 3737
rect 9815 3711 9841 3737
rect 10375 3711 10401 3737
rect 10487 3711 10513 3737
rect 11551 3711 11577 3737
rect 12447 3711 12473 3737
rect 13119 3711 13145 3737
rect 13287 3711 13313 3737
rect 13567 3711 13593 3737
rect 14519 3711 14545 3737
rect 15359 3711 15385 3737
rect 17879 3711 17905 3737
rect 18831 3711 18857 3737
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 911 3319 937 3345
rect 2087 3319 2113 3345
rect 3823 3319 3849 3345
rect 4999 3319 5025 3345
rect 5559 3319 5585 3345
rect 5839 3319 5865 3345
rect 5951 3319 5977 3345
rect 7799 3319 7825 3345
rect 8807 3319 8833 3345
rect 9255 3319 9281 3345
rect 9759 3319 9785 3345
rect 9927 3319 9953 3345
rect 11103 3319 11129 3345
rect 11383 3319 11409 3345
rect 11495 3319 11521 3345
rect 12559 3319 12585 3345
rect 12727 3319 12753 3345
rect 12951 3319 12977 3345
rect 16255 3319 16281 3345
rect 16367 3319 16393 3345
rect 16927 3319 16953 3345
rect 17711 3319 17737 3345
rect 17823 3319 17849 3345
rect 18383 3319 18409 3345
rect 2087 3263 2113 3289
rect 3823 3263 3849 3289
rect 8807 3263 8833 3289
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2031 2983 2057 3009
rect 11719 2983 11745 3009
rect 14015 2983 14041 3009
rect 15247 2983 15273 3009
rect 17991 2983 18017 3009
rect 911 2927 937 2953
rect 2031 2927 2057 2953
rect 3823 2927 3849 2953
rect 3935 2927 3961 2953
rect 4495 2927 4521 2953
rect 6119 2927 6145 2953
rect 6287 2927 6313 2953
rect 6511 2927 6537 2953
rect 7519 2927 7545 2953
rect 7743 2927 7769 2953
rect 7967 2927 7993 2953
rect 9311 2927 9337 2953
rect 9759 2927 9785 2953
rect 9983 2927 10009 2953
rect 11047 2927 11073 2953
rect 11663 2927 11689 2953
rect 13119 2927 13145 2953
rect 14015 2927 14041 2953
rect 14351 2927 14377 2953
rect 15135 2927 15161 2953
rect 17991 2927 18017 2953
rect 18775 2927 18801 2953
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 911 2535 937 2561
rect 2031 2535 2057 2561
rect 3991 2535 4017 2561
rect 4999 2535 5025 2561
rect 5559 2535 5585 2561
rect 6455 2535 6481 2561
rect 8079 2535 8105 2561
rect 8247 2535 8273 2561
rect 8471 2535 8497 2561
rect 9255 2535 9281 2561
rect 10431 2535 10457 2561
rect 11047 2535 11073 2561
rect 11663 2535 11689 2561
rect 12559 2535 12585 2561
rect 13455 2535 13481 2561
rect 14799 2535 14825 2561
rect 15247 2535 15273 2561
rect 15471 2535 15497 2561
rect 17487 2535 17513 2561
rect 17767 2535 17793 2561
rect 17879 2535 17905 2561
rect 2031 2479 2057 2505
rect 3991 2479 4017 2505
rect 6455 2479 6481 2505
rect 10431 2479 10457 2505
rect 11775 2479 11801 2505
rect 13399 2479 13425 2505
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 2031 2199 2057 2225
rect 7015 2199 7041 2225
rect 8359 2199 8385 2225
rect 10431 2199 10457 2225
rect 13791 2199 13817 2225
rect 15247 2199 15273 2225
rect 17879 2199 17905 2225
rect 911 2143 937 2169
rect 2031 2143 2057 2169
rect 3823 2143 3849 2169
rect 3935 2143 3961 2169
rect 4495 2143 4521 2169
rect 6119 2143 6145 2169
rect 7015 2143 7041 2169
rect 7519 2143 7545 2169
rect 8359 2143 8385 2169
rect 9255 2143 9281 2169
rect 10431 2143 10457 2169
rect 10879 2143 10905 2169
rect 11159 2143 11185 2169
rect 11383 2143 11409 2169
rect 12839 2143 12865 2169
rect 13623 2143 13649 2169
rect 14295 2143 14321 2169
rect 15247 2143 15273 2169
rect 17879 2143 17905 2169
rect 18775 2143 18801 2169
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 967 1751 993 1777
rect 2087 1751 2113 1777
rect 2871 1751 2897 1777
rect 3823 1751 3849 1777
rect 5223 1751 5249 1777
rect 5783 1751 5809 1777
rect 5895 1751 5921 1777
rect 7463 1751 7489 1777
rect 7631 1751 7657 1777
rect 7855 1751 7881 1777
rect 9423 1751 9449 1777
rect 9591 1751 9617 1777
rect 9815 1751 9841 1777
rect 10879 1751 10905 1777
rect 11663 1751 11689 1777
rect 12671 1751 12697 1777
rect 13623 1751 13649 1777
rect 14743 1751 14769 1777
rect 15527 1751 15553 1777
rect 2087 1695 2113 1721
rect 3823 1695 3849 1721
rect 11663 1695 11689 1721
rect 13623 1695 13649 1721
rect 14743 1695 14769 1721
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 1344 29600 1400 30000
rect 3808 29600 3864 30000
rect 6272 29600 6328 30000
rect 8736 29600 8792 30000
rect 11200 29600 11256 30000
rect 13664 29600 13720 30000
rect 16128 29600 16184 30000
rect 18592 29600 18648 30000
rect 1358 26922 1386 29600
rect 1358 26889 1386 26894
rect 1750 27930 1778 27935
rect 1638 25689 1666 25695
rect 1638 25663 1639 25689
rect 1665 25663 1666 25689
rect 1582 25298 1610 25303
rect 1638 25298 1666 25663
rect 1582 25297 1722 25298
rect 1582 25271 1583 25297
rect 1609 25271 1722 25297
rect 1582 25270 1722 25271
rect 1582 24906 1610 25270
rect 1694 25242 1722 25270
rect 1694 25209 1722 25214
rect 1638 24906 1666 24911
rect 1582 24905 1666 24906
rect 1582 24879 1639 24905
rect 1665 24879 1666 24905
rect 1582 24878 1666 24879
rect 1582 24513 1610 24878
rect 1638 24873 1666 24878
rect 1582 24487 1583 24513
rect 1609 24487 1610 24513
rect 1582 23730 1610 24487
rect 1582 23683 1610 23702
rect 1414 22945 1442 22951
rect 1414 22919 1415 22945
rect 1441 22919 1442 22945
rect 1414 22161 1442 22919
rect 1414 22135 1415 22161
rect 1441 22135 1442 22161
rect 1414 21378 1442 22135
rect 1582 21378 1610 21383
rect 1414 21377 1610 21378
rect 1414 21351 1583 21377
rect 1609 21351 1610 21377
rect 1414 21350 1610 21351
rect 1582 20593 1610 21350
rect 1582 20567 1583 20593
rect 1609 20567 1610 20593
rect 1582 19809 1610 20567
rect 1582 19783 1583 19809
rect 1609 19783 1610 19809
rect 1582 19025 1610 19783
rect 1582 18999 1583 19025
rect 1609 18999 1610 19025
rect 1582 18241 1610 18999
rect 1582 18215 1583 18241
rect 1609 18215 1610 18241
rect 1582 17682 1610 18215
rect 1582 17457 1610 17654
rect 1582 17431 1583 17457
rect 1609 17431 1610 17457
rect 1582 17425 1610 17431
rect 1582 16674 1610 16679
rect 1750 16674 1778 27902
rect 2238 27846 2370 27851
rect 2266 27818 2290 27846
rect 2318 27818 2342 27846
rect 2238 27813 2370 27818
rect 2238 27062 2370 27067
rect 2266 27034 2290 27062
rect 2318 27034 2342 27062
rect 2238 27029 2370 27034
rect 2086 26922 2114 26927
rect 2086 24906 2114 26894
rect 3374 26865 3402 26871
rect 3374 26839 3375 26865
rect 3401 26839 3402 26865
rect 3318 26474 3346 26479
rect 3374 26474 3402 26839
rect 3822 26866 3850 29600
rect 3822 26800 3850 26838
rect 4494 26866 4522 26871
rect 3318 26473 3402 26474
rect 3318 26447 3319 26473
rect 3345 26447 3402 26473
rect 3318 26446 3402 26447
rect 4494 26529 4522 26838
rect 4494 26503 4495 26529
rect 4521 26503 4522 26529
rect 4494 26474 4522 26503
rect 5838 26529 5866 26535
rect 5838 26503 5839 26529
rect 5865 26503 5866 26529
rect 2814 26418 2842 26423
rect 2238 26278 2370 26283
rect 2266 26250 2290 26278
rect 2318 26250 2342 26278
rect 2238 26245 2370 26250
rect 2814 25745 2842 26390
rect 2814 25719 2815 25745
rect 2841 25719 2842 25745
rect 2814 25689 2842 25719
rect 2814 25663 2815 25689
rect 2841 25663 2842 25689
rect 2238 25494 2370 25499
rect 2266 25466 2290 25494
rect 2318 25466 2342 25494
rect 2238 25461 2370 25466
rect 2478 25298 2506 25303
rect 2478 25241 2506 25270
rect 2814 25298 2842 25663
rect 2814 25265 2842 25270
rect 3094 26082 3122 26087
rect 3318 26082 3346 26446
rect 4494 26427 4522 26446
rect 5166 26473 5194 26479
rect 5166 26447 5167 26473
rect 5193 26447 5194 26473
rect 3094 26081 3318 26082
rect 3094 26055 3095 26081
rect 3121 26055 3318 26081
rect 3094 26054 3318 26055
rect 3094 25689 3122 26054
rect 3318 26016 3346 26054
rect 3542 26081 3570 26087
rect 3542 26055 3543 26081
rect 3569 26055 3570 26081
rect 3094 25663 3095 25689
rect 3121 25663 3122 25689
rect 3094 25297 3122 25663
rect 3094 25271 3095 25297
rect 3121 25271 3122 25297
rect 2478 25215 2479 25241
rect 2505 25215 2506 25241
rect 2478 25209 2506 25215
rect 3094 25242 3122 25271
rect 2310 24906 2338 24911
rect 2086 24905 2338 24906
rect 2086 24879 2087 24905
rect 2113 24879 2311 24905
rect 2337 24879 2338 24905
rect 2086 24878 2338 24879
rect 2086 24873 2114 24878
rect 2142 24514 2170 24878
rect 2310 24873 2338 24878
rect 3094 24905 3122 25214
rect 3094 24879 3095 24905
rect 3121 24879 3122 24905
rect 2238 24710 2370 24715
rect 2266 24682 2290 24710
rect 2318 24682 2342 24710
rect 2238 24677 2370 24682
rect 2142 24513 2282 24514
rect 2142 24487 2143 24513
rect 2169 24487 2282 24513
rect 2142 24486 2282 24487
rect 2142 24481 2170 24486
rect 2254 24458 2282 24486
rect 3094 24513 3122 24879
rect 3094 24487 3095 24513
rect 3121 24487 3122 24513
rect 3094 24481 3122 24487
rect 3542 25689 3570 26055
rect 3542 25663 3543 25689
rect 3569 25663 3570 25689
rect 3542 25297 3570 25663
rect 3542 25271 3543 25297
rect 3569 25271 3570 25297
rect 3542 24905 3570 25271
rect 3542 24879 3543 24905
rect 3569 24879 3570 24905
rect 3542 24513 3570 24879
rect 3542 24487 3543 24513
rect 3569 24487 3570 24513
rect 2254 24457 2338 24458
rect 2254 24431 2255 24457
rect 2281 24431 2338 24457
rect 2254 24430 2338 24431
rect 2254 24425 2282 24430
rect 1918 24234 1946 24239
rect 1862 24122 1890 24127
rect 1806 24121 1890 24122
rect 1806 24095 1863 24121
rect 1889 24095 1890 24121
rect 1806 24094 1890 24095
rect 1806 23730 1834 24094
rect 1862 24089 1890 24094
rect 1806 20538 1834 23702
rect 1918 23730 1946 24206
rect 2310 24122 2338 24430
rect 2534 24122 2562 24127
rect 2310 24121 2534 24122
rect 2310 24095 2311 24121
rect 2337 24095 2534 24121
rect 2310 24094 2534 24095
rect 2310 24089 2338 24094
rect 2238 23926 2370 23931
rect 2266 23898 2290 23926
rect 2318 23898 2342 23926
rect 2238 23893 2370 23898
rect 1918 23337 1946 23702
rect 2478 23729 2506 24094
rect 2534 24056 2562 24094
rect 3318 24121 3346 24127
rect 3318 24095 3319 24121
rect 3345 24095 3346 24121
rect 2478 23703 2479 23729
rect 2505 23703 2506 23729
rect 2478 23673 2506 23703
rect 3150 23730 3178 23735
rect 3150 23683 3178 23702
rect 3318 23730 3346 24095
rect 3542 24122 3570 24487
rect 3542 23730 3570 24094
rect 3766 26081 3794 26087
rect 3766 26055 3767 26081
rect 3793 26055 3794 26081
rect 3766 25689 3794 26055
rect 4830 26082 4858 26087
rect 4830 26035 4858 26054
rect 5166 26082 5194 26447
rect 3766 25663 3767 25689
rect 3793 25663 3794 25689
rect 3766 25297 3794 25663
rect 5166 25689 5194 26054
rect 5166 25663 5167 25689
rect 5193 25663 5194 25689
rect 3766 25271 3767 25297
rect 3793 25271 3794 25297
rect 3766 24905 3794 25271
rect 3766 24879 3767 24905
rect 3793 24879 3794 24905
rect 3766 24513 3794 24879
rect 3766 24487 3767 24513
rect 3793 24487 3794 24513
rect 3766 24122 3794 24487
rect 4886 25297 4914 25303
rect 4886 25271 4887 25297
rect 4913 25271 4914 25297
rect 4886 24905 4914 25271
rect 4886 24879 4887 24905
rect 4913 24879 4914 24905
rect 4886 24513 4914 24879
rect 5166 24906 5194 25663
rect 5726 26474 5754 26479
rect 5838 26474 5866 26503
rect 5754 26446 5866 26474
rect 5726 26081 5754 26446
rect 5726 26055 5727 26081
rect 5753 26055 5754 26081
rect 5726 26025 5754 26055
rect 5726 25999 5727 26025
rect 5753 25999 5754 26025
rect 5726 25690 5754 25999
rect 5838 25745 5866 25751
rect 5838 25719 5839 25745
rect 5865 25719 5866 25745
rect 5838 25690 5866 25719
rect 5726 25689 5866 25690
rect 5726 25663 5727 25689
rect 5753 25663 5866 25689
rect 5726 25662 5866 25663
rect 5726 24962 5754 25662
rect 5782 25297 5810 25303
rect 5782 25271 5783 25297
rect 5809 25271 5810 25297
rect 5782 25242 5810 25271
rect 6286 25242 6314 29600
rect 5782 25241 5866 25242
rect 5782 25215 5783 25241
rect 5809 25215 5866 25241
rect 5782 25214 5866 25215
rect 5782 25209 5810 25214
rect 5726 24929 5754 24934
rect 5838 24961 5866 25214
rect 6286 25209 6314 25214
rect 7126 25297 7154 25303
rect 7126 25271 7127 25297
rect 7153 25271 7154 25297
rect 5838 24935 5839 24961
rect 5865 24935 5866 24961
rect 5166 24873 5194 24878
rect 5838 24905 5866 24935
rect 5838 24879 5839 24905
rect 5865 24879 5866 24905
rect 4886 24487 4887 24513
rect 4913 24487 4914 24513
rect 3990 24122 4018 24127
rect 3794 24094 3850 24122
rect 3766 24075 3794 24094
rect 3598 23730 3626 23735
rect 3542 23729 3626 23730
rect 3542 23703 3599 23729
rect 3625 23703 3626 23729
rect 3542 23702 3626 23703
rect 3318 23697 3346 23702
rect 3598 23697 3626 23702
rect 3822 23729 3850 24094
rect 3990 24075 4018 24094
rect 4886 24122 4914 24487
rect 5782 24513 5810 24519
rect 5782 24487 5783 24513
rect 5809 24487 5810 24513
rect 5782 24458 5810 24487
rect 5838 24458 5866 24879
rect 5782 24457 5866 24458
rect 5782 24431 5783 24457
rect 5809 24431 5866 24457
rect 5782 24430 5866 24431
rect 5782 24425 5810 24430
rect 5838 24178 5866 24430
rect 6622 24906 6650 24911
rect 6622 24402 6650 24878
rect 6622 24369 6650 24374
rect 7070 24513 7098 24519
rect 7070 24487 7071 24513
rect 7097 24487 7098 24513
rect 7070 24402 7098 24487
rect 7126 24514 7154 25271
rect 8022 25297 8050 25303
rect 8022 25271 8023 25297
rect 8049 25271 8050 25297
rect 8022 25241 8050 25271
rect 8022 25215 8023 25241
rect 8049 25215 8050 25241
rect 7126 24481 7154 24486
rect 7518 24962 7546 24967
rect 7518 24905 7546 24934
rect 7518 24879 7519 24905
rect 7545 24879 7546 24905
rect 7518 24458 7546 24879
rect 7518 24425 7546 24430
rect 7966 24513 7994 24519
rect 7966 24487 7967 24513
rect 7993 24487 7994 24513
rect 7966 24458 7994 24487
rect 7966 24411 7994 24430
rect 7070 24369 7098 24374
rect 3822 23703 3823 23729
rect 3849 23703 3850 23729
rect 2478 23647 2479 23673
rect 2505 23647 2506 23673
rect 1918 23311 1919 23337
rect 1945 23311 1946 23337
rect 1918 22554 1946 23311
rect 2422 23338 2450 23343
rect 2478 23338 2506 23647
rect 3822 23674 3850 23703
rect 4886 23730 4914 24094
rect 5166 24122 5194 24127
rect 5166 24075 5194 24094
rect 5838 24121 5866 24150
rect 7518 24177 7546 24183
rect 7518 24151 7519 24177
rect 7545 24151 7546 24177
rect 5838 24095 5839 24121
rect 5865 24095 5866 24121
rect 4886 23664 4914 23702
rect 5782 23730 5810 23735
rect 5838 23730 5866 24095
rect 5782 23729 5866 23730
rect 5782 23703 5783 23729
rect 5809 23703 5866 23729
rect 5782 23702 5866 23703
rect 6062 24122 6090 24127
rect 5782 23674 5810 23702
rect 3822 23641 3850 23646
rect 5782 23608 5810 23646
rect 4438 23393 4466 23399
rect 4438 23367 4439 23393
rect 4465 23367 4466 23393
rect 2534 23338 2562 23343
rect 2422 23337 2562 23338
rect 2422 23311 2423 23337
rect 2449 23311 2535 23337
rect 2561 23311 2562 23337
rect 2422 23310 2562 23311
rect 2422 23305 2450 23310
rect 2238 23142 2370 23147
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2238 23109 2370 23114
rect 2478 22945 2506 23310
rect 2534 23305 2562 23310
rect 3598 23337 3626 23343
rect 3598 23311 3599 23337
rect 3625 23311 3626 23337
rect 2478 22919 2479 22945
rect 2505 22919 2506 22945
rect 2478 22889 2506 22919
rect 2478 22863 2479 22889
rect 2505 22863 2506 22889
rect 2422 22554 2450 22559
rect 2478 22554 2506 22863
rect 2534 22554 2562 22559
rect 1918 22553 2170 22554
rect 1918 22527 1919 22553
rect 1945 22527 2170 22553
rect 1918 22526 2170 22527
rect 1918 22521 1946 22526
rect 2142 21854 2170 22526
rect 2422 22553 3066 22554
rect 2422 22527 2423 22553
rect 2449 22527 2535 22553
rect 2561 22527 3066 22553
rect 2422 22526 3066 22527
rect 2422 22521 2450 22526
rect 2534 22521 2562 22526
rect 2238 22358 2370 22363
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2238 22325 2370 22330
rect 1806 20505 1834 20510
rect 1862 21826 2170 21854
rect 2254 22161 2282 22167
rect 2254 22135 2255 22161
rect 2281 22135 2282 22161
rect 2254 22105 2282 22135
rect 2254 22079 2255 22105
rect 2281 22079 2282 22105
rect 1862 21769 1890 21826
rect 1862 21743 1863 21769
rect 1889 21743 1890 21769
rect 1862 20985 1890 21743
rect 2254 21770 2282 22079
rect 2254 21737 2282 21742
rect 3038 21825 3066 22526
rect 3038 21799 3039 21825
rect 3065 21799 3066 21825
rect 3038 21770 3066 21799
rect 3598 22553 3626 23311
rect 4438 23337 4466 23367
rect 4438 23311 4439 23337
rect 4465 23311 4466 23337
rect 3598 22527 3599 22553
rect 3625 22527 3626 22553
rect 2238 21574 2370 21579
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2238 21541 2370 21546
rect 1862 20959 1863 20985
rect 1889 20959 1890 20985
rect 1862 20201 1890 20959
rect 2478 21377 2506 21383
rect 2478 21351 2479 21377
rect 2505 21351 2506 21377
rect 2478 21322 2506 21351
rect 2238 20790 2370 20795
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2238 20757 2370 20762
rect 2478 20593 2506 21294
rect 3038 21322 3066 21742
rect 3038 21041 3066 21294
rect 3038 21015 3039 21041
rect 3065 21015 3066 21041
rect 3038 20985 3066 21015
rect 3038 20959 3039 20985
rect 3065 20959 3066 20985
rect 3038 20953 3066 20959
rect 3374 21770 3402 21775
rect 3598 21770 3626 22527
rect 3934 22945 3962 22951
rect 3934 22919 3935 22945
rect 3961 22919 3962 22945
rect 3934 22161 3962 22919
rect 4382 22946 4410 22951
rect 4438 22946 4466 23311
rect 6062 23337 6090 24094
rect 6342 24122 6370 24127
rect 6342 24075 6370 24094
rect 7518 24122 7546 24151
rect 7518 24075 7546 24094
rect 8022 24122 8050 25215
rect 8582 24514 8610 24519
rect 8582 24467 8610 24486
rect 8358 24458 8386 24463
rect 8358 24402 8386 24430
rect 8750 24458 8778 29600
rect 9918 28238 10050 28243
rect 9946 28210 9970 28238
rect 9998 28210 10022 28238
rect 9918 28205 10050 28210
rect 11214 27734 11242 29600
rect 11046 27706 11242 27734
rect 9918 27454 10050 27459
rect 9946 27426 9970 27454
rect 9998 27426 10022 27454
rect 9918 27421 10050 27426
rect 9918 26670 10050 26675
rect 9946 26642 9970 26670
rect 9998 26642 10022 26670
rect 9918 26637 10050 26642
rect 9918 25886 10050 25891
rect 9946 25858 9970 25886
rect 9998 25858 10022 25886
rect 9918 25853 10050 25858
rect 9918 25102 10050 25107
rect 9946 25074 9970 25102
rect 9998 25074 10022 25102
rect 9918 25069 10050 25074
rect 8750 24425 8778 24430
rect 9142 24514 9170 24519
rect 8582 24402 8610 24407
rect 8358 24374 8442 24402
rect 7126 23729 7154 23735
rect 7126 23703 7127 23729
rect 7153 23703 7154 23729
rect 6062 23311 6063 23337
rect 6089 23311 6090 23337
rect 4494 22946 4522 22951
rect 4382 22945 4522 22946
rect 4382 22919 4383 22945
rect 4409 22919 4495 22945
rect 4521 22919 4522 22945
rect 4382 22918 4522 22919
rect 4382 22913 4410 22918
rect 3934 22135 3935 22161
rect 3961 22135 3962 22161
rect 3934 21854 3962 22135
rect 4438 22609 4466 22918
rect 4494 22913 4522 22918
rect 5278 22945 5306 22951
rect 5278 22919 5279 22945
rect 5305 22919 5306 22945
rect 4438 22583 4439 22609
rect 4465 22583 4466 22609
rect 4438 22553 4466 22583
rect 4438 22527 4439 22553
rect 4465 22527 4466 22553
rect 4438 21854 4466 22527
rect 4774 22161 4802 22167
rect 4774 22135 4775 22161
rect 4801 22135 4802 22161
rect 4774 22105 4802 22135
rect 4774 22079 4775 22105
rect 4801 22079 4802 22105
rect 4774 21854 4802 22079
rect 3374 21769 3626 21770
rect 3374 21743 3375 21769
rect 3401 21743 3626 21769
rect 3374 21742 3626 21743
rect 3822 21826 3962 21854
rect 4270 21826 4802 21854
rect 5278 22161 5306 22919
rect 5278 22135 5279 22161
rect 5305 22135 5306 22161
rect 3374 20985 3402 21742
rect 3374 20959 3375 20985
rect 3401 20959 3402 20985
rect 2478 20567 2479 20593
rect 2505 20567 2506 20593
rect 2478 20537 2506 20567
rect 2478 20511 2479 20537
rect 2505 20511 2506 20537
rect 2478 20505 2506 20511
rect 1862 20175 1863 20201
rect 1889 20175 1890 20201
rect 1862 19417 1890 20175
rect 2422 20202 2450 20207
rect 2534 20202 2562 20207
rect 2422 20201 2562 20202
rect 2422 20175 2423 20201
rect 2449 20175 2535 20201
rect 2561 20175 2562 20201
rect 2422 20174 2562 20175
rect 2238 20006 2370 20011
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2238 19973 2370 19978
rect 1862 19391 1863 19417
rect 1889 19391 1890 19417
rect 1862 18633 1890 19391
rect 2422 19809 2450 20174
rect 2534 20169 2562 20174
rect 3374 20201 3402 20959
rect 3374 20175 3375 20201
rect 3401 20175 3402 20201
rect 2422 19783 2423 19809
rect 2449 19783 2450 19809
rect 2422 19753 2450 19783
rect 2422 19727 2423 19753
rect 2449 19727 2450 19753
rect 2422 19418 2450 19727
rect 2534 19418 2562 19423
rect 2422 19417 2562 19418
rect 2422 19391 2423 19417
rect 2449 19391 2535 19417
rect 2561 19391 2562 19417
rect 2422 19390 2562 19391
rect 2422 19385 2450 19390
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 1862 18607 1863 18633
rect 1889 18607 1890 18633
rect 1862 17906 1890 18607
rect 2478 19026 2506 19031
rect 2534 19026 2562 19390
rect 2478 19025 2562 19026
rect 2478 18999 2479 19025
rect 2505 18999 2562 19025
rect 2478 18998 2562 18999
rect 3374 19417 3402 20175
rect 3374 19391 3375 19417
rect 3401 19391 3402 19417
rect 2478 18969 2506 18998
rect 2478 18943 2479 18969
rect 2505 18943 2506 18969
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2478 18242 2506 18943
rect 2478 18185 2506 18214
rect 2478 18159 2479 18185
rect 2505 18159 2506 18185
rect 2478 18153 2506 18159
rect 3038 18689 3066 18695
rect 3038 18663 3039 18689
rect 3065 18663 3066 18689
rect 3038 18633 3066 18663
rect 3038 18607 3039 18633
rect 3065 18607 3066 18633
rect 3038 18242 3066 18607
rect 1862 17849 1890 17878
rect 1862 17823 1863 17849
rect 1889 17823 1890 17849
rect 1862 17682 1890 17823
rect 3038 17905 3066 18214
rect 3038 17879 3039 17905
rect 3065 17879 3066 17905
rect 3038 17850 3066 17879
rect 3038 17803 3066 17822
rect 3374 18633 3402 19391
rect 3374 18607 3375 18633
rect 3401 18607 3402 18633
rect 3374 18242 3402 18607
rect 3822 21377 3850 21826
rect 4214 21825 4298 21826
rect 4214 21799 4271 21825
rect 4297 21799 4298 21825
rect 4214 21798 4298 21799
rect 4214 21770 4242 21798
rect 4270 21793 4298 21798
rect 4214 21723 4242 21742
rect 3822 21351 3823 21377
rect 3849 21351 3850 21377
rect 3822 20593 3850 21351
rect 4774 21377 4802 21383
rect 4774 21351 4775 21377
rect 4801 21351 4802 21377
rect 4774 21321 4802 21351
rect 4774 21295 4775 21321
rect 4801 21295 4802 21321
rect 4494 21042 4522 21047
rect 4774 21042 4802 21295
rect 4494 21041 4802 21042
rect 4494 21015 4495 21041
rect 4521 21015 4802 21041
rect 4494 21014 4802 21015
rect 5278 21377 5306 22135
rect 5278 21351 5279 21377
rect 5305 21351 5306 21377
rect 4494 20985 4522 21014
rect 4494 20959 4495 20985
rect 4521 20959 4522 20985
rect 3822 20567 3823 20593
rect 3849 20567 3850 20593
rect 3822 19809 3850 20567
rect 4382 20594 4410 20599
rect 4494 20594 4522 20959
rect 4382 20593 4522 20594
rect 4382 20567 4383 20593
rect 4409 20567 4495 20593
rect 4521 20567 4522 20593
rect 4382 20566 4522 20567
rect 4382 20561 4410 20566
rect 4438 20257 4466 20566
rect 4494 20561 4522 20566
rect 5278 20593 5306 21351
rect 5278 20567 5279 20593
rect 5305 20567 5306 20593
rect 4438 20231 4439 20257
rect 4465 20231 4466 20257
rect 4438 20201 4466 20231
rect 4438 20175 4439 20201
rect 4465 20175 4466 20201
rect 3822 19783 3823 19809
rect 3849 19783 3850 19809
rect 3822 19026 3850 19783
rect 4382 19810 4410 19815
rect 4438 19810 4466 20175
rect 4494 19810 4522 19815
rect 4382 19809 4522 19810
rect 4382 19783 4383 19809
rect 4409 19783 4495 19809
rect 4521 19783 4522 19809
rect 4382 19782 4522 19783
rect 4382 19777 4410 19782
rect 4438 19473 4466 19782
rect 4494 19777 4522 19782
rect 5278 19809 5306 20567
rect 6062 22553 6090 23311
rect 6062 22527 6063 22553
rect 6089 22527 6090 22553
rect 6062 21769 6090 22527
rect 6342 23338 6370 23343
rect 6454 23338 6482 23343
rect 6342 23337 6482 23338
rect 6342 23311 6343 23337
rect 6369 23311 6455 23337
rect 6481 23311 6482 23337
rect 6342 23310 6482 23311
rect 6342 22945 6370 23310
rect 6454 23305 6482 23310
rect 7126 23338 7154 23703
rect 8022 23729 8050 24094
rect 8022 23703 8023 23729
rect 8049 23703 8050 23729
rect 8022 23673 8050 23703
rect 8414 23730 8442 24374
rect 8414 23697 8442 23702
rect 8582 23729 8610 24374
rect 8582 23703 8583 23729
rect 8609 23703 8610 23729
rect 8022 23647 8023 23673
rect 8049 23647 8050 23673
rect 7238 23338 7266 23343
rect 7126 23337 7266 23338
rect 7126 23311 7239 23337
rect 7265 23311 7266 23337
rect 7126 23310 7266 23311
rect 6342 22919 6343 22945
rect 6369 22919 6370 22945
rect 6342 22889 6370 22919
rect 6342 22863 6343 22889
rect 6369 22863 6370 22889
rect 6342 22554 6370 22863
rect 7126 22945 7154 23310
rect 7238 23305 7266 23310
rect 8022 23338 8050 23647
rect 8190 23393 8218 23399
rect 8190 23367 8191 23393
rect 8217 23367 8218 23393
rect 8190 23338 8218 23367
rect 8022 23337 8218 23338
rect 8022 23311 8023 23337
rect 8049 23311 8218 23337
rect 8022 23310 8218 23311
rect 7126 22919 7127 22945
rect 7153 22919 7154 22945
rect 6454 22554 6482 22559
rect 6342 22553 6482 22554
rect 6342 22527 6343 22553
rect 6369 22527 6455 22553
rect 6481 22527 6482 22553
rect 6342 22526 6482 22527
rect 6342 22161 6370 22526
rect 6454 22521 6482 22526
rect 6342 22135 6343 22161
rect 6369 22135 6370 22161
rect 6342 22106 6370 22135
rect 7126 22161 7154 22919
rect 8022 22945 8050 23310
rect 8582 23282 8610 23703
rect 9142 24121 9170 24486
rect 9478 24513 9506 24519
rect 9478 24487 9479 24513
rect 9505 24487 9506 24513
rect 9478 24457 9506 24487
rect 9478 24431 9479 24457
rect 9505 24431 9506 24457
rect 9478 24178 9506 24431
rect 9918 24318 10050 24323
rect 9946 24290 9970 24318
rect 9998 24290 10022 24318
rect 9918 24285 10050 24290
rect 9814 24178 9842 24183
rect 9478 24177 9842 24178
rect 9478 24151 9815 24177
rect 9841 24151 9842 24177
rect 9478 24150 9842 24151
rect 9142 24095 9143 24121
rect 9169 24095 9170 24121
rect 8582 23249 8610 23254
rect 9086 23337 9114 23343
rect 9086 23311 9087 23337
rect 9113 23311 9114 23337
rect 9086 23282 9114 23311
rect 9142 23338 9170 24095
rect 9814 24121 9842 24150
rect 9814 24095 9815 24121
rect 9841 24095 9842 24121
rect 9142 23305 9170 23310
rect 9422 23730 9450 23735
rect 9422 23673 9450 23702
rect 9422 23647 9423 23673
rect 9449 23647 9450 23673
rect 9422 23338 9450 23647
rect 9534 23338 9562 23343
rect 9422 23337 9562 23338
rect 9422 23311 9423 23337
rect 9449 23311 9535 23337
rect 9561 23311 9562 23337
rect 9422 23310 9562 23311
rect 9086 23249 9114 23254
rect 8022 22919 8023 22945
rect 8049 22919 8050 22945
rect 8022 22889 8050 22919
rect 8022 22863 8023 22889
rect 8049 22863 8050 22889
rect 7126 22135 7127 22161
rect 7153 22135 7154 22161
rect 6342 22105 6706 22106
rect 6342 22079 6343 22105
rect 6369 22079 6706 22105
rect 6342 22078 6706 22079
rect 6342 22073 6370 22078
rect 6678 21854 6706 22078
rect 6454 21826 6706 21854
rect 6062 21743 6063 21769
rect 6089 21743 6090 21769
rect 6062 21042 6090 21743
rect 6342 21770 6370 21775
rect 6454 21770 6482 21826
rect 6342 21769 6482 21770
rect 6342 21743 6343 21769
rect 6369 21743 6455 21769
rect 6481 21743 6482 21769
rect 6342 21742 6482 21743
rect 6342 21737 6370 21742
rect 6062 20985 6090 21014
rect 6454 21377 6482 21742
rect 6454 21351 6455 21377
rect 6481 21351 6482 21377
rect 6454 21321 6482 21351
rect 6454 21295 6455 21321
rect 6481 21295 6482 21321
rect 6062 20959 6063 20985
rect 6089 20959 6090 20985
rect 6062 20201 6090 20959
rect 6342 20986 6370 20991
rect 6454 20986 6482 21295
rect 6342 20985 6482 20986
rect 6342 20959 6343 20985
rect 6369 20959 6455 20985
rect 6481 20959 6482 20985
rect 6342 20958 6482 20959
rect 6342 20953 6370 20958
rect 6454 20593 6482 20958
rect 6454 20567 6455 20593
rect 6481 20567 6482 20593
rect 6454 20537 6482 20567
rect 7126 21377 7154 22135
rect 7126 21351 7127 21377
rect 7153 21351 7154 21377
rect 7126 21042 7154 21351
rect 7126 20594 7154 21014
rect 7462 22553 7490 22559
rect 7462 22527 7463 22553
rect 7489 22527 7490 22553
rect 7462 21769 7490 22527
rect 8022 22554 8050 22863
rect 8414 22945 8442 22951
rect 8414 22919 8415 22945
rect 8441 22919 8442 22945
rect 8022 22521 8050 22526
rect 8358 22609 8386 22615
rect 8358 22583 8359 22609
rect 8385 22583 8386 22609
rect 8358 22554 8386 22583
rect 8358 22507 8386 22526
rect 7798 22161 7826 22167
rect 7798 22135 7799 22161
rect 7825 22135 7826 22161
rect 7798 22105 7826 22135
rect 8414 22162 8442 22919
rect 9142 22553 9170 22559
rect 9142 22527 9143 22553
rect 9169 22527 9170 22553
rect 8414 22161 8610 22162
rect 8414 22135 8415 22161
rect 8441 22135 8610 22161
rect 8414 22134 8610 22135
rect 8414 22129 8442 22134
rect 7798 22079 7799 22105
rect 7825 22079 7826 22105
rect 7798 21854 7826 22079
rect 7462 21743 7463 21769
rect 7489 21743 7490 21769
rect 7462 20986 7490 21743
rect 7686 21826 7826 21854
rect 7686 21769 7714 21826
rect 7686 21743 7687 21769
rect 7713 21743 7714 21769
rect 7574 21377 7602 21383
rect 7574 21351 7575 21377
rect 7601 21351 7602 21377
rect 7574 21322 7602 21351
rect 7686 21322 7714 21743
rect 7798 21770 7826 21826
rect 7910 21770 7938 21775
rect 7798 21769 7938 21770
rect 7798 21743 7911 21769
rect 7937 21743 7938 21769
rect 7798 21742 7938 21743
rect 7910 21737 7938 21742
rect 8582 21377 8610 22134
rect 9142 21769 9170 22527
rect 9142 21743 9143 21769
rect 9169 21743 9170 21769
rect 8582 21351 8583 21377
rect 8609 21351 8610 21377
rect 7798 21322 7826 21327
rect 7574 21321 7826 21322
rect 7574 21295 7799 21321
rect 7825 21295 7826 21321
rect 7574 21294 7826 21295
rect 7518 21042 7546 21047
rect 7518 20986 7546 21014
rect 7462 20985 7546 20986
rect 7462 20959 7519 20985
rect 7545 20959 7546 20985
rect 7462 20958 7546 20959
rect 7462 20594 7490 20958
rect 7518 20953 7546 20958
rect 7126 20593 7490 20594
rect 7126 20567 7127 20593
rect 7153 20567 7490 20593
rect 7126 20566 7490 20567
rect 7126 20561 7154 20566
rect 6454 20511 6455 20537
rect 6481 20511 6482 20537
rect 6062 20175 6063 20201
rect 6089 20175 6090 20201
rect 6062 20169 6090 20175
rect 6342 20202 6370 20207
rect 6454 20202 6482 20511
rect 6342 20201 6482 20202
rect 6342 20175 6343 20201
rect 6369 20175 6455 20201
rect 6481 20175 6482 20201
rect 6342 20174 6482 20175
rect 6342 20169 6370 20174
rect 5278 19783 5279 19809
rect 5305 19783 5306 19809
rect 4438 19447 4439 19473
rect 4465 19447 4466 19473
rect 4438 19417 4466 19447
rect 4438 19391 4439 19417
rect 4465 19391 4466 19417
rect 3822 18242 3850 18998
rect 4382 19026 4410 19031
rect 4438 19026 4466 19391
rect 5278 19417 5306 19783
rect 5278 19391 5279 19417
rect 5305 19391 5306 19417
rect 4494 19026 4522 19031
rect 4382 19025 4522 19026
rect 4382 18999 4383 19025
rect 4409 18999 4495 19025
rect 4521 18999 4522 19025
rect 4382 18998 4522 18999
rect 4382 18993 4410 18998
rect 4438 18689 4466 18998
rect 4494 18993 4522 18998
rect 5278 19026 5306 19391
rect 5278 18979 5306 18998
rect 6398 19809 6426 20174
rect 6454 20169 6482 20174
rect 7462 20201 7490 20566
rect 7462 20175 7463 20201
rect 7489 20175 7490 20201
rect 7462 20169 7490 20175
rect 7574 20593 7602 21294
rect 7686 20986 7714 21294
rect 7798 21289 7826 21294
rect 8582 21042 8610 21351
rect 7910 20986 7938 20991
rect 7686 20985 7938 20986
rect 7686 20959 7687 20985
rect 7713 20959 7911 20985
rect 7937 20959 7938 20985
rect 7686 20958 7938 20959
rect 7686 20953 7714 20958
rect 7910 20953 7938 20958
rect 7574 20567 7575 20593
rect 7601 20567 7602 20593
rect 7574 20538 7602 20567
rect 8582 20593 8610 21014
rect 8582 20567 8583 20593
rect 8609 20567 8610 20593
rect 7798 20538 7826 20543
rect 7574 20537 7826 20538
rect 7574 20511 7799 20537
rect 7825 20511 7826 20537
rect 7574 20510 7826 20511
rect 6398 19783 6399 19809
rect 6425 19783 6426 19809
rect 6398 19753 6426 19783
rect 6398 19727 6399 19753
rect 6425 19727 6426 19753
rect 6398 19473 6426 19727
rect 6398 19447 6399 19473
rect 6425 19447 6426 19473
rect 6398 19417 6426 19447
rect 6398 19391 6399 19417
rect 6425 19391 6426 19417
rect 6398 19025 6426 19391
rect 6398 18999 6399 19025
rect 6425 18999 6426 19025
rect 4438 18663 4439 18689
rect 4465 18663 4466 18689
rect 4438 18633 4466 18663
rect 6398 18969 6426 18999
rect 6398 18943 6399 18969
rect 6425 18943 6426 18969
rect 6398 18689 6426 18943
rect 6398 18663 6399 18689
rect 6425 18663 6426 18689
rect 4438 18607 4439 18633
rect 4465 18607 4466 18633
rect 3374 18241 3850 18242
rect 3374 18215 3823 18241
rect 3849 18215 3850 18241
rect 3374 18214 3850 18215
rect 3374 17906 3402 18214
rect 3822 18209 3850 18214
rect 4382 18242 4410 18247
rect 4438 18242 4466 18607
rect 5278 18633 5306 18639
rect 5278 18607 5279 18633
rect 5305 18607 5306 18633
rect 4494 18242 4522 18247
rect 4382 18241 4522 18242
rect 4382 18215 4383 18241
rect 4409 18215 4495 18241
rect 4521 18215 4522 18241
rect 4382 18214 4522 18215
rect 4382 18209 4410 18214
rect 3374 17849 3402 17878
rect 3374 17823 3375 17849
rect 3401 17823 3402 17849
rect 3374 17817 3402 17823
rect 4438 17905 4466 18214
rect 4494 18209 4522 18214
rect 5278 18241 5306 18607
rect 5278 18215 5279 18241
rect 5305 18215 5306 18241
rect 4438 17879 4439 17905
rect 4465 17879 4466 17905
rect 4438 17850 4466 17879
rect 1862 17065 1890 17654
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 1862 17039 1863 17065
rect 1889 17039 1890 17065
rect 1862 17033 1890 17039
rect 2422 17457 2450 17463
rect 2422 17431 2423 17457
rect 2449 17431 2450 17457
rect 2422 17401 2450 17431
rect 2422 17375 2423 17401
rect 2449 17375 2450 17401
rect 2422 17066 2450 17375
rect 3878 17457 3906 17463
rect 3878 17431 3879 17457
rect 3905 17431 3906 17457
rect 2590 17066 2618 17071
rect 2422 17065 2618 17066
rect 2422 17039 2423 17065
rect 2449 17039 2591 17065
rect 2617 17039 2618 17065
rect 2422 17038 2618 17039
rect 2422 17033 2450 17038
rect 2238 16870 2370 16875
rect 1582 16673 1778 16674
rect 1582 16647 1583 16673
rect 1609 16647 1778 16673
rect 1582 16646 1778 16647
rect 1358 15890 1386 15895
rect 1582 15890 1610 16646
rect 1750 16282 1778 16646
rect 2086 16842 2114 16847
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 1862 16282 1890 16287
rect 1750 16281 1890 16282
rect 1750 16255 1863 16281
rect 1889 16255 1890 16281
rect 1750 16254 1890 16255
rect 1358 15889 1610 15890
rect 1358 15863 1359 15889
rect 1385 15863 1610 15889
rect 1358 15862 1610 15863
rect 1358 15105 1386 15862
rect 1358 15079 1359 15105
rect 1385 15079 1386 15105
rect 1358 14321 1386 15079
rect 1358 14295 1359 14321
rect 1385 14295 1386 14321
rect 1358 13537 1386 14295
rect 1358 13511 1359 13537
rect 1385 13511 1386 13537
rect 1358 12753 1386 13511
rect 1862 15497 1890 16254
rect 1862 15471 1863 15497
rect 1889 15471 1890 15497
rect 1862 14713 1890 15471
rect 1862 14687 1863 14713
rect 1889 14687 1890 14713
rect 1862 13929 1890 14687
rect 1862 13903 1863 13929
rect 1889 13903 1890 13929
rect 1358 12727 1359 12753
rect 1385 12727 1386 12753
rect 1358 11969 1386 12727
rect 1358 11943 1359 11969
rect 1385 11943 1386 11969
rect 1358 11937 1386 11943
rect 1694 13146 1722 13151
rect 1414 11185 1442 11191
rect 1414 11159 1415 11185
rect 1441 11159 1442 11185
rect 1414 10401 1442 11159
rect 1414 10375 1415 10401
rect 1441 10375 1442 10401
rect 1414 9618 1442 10375
rect 1582 9618 1610 9623
rect 1414 9617 1610 9618
rect 1414 9591 1583 9617
rect 1609 9591 1610 9617
rect 1414 9590 1610 9591
rect 910 9450 938 9455
rect 910 4129 938 9422
rect 1582 9282 1610 9590
rect 1582 9249 1610 9254
rect 1582 8833 1610 8839
rect 1582 8807 1583 8833
rect 1609 8807 1610 8833
rect 1582 8050 1610 8807
rect 1582 8003 1610 8022
rect 1582 7266 1610 7271
rect 1582 6481 1610 7238
rect 1582 6455 1583 6481
rect 1609 6455 1610 6481
rect 1582 6449 1610 6455
rect 1638 6090 1666 6095
rect 1694 6090 1722 13118
rect 1862 13145 1890 13903
rect 1862 13119 1863 13145
rect 1889 13119 1890 13145
rect 1862 12361 1890 13119
rect 1862 12335 1863 12361
rect 1889 12335 1890 12361
rect 1862 11578 1890 12335
rect 1862 11512 1890 11550
rect 1918 10793 1946 10799
rect 1918 10767 1919 10793
rect 1945 10767 1946 10793
rect 1918 10009 1946 10767
rect 1918 9983 1919 10009
rect 1945 9983 1946 10009
rect 1918 9282 1946 9983
rect 1918 9225 1946 9254
rect 1918 9199 1919 9225
rect 1945 9199 1946 9225
rect 1918 9193 1946 9199
rect 2086 8498 2114 16814
rect 2310 16673 2338 16679
rect 2310 16647 2311 16673
rect 2337 16647 2338 16673
rect 2310 16617 2338 16647
rect 2310 16591 2311 16617
rect 2337 16591 2338 16617
rect 2310 16282 2338 16591
rect 2534 16282 2562 16287
rect 2310 16281 2562 16282
rect 2310 16255 2311 16281
rect 2337 16255 2535 16281
rect 2561 16255 2562 16281
rect 2310 16254 2562 16255
rect 2310 16249 2338 16254
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2478 15889 2506 16254
rect 2534 16249 2562 16254
rect 2590 15974 2618 17038
rect 2478 15863 2479 15889
rect 2505 15863 2506 15889
rect 2478 15834 2506 15863
rect 2142 15833 2506 15834
rect 2142 15807 2479 15833
rect 2505 15807 2506 15833
rect 2142 15806 2506 15807
rect 2142 13538 2170 15806
rect 2478 15801 2506 15806
rect 2534 15946 2618 15974
rect 3430 17065 3458 17071
rect 3430 17039 3431 17065
rect 3457 17039 3458 17065
rect 3430 16281 3458 17039
rect 3430 16255 3431 16281
rect 3457 16255 3458 16281
rect 3430 15974 3458 16255
rect 3878 16673 3906 17431
rect 4382 17458 4410 17463
rect 4438 17458 4466 17822
rect 5278 17849 5306 18215
rect 5278 17823 5279 17849
rect 5305 17823 5306 17849
rect 4494 17458 4522 17463
rect 4382 17457 4522 17458
rect 4382 17431 4383 17457
rect 4409 17431 4495 17457
rect 4521 17431 4522 17457
rect 4382 17430 4522 17431
rect 4382 17425 4410 17430
rect 4438 17121 4466 17430
rect 4494 17425 4522 17430
rect 5278 17457 5306 17823
rect 5278 17431 5279 17457
rect 5305 17431 5306 17457
rect 4438 17095 4439 17121
rect 4465 17095 4466 17121
rect 4438 17066 4466 17095
rect 3878 16647 3879 16673
rect 3905 16647 3906 16673
rect 3878 15974 3906 16647
rect 4382 17065 4466 17066
rect 4382 17039 4439 17065
rect 4465 17039 4466 17065
rect 4382 17038 4466 17039
rect 4382 16674 4410 17038
rect 4438 17033 4466 17038
rect 5278 17065 5306 17431
rect 5278 17039 5279 17065
rect 5305 17039 5306 17065
rect 4494 16674 4522 16679
rect 4382 16673 4522 16674
rect 4382 16647 4383 16673
rect 4409 16647 4495 16673
rect 4521 16647 4522 16673
rect 4382 16646 4522 16647
rect 4382 16641 4410 16646
rect 4438 16337 4466 16646
rect 4494 16641 4522 16646
rect 5278 16673 5306 17039
rect 5278 16647 5279 16673
rect 5305 16647 5306 16673
rect 4438 16311 4439 16337
rect 4465 16311 4466 16337
rect 4438 16281 4466 16311
rect 4438 16255 4439 16281
rect 4465 16255 4466 16281
rect 4438 15974 4466 16255
rect 3430 15946 3626 15974
rect 3878 15946 4074 15974
rect 2422 15498 2450 15503
rect 2534 15498 2562 15946
rect 2422 15497 2562 15498
rect 2422 15471 2423 15497
rect 2449 15471 2535 15497
rect 2561 15471 2562 15497
rect 2422 15470 2562 15471
rect 2422 15465 2450 15470
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2478 15106 2506 15111
rect 2534 15106 2562 15470
rect 2478 15105 2562 15106
rect 2478 15079 2479 15105
rect 2505 15079 2562 15105
rect 2478 15078 2562 15079
rect 3598 15497 3626 15946
rect 3598 15471 3599 15497
rect 3625 15471 3626 15497
rect 2478 15049 2506 15078
rect 2478 15023 2479 15049
rect 2505 15023 2506 15049
rect 2422 14714 2450 14719
rect 2478 14714 2506 15023
rect 2534 14714 2562 14719
rect 2422 14713 2562 14714
rect 2422 14687 2423 14713
rect 2449 14687 2535 14713
rect 2561 14687 2562 14713
rect 2422 14686 2562 14687
rect 2422 14681 2450 14686
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2478 14322 2506 14327
rect 2534 14322 2562 14686
rect 2478 14321 2534 14322
rect 2478 14295 2479 14321
rect 2505 14295 2534 14321
rect 2478 14294 2534 14295
rect 2478 14265 2506 14294
rect 2478 14239 2479 14265
rect 2505 14239 2506 14265
rect 2534 14256 2562 14294
rect 3598 14713 3626 15471
rect 3598 14687 3599 14713
rect 3625 14687 3626 14713
rect 2422 13930 2450 13935
rect 2478 13930 2506 14239
rect 2590 13930 2618 13935
rect 2422 13929 2618 13930
rect 2422 13903 2423 13929
rect 2449 13903 2591 13929
rect 2617 13903 2618 13929
rect 2422 13902 2618 13903
rect 2422 13897 2450 13902
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2142 13537 2282 13538
rect 2142 13511 2143 13537
rect 2169 13511 2282 13537
rect 2142 13510 2282 13511
rect 2142 13505 2170 13510
rect 2254 13482 2282 13510
rect 2254 13481 2338 13482
rect 2254 13455 2255 13481
rect 2281 13455 2338 13481
rect 2254 13454 2338 13455
rect 2254 13449 2282 13454
rect 2310 13146 2338 13454
rect 2534 13146 2562 13151
rect 2310 13145 2562 13146
rect 2310 13119 2311 13145
rect 2337 13119 2535 13145
rect 2561 13119 2562 13145
rect 2310 13118 2562 13119
rect 2310 13113 2338 13118
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2478 12753 2506 13118
rect 2534 13113 2562 13118
rect 2478 12727 2479 12753
rect 2505 12727 2506 12753
rect 2478 12697 2506 12727
rect 2478 12671 2479 12697
rect 2505 12671 2506 12697
rect 2422 12362 2450 12367
rect 2478 12362 2506 12671
rect 2534 12362 2562 12367
rect 2422 12361 2534 12362
rect 2422 12335 2423 12361
rect 2449 12335 2534 12361
rect 2422 12334 2534 12335
rect 2422 12329 2450 12334
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2478 11969 2506 12334
rect 2534 12296 2562 12334
rect 2478 11943 2479 11969
rect 2505 11943 2506 11969
rect 2478 11913 2506 11943
rect 2478 11887 2479 11913
rect 2505 11887 2506 11913
rect 2422 11578 2450 11583
rect 2478 11578 2506 11887
rect 2534 11578 2562 11583
rect 2422 11577 2562 11578
rect 2422 11551 2423 11577
rect 2449 11551 2535 11577
rect 2561 11551 2562 11577
rect 2422 11550 2562 11551
rect 2422 11545 2450 11550
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2478 11185 2506 11550
rect 2534 11545 2562 11550
rect 2478 11159 2479 11185
rect 2505 11159 2506 11185
rect 2478 11130 2506 11159
rect 2478 11129 2562 11130
rect 2478 11103 2479 11129
rect 2505 11103 2562 11129
rect 2478 11102 2562 11103
rect 2478 11097 2506 11102
rect 2422 10794 2450 10799
rect 2534 10794 2562 11102
rect 2422 10793 2562 10794
rect 2422 10767 2423 10793
rect 2449 10767 2535 10793
rect 2561 10767 2562 10793
rect 2422 10766 2562 10767
rect 2422 10761 2450 10766
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2478 10401 2506 10766
rect 2534 10761 2562 10766
rect 2478 10375 2479 10401
rect 2505 10375 2506 10401
rect 2478 10345 2506 10375
rect 2478 10319 2479 10345
rect 2505 10319 2506 10345
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 2478 9617 2506 10319
rect 2478 9591 2479 9617
rect 2505 9591 2506 9617
rect 2478 9561 2506 9591
rect 2478 9535 2479 9561
rect 2505 9535 2506 9561
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 1918 8441 1946 8447
rect 1918 8415 1919 8441
rect 1945 8415 1946 8441
rect 1918 8050 1946 8415
rect 1918 7658 1946 8022
rect 1918 7625 1946 7630
rect 2086 7266 2114 8470
rect 2478 8833 2506 9535
rect 2478 8807 2479 8833
rect 2505 8807 2506 8833
rect 2478 8777 2506 8807
rect 2478 8751 2479 8777
rect 2505 8751 2506 8777
rect 2478 8442 2506 8751
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 2478 8049 2506 8414
rect 2478 8023 2479 8049
rect 2505 8023 2506 8049
rect 2478 7993 2506 8023
rect 2478 7967 2479 7993
rect 2505 7967 2506 7993
rect 2478 7961 2506 7967
rect 2142 7658 2170 7663
rect 2142 7611 2170 7630
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 2086 6873 2114 7238
rect 2478 7266 2506 7271
rect 2590 7266 2618 13902
rect 3598 13929 3626 14687
rect 3598 13903 3599 13929
rect 3625 13903 3626 13929
rect 3598 13145 3626 13903
rect 3598 13119 3599 13145
rect 3625 13119 3626 13145
rect 3598 12474 3626 13119
rect 4046 15889 4074 15946
rect 4046 15863 4047 15889
rect 4073 15863 4074 15889
rect 4046 15105 4074 15863
rect 4270 15946 4466 15974
rect 5278 16281 5306 16647
rect 5278 16255 5279 16281
rect 5305 16255 5306 16281
rect 4270 15890 4298 15946
rect 4494 15890 4522 15895
rect 4270 15889 4522 15890
rect 4270 15863 4271 15889
rect 4297 15863 4495 15889
rect 4521 15863 4522 15889
rect 4270 15862 4522 15863
rect 4270 15857 4298 15862
rect 4494 15553 4522 15862
rect 4494 15527 4495 15553
rect 4521 15527 4522 15553
rect 4494 15497 4522 15527
rect 4494 15471 4495 15497
rect 4521 15471 4522 15497
rect 4046 15079 4047 15105
rect 4073 15079 4074 15105
rect 4046 14321 4074 15079
rect 4382 15106 4410 15111
rect 4494 15106 4522 15471
rect 4382 15105 4522 15106
rect 4382 15079 4383 15105
rect 4409 15079 4495 15105
rect 4521 15079 4522 15105
rect 4382 15078 4522 15079
rect 4382 15073 4410 15078
rect 4494 14769 4522 15078
rect 4494 14743 4495 14769
rect 4521 14743 4522 14769
rect 4494 14713 4522 14743
rect 5278 15889 5306 16255
rect 6398 18633 6426 18663
rect 6398 18607 6399 18633
rect 6425 18607 6426 18633
rect 6398 18241 6426 18607
rect 6958 19809 6986 19815
rect 6958 19783 6959 19809
rect 6985 19783 6986 19809
rect 6958 19417 6986 19783
rect 7350 19810 7378 19815
rect 7574 19810 7602 20510
rect 7686 20202 7714 20510
rect 7798 20505 7826 20510
rect 7910 20202 7938 20207
rect 7686 20201 7938 20202
rect 7686 20175 7687 20201
rect 7713 20175 7911 20201
rect 7937 20175 7938 20201
rect 7686 20174 7938 20175
rect 7686 20169 7714 20174
rect 7910 20169 7938 20174
rect 7350 19809 7602 19810
rect 7350 19783 7351 19809
rect 7377 19783 7575 19809
rect 7601 19783 7602 19809
rect 7350 19782 7602 19783
rect 6958 19391 6959 19417
rect 6985 19391 6986 19417
rect 6958 18634 6986 19391
rect 7238 19418 7266 19423
rect 7350 19418 7378 19782
rect 7238 19417 7378 19418
rect 7238 19391 7239 19417
rect 7265 19391 7351 19417
rect 7377 19391 7378 19417
rect 7238 19390 7378 19391
rect 7238 19385 7266 19390
rect 7126 19025 7154 19031
rect 7126 18999 7127 19025
rect 7153 18999 7154 19025
rect 7126 18634 7154 18999
rect 7350 19025 7378 19390
rect 7350 18999 7351 19025
rect 7377 18999 7378 19025
rect 6958 18633 7154 18634
rect 6958 18607 6959 18633
rect 6985 18607 7154 18633
rect 6958 18606 7154 18607
rect 6958 18601 6986 18606
rect 6398 18215 6399 18241
rect 6425 18215 6426 18241
rect 6398 18185 6426 18215
rect 6398 18159 6399 18185
rect 6425 18159 6426 18185
rect 6398 17905 6426 18159
rect 6398 17879 6399 17905
rect 6425 17879 6426 17905
rect 6398 17850 6426 17879
rect 7126 18241 7154 18606
rect 7238 18634 7266 18639
rect 7350 18634 7378 18999
rect 7574 19025 7602 19782
rect 8582 19810 8610 20567
rect 8582 19763 8610 19782
rect 8750 21378 8778 21383
rect 8974 21378 9002 21383
rect 8750 21377 9002 21378
rect 8750 21351 8751 21377
rect 8777 21351 8975 21377
rect 9001 21351 9002 21377
rect 8750 21350 9002 21351
rect 8750 20594 8778 21350
rect 8974 21345 9002 21350
rect 9142 20985 9170 21743
rect 9142 20959 9143 20985
rect 9169 20959 9170 20985
rect 8974 20594 9002 20599
rect 8750 20593 9002 20594
rect 8750 20567 8751 20593
rect 8777 20567 8975 20593
rect 9001 20567 9002 20593
rect 8750 20566 9002 20567
rect 8750 19810 8778 20566
rect 8974 20561 9002 20566
rect 9142 20201 9170 20959
rect 9142 20175 9143 20201
rect 9169 20175 9170 20201
rect 8974 19810 9002 19815
rect 8750 19809 9002 19810
rect 8750 19783 8751 19809
rect 8777 19783 8975 19809
rect 9001 19783 9002 19809
rect 8750 19782 9002 19783
rect 7574 18999 7575 19025
rect 7601 18999 7602 19025
rect 7574 18993 7602 18999
rect 8414 19025 8442 19031
rect 8414 18999 8415 19025
rect 8441 18999 8442 19025
rect 7238 18633 7378 18634
rect 7238 18607 7239 18633
rect 7265 18607 7351 18633
rect 7377 18607 7378 18633
rect 7238 18606 7378 18607
rect 7238 18601 7266 18606
rect 7126 18215 7127 18241
rect 7153 18215 7154 18241
rect 6398 17457 6426 17822
rect 6958 17850 6986 17855
rect 7126 17850 7154 18215
rect 7350 18242 7378 18606
rect 7574 18242 7602 18247
rect 7350 18241 7574 18242
rect 7350 18215 7351 18241
rect 7377 18215 7574 18241
rect 7350 18214 7574 18215
rect 6958 17849 7154 17850
rect 6958 17823 6959 17849
rect 6985 17823 7154 17849
rect 6958 17822 7154 17823
rect 6958 17817 6986 17822
rect 6398 17431 6399 17457
rect 6425 17431 6426 17457
rect 6398 17401 6426 17431
rect 6398 17375 6399 17401
rect 6425 17375 6426 17401
rect 6398 17121 6426 17375
rect 6398 17095 6399 17121
rect 6425 17095 6426 17121
rect 6398 17065 6426 17095
rect 7126 17457 7154 17822
rect 7182 17850 7210 17855
rect 7350 17850 7378 18214
rect 7574 18176 7602 18214
rect 8414 18241 8442 18999
rect 8414 18215 8415 18241
rect 8441 18215 8442 18241
rect 7210 17849 7378 17850
rect 7210 17823 7351 17849
rect 7377 17823 7378 17849
rect 7210 17822 7378 17823
rect 7182 17803 7210 17822
rect 7350 17817 7378 17822
rect 8414 17850 8442 18215
rect 8750 19026 8778 19782
rect 8974 19777 9002 19782
rect 9142 19810 9170 20175
rect 9142 19418 9170 19782
rect 9142 19371 9170 19390
rect 9310 20986 9338 20991
rect 9422 20986 9450 23310
rect 9534 23305 9562 23310
rect 9478 22945 9506 22951
rect 9478 22919 9479 22945
rect 9505 22919 9506 22945
rect 9478 22889 9506 22919
rect 9478 22863 9479 22889
rect 9505 22863 9506 22889
rect 9478 22554 9506 22863
rect 9478 22162 9506 22526
rect 9478 22105 9506 22134
rect 9478 22079 9479 22105
rect 9505 22079 9506 22105
rect 9478 22073 9506 22079
rect 9814 22609 9842 24095
rect 9918 23534 10050 23539
rect 9946 23506 9970 23534
rect 9998 23506 10022 23534
rect 9918 23501 10050 23506
rect 10598 23338 10626 23343
rect 10374 23282 10402 23287
rect 9918 22750 10050 22755
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 9918 22717 10050 22722
rect 9814 22583 9815 22609
rect 9841 22583 9842 22609
rect 9814 22553 9842 22583
rect 9814 22527 9815 22553
rect 9841 22527 9842 22553
rect 9814 22162 9842 22527
rect 9814 21882 9842 22134
rect 10374 22553 10402 23254
rect 10598 22946 10626 23310
rect 10598 22913 10626 22918
rect 10374 22527 10375 22553
rect 10401 22527 10402 22553
rect 9918 21966 10050 21971
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 9918 21933 10050 21938
rect 10038 21882 10066 21887
rect 9814 21849 9842 21854
rect 9982 21826 10066 21854
rect 9982 21825 10010 21826
rect 9982 21799 9983 21825
rect 10009 21799 10010 21825
rect 9982 21769 10010 21799
rect 9982 21743 9983 21769
rect 10009 21743 10010 21769
rect 9982 21737 10010 21743
rect 10374 21770 10402 22527
rect 10374 21737 10402 21742
rect 10598 21770 10626 21775
rect 10598 21723 10626 21742
rect 9918 21182 10050 21187
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 9918 21149 10050 21154
rect 9534 21042 9562 21047
rect 9534 20986 9562 21014
rect 9310 20985 9562 20986
rect 9310 20959 9311 20985
rect 9337 20959 9535 20985
rect 9561 20959 9562 20985
rect 9310 20958 9562 20959
rect 9310 20202 9338 20958
rect 9534 20953 9562 20958
rect 10598 20985 10626 20991
rect 10598 20959 10599 20985
rect 10625 20959 10626 20985
rect 9918 20398 10050 20403
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 9918 20365 10050 20370
rect 9534 20202 9562 20207
rect 9310 20201 9562 20202
rect 9310 20175 9311 20201
rect 9337 20175 9535 20201
rect 9561 20175 9562 20201
rect 9310 20174 9562 20175
rect 9310 19418 9338 20174
rect 9534 20169 9562 20174
rect 10598 20201 10626 20959
rect 10598 20175 10599 20201
rect 10625 20175 10626 20201
rect 9918 19614 10050 19619
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 9918 19581 10050 19586
rect 9534 19418 9562 19423
rect 9310 19417 9562 19418
rect 9310 19391 9311 19417
rect 9337 19391 9535 19417
rect 9561 19391 9562 19417
rect 9310 19390 9562 19391
rect 8974 19026 9002 19031
rect 8750 19025 9002 19026
rect 8750 18999 8751 19025
rect 8777 18999 8975 19025
rect 9001 18999 9002 19025
rect 8750 18998 9002 18999
rect 8750 18242 8778 18998
rect 8974 18993 9002 18998
rect 8750 18195 8778 18214
rect 8862 18633 8890 18639
rect 8862 18607 8863 18633
rect 8889 18607 8890 18633
rect 8862 17850 8890 18607
rect 9310 18634 9338 19390
rect 9534 19385 9562 19390
rect 10598 19418 10626 20175
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9534 18634 9562 18639
rect 9310 18633 9562 18634
rect 9310 18607 9311 18633
rect 9337 18607 9535 18633
rect 9561 18607 9562 18633
rect 9310 18606 9562 18607
rect 8974 18242 9002 18247
rect 8974 18195 9002 18214
rect 9310 18242 9338 18606
rect 9534 18601 9562 18606
rect 10598 18633 10626 19390
rect 10598 18607 10599 18633
rect 10625 18607 10626 18633
rect 8414 17849 8890 17850
rect 8414 17823 8863 17849
rect 8889 17823 8890 17849
rect 8414 17822 8890 17823
rect 7126 17431 7127 17457
rect 7153 17431 7154 17457
rect 6398 17039 6399 17065
rect 6425 17039 6426 17065
rect 6398 16673 6426 17039
rect 6958 17066 6986 17071
rect 7126 17066 7154 17431
rect 6958 17065 7154 17066
rect 6958 17039 6959 17065
rect 6985 17039 7154 17065
rect 6958 17038 7154 17039
rect 6958 17033 6986 17038
rect 6398 16647 6399 16673
rect 6425 16647 6426 16673
rect 6398 16617 6426 16647
rect 6398 16591 6399 16617
rect 6425 16591 6426 16617
rect 6398 16337 6426 16591
rect 6398 16311 6399 16337
rect 6425 16311 6426 16337
rect 6398 16281 6426 16311
rect 7126 16673 7154 17038
rect 7126 16647 7127 16673
rect 7153 16647 7154 16673
rect 6398 16255 6399 16281
rect 6425 16255 6426 16281
rect 6398 15974 6426 16255
rect 6958 16282 6986 16287
rect 7126 16282 7154 16647
rect 6958 16281 7154 16282
rect 6958 16255 6959 16281
rect 6985 16255 7154 16281
rect 6958 16254 7154 16255
rect 6958 16249 6986 16254
rect 6230 15946 6426 15974
rect 7126 16002 7154 16254
rect 5278 15863 5279 15889
rect 5305 15863 5306 15889
rect 5278 15497 5306 15863
rect 5278 15471 5279 15497
rect 5305 15471 5306 15497
rect 5278 15105 5306 15471
rect 5278 15079 5279 15105
rect 5305 15079 5306 15105
rect 4494 14687 4495 14713
rect 4521 14687 4522 14713
rect 4046 14295 4047 14321
rect 4073 14295 4074 14321
rect 4046 13537 4074 14295
rect 4382 14322 4410 14327
rect 4494 14322 4522 14687
rect 4410 14321 4522 14322
rect 4410 14295 4495 14321
rect 4521 14295 4522 14321
rect 4410 14294 4522 14295
rect 4382 14256 4410 14294
rect 4494 13985 4522 14294
rect 4494 13959 4495 13985
rect 4521 13959 4522 13985
rect 4494 13929 4522 13959
rect 4494 13903 4495 13929
rect 4521 13903 4522 13929
rect 4046 13511 4047 13537
rect 4073 13511 4074 13537
rect 4046 12753 4074 13511
rect 4382 13538 4410 13543
rect 4494 13538 4522 13903
rect 4382 13537 4522 13538
rect 4382 13511 4383 13537
rect 4409 13511 4495 13537
rect 4521 13511 4522 13537
rect 4382 13510 4522 13511
rect 4382 13505 4410 13510
rect 4494 13201 4522 13510
rect 4494 13175 4495 13201
rect 4521 13175 4522 13201
rect 4494 13145 4522 13175
rect 4494 13119 4495 13145
rect 4521 13119 4522 13145
rect 4046 12727 4047 12753
rect 4073 12727 4074 12753
rect 4046 12474 4074 12727
rect 4382 12754 4410 12759
rect 4494 12754 4522 13119
rect 4382 12753 4522 12754
rect 4382 12727 4383 12753
rect 4409 12727 4495 12753
rect 4521 12727 4522 12753
rect 4382 12726 4522 12727
rect 4382 12721 4410 12726
rect 4494 12721 4522 12726
rect 5222 14714 5250 14719
rect 5278 14714 5306 15079
rect 6174 15889 6202 15895
rect 6174 15863 6175 15889
rect 6201 15863 6202 15889
rect 6174 15834 6202 15863
rect 6230 15834 6258 15946
rect 6174 15833 6258 15834
rect 6174 15807 6231 15833
rect 6257 15807 6258 15833
rect 6174 15806 6258 15807
rect 6174 15553 6202 15806
rect 6230 15801 6258 15806
rect 7126 15889 7154 15974
rect 7798 17457 7826 17463
rect 7798 17431 7799 17457
rect 7825 17431 7826 17457
rect 7798 17401 7826 17431
rect 7798 17375 7799 17401
rect 7825 17375 7826 17401
rect 7798 17121 7826 17375
rect 7798 17095 7799 17121
rect 7825 17095 7826 17121
rect 7798 17065 7826 17095
rect 7798 17039 7799 17065
rect 7825 17039 7826 17065
rect 7798 16673 7826 17039
rect 7798 16647 7799 16673
rect 7825 16647 7826 16673
rect 7798 16617 7826 16647
rect 7798 16591 7799 16617
rect 7825 16591 7826 16617
rect 7798 16337 7826 16591
rect 7798 16311 7799 16337
rect 7825 16311 7826 16337
rect 7798 16281 7826 16311
rect 7798 16255 7799 16281
rect 7825 16255 7826 16281
rect 7126 15863 7127 15889
rect 7153 15863 7154 15889
rect 6174 15527 6175 15553
rect 6201 15527 6202 15553
rect 6174 15497 6202 15527
rect 6174 15471 6175 15497
rect 6201 15471 6202 15497
rect 6174 15105 6202 15471
rect 6174 15079 6175 15105
rect 6201 15079 6202 15105
rect 6174 15050 6202 15079
rect 6958 15498 6986 15503
rect 7126 15498 7154 15863
rect 6958 15497 7154 15498
rect 6958 15471 6959 15497
rect 6985 15471 7154 15497
rect 6958 15470 7154 15471
rect 7630 15889 7658 15895
rect 7630 15863 7631 15889
rect 7657 15863 7658 15889
rect 7630 15834 7658 15863
rect 7798 15834 7826 16255
rect 7630 15833 7826 15834
rect 7630 15807 7799 15833
rect 7825 15807 7826 15833
rect 7630 15806 7826 15807
rect 7630 15553 7658 15806
rect 7798 15801 7826 15806
rect 8414 17457 8442 17822
rect 8862 17817 8890 17822
rect 9310 17850 9338 18214
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9534 17850 9562 17855
rect 9310 17849 9562 17850
rect 9310 17823 9311 17849
rect 9337 17823 9535 17849
rect 9561 17823 9562 17849
rect 9310 17822 9562 17823
rect 9310 17817 9338 17822
rect 9534 17817 9562 17822
rect 10598 17850 10626 18607
rect 10598 17803 10626 17822
rect 8414 17431 8415 17457
rect 8441 17431 8442 17457
rect 8414 16673 8442 17431
rect 9310 17457 9338 17463
rect 9310 17431 9311 17457
rect 9337 17431 9338 17457
rect 9310 17401 9338 17431
rect 9310 17375 9311 17401
rect 9337 17375 9338 17401
rect 8414 16647 8415 16673
rect 8441 16647 8442 16673
rect 8414 16002 8442 16647
rect 8414 15889 8442 15974
rect 8862 17065 8890 17071
rect 8862 17039 8863 17065
rect 8889 17039 8890 17065
rect 8862 16281 8890 17039
rect 8862 16255 8863 16281
rect 8889 16255 8890 16281
rect 8414 15863 8415 15889
rect 8441 15863 8442 15889
rect 7630 15527 7631 15553
rect 7657 15527 7658 15553
rect 7630 15497 7658 15527
rect 7630 15471 7631 15497
rect 7657 15471 7658 15497
rect 6958 15105 6986 15470
rect 6958 15079 6959 15105
rect 6985 15079 6986 15105
rect 6230 15050 6258 15055
rect 6174 15049 6258 15050
rect 6174 15023 6231 15049
rect 6257 15023 6258 15049
rect 6174 15022 6258 15023
rect 6174 14769 6202 15022
rect 6230 15017 6258 15022
rect 6174 14743 6175 14769
rect 6201 14743 6202 14769
rect 5222 14713 5306 14714
rect 5222 14687 5223 14713
rect 5249 14687 5306 14713
rect 5222 14686 5306 14687
rect 5950 14714 5978 14719
rect 6174 14714 6202 14743
rect 5950 14713 6202 14714
rect 5950 14687 5951 14713
rect 5977 14687 6202 14713
rect 5950 14686 6202 14687
rect 6958 14713 6986 15079
rect 6958 14687 6959 14713
rect 6985 14687 6986 14713
rect 5222 14322 5250 14686
rect 5278 14322 5306 14327
rect 5222 14321 5306 14322
rect 5222 14295 5279 14321
rect 5305 14295 5306 14321
rect 5222 14294 5306 14295
rect 5222 13929 5250 14294
rect 5278 14289 5306 14294
rect 5838 14322 5866 14327
rect 5894 14322 5922 14327
rect 5950 14322 5978 14686
rect 5838 14321 5894 14322
rect 5838 14295 5839 14321
rect 5865 14295 5894 14321
rect 5838 14294 5894 14295
rect 5922 14321 5978 14322
rect 5922 14295 5951 14321
rect 5977 14295 5978 14321
rect 5922 14294 5978 14295
rect 5838 14289 5866 14294
rect 5222 13903 5223 13929
rect 5249 13903 5250 13929
rect 5222 13538 5250 13903
rect 5782 13930 5810 13935
rect 5894 13930 5922 14294
rect 5950 14289 5978 14294
rect 6958 14321 6986 14687
rect 6958 14295 6959 14321
rect 6985 14295 6986 14321
rect 5782 13929 5922 13930
rect 5782 13903 5783 13929
rect 5809 13903 5895 13929
rect 5921 13903 5922 13929
rect 5782 13902 5922 13903
rect 5782 13897 5810 13902
rect 5278 13538 5306 13543
rect 5222 13537 5306 13538
rect 5222 13511 5279 13537
rect 5305 13511 5306 13537
rect 5222 13510 5306 13511
rect 5222 13145 5250 13510
rect 5278 13505 5306 13510
rect 5838 13538 5866 13543
rect 5894 13538 5922 13902
rect 6958 13929 6986 14295
rect 6958 13903 6959 13929
rect 6985 13903 6986 13929
rect 5950 13538 5978 13543
rect 5838 13537 5978 13538
rect 5838 13511 5839 13537
rect 5865 13511 5951 13537
rect 5977 13511 5978 13537
rect 5838 13510 5978 13511
rect 5838 13505 5866 13510
rect 5222 13119 5223 13145
rect 5249 13119 5250 13145
rect 5222 12754 5250 13119
rect 5782 13146 5810 13151
rect 5894 13146 5922 13510
rect 5950 13505 5978 13510
rect 6958 13537 6986 13903
rect 6958 13511 6959 13537
rect 6985 13511 6986 13537
rect 5782 13145 5922 13146
rect 5782 13119 5783 13145
rect 5809 13119 5895 13145
rect 5921 13119 5922 13145
rect 5782 13118 5922 13119
rect 5782 13113 5810 13118
rect 5278 12754 5306 12759
rect 5222 12753 5306 12754
rect 5222 12727 5279 12753
rect 5305 12727 5306 12753
rect 5222 12726 5306 12727
rect 3598 12446 4074 12474
rect 3598 12361 3626 12446
rect 3598 12335 3599 12361
rect 3625 12335 3626 12361
rect 3598 12329 3626 12335
rect 3766 12362 3794 12367
rect 3766 12315 3794 12334
rect 3990 12362 4018 12367
rect 3990 12315 4018 12334
rect 4046 11970 4074 12446
rect 4158 12362 4186 12367
rect 4186 12334 4802 12362
rect 4158 12329 4186 12334
rect 4102 11970 4130 11975
rect 4046 11942 4102 11970
rect 4102 11923 4130 11942
rect 4214 11970 4242 11975
rect 3318 11578 3346 11583
rect 3318 11186 3346 11550
rect 3878 11578 3906 11583
rect 3990 11578 4018 11583
rect 3878 11577 4018 11578
rect 3878 11551 3879 11577
rect 3905 11551 3991 11577
rect 4017 11551 4018 11577
rect 3878 11550 4018 11551
rect 3878 11545 3906 11550
rect 3318 11185 3402 11186
rect 3318 11159 3319 11185
rect 3345 11159 3402 11185
rect 3318 11158 3402 11159
rect 3318 11153 3346 11158
rect 3374 11130 3402 11158
rect 3374 10793 3402 11102
rect 3990 11185 4018 11550
rect 3990 11159 3991 11185
rect 4017 11159 4018 11185
rect 3990 11130 4018 11159
rect 4102 11186 4130 11191
rect 4102 11130 4130 11158
rect 3990 11129 4130 11130
rect 3990 11103 4103 11129
rect 4129 11103 4130 11129
rect 3990 11102 4130 11103
rect 3374 10767 3375 10793
rect 3401 10767 3402 10793
rect 3374 10401 3402 10767
rect 3878 10794 3906 10799
rect 3990 10794 4018 11102
rect 4102 11097 4130 11102
rect 4214 11130 4242 11942
rect 4774 11969 4802 12334
rect 4774 11943 4775 11969
rect 4801 11943 4802 11969
rect 4774 11913 4802 11943
rect 4774 11887 4775 11913
rect 4801 11887 4802 11913
rect 4774 11881 4802 11887
rect 5222 12361 5250 12726
rect 5278 12721 5306 12726
rect 5838 12754 5866 12759
rect 5894 12754 5922 13118
rect 6958 13145 6986 13511
rect 6958 13119 6959 13145
rect 6985 13119 6986 13145
rect 5950 12754 5978 12759
rect 5838 12753 5978 12754
rect 5838 12727 5839 12753
rect 5865 12727 5951 12753
rect 5977 12727 5978 12753
rect 5838 12726 5978 12727
rect 5838 12721 5866 12726
rect 5222 12335 5223 12361
rect 5249 12335 5250 12361
rect 5222 11970 5250 12335
rect 5950 12418 5978 12726
rect 6958 12753 6986 13119
rect 6958 12727 6959 12753
rect 6985 12727 6986 12753
rect 6174 12418 6202 12423
rect 5950 12417 6202 12418
rect 5950 12391 6175 12417
rect 6201 12391 6202 12417
rect 5950 12390 6202 12391
rect 5950 12361 5978 12390
rect 6174 12385 6202 12390
rect 5950 12335 5951 12361
rect 5977 12335 5978 12361
rect 5278 11970 5306 11975
rect 5222 11969 5306 11970
rect 5222 11943 5279 11969
rect 5305 11943 5306 11969
rect 5222 11942 5306 11943
rect 5222 11577 5250 11942
rect 5278 11937 5306 11942
rect 5838 11970 5866 11975
rect 5950 11970 5978 12335
rect 5838 11969 5978 11970
rect 5838 11943 5839 11969
rect 5865 11943 5951 11969
rect 5977 11943 5978 11969
rect 5838 11942 5978 11943
rect 5838 11937 5866 11942
rect 5222 11551 5223 11577
rect 5249 11551 5250 11577
rect 4214 11097 4242 11102
rect 4662 11185 4690 11191
rect 4662 11159 4663 11185
rect 4689 11159 4690 11185
rect 4662 11130 4690 11159
rect 5054 11186 5082 11191
rect 5054 11139 5082 11158
rect 3878 10793 4018 10794
rect 3878 10767 3879 10793
rect 3905 10767 3991 10793
rect 4017 10767 4018 10793
rect 3878 10766 4018 10767
rect 3878 10761 3906 10766
rect 3374 10375 3375 10401
rect 3401 10375 3402 10401
rect 3038 10065 3066 10071
rect 3038 10039 3039 10065
rect 3065 10039 3066 10065
rect 3038 10010 3066 10039
rect 3038 9963 3066 9982
rect 3374 10009 3402 10375
rect 3374 9983 3375 10009
rect 3401 9983 3402 10009
rect 3374 9977 3402 9983
rect 3766 10401 3794 10407
rect 3766 10375 3767 10401
rect 3793 10375 3794 10401
rect 3766 10010 3794 10375
rect 3990 10401 4018 10766
rect 3990 10375 3991 10401
rect 4017 10375 4018 10401
rect 3990 10010 4018 10375
rect 4662 10401 4690 11102
rect 5222 11130 5250 11551
rect 5950 11634 5978 11942
rect 6342 12362 6370 12367
rect 6174 11802 6202 11807
rect 6174 11634 6202 11774
rect 5950 11633 6202 11634
rect 5950 11607 6175 11633
rect 6201 11607 6202 11633
rect 5950 11606 6202 11607
rect 5950 11577 5978 11606
rect 6174 11601 6202 11606
rect 5950 11551 5951 11577
rect 5977 11551 5978 11577
rect 5950 11545 5978 11551
rect 5278 11186 5306 11191
rect 5278 11139 5306 11158
rect 5222 11097 5250 11102
rect 5838 10849 5866 10855
rect 5838 10823 5839 10849
rect 5865 10823 5866 10849
rect 4662 10375 4663 10401
rect 4689 10375 4690 10401
rect 4662 10094 4690 10375
rect 4886 10793 4914 10799
rect 4886 10767 4887 10793
rect 4913 10767 4914 10793
rect 4886 10094 4914 10767
rect 5838 10793 5866 10823
rect 5838 10767 5839 10793
rect 5865 10767 5866 10793
rect 5110 10401 5138 10407
rect 5838 10402 5866 10767
rect 5110 10375 5111 10401
rect 5137 10375 5138 10401
rect 4662 10066 5026 10094
rect 3794 10009 4018 10010
rect 3794 9983 3991 10009
rect 4017 9983 4018 10009
rect 3794 9982 4018 9983
rect 3318 9617 3346 9623
rect 3318 9591 3319 9617
rect 3345 9591 3346 9617
rect 3318 9562 3346 9591
rect 3654 9618 3682 9623
rect 3766 9618 3794 9982
rect 3990 9977 4018 9982
rect 4998 10009 5026 10066
rect 4998 9983 4999 10009
rect 5025 9983 5026 10009
rect 3654 9617 3794 9618
rect 3654 9591 3655 9617
rect 3681 9591 3767 9617
rect 3793 9591 3794 9617
rect 3654 9590 3794 9591
rect 3654 9585 3682 9590
rect 2814 9281 2842 9287
rect 2814 9255 2815 9281
rect 2841 9255 2842 9281
rect 2814 9225 2842 9255
rect 2814 9199 2815 9225
rect 2841 9199 2842 9225
rect 2814 8497 2842 9199
rect 2814 8471 2815 8497
rect 2841 8471 2842 8497
rect 2814 8442 2842 8471
rect 3318 9282 3346 9534
rect 3318 9225 3346 9254
rect 3766 9282 3794 9590
rect 4942 9618 4970 9623
rect 4998 9618 5026 9983
rect 4942 9617 5026 9618
rect 4942 9591 4943 9617
rect 4969 9591 5026 9617
rect 4942 9590 5026 9591
rect 4942 9585 4970 9590
rect 3318 9199 3319 9225
rect 3345 9199 3346 9225
rect 3318 8833 3346 9199
rect 3318 8807 3319 8833
rect 3345 8807 3346 8833
rect 2814 8395 2842 8414
rect 3038 8442 3066 8447
rect 3038 7713 3066 8414
rect 3318 8441 3346 8807
rect 3318 8415 3319 8441
rect 3345 8415 3346 8441
rect 3318 8049 3346 8415
rect 3654 9226 3682 9231
rect 3766 9226 3794 9254
rect 3654 9225 3794 9226
rect 3654 9199 3655 9225
rect 3681 9199 3767 9225
rect 3793 9199 3794 9225
rect 3654 9198 3794 9199
rect 3654 8834 3682 9198
rect 3766 9193 3794 9198
rect 4998 9225 5026 9590
rect 4998 9199 4999 9225
rect 5025 9199 5026 9225
rect 3766 8834 3794 8839
rect 3654 8833 3794 8834
rect 3654 8807 3655 8833
rect 3681 8807 3767 8833
rect 3793 8807 3794 8833
rect 3654 8806 3794 8807
rect 3654 8442 3682 8806
rect 3766 8801 3794 8806
rect 4942 8834 4970 8839
rect 4998 8834 5026 9199
rect 4942 8833 5026 8834
rect 4942 8807 4943 8833
rect 4969 8807 5026 8833
rect 4942 8806 5026 8807
rect 4942 8801 4970 8806
rect 3766 8442 3794 8447
rect 3682 8441 3794 8442
rect 3682 8415 3767 8441
rect 3793 8415 3794 8441
rect 3682 8414 3794 8415
rect 3318 8023 3319 8049
rect 3345 8023 3346 8049
rect 3318 8017 3346 8023
rect 3598 8386 3626 8391
rect 3038 7687 3039 7713
rect 3065 7687 3066 7713
rect 3038 7657 3066 7687
rect 3038 7631 3039 7657
rect 3065 7631 3066 7657
rect 3038 7625 3066 7631
rect 3598 7658 3626 8358
rect 3654 8050 3682 8414
rect 3766 8409 3794 8414
rect 4998 8441 5026 8806
rect 5110 9617 5138 10375
rect 5334 10401 5866 10402
rect 5334 10375 5839 10401
rect 5865 10375 5866 10401
rect 5334 10374 5866 10375
rect 5334 10094 5362 10374
rect 5838 10369 5866 10374
rect 5334 10066 5474 10094
rect 5446 10010 5474 10066
rect 5558 10010 5586 10015
rect 5446 10009 5586 10010
rect 5446 9983 5447 10009
rect 5473 9983 5559 10009
rect 5585 9983 5586 10009
rect 5446 9982 5586 9983
rect 5446 9977 5474 9982
rect 5110 9591 5111 9617
rect 5137 9591 5138 9617
rect 5110 9282 5138 9591
rect 5110 8833 5138 9254
rect 5558 9617 5586 9982
rect 5558 9591 5559 9617
rect 5585 9591 5586 9617
rect 5446 9226 5474 9231
rect 5558 9226 5586 9591
rect 6342 10009 6370 12334
rect 6958 12361 6986 12727
rect 7630 15105 7658 15471
rect 7630 15079 7631 15105
rect 7657 15079 7658 15105
rect 7630 15050 7658 15079
rect 8414 15105 8442 15863
rect 8414 15079 8415 15105
rect 8441 15079 8442 15105
rect 7798 15050 7826 15055
rect 7630 15049 7826 15050
rect 7630 15023 7799 15049
rect 7825 15023 7826 15049
rect 7630 15022 7826 15023
rect 7630 14769 7658 15022
rect 7798 15017 7826 15022
rect 7630 14743 7631 14769
rect 7657 14743 7658 14769
rect 7630 14713 7658 14743
rect 7630 14687 7631 14713
rect 7657 14687 7658 14713
rect 7630 14321 7658 14687
rect 7630 14295 7631 14321
rect 7657 14295 7658 14321
rect 7630 14266 7658 14295
rect 8414 14321 8442 15079
rect 8414 14295 8415 14321
rect 8441 14295 8442 14321
rect 7798 14266 7826 14271
rect 7630 14265 7826 14266
rect 7630 14239 7799 14265
rect 7825 14239 7826 14265
rect 7630 14238 7826 14239
rect 7630 13985 7658 14238
rect 7798 14233 7826 14238
rect 7630 13959 7631 13985
rect 7657 13959 7658 13985
rect 7630 13929 7658 13959
rect 7630 13903 7631 13929
rect 7657 13903 7658 13929
rect 7630 13537 7658 13903
rect 7630 13511 7631 13537
rect 7657 13511 7658 13537
rect 7630 13482 7658 13511
rect 8414 13537 8442 14295
rect 8414 13511 8415 13537
rect 8441 13511 8442 13537
rect 7798 13482 7826 13487
rect 7630 13481 7826 13482
rect 7630 13455 7799 13481
rect 7825 13455 7826 13481
rect 7630 13454 7826 13455
rect 7630 13201 7658 13454
rect 7798 13449 7826 13454
rect 7630 13175 7631 13201
rect 7657 13175 7658 13201
rect 7630 13145 7658 13175
rect 7630 13119 7631 13145
rect 7657 13119 7658 13145
rect 7630 12753 7658 13119
rect 7630 12727 7631 12753
rect 7657 12727 7658 12753
rect 7630 12698 7658 12727
rect 8414 12753 8442 13511
rect 8414 12727 8415 12753
rect 8441 12727 8442 12753
rect 7798 12698 7826 12703
rect 7630 12697 7826 12698
rect 7630 12671 7799 12697
rect 7825 12671 7826 12697
rect 7630 12670 7826 12671
rect 7630 12417 7658 12670
rect 7798 12665 7826 12670
rect 7630 12391 7631 12417
rect 7657 12391 7658 12417
rect 6958 12335 6959 12361
rect 6985 12335 6986 12361
rect 6958 11969 6986 12335
rect 6958 11943 6959 11969
rect 6985 11943 6986 11969
rect 6958 11577 6986 11943
rect 6958 11551 6959 11577
rect 6985 11551 6986 11577
rect 6958 11185 6986 11551
rect 6958 11159 6959 11185
rect 6985 11159 6986 11185
rect 6958 10793 6986 11159
rect 7574 12362 7602 12367
rect 7630 12362 7658 12391
rect 7574 12361 7658 12362
rect 7574 12335 7575 12361
rect 7601 12335 7658 12361
rect 7574 12334 7658 12335
rect 7574 11969 7602 12334
rect 7574 11943 7575 11969
rect 7601 11943 7602 11969
rect 7574 11802 7602 11943
rect 8414 12306 8442 12727
rect 8414 11969 8442 12278
rect 8806 15889 8834 15895
rect 8806 15863 8807 15889
rect 8833 15863 8834 15889
rect 8806 15105 8834 15863
rect 8806 15079 8807 15105
rect 8833 15079 8834 15105
rect 8806 14321 8834 15079
rect 8806 14295 8807 14321
rect 8833 14295 8834 14321
rect 8806 14266 8834 14295
rect 8806 13537 8834 14238
rect 8806 13511 8807 13537
rect 8833 13511 8834 13537
rect 8806 13482 8834 13511
rect 8806 12753 8834 13454
rect 8806 12727 8807 12753
rect 8833 12727 8834 12753
rect 8414 11943 8415 11969
rect 8441 11943 8442 11969
rect 7574 11634 7602 11774
rect 7798 11913 7826 11919
rect 7798 11887 7799 11913
rect 7825 11887 7826 11913
rect 7798 11802 7826 11887
rect 7630 11634 7658 11639
rect 7574 11633 7658 11634
rect 7574 11607 7631 11633
rect 7657 11607 7658 11633
rect 7574 11606 7658 11607
rect 7574 11577 7602 11606
rect 7630 11601 7658 11606
rect 7574 11551 7575 11577
rect 7601 11551 7602 11577
rect 7574 11185 7602 11551
rect 7574 11159 7575 11185
rect 7601 11159 7602 11185
rect 7574 11153 7602 11159
rect 6958 10767 6959 10793
rect 6985 10767 6986 10793
rect 6958 10402 6986 10767
rect 6342 9983 6343 10009
rect 6369 9983 6370 10009
rect 6342 9562 6370 9983
rect 6342 9529 6370 9534
rect 6846 10401 6986 10402
rect 6846 10375 6959 10401
rect 6985 10375 6986 10401
rect 6846 10374 6986 10375
rect 6846 9617 6874 10374
rect 6958 10369 6986 10374
rect 7798 11129 7826 11774
rect 7798 11103 7799 11129
rect 7825 11103 7826 11129
rect 7798 10849 7826 11103
rect 7798 10823 7799 10849
rect 7825 10823 7826 10849
rect 7798 10793 7826 10823
rect 7798 10767 7799 10793
rect 7825 10767 7826 10793
rect 7798 10401 7826 10767
rect 7798 10375 7799 10401
rect 7825 10375 7826 10401
rect 7798 10345 7826 10375
rect 7798 10319 7799 10345
rect 7825 10319 7826 10345
rect 7798 10313 7826 10319
rect 8414 11185 8442 11943
rect 8414 11159 8415 11185
rect 8441 11159 8442 11185
rect 8414 10401 8442 11159
rect 8750 11970 8778 11975
rect 8806 11970 8834 12727
rect 8862 15497 8890 16255
rect 9310 17066 9338 17375
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9534 17066 9562 17071
rect 9310 17065 9562 17066
rect 9310 17039 9311 17065
rect 9337 17039 9535 17065
rect 9561 17039 9562 17065
rect 9310 17038 9562 17039
rect 9310 16673 9338 17038
rect 9534 17033 9562 17038
rect 10598 17065 10626 17071
rect 10598 17039 10599 17065
rect 10625 17039 10626 17065
rect 9310 16647 9311 16673
rect 9337 16647 9338 16673
rect 9310 16617 9338 16647
rect 9310 16591 9311 16617
rect 9337 16591 9338 16617
rect 9310 16282 9338 16591
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9534 16282 9562 16287
rect 9310 16281 9562 16282
rect 9310 16255 9311 16281
rect 9337 16255 9535 16281
rect 9561 16255 9562 16281
rect 9310 16254 9562 16255
rect 8862 15471 8863 15497
rect 8889 15471 8890 15497
rect 8862 14713 8890 15471
rect 8862 14687 8863 14713
rect 8889 14687 8890 14713
rect 8862 13929 8890 14687
rect 8974 15889 9002 15895
rect 8974 15863 8975 15889
rect 9001 15863 9002 15889
rect 8974 15105 9002 15863
rect 8974 15079 8975 15105
rect 9001 15079 9002 15105
rect 8974 14321 9002 15079
rect 8974 14295 8975 14321
rect 9001 14295 9002 14321
rect 8974 14266 9002 14295
rect 8974 14233 9002 14238
rect 9310 15497 9338 16254
rect 9310 15471 9311 15497
rect 9337 15471 9338 15497
rect 9310 14714 9338 15471
rect 9478 15498 9506 16254
rect 9534 16249 9562 16254
rect 10598 16282 10626 17039
rect 10822 16673 10850 16679
rect 10822 16647 10823 16673
rect 10849 16647 10850 16673
rect 10822 16282 10850 16647
rect 10598 16281 10850 16282
rect 10598 16255 10599 16281
rect 10625 16255 10850 16281
rect 10598 16254 10850 16255
rect 10598 16249 10626 16254
rect 10822 15889 10850 16254
rect 10822 15863 10823 15889
rect 10849 15863 10850 15889
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9534 15498 9562 15503
rect 9478 15497 9562 15498
rect 9478 15471 9535 15497
rect 9561 15471 9562 15497
rect 9478 15470 9562 15471
rect 9534 15465 9562 15470
rect 10374 15497 10402 15503
rect 10374 15471 10375 15497
rect 10401 15471 10402 15497
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9534 14714 9562 14719
rect 9310 14713 9562 14714
rect 9310 14687 9311 14713
rect 9337 14687 9535 14713
rect 9561 14687 9562 14713
rect 9310 14686 9562 14687
rect 8862 13903 8863 13929
rect 8889 13903 8890 13929
rect 8862 13538 8890 13903
rect 9310 13930 9338 14686
rect 9534 14681 9562 14686
rect 10374 14713 10402 15471
rect 10374 14687 10375 14713
rect 10401 14687 10402 14713
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9534 13930 9562 13935
rect 9310 13929 9534 13930
rect 9310 13903 9311 13929
rect 9337 13903 9534 13929
rect 9310 13902 9534 13903
rect 8862 13145 8890 13510
rect 8974 13537 9002 13543
rect 8974 13511 8975 13537
rect 9001 13511 9002 13537
rect 8974 13482 9002 13511
rect 8974 13449 9002 13454
rect 8862 13119 8863 13145
rect 8889 13119 8890 13145
rect 8862 12361 8890 13119
rect 9310 13146 9338 13902
rect 9534 13864 9562 13902
rect 10374 13929 10402 14687
rect 10374 13903 10375 13929
rect 10401 13903 10402 13929
rect 10374 13538 10402 13903
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9534 13146 9562 13151
rect 9310 13145 9562 13146
rect 9310 13119 9311 13145
rect 9337 13119 9535 13145
rect 9561 13119 9562 13145
rect 9310 13118 9562 13119
rect 8862 12335 8863 12361
rect 8889 12335 8890 12361
rect 8862 12306 8890 12335
rect 8862 12273 8890 12278
rect 8974 12753 9002 12759
rect 8974 12727 8975 12753
rect 9001 12727 9002 12753
rect 8974 11970 9002 12727
rect 9310 12362 9338 13118
rect 9534 13113 9562 13118
rect 10374 13145 10402 13510
rect 10822 15105 10850 15863
rect 10822 15079 10823 15105
rect 10849 15079 10850 15105
rect 10822 14321 10850 15079
rect 10822 14295 10823 14321
rect 10849 14295 10850 14321
rect 10822 13538 10850 14295
rect 10822 13491 10850 13510
rect 10934 15498 10962 15503
rect 10374 13119 10375 13145
rect 10401 13119 10402 13145
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9534 12362 9562 12367
rect 9310 12361 9562 12362
rect 9310 12335 9311 12361
rect 9337 12335 9535 12361
rect 9561 12335 9562 12361
rect 9310 12334 9562 12335
rect 9310 11970 9338 12334
rect 9534 12329 9562 12334
rect 10318 12362 10346 12367
rect 10318 12315 10346 12334
rect 8750 11969 9338 11970
rect 8750 11943 8751 11969
rect 8777 11943 8975 11969
rect 9001 11943 9338 11969
rect 8750 11942 9338 11943
rect 8750 11802 8778 11942
rect 8974 11937 9002 11942
rect 8750 11298 8778 11774
rect 9030 11577 9058 11583
rect 9030 11551 9031 11577
rect 9057 11551 9058 11577
rect 8750 11270 9002 11298
rect 8750 11185 8778 11270
rect 8750 11159 8751 11185
rect 8777 11159 8778 11185
rect 8750 11153 8778 11159
rect 8974 11185 9002 11270
rect 8974 11159 8975 11185
rect 9001 11159 9002 11185
rect 8974 11153 9002 11159
rect 8414 10375 8415 10401
rect 8441 10375 8442 10401
rect 6846 9591 6847 9617
rect 6873 9591 6874 9617
rect 5446 9225 5586 9226
rect 5446 9199 5447 9225
rect 5473 9199 5559 9225
rect 5585 9199 5586 9225
rect 5446 9198 5586 9199
rect 5446 9193 5474 9198
rect 5110 8807 5111 8833
rect 5137 8807 5138 8833
rect 5110 8801 5138 8807
rect 5558 8833 5586 9198
rect 5558 8807 5559 8833
rect 5585 8807 5586 8833
rect 4998 8415 4999 8441
rect 5025 8415 5026 8441
rect 4998 8386 5026 8415
rect 5446 8442 5474 8447
rect 5558 8442 5586 8807
rect 5446 8441 5586 8442
rect 5446 8415 5447 8441
rect 5473 8415 5559 8441
rect 5585 8415 5586 8441
rect 5446 8414 5586 8415
rect 5446 8409 5474 8414
rect 3822 8050 3850 8055
rect 3654 8049 3850 8050
rect 3654 8023 3655 8049
rect 3681 8023 3823 8049
rect 3849 8023 3850 8049
rect 3654 8022 3850 8023
rect 3654 8017 3682 8022
rect 2478 7265 2618 7266
rect 2478 7239 2479 7265
rect 2505 7239 2618 7265
rect 2478 7238 2618 7239
rect 3542 7266 3570 7271
rect 3598 7266 3626 7630
rect 3542 7265 3626 7266
rect 3542 7239 3543 7265
rect 3569 7239 3626 7265
rect 3542 7238 3626 7239
rect 3822 7658 3850 8022
rect 4998 8049 5026 8358
rect 4998 8023 4999 8049
rect 5025 8023 5026 8049
rect 3990 7658 4018 7663
rect 3822 7657 4018 7658
rect 3822 7631 3823 7657
rect 3849 7631 3991 7657
rect 4017 7631 4018 7657
rect 3822 7630 4018 7631
rect 3822 7266 3850 7630
rect 3990 7625 4018 7630
rect 4998 7657 5026 8023
rect 5558 8049 5586 8414
rect 5558 8023 5559 8049
rect 5585 8023 5586 8049
rect 5558 7994 5586 8023
rect 6342 9225 6370 9231
rect 6342 9199 6343 9225
rect 6369 9199 6370 9225
rect 6342 8441 6370 9199
rect 6342 8415 6343 8441
rect 6369 8415 6370 8441
rect 5670 7994 5698 7999
rect 5558 7993 5698 7994
rect 5558 7967 5671 7993
rect 5697 7967 5698 7993
rect 5558 7966 5698 7967
rect 4998 7631 4999 7657
rect 5025 7631 5026 7657
rect 4998 7602 5026 7631
rect 5446 7658 5474 7663
rect 5558 7658 5586 7966
rect 5670 7961 5698 7966
rect 5446 7657 5586 7658
rect 5446 7631 5447 7657
rect 5473 7631 5559 7657
rect 5585 7631 5586 7657
rect 5446 7630 5586 7631
rect 5446 7625 5474 7630
rect 3934 7266 3962 7271
rect 3822 7265 3962 7266
rect 3822 7239 3823 7265
rect 3849 7239 3935 7265
rect 3961 7239 3962 7265
rect 3822 7238 3962 7239
rect 2478 7209 2506 7238
rect 2478 7183 2479 7209
rect 2505 7183 2506 7209
rect 2478 7177 2506 7183
rect 2086 6847 2087 6873
rect 2113 6847 2114 6873
rect 2086 6841 2114 6847
rect 2422 6874 2450 6879
rect 2534 6874 2562 7238
rect 2422 6873 2562 6874
rect 2422 6847 2423 6873
rect 2449 6847 2535 6873
rect 2561 6847 2562 6873
rect 2422 6846 2562 6847
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 1638 6089 1722 6090
rect 1638 6063 1639 6089
rect 1665 6063 1722 6089
rect 1638 6062 1722 6063
rect 2422 6481 2450 6846
rect 2534 6841 2562 6846
rect 3542 6873 3570 7238
rect 3542 6847 3543 6873
rect 3569 6847 3570 6873
rect 2422 6455 2423 6481
rect 2449 6455 2450 6481
rect 2422 6425 2450 6455
rect 2422 6399 2423 6425
rect 2449 6399 2450 6425
rect 2422 6145 2450 6399
rect 2422 6119 2423 6145
rect 2449 6119 2450 6145
rect 2422 6089 2450 6119
rect 2422 6063 2423 6089
rect 2449 6063 2450 6089
rect 910 4103 911 4129
rect 937 4103 938 4129
rect 910 3737 938 4103
rect 910 3711 911 3737
rect 937 3711 938 3737
rect 910 3345 938 3711
rect 910 3319 911 3345
rect 937 3319 938 3345
rect 910 2953 938 3319
rect 910 2927 911 2953
rect 937 2927 938 2953
rect 910 2561 938 2927
rect 910 2535 911 2561
rect 937 2535 938 2561
rect 910 2169 938 2535
rect 910 2143 911 2169
rect 937 2143 938 2169
rect 910 2137 938 2143
rect 966 5754 994 5759
rect 966 1834 994 5726
rect 1582 5698 1610 5703
rect 1638 5698 1666 6062
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 1582 5697 1666 5698
rect 1582 5671 1583 5697
rect 1609 5671 1666 5697
rect 1582 5670 1666 5671
rect 1582 5665 1610 5670
rect 1638 5306 1666 5670
rect 1582 5305 1666 5306
rect 1582 5279 1639 5305
rect 1665 5279 1666 5305
rect 1582 5278 1666 5279
rect 1582 5194 1610 5278
rect 1638 5273 1666 5278
rect 2422 5698 2450 6063
rect 3542 6481 3570 6847
rect 3542 6455 3543 6481
rect 3569 6455 3570 6481
rect 3542 6089 3570 6455
rect 3822 6874 3850 7238
rect 3934 7233 3962 7238
rect 4998 7265 5026 7574
rect 4998 7239 4999 7265
rect 5025 7239 5026 7265
rect 3990 6874 4018 6879
rect 3822 6873 4018 6874
rect 3822 6847 3823 6873
rect 3849 6847 3991 6873
rect 4017 6847 4018 6873
rect 3822 6846 4018 6847
rect 3822 6482 3850 6846
rect 3990 6762 4018 6846
rect 3990 6729 4018 6734
rect 4998 6873 5026 7239
rect 5558 7265 5586 7630
rect 5558 7239 5559 7265
rect 5585 7239 5586 7265
rect 5558 7210 5586 7239
rect 6342 7657 6370 8415
rect 6342 7631 6343 7657
rect 6369 7631 6370 7657
rect 6342 7602 6370 7631
rect 5670 7210 5698 7215
rect 5558 7209 5698 7210
rect 5558 7183 5671 7209
rect 5697 7183 5698 7209
rect 5558 7182 5698 7183
rect 4998 6847 4999 6873
rect 5025 6847 5026 6873
rect 3934 6482 3962 6487
rect 3822 6481 3962 6482
rect 3822 6455 3823 6481
rect 3849 6455 3935 6481
rect 3961 6455 3962 6481
rect 3822 6454 3962 6455
rect 3822 6449 3850 6454
rect 3542 6063 3543 6089
rect 3569 6063 3570 6089
rect 3542 6057 3570 6063
rect 3878 6090 3906 6095
rect 3934 6090 3962 6454
rect 4998 6481 5026 6847
rect 5446 6874 5474 6879
rect 5558 6874 5586 7182
rect 5670 7177 5698 7182
rect 5446 6873 5586 6874
rect 5446 6847 5447 6873
rect 5473 6847 5559 6873
rect 5585 6847 5586 6873
rect 5446 6846 5586 6847
rect 5446 6841 5474 6846
rect 4998 6455 4999 6481
rect 5025 6455 5026 6481
rect 3990 6090 4018 6095
rect 3878 6089 4018 6090
rect 3878 6063 3879 6089
rect 3905 6063 3991 6089
rect 4017 6063 4018 6089
rect 3878 6062 4018 6063
rect 3878 6057 3906 6062
rect 3990 6057 4018 6062
rect 4998 6089 5026 6455
rect 5558 6762 5586 6846
rect 5558 6481 5586 6734
rect 5558 6455 5559 6481
rect 5585 6455 5586 6481
rect 5558 6426 5586 6455
rect 6342 6873 6370 7574
rect 6342 6847 6343 6873
rect 6369 6847 6370 6873
rect 6342 6482 6370 6847
rect 6846 8833 6874 9591
rect 6846 8807 6847 8833
rect 6873 8807 6874 8833
rect 6846 8049 6874 8807
rect 6846 8023 6847 8049
rect 6873 8023 6874 8049
rect 6846 7265 6874 8023
rect 6846 7239 6847 7265
rect 6873 7239 6874 7265
rect 6846 6482 6874 7239
rect 6342 6481 6874 6482
rect 6342 6455 6847 6481
rect 6873 6455 6874 6481
rect 6342 6454 6874 6455
rect 5670 6426 5698 6431
rect 5558 6425 5698 6426
rect 5558 6399 5671 6425
rect 5697 6399 5698 6425
rect 5558 6398 5698 6399
rect 4998 6063 4999 6089
rect 5025 6063 5026 6089
rect 2422 5641 2450 5670
rect 2422 5615 2423 5641
rect 2449 5615 2450 5641
rect 2422 5361 2450 5615
rect 2422 5335 2423 5361
rect 2449 5335 2450 5361
rect 2422 5305 2450 5335
rect 2422 5279 2423 5305
rect 2449 5279 2450 5305
rect 1582 4913 1610 5166
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 1582 4887 1583 4913
rect 1609 4887 1610 4913
rect 1582 4521 1610 4887
rect 2422 4913 2450 5279
rect 2422 4887 2423 4913
rect 2449 4887 2450 4913
rect 2422 4857 2450 4887
rect 2422 4831 2423 4857
rect 2449 4831 2450 4857
rect 2422 4577 2450 4831
rect 2422 4551 2423 4577
rect 2449 4551 2450 4577
rect 1582 4495 1583 4521
rect 1609 4495 1610 4521
rect 1582 4489 1610 4495
rect 2030 4522 2058 4527
rect 2030 3009 2058 4494
rect 2422 4521 2450 4551
rect 2422 4495 2423 4521
rect 2449 4495 2450 4521
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2422 4214 2450 4495
rect 2870 5697 2898 5703
rect 2870 5671 2871 5697
rect 2897 5671 2898 5697
rect 2870 5305 2898 5671
rect 3374 5698 3402 5703
rect 3542 5698 3570 5703
rect 3402 5697 3570 5698
rect 3402 5671 3543 5697
rect 3569 5671 3570 5697
rect 3402 5670 3570 5671
rect 3374 5651 3402 5670
rect 3542 5665 3570 5670
rect 4998 5697 5026 6063
rect 5446 6090 5474 6095
rect 5558 6090 5586 6398
rect 5670 6393 5698 6398
rect 5446 6089 5558 6090
rect 5446 6063 5447 6089
rect 5473 6063 5558 6089
rect 5446 6062 5558 6063
rect 5446 6057 5474 6062
rect 4998 5671 4999 5697
rect 5025 5671 5026 5697
rect 2870 5279 2871 5305
rect 2897 5279 2898 5305
rect 2870 5194 2898 5279
rect 2870 4913 2898 5166
rect 2870 4887 2871 4913
rect 2897 4887 2898 4913
rect 2870 4521 2898 4887
rect 3430 5306 3458 5311
rect 3542 5306 3570 5311
rect 3430 5305 3570 5306
rect 3430 5279 3431 5305
rect 3457 5279 3543 5305
rect 3569 5279 3570 5305
rect 3430 5278 3570 5279
rect 3430 4914 3458 5278
rect 3542 5273 3570 5278
rect 4998 5305 5026 5671
rect 5558 5697 5586 6062
rect 6342 6089 6370 6454
rect 6846 6449 6874 6454
rect 6902 10010 6930 10015
rect 7014 10010 7042 10015
rect 6902 10009 7042 10010
rect 6902 9983 6903 10009
rect 6929 9983 7015 10009
rect 7041 9983 7042 10009
rect 6902 9982 7042 9983
rect 6902 9226 6930 9982
rect 7014 9977 7042 9982
rect 7294 9618 7322 9623
rect 7518 9618 7546 9623
rect 7294 9617 7546 9618
rect 7294 9591 7295 9617
rect 7321 9591 7519 9617
rect 7545 9591 7546 9617
rect 7294 9590 7546 9591
rect 7014 9226 7042 9231
rect 6902 9225 7042 9226
rect 6902 9199 6903 9225
rect 6929 9199 7015 9225
rect 7041 9199 7042 9225
rect 6902 9198 7042 9199
rect 6902 8442 6930 9198
rect 7014 9193 7042 9198
rect 7294 8834 7322 9590
rect 7518 9585 7546 9590
rect 8414 9617 8442 10375
rect 9030 10793 9058 11551
rect 9310 11578 9338 11942
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9534 11578 9562 11583
rect 9310 11577 9562 11578
rect 9310 11551 9311 11577
rect 9337 11551 9535 11577
rect 9561 11551 9562 11577
rect 9310 11550 9562 11551
rect 9310 11545 9338 11550
rect 9534 11545 9562 11550
rect 10318 11578 10346 11583
rect 10374 11578 10402 13119
rect 10934 12753 10962 15470
rect 10934 12727 10935 12753
rect 10961 12727 10962 12753
rect 10934 12362 10962 12727
rect 10934 12329 10962 12334
rect 10318 11577 10402 11578
rect 10318 11551 10319 11577
rect 10345 11551 10402 11577
rect 10318 11550 10402 11551
rect 10934 11969 10962 11975
rect 10934 11943 10935 11969
rect 10961 11943 10962 11969
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10850 9842 10855
rect 9030 10767 9031 10793
rect 9057 10767 9058 10793
rect 9030 10010 9058 10767
rect 9758 10849 9842 10850
rect 9758 10823 9815 10849
rect 9841 10823 9842 10849
rect 9758 10822 9842 10823
rect 9758 10793 9786 10822
rect 9814 10817 9842 10822
rect 9758 10767 9759 10793
rect 9785 10767 9786 10793
rect 9254 10401 9282 10407
rect 9254 10375 9255 10401
rect 9281 10375 9282 10401
rect 9254 10345 9282 10375
rect 9254 10319 9255 10345
rect 9281 10319 9282 10345
rect 9086 10010 9114 10015
rect 9030 10009 9114 10010
rect 9030 9983 9087 10009
rect 9113 9983 9114 10009
rect 9030 9982 9114 9983
rect 8414 9591 8415 9617
rect 8441 9591 8442 9617
rect 7518 8834 7546 8839
rect 7294 8833 7546 8834
rect 7294 8807 7295 8833
rect 7321 8807 7519 8833
rect 7545 8807 7546 8833
rect 7294 8806 7546 8807
rect 7014 8442 7042 8447
rect 6902 8441 7042 8442
rect 6902 8415 6903 8441
rect 6929 8415 7015 8441
rect 7041 8415 7042 8441
rect 6902 8414 7042 8415
rect 6902 7658 6930 8414
rect 7014 8409 7042 8414
rect 7294 8050 7322 8806
rect 7518 8801 7546 8806
rect 8414 8833 8442 9591
rect 8414 8807 8415 8833
rect 8441 8807 8442 8833
rect 7518 8050 7546 8055
rect 7294 8049 7546 8050
rect 7294 8023 7295 8049
rect 7321 8023 7519 8049
rect 7545 8023 7546 8049
rect 7294 8022 7546 8023
rect 7014 7658 7042 7663
rect 6902 7657 7042 7658
rect 6902 7631 6903 7657
rect 6929 7631 7015 7657
rect 7041 7631 7042 7657
rect 6902 7630 7042 7631
rect 6902 6874 6930 7630
rect 7014 7625 7042 7630
rect 7294 7266 7322 8022
rect 7518 8017 7546 8022
rect 8414 8049 8442 8807
rect 8414 8023 8415 8049
rect 8441 8023 8442 8049
rect 7518 7266 7546 7271
rect 7294 7265 7518 7266
rect 7294 7239 7295 7265
rect 7321 7239 7518 7265
rect 7294 7238 7518 7239
rect 7014 6874 7042 6879
rect 6902 6873 7042 6874
rect 6902 6847 6903 6873
rect 6929 6847 7015 6873
rect 7041 6847 7042 6873
rect 6902 6846 7042 6847
rect 6902 6482 6930 6846
rect 7014 6841 7042 6846
rect 7294 6482 7322 7238
rect 7518 7200 7546 7238
rect 8414 7265 8442 8023
rect 8414 7239 8415 7265
rect 8441 7239 8442 7265
rect 8414 7233 8442 7239
rect 8750 9618 8778 9623
rect 8974 9618 9002 9623
rect 8750 9617 8974 9618
rect 8750 9591 8751 9617
rect 8777 9591 8974 9617
rect 8750 9590 8974 9591
rect 8750 8834 8778 9590
rect 8974 9552 9002 9590
rect 9086 9226 9114 9982
rect 9254 10010 9282 10319
rect 9758 10094 9786 10767
rect 10318 10793 10346 11550
rect 10318 10767 10319 10793
rect 10345 10767 10346 10793
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9534 10066 9786 10094
rect 10318 10122 10346 10767
rect 9310 10010 9338 10015
rect 9534 10010 9562 10066
rect 9254 10009 9562 10010
rect 9254 9983 9311 10009
rect 9337 9983 9535 10009
rect 9561 9983 9562 10009
rect 9254 9982 9562 9983
rect 9254 9618 9282 9982
rect 9310 9977 9338 9982
rect 9534 9977 9562 9982
rect 10318 10009 10346 10094
rect 10318 9983 10319 10009
rect 10345 9983 10346 10009
rect 9282 9590 9338 9618
rect 9254 9585 9282 9590
rect 8974 8834 9002 8839
rect 8750 8833 9002 8834
rect 8750 8807 8751 8833
rect 8777 8807 8975 8833
rect 9001 8807 9002 8833
rect 8750 8806 9002 8807
rect 8750 8050 8778 8806
rect 8974 8801 9002 8806
rect 9086 8441 9114 9198
rect 9310 9226 9338 9590
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9534 9282 9562 9287
rect 9534 9226 9562 9254
rect 9310 9225 9562 9226
rect 9310 9199 9311 9225
rect 9337 9199 9535 9225
rect 9561 9199 9562 9225
rect 9310 9198 9562 9199
rect 9310 9193 9338 9198
rect 9534 9193 9562 9198
rect 10318 9226 10346 9983
rect 10822 11186 10850 11191
rect 10934 11186 10962 11943
rect 10822 11185 10962 11186
rect 10822 11159 10823 11185
rect 10849 11159 10962 11185
rect 10822 11158 10962 11159
rect 10822 10402 10850 11158
rect 10822 10122 10850 10374
rect 10822 9617 10850 10094
rect 11046 10010 11074 27706
rect 11494 23393 11522 23399
rect 11494 23367 11495 23393
rect 11521 23367 11522 23393
rect 11494 23337 11522 23367
rect 11494 23311 11495 23337
rect 11521 23311 11522 23337
rect 11102 22946 11130 22951
rect 11102 22899 11130 22918
rect 11382 22946 11410 22951
rect 11494 22946 11522 23311
rect 11382 22945 11522 22946
rect 11382 22919 11383 22945
rect 11409 22919 11495 22945
rect 11521 22919 11522 22945
rect 11382 22918 11522 22919
rect 11270 22609 11298 22615
rect 11270 22583 11271 22609
rect 11297 22583 11298 22609
rect 11270 22553 11298 22583
rect 11270 22527 11271 22553
rect 11297 22527 11298 22553
rect 11102 22161 11130 22167
rect 11102 22135 11103 22161
rect 11129 22135 11130 22161
rect 11102 21770 11130 22135
rect 11270 22161 11298 22527
rect 11270 22135 11271 22161
rect 11297 22135 11298 22161
rect 11270 21826 11298 22135
rect 11382 22162 11410 22918
rect 11494 22913 11522 22918
rect 12278 22946 12306 22951
rect 11382 21882 11410 22134
rect 11270 21793 11298 21798
rect 11326 21826 11410 21854
rect 11494 22161 11522 22167
rect 11494 22135 11495 22161
rect 11521 22135 11522 22161
rect 11494 21826 11522 22135
rect 11102 21377 11130 21742
rect 11102 21351 11103 21377
rect 11129 21351 11130 21377
rect 11102 20706 11130 21351
rect 11102 20673 11130 20678
rect 11326 21041 11354 21826
rect 11494 21769 11522 21798
rect 11494 21743 11495 21769
rect 11521 21743 11522 21769
rect 11382 21378 11410 21383
rect 11494 21378 11522 21743
rect 11550 21378 11578 21383
rect 11382 21377 11578 21378
rect 11382 21351 11383 21377
rect 11409 21351 11551 21377
rect 11577 21351 11578 21377
rect 11382 21350 11578 21351
rect 12278 21378 12306 22918
rect 12558 22162 12586 22167
rect 12838 22162 12866 22167
rect 12558 22161 12810 22162
rect 12558 22135 12559 22161
rect 12585 22135 12810 22161
rect 12558 22134 12810 22135
rect 12558 22129 12586 22134
rect 12782 21854 12810 22134
rect 12838 22115 12866 22134
rect 12950 22162 12978 22167
rect 12950 22115 12978 22134
rect 12670 21826 12810 21854
rect 12558 21378 12586 21383
rect 12278 21377 12586 21378
rect 12278 21351 12559 21377
rect 12585 21351 12586 21377
rect 12278 21350 12586 21351
rect 11382 21345 11410 21350
rect 11326 21015 11327 21041
rect 11353 21015 11354 21041
rect 11326 20985 11354 21015
rect 11326 20959 11327 20985
rect 11353 20959 11354 20985
rect 11102 20593 11130 20599
rect 11102 20567 11103 20593
rect 11129 20567 11130 20593
rect 11102 19809 11130 20567
rect 11326 20594 11354 20959
rect 11550 21042 11578 21350
rect 11494 20594 11522 20599
rect 11326 20593 11522 20594
rect 11326 20567 11327 20593
rect 11353 20567 11495 20593
rect 11521 20567 11522 20593
rect 11326 20566 11522 20567
rect 11326 20561 11354 20566
rect 11494 20257 11522 20566
rect 11494 20231 11495 20257
rect 11521 20231 11522 20257
rect 11494 20201 11522 20231
rect 11494 20175 11495 20201
rect 11521 20175 11522 20201
rect 11102 19783 11103 19809
rect 11129 19783 11130 19809
rect 11102 19025 11130 19783
rect 11382 19810 11410 19815
rect 11494 19810 11522 20175
rect 11382 19809 11494 19810
rect 11382 19783 11383 19809
rect 11409 19783 11494 19809
rect 11382 19782 11494 19783
rect 11382 19777 11410 19782
rect 11494 19744 11522 19782
rect 11494 19474 11522 19479
rect 11550 19474 11578 21014
rect 12558 20986 12586 21350
rect 12558 20953 12586 20958
rect 12558 20706 12586 20711
rect 12558 20593 12586 20678
rect 12558 20567 12559 20593
rect 12585 20567 12586 20593
rect 12558 20258 12586 20567
rect 12558 20225 12586 20230
rect 11494 19473 11578 19474
rect 11494 19447 11495 19473
rect 11521 19447 11578 19473
rect 11494 19446 11578 19447
rect 12558 19809 12586 19815
rect 12558 19783 12559 19809
rect 12585 19783 12586 19809
rect 11494 19417 11522 19446
rect 11494 19391 11495 19417
rect 11521 19391 11522 19417
rect 11102 18999 11103 19025
rect 11129 18999 11130 19025
rect 11102 18241 11130 18999
rect 11382 19026 11410 19031
rect 11494 19026 11522 19391
rect 11382 19025 11522 19026
rect 11382 18999 11383 19025
rect 11409 18999 11495 19025
rect 11521 18999 11522 19025
rect 11382 18998 11522 18999
rect 11382 18993 11410 18998
rect 11494 18689 11522 18998
rect 11494 18663 11495 18689
rect 11521 18663 11522 18689
rect 11494 18633 11522 18663
rect 11494 18607 11495 18633
rect 11521 18607 11522 18633
rect 11102 18215 11103 18241
rect 11129 18215 11130 18241
rect 11102 17850 11130 18215
rect 11382 18242 11410 18247
rect 11494 18242 11522 18607
rect 11382 18241 11522 18242
rect 11382 18215 11383 18241
rect 11409 18215 11495 18241
rect 11521 18215 11522 18241
rect 11382 18214 11522 18215
rect 11382 18209 11410 18214
rect 11102 17458 11130 17822
rect 11494 17905 11522 18214
rect 11494 17879 11495 17905
rect 11521 17879 11522 17905
rect 11494 17849 11522 17879
rect 11494 17823 11495 17849
rect 11521 17823 11522 17849
rect 11494 17817 11522 17823
rect 12558 19025 12586 19783
rect 12670 19586 12698 21826
rect 12782 21770 12810 21826
rect 12838 21770 12866 21775
rect 12782 21769 12866 21770
rect 12782 21743 12839 21769
rect 12865 21743 12866 21769
rect 12782 21742 12866 21743
rect 12838 21737 12866 21742
rect 13398 21770 13426 21775
rect 13566 21770 13594 21775
rect 13398 21769 13594 21770
rect 13398 21743 13399 21769
rect 13425 21743 13567 21769
rect 13593 21743 13594 21769
rect 13398 21742 13594 21743
rect 13398 21737 13426 21742
rect 12726 21378 12754 21383
rect 12950 21378 12978 21383
rect 12726 21377 12978 21378
rect 12726 21351 12727 21377
rect 12753 21351 12951 21377
rect 12977 21351 12978 21377
rect 12726 21350 12978 21351
rect 12726 21042 12754 21350
rect 12950 21345 12978 21350
rect 12726 20594 12754 21014
rect 13286 21042 13314 21047
rect 13118 20986 13146 20991
rect 12950 20594 12978 20599
rect 12726 20593 12978 20594
rect 12726 20567 12727 20593
rect 12753 20567 12951 20593
rect 12977 20567 12978 20593
rect 12726 20566 12978 20567
rect 12726 20561 12754 20566
rect 12950 20561 12978 20566
rect 13062 20258 13090 20263
rect 13062 20201 13090 20230
rect 13062 20175 13063 20201
rect 13089 20175 13090 20201
rect 13062 20169 13090 20175
rect 13118 20202 13146 20958
rect 13118 20169 13146 20174
rect 13286 20985 13314 21014
rect 13286 20959 13287 20985
rect 13313 20959 13314 20985
rect 13286 20202 13314 20959
rect 13510 21042 13538 21047
rect 13510 20985 13538 21014
rect 13510 20959 13511 20985
rect 13537 20959 13538 20985
rect 13510 20953 13538 20959
rect 13510 20202 13538 20207
rect 13286 20201 13538 20202
rect 13286 20175 13287 20201
rect 13313 20175 13511 20201
rect 13537 20175 13538 20201
rect 13286 20174 13538 20175
rect 13286 20169 13314 20174
rect 13510 20169 13538 20174
rect 12726 19810 12754 19815
rect 12726 19763 12754 19782
rect 12950 19810 12978 19815
rect 12950 19763 12978 19782
rect 13566 19810 13594 21742
rect 12670 19558 12810 19586
rect 12558 18999 12559 19025
rect 12585 18999 12586 19025
rect 12558 18241 12586 18999
rect 12558 18215 12559 18241
rect 12585 18215 12586 18241
rect 11102 17411 11130 17430
rect 11382 17458 11410 17463
rect 11494 17458 11522 17463
rect 11382 17457 11522 17458
rect 11382 17431 11383 17457
rect 11409 17431 11495 17457
rect 11521 17431 11522 17457
rect 11382 17430 11522 17431
rect 11270 17121 11298 17127
rect 11270 17095 11271 17121
rect 11297 17095 11298 17121
rect 11270 17065 11298 17095
rect 11270 17039 11271 17065
rect 11297 17039 11298 17065
rect 11270 16674 11298 17039
rect 11270 16337 11298 16646
rect 11270 16311 11271 16337
rect 11297 16311 11298 16337
rect 11270 16281 11298 16311
rect 11270 16255 11271 16281
rect 11297 16255 11298 16281
rect 11270 15554 11298 16255
rect 11382 15974 11410 17430
rect 11494 17425 11522 17430
rect 12558 17458 12586 18215
rect 11326 15946 11410 15974
rect 11494 16674 11522 16679
rect 11326 15913 11354 15918
rect 11494 15889 11522 16646
rect 12558 16673 12586 17430
rect 12558 16647 12559 16673
rect 12585 16647 12586 16673
rect 12558 16641 12586 16647
rect 12782 19026 12810 19558
rect 12726 15946 12754 15951
rect 11494 15863 11495 15889
rect 11521 15863 11522 15889
rect 11438 15554 11466 15559
rect 11270 15553 11466 15554
rect 11270 15527 11439 15553
rect 11465 15527 11466 15553
rect 11270 15526 11466 15527
rect 11438 15497 11466 15526
rect 11438 15471 11439 15497
rect 11465 15471 11466 15497
rect 11438 14769 11466 15471
rect 11438 14743 11439 14769
rect 11465 14743 11466 14769
rect 11438 14713 11466 14743
rect 11438 14687 11439 14713
rect 11465 14687 11466 14713
rect 11438 13986 11466 14687
rect 11494 15105 11522 15863
rect 12278 15889 12306 15895
rect 12278 15863 12279 15889
rect 12305 15863 12306 15889
rect 11774 15834 11802 15839
rect 11494 15079 11495 15105
rect 11521 15079 11522 15105
rect 11494 14321 11522 15079
rect 11494 14295 11495 14321
rect 11521 14295 11522 14321
rect 11494 14289 11522 14295
rect 11718 15833 11802 15834
rect 11718 15807 11775 15833
rect 11801 15807 11802 15833
rect 11718 15806 11802 15807
rect 11718 15050 11746 15806
rect 11774 15801 11802 15806
rect 12278 15105 12306 15863
rect 12726 15889 12754 15918
rect 12726 15863 12727 15889
rect 12753 15863 12754 15889
rect 12726 15857 12754 15863
rect 12278 15079 12279 15105
rect 12305 15079 12306 15105
rect 11774 15050 11802 15055
rect 11718 15049 11802 15050
rect 11718 15023 11775 15049
rect 11801 15023 11802 15049
rect 11718 15022 11802 15023
rect 11718 14266 11746 15022
rect 11774 15017 11802 15022
rect 12278 14321 12306 15079
rect 12278 14295 12279 14321
rect 12305 14295 12306 14321
rect 11774 14266 11802 14271
rect 11746 14265 11802 14266
rect 11746 14239 11775 14265
rect 11801 14239 11802 14265
rect 11746 14238 11802 14239
rect 11494 13986 11522 13991
rect 11438 13985 11522 13986
rect 11438 13959 11495 13985
rect 11521 13959 11522 13985
rect 11438 13958 11522 13959
rect 11494 13930 11522 13958
rect 11718 13930 11746 14238
rect 11774 14233 11802 14238
rect 11522 13902 11746 13930
rect 11494 13864 11522 13902
rect 11718 13537 11746 13902
rect 11718 13511 11719 13537
rect 11745 13511 11746 13537
rect 11718 13482 11746 13511
rect 12278 13537 12306 14295
rect 12278 13511 12279 13537
rect 12305 13511 12306 13537
rect 11774 13482 11802 13487
rect 11718 13481 11802 13482
rect 11718 13455 11775 13481
rect 11801 13455 11802 13481
rect 11718 13454 11802 13455
rect 11494 13201 11522 13207
rect 11494 13175 11495 13201
rect 11521 13175 11522 13201
rect 11494 13146 11522 13175
rect 11718 13146 11746 13454
rect 11774 13449 11802 13454
rect 11494 13145 11746 13146
rect 11494 13119 11495 13145
rect 11521 13119 11746 13145
rect 11494 13118 11746 13119
rect 11494 13113 11522 13118
rect 11718 12753 11746 13118
rect 11718 12727 11719 12753
rect 11745 12727 11746 12753
rect 11718 12698 11746 12727
rect 12278 12753 12306 13511
rect 12782 13034 12810 18998
rect 13118 19417 13146 19423
rect 13118 19391 13119 19417
rect 13145 19391 13146 19417
rect 13118 18633 13146 19391
rect 13118 18607 13119 18633
rect 13145 18607 13146 18633
rect 13118 17849 13146 18607
rect 13118 17823 13119 17849
rect 13145 17823 13146 17849
rect 13118 17458 13146 17823
rect 13118 17066 13146 17430
rect 13118 16281 13146 17038
rect 13118 16255 13119 16281
rect 13145 16255 13146 16281
rect 13118 16249 13146 16255
rect 13398 19418 13426 19423
rect 13566 19418 13594 19782
rect 13398 19417 13594 19418
rect 13398 19391 13399 19417
rect 13425 19391 13567 19417
rect 13593 19391 13594 19417
rect 13398 19390 13594 19391
rect 13398 19025 13426 19390
rect 13566 19385 13594 19390
rect 13398 18999 13399 19025
rect 13425 18999 13426 19025
rect 13398 18969 13426 18999
rect 13398 18943 13399 18969
rect 13425 18943 13426 18969
rect 13398 18634 13426 18943
rect 13510 18634 13538 18639
rect 13398 18633 13538 18634
rect 13398 18607 13399 18633
rect 13425 18607 13511 18633
rect 13537 18607 13538 18633
rect 13398 18606 13538 18607
rect 13398 18241 13426 18606
rect 13510 18601 13538 18606
rect 13398 18215 13399 18241
rect 13425 18215 13426 18241
rect 13398 18185 13426 18215
rect 13398 18159 13399 18185
rect 13425 18159 13426 18185
rect 13398 17850 13426 18159
rect 13510 17850 13538 17855
rect 13398 17849 13538 17850
rect 13398 17823 13399 17849
rect 13425 17823 13511 17849
rect 13537 17823 13538 17849
rect 13398 17822 13538 17823
rect 13398 17457 13426 17822
rect 13510 17817 13538 17822
rect 13398 17431 13399 17457
rect 13425 17431 13426 17457
rect 13398 17401 13426 17431
rect 13398 17375 13399 17401
rect 13425 17375 13426 17401
rect 13398 17066 13426 17375
rect 13510 17066 13538 17071
rect 13398 17065 13538 17066
rect 13398 17039 13399 17065
rect 13425 17039 13511 17065
rect 13537 17039 13538 17065
rect 13398 17038 13538 17039
rect 13398 16673 13426 17038
rect 13510 17033 13538 17038
rect 13398 16647 13399 16673
rect 13425 16647 13426 16673
rect 13398 16617 13426 16647
rect 13398 16591 13399 16617
rect 13425 16591 13426 16617
rect 13398 16282 13426 16591
rect 13510 16282 13538 16287
rect 13398 16281 13538 16282
rect 13398 16255 13399 16281
rect 13425 16255 13511 16281
rect 13537 16255 13538 16281
rect 13398 16254 13538 16255
rect 13398 16249 13426 16254
rect 12950 15946 12978 15951
rect 12950 15889 12978 15918
rect 12950 15863 12951 15889
rect 12977 15863 12978 15889
rect 12950 15857 12978 15863
rect 13454 15946 13482 16254
rect 13510 16249 13538 16254
rect 12782 13001 12810 13006
rect 12838 15497 12866 15503
rect 12838 15471 12839 15497
rect 12865 15471 12866 15497
rect 12838 14713 12866 15471
rect 13398 15498 13426 15503
rect 13454 15498 13482 15918
rect 13510 15498 13538 15503
rect 13398 15497 13538 15498
rect 13398 15471 13399 15497
rect 13425 15471 13511 15497
rect 13537 15471 13538 15497
rect 13398 15470 13538 15471
rect 13398 15465 13426 15470
rect 12838 14687 12839 14713
rect 12865 14687 12866 14713
rect 12838 13929 12866 14687
rect 13342 15105 13370 15111
rect 13342 15079 13343 15105
rect 13369 15079 13370 15105
rect 13342 15049 13370 15079
rect 13342 15023 13343 15049
rect 13369 15023 13370 15049
rect 13342 14322 13370 15023
rect 13398 14714 13426 14719
rect 13510 14714 13538 15470
rect 13398 14713 13538 14714
rect 13398 14687 13399 14713
rect 13425 14687 13511 14713
rect 13537 14687 13538 14713
rect 13398 14686 13538 14687
rect 13398 14681 13426 14686
rect 13398 14322 13426 14327
rect 13342 14321 13426 14322
rect 13342 14295 13399 14321
rect 13425 14295 13426 14321
rect 13342 14294 13426 14295
rect 13398 14266 13426 14294
rect 13398 14219 13426 14238
rect 12838 13903 12839 13929
rect 12865 13903 12866 13929
rect 12838 13145 12866 13903
rect 13398 13930 13426 13935
rect 13510 13930 13538 14686
rect 13398 13929 13538 13930
rect 13398 13903 13399 13929
rect 13425 13903 13511 13929
rect 13537 13903 13538 13929
rect 13398 13902 13538 13903
rect 13398 13897 13426 13902
rect 13454 13537 13482 13902
rect 13510 13897 13538 13902
rect 13454 13511 13455 13537
rect 13481 13511 13482 13537
rect 13454 13481 13482 13511
rect 13454 13455 13455 13481
rect 13481 13455 13482 13481
rect 12838 13119 12839 13145
rect 12865 13119 12866 13145
rect 12278 12727 12279 12753
rect 12305 12727 12306 12753
rect 11774 12698 11802 12703
rect 11718 12697 11802 12698
rect 11718 12671 11775 12697
rect 11801 12671 11802 12697
rect 11718 12670 11802 12671
rect 11494 12417 11522 12423
rect 11494 12391 11495 12417
rect 11521 12391 11522 12417
rect 11494 12362 11522 12391
rect 11718 12362 11746 12670
rect 11774 12665 11802 12670
rect 11494 12361 11746 12362
rect 11494 12335 11495 12361
rect 11521 12335 11746 12361
rect 11494 12334 11746 12335
rect 11494 12329 11522 12334
rect 11382 11970 11410 11975
rect 11494 11970 11522 11975
rect 11382 11969 11522 11970
rect 11382 11943 11383 11969
rect 11409 11943 11495 11969
rect 11521 11943 11522 11969
rect 11382 11942 11522 11943
rect 11382 11937 11410 11942
rect 11494 11633 11522 11942
rect 11494 11607 11495 11633
rect 11521 11607 11522 11633
rect 11494 11578 11522 11607
rect 11382 11186 11410 11191
rect 11494 11186 11522 11550
rect 11382 11185 11522 11186
rect 11382 11159 11383 11185
rect 11409 11159 11495 11185
rect 11521 11159 11522 11185
rect 11382 11158 11522 11159
rect 11382 11153 11410 11158
rect 11494 10849 11522 11158
rect 11494 10823 11495 10849
rect 11521 10823 11522 10849
rect 11494 10793 11522 10823
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11382 10402 11410 10407
rect 11494 10402 11522 10767
rect 11382 10401 11522 10402
rect 11382 10375 11383 10401
rect 11409 10375 11495 10401
rect 11521 10375 11522 10401
rect 11382 10374 11522 10375
rect 11382 10094 11410 10374
rect 11494 10369 11522 10374
rect 12278 11969 12306 12727
rect 12278 11943 12279 11969
rect 12305 11943 12306 11969
rect 12278 11185 12306 11943
rect 12278 11159 12279 11185
rect 12305 11159 12306 11185
rect 12278 10794 12306 11159
rect 12278 10402 12306 10766
rect 12838 12362 12866 13119
rect 13398 13146 13426 13151
rect 13454 13146 13482 13455
rect 13510 13146 13538 13151
rect 13398 13145 13538 13146
rect 13398 13119 13399 13145
rect 13425 13119 13511 13145
rect 13537 13119 13538 13145
rect 13398 13118 13538 13119
rect 13398 13113 13426 13118
rect 13454 12753 13482 13118
rect 13510 13113 13538 13118
rect 13454 12727 13455 12753
rect 13481 12727 13482 12753
rect 13454 12698 13482 12727
rect 13454 12697 13538 12698
rect 13454 12671 13455 12697
rect 13481 12671 13538 12697
rect 13454 12670 13538 12671
rect 13454 12665 13482 12670
rect 12838 11577 12866 12334
rect 12838 11551 12839 11577
rect 12865 11551 12866 11577
rect 12838 10794 12866 11551
rect 13398 12362 13426 12367
rect 13510 12362 13538 12670
rect 13398 12361 13538 12362
rect 13398 12335 13399 12361
rect 13425 12335 13511 12361
rect 13537 12335 13538 12361
rect 13398 12334 13538 12335
rect 13398 11969 13426 12334
rect 13510 12329 13538 12334
rect 13398 11943 13399 11969
rect 13425 11943 13426 11969
rect 13398 11913 13426 11943
rect 13398 11887 13399 11913
rect 13425 11887 13426 11913
rect 13398 11578 13426 11887
rect 13510 11578 13538 11583
rect 13426 11577 13538 11578
rect 13426 11551 13511 11577
rect 13537 11551 13538 11577
rect 13426 11550 13538 11551
rect 13398 11512 13426 11550
rect 13454 11185 13482 11550
rect 13510 11545 13538 11550
rect 13454 11159 13455 11185
rect 13481 11159 13482 11185
rect 13454 11129 13482 11159
rect 13454 11103 13455 11129
rect 13481 11103 13482 11129
rect 12838 10747 12866 10766
rect 13398 10794 13426 10799
rect 13454 10794 13482 11103
rect 13510 10794 13538 10799
rect 13398 10793 13538 10794
rect 13398 10767 13399 10793
rect 13425 10767 13511 10793
rect 13537 10767 13538 10793
rect 13398 10766 13538 10767
rect 13398 10761 13426 10766
rect 12278 10355 12306 10374
rect 13454 10401 13482 10766
rect 13510 10761 13538 10766
rect 13454 10375 13455 10401
rect 13481 10375 13482 10401
rect 13454 10345 13482 10375
rect 13454 10319 13455 10345
rect 13481 10319 13482 10345
rect 13454 10234 13482 10319
rect 13454 10206 13650 10234
rect 11046 9977 11074 9982
rect 11270 10066 11410 10094
rect 13566 10122 13594 10127
rect 11270 10065 11298 10066
rect 11270 10039 11271 10065
rect 11297 10039 11298 10065
rect 11270 10009 11298 10039
rect 11270 9983 11271 10009
rect 11297 9983 11298 10009
rect 10822 9591 10823 9617
rect 10849 9591 10850 9617
rect 10822 9585 10850 9591
rect 11270 9618 11298 9983
rect 12838 10009 12866 10015
rect 12838 9983 12839 10009
rect 12865 9983 12866 10009
rect 11494 9618 11522 9623
rect 11270 9617 11522 9618
rect 11270 9591 11271 9617
rect 11297 9591 11495 9617
rect 11521 9591 11522 9617
rect 11270 9590 11522 9591
rect 10318 9179 10346 9198
rect 10990 9282 11018 9287
rect 10990 9225 11018 9254
rect 10990 9199 10991 9225
rect 11017 9199 11018 9225
rect 10990 9193 11018 9199
rect 11270 9282 11298 9590
rect 11494 9585 11522 9590
rect 12558 9618 12586 9623
rect 12558 9571 12586 9590
rect 12838 9618 12866 9983
rect 13398 10010 13426 10015
rect 10598 8834 10626 8839
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9086 8415 9087 8441
rect 9113 8415 9114 8441
rect 8974 8050 9002 8055
rect 8750 8049 9002 8050
rect 8750 8023 8751 8049
rect 8777 8023 8975 8049
rect 9001 8023 9002 8049
rect 8750 8022 9002 8023
rect 8750 7266 8778 8022
rect 8974 8017 9002 8022
rect 9086 7657 9114 8415
rect 9086 7631 9087 7657
rect 9113 7631 9114 7657
rect 9086 7625 9114 7631
rect 9310 8442 9338 8447
rect 9534 8442 9562 8447
rect 9310 8441 9562 8442
rect 9310 8415 9311 8441
rect 9337 8415 9535 8441
rect 9561 8415 9562 8441
rect 9310 8414 9562 8415
rect 9310 7658 9338 8414
rect 9534 8409 9562 8414
rect 10598 8442 10626 8806
rect 11102 8834 11130 8839
rect 11102 8787 11130 8806
rect 11270 8834 11298 9254
rect 12838 9226 12866 9590
rect 12838 9160 12866 9198
rect 13342 9617 13370 9623
rect 13342 9591 13343 9617
rect 13369 9591 13370 9617
rect 13342 9561 13370 9591
rect 13342 9535 13343 9561
rect 13369 9535 13370 9561
rect 13342 9338 13370 9535
rect 13342 9225 13370 9310
rect 13342 9199 13343 9225
rect 13369 9199 13370 9225
rect 11494 8834 11522 8839
rect 11270 8833 11522 8834
rect 11270 8807 11271 8833
rect 11297 8807 11495 8833
rect 11521 8807 11522 8833
rect 11270 8806 11522 8807
rect 10598 8376 10626 8414
rect 11270 8497 11298 8806
rect 11494 8801 11522 8806
rect 12278 8833 12306 8839
rect 12278 8807 12279 8833
rect 12305 8807 12306 8833
rect 11270 8471 11271 8497
rect 11297 8471 11298 8497
rect 11270 8441 11298 8471
rect 11270 8415 11271 8441
rect 11297 8415 11298 8441
rect 11270 8409 11298 8415
rect 11102 8049 11130 8055
rect 11102 8023 11103 8049
rect 11129 8023 11130 8049
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9534 7658 9562 7663
rect 9310 7657 9562 7658
rect 9310 7631 9311 7657
rect 9337 7631 9535 7657
rect 9561 7631 9562 7657
rect 9310 7630 9562 7631
rect 9310 7602 9338 7630
rect 9534 7625 9562 7630
rect 10598 7658 10626 7663
rect 10598 7611 10626 7630
rect 11102 7658 11130 8023
rect 11998 8049 12026 8055
rect 11998 8023 11999 8049
rect 12025 8023 12026 8049
rect 11998 7993 12026 8023
rect 11998 7967 11999 7993
rect 12025 7967 12026 7993
rect 9198 7574 9338 7602
rect 8750 7219 8778 7238
rect 8974 7266 9002 7271
rect 9198 7266 9226 7574
rect 9002 7238 9226 7266
rect 11102 7265 11130 7630
rect 11494 7713 11522 7719
rect 11494 7687 11495 7713
rect 11521 7687 11522 7713
rect 11494 7657 11522 7687
rect 11494 7631 11495 7657
rect 11521 7631 11522 7657
rect 11494 7546 11522 7631
rect 11998 7546 12026 7967
rect 11494 7518 12026 7546
rect 11102 7239 11103 7265
rect 11129 7239 11130 7265
rect 8974 7219 9002 7238
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10990 6929 11018 6935
rect 10990 6903 10991 6929
rect 11017 6903 11018 6929
rect 9814 6873 9842 6879
rect 9814 6847 9815 6873
rect 9841 6847 9842 6873
rect 9814 6538 9842 6847
rect 7518 6482 7546 6487
rect 6902 6481 7546 6482
rect 6902 6455 7295 6481
rect 7321 6455 7519 6481
rect 7545 6455 7546 6481
rect 6902 6454 7546 6455
rect 6342 6063 6343 6089
rect 6369 6063 6370 6089
rect 6342 6057 6370 6063
rect 6790 6090 6818 6095
rect 6902 6090 6930 6454
rect 7294 6449 7322 6454
rect 7518 6449 7546 6454
rect 9534 6481 9562 6487
rect 9534 6455 9535 6481
rect 9561 6455 9562 6481
rect 7014 6090 7042 6095
rect 6818 6089 7042 6090
rect 6818 6063 7015 6089
rect 7041 6063 7042 6089
rect 6818 6062 7042 6063
rect 6790 6043 6818 6062
rect 7014 6057 7042 6062
rect 5558 5671 5559 5697
rect 5585 5671 5586 5697
rect 5558 5642 5586 5671
rect 8302 5698 8330 5703
rect 8414 5698 8442 5703
rect 8302 5697 8442 5698
rect 8302 5671 8303 5697
rect 8329 5671 8415 5697
rect 8441 5671 8442 5697
rect 8302 5670 8442 5671
rect 5670 5642 5698 5647
rect 5558 5641 5698 5642
rect 5558 5615 5671 5641
rect 5697 5615 5698 5641
rect 5558 5614 5698 5615
rect 4998 5279 4999 5305
rect 5025 5279 5026 5305
rect 3542 4914 3570 4919
rect 3430 4913 3542 4914
rect 3430 4887 3431 4913
rect 3457 4887 3542 4913
rect 3430 4886 3542 4887
rect 2870 4495 2871 4521
rect 2897 4495 2898 4521
rect 2870 4489 2898 4495
rect 3374 4522 3402 4527
rect 3430 4522 3458 4886
rect 3542 4848 3570 4886
rect 4998 4913 5026 5279
rect 5390 5306 5418 5311
rect 5558 5306 5586 5614
rect 5670 5609 5698 5614
rect 5390 5305 5586 5306
rect 5390 5279 5391 5305
rect 5417 5279 5559 5305
rect 5585 5279 5586 5305
rect 5390 5278 5586 5279
rect 4998 4887 4999 4913
rect 5025 4887 5026 4913
rect 4998 4881 5026 4887
rect 5166 4914 5194 4919
rect 5166 4867 5194 4886
rect 5390 4914 5418 5278
rect 5558 5273 5586 5278
rect 7518 5305 7546 5311
rect 7518 5279 7519 5305
rect 7545 5279 7546 5305
rect 5390 4867 5418 4886
rect 6062 4577 6090 4583
rect 6062 4551 6063 4577
rect 6089 4551 6090 4577
rect 3542 4522 3570 4527
rect 3402 4521 3570 4522
rect 3402 4495 3543 4521
rect 3569 4495 3570 4521
rect 3402 4494 3570 4495
rect 3374 4475 3402 4494
rect 3542 4489 3570 4494
rect 6062 4521 6090 4551
rect 6062 4495 6063 4521
rect 6089 4495 6090 4521
rect 2030 2983 2031 3009
rect 2057 2983 2058 3009
rect 2030 2953 2058 2983
rect 2030 2927 2031 2953
rect 2057 2927 2058 2953
rect 2030 2561 2058 2927
rect 2030 2535 2031 2561
rect 2057 2535 2058 2561
rect 2030 2505 2058 2535
rect 2030 2479 2031 2505
rect 2057 2479 2058 2505
rect 2030 2225 2058 2479
rect 2030 2199 2031 2225
rect 2057 2199 2058 2225
rect 2030 2169 2058 2199
rect 2030 2143 2031 2169
rect 2057 2143 2058 2169
rect 2030 2137 2058 2143
rect 2086 4186 2450 4214
rect 6062 4214 6090 4495
rect 7014 4522 7042 4527
rect 7014 4475 7042 4494
rect 7518 4522 7546 5279
rect 7798 4913 7826 4919
rect 7798 4887 7799 4913
rect 7825 4887 7826 4913
rect 7574 4522 7602 4527
rect 7798 4522 7826 4887
rect 7546 4521 7826 4522
rect 7546 4495 7575 4521
rect 7601 4495 7826 4521
rect 7546 4494 7826 4495
rect 7518 4456 7546 4494
rect 7574 4214 7602 4494
rect 5782 4186 5810 4191
rect 2086 4129 2114 4186
rect 2086 4103 2087 4129
rect 2113 4103 2114 4129
rect 2086 4073 2114 4103
rect 2086 4047 2087 4073
rect 2113 4047 2114 4073
rect 2086 3793 2114 4047
rect 3878 4129 3906 4135
rect 3878 4103 3879 4129
rect 3905 4103 3906 4129
rect 3878 4074 3906 4103
rect 4046 4130 4074 4135
rect 3878 4073 4018 4074
rect 3878 4047 3879 4073
rect 3905 4047 4018 4073
rect 3878 4046 4018 4047
rect 3878 4041 3906 4046
rect 2086 3767 2087 3793
rect 2113 3767 2114 3793
rect 2086 3737 2114 3767
rect 2086 3711 2087 3737
rect 2113 3711 2114 3737
rect 2086 3345 2114 3711
rect 3822 3738 3850 3743
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2086 3319 2087 3345
rect 2113 3319 2114 3345
rect 2086 3289 2114 3319
rect 2086 3263 2087 3289
rect 2113 3263 2114 3289
rect 966 1777 994 1806
rect 966 1751 967 1777
rect 993 1751 994 1777
rect 966 1745 994 1751
rect 1694 2058 1722 2063
rect 1694 400 1722 2030
rect 2086 1778 2114 3263
rect 3822 3345 3850 3710
rect 3822 3319 3823 3345
rect 3849 3319 3850 3345
rect 3822 3289 3850 3319
rect 3822 3263 3823 3289
rect 3849 3263 3850 3289
rect 3822 2954 3850 3263
rect 3934 2954 3962 2959
rect 3822 2953 3962 2954
rect 3822 2927 3823 2953
rect 3849 2927 3935 2953
rect 3961 2927 3962 2953
rect 3822 2926 3962 2927
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 3822 2170 3850 2926
rect 3934 2921 3962 2926
rect 3990 2562 4018 4046
rect 4046 3738 4074 4102
rect 4998 4129 5026 4135
rect 4998 4103 4999 4129
rect 5025 4103 5026 4129
rect 4046 3672 4074 3710
rect 4494 3737 4522 3743
rect 4494 3711 4495 3737
rect 4521 3711 4522 3737
rect 4494 3346 4522 3711
rect 4494 3313 4522 3318
rect 4998 3346 5026 4103
rect 5782 4129 5810 4158
rect 5782 4103 5783 4129
rect 5809 4103 5810 4129
rect 5782 4097 5810 4103
rect 6006 4186 6034 4191
rect 6062 4186 6594 4214
rect 6006 4129 6034 4158
rect 6006 4103 6007 4129
rect 6033 4103 6034 4129
rect 6006 4097 6034 4103
rect 6454 4130 6482 4135
rect 6454 4083 6482 4102
rect 6342 3738 6370 3743
rect 6566 3738 6594 4158
rect 7518 4186 7602 4214
rect 6342 3737 6594 3738
rect 6342 3711 6343 3737
rect 6369 3711 6567 3737
rect 6593 3711 6594 3737
rect 6342 3710 6594 3711
rect 6342 3705 6370 3710
rect 4998 3299 5026 3318
rect 5558 3346 5586 3351
rect 3990 2505 4018 2534
rect 3990 2479 3991 2505
rect 4017 2479 4018 2505
rect 3990 2473 4018 2479
rect 4494 2953 4522 2959
rect 4494 2927 4495 2953
rect 4521 2927 4522 2953
rect 3934 2170 3962 2175
rect 3822 2169 3962 2170
rect 3822 2143 3823 2169
rect 3849 2143 3935 2169
rect 3961 2143 3962 2169
rect 3822 2142 3962 2143
rect 3822 2137 3850 2142
rect 3934 2137 3962 2142
rect 4494 2170 4522 2927
rect 4494 2123 4522 2142
rect 4998 2561 5026 2567
rect 4998 2535 4999 2561
rect 5025 2535 5026 2561
rect 4998 2170 5026 2535
rect 5558 2562 5586 3318
rect 5838 3346 5866 3351
rect 5950 3346 5978 3351
rect 5838 3345 5978 3346
rect 5838 3319 5839 3345
rect 5865 3319 5951 3345
rect 5977 3319 5978 3345
rect 5838 3318 5978 3319
rect 5838 3313 5866 3318
rect 5558 2515 5586 2534
rect 5894 2954 5922 3318
rect 5950 3313 5978 3318
rect 5894 2618 5922 2926
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 2086 1721 2114 1750
rect 2870 1834 2898 1839
rect 2870 1777 2898 1806
rect 2870 1751 2871 1777
rect 2897 1751 2898 1777
rect 2870 1745 2898 1751
rect 3822 1778 3850 1783
rect 2086 1695 2087 1721
rect 2113 1695 2114 1721
rect 2086 1689 2114 1695
rect 3822 1721 3850 1750
rect 3822 1695 3823 1721
rect 3849 1695 3850 1721
rect 3822 1689 3850 1695
rect 4998 1778 5026 2142
rect 5222 1778 5250 1783
rect 4998 1777 5250 1778
rect 4998 1751 5223 1777
rect 5249 1751 5250 1777
rect 4998 1750 5250 1751
rect 4998 400 5026 1750
rect 5222 1745 5250 1750
rect 5782 1778 5810 1783
rect 5894 1778 5922 2590
rect 5782 1777 5922 1778
rect 5782 1751 5783 1777
rect 5809 1751 5895 1777
rect 5921 1751 5922 1777
rect 5782 1750 5922 1751
rect 5782 1745 5810 1750
rect 5894 1745 5922 1750
rect 6118 2953 6146 2959
rect 6118 2927 6119 2953
rect 6145 2927 6146 2953
rect 6118 2562 6146 2927
rect 6286 2954 6314 2959
rect 6286 2907 6314 2926
rect 6510 2954 6538 2959
rect 6510 2907 6538 2926
rect 6118 2169 6146 2534
rect 6454 2562 6482 2567
rect 6566 2562 6594 3710
rect 7014 4130 7042 4135
rect 7014 3737 7042 4102
rect 7014 3711 7015 3737
rect 7041 3711 7042 3737
rect 7014 3402 7042 3711
rect 7518 3737 7546 4186
rect 7518 3711 7519 3737
rect 7545 3711 7546 3737
rect 7518 3705 7546 3711
rect 7798 4129 7826 4494
rect 8302 4214 8330 5670
rect 8414 5665 8442 5670
rect 8974 5698 9002 5703
rect 8974 5651 9002 5670
rect 9534 5698 9562 6455
rect 8358 5361 8386 5367
rect 8358 5335 8359 5361
rect 8385 5335 8386 5361
rect 8358 5305 8386 5335
rect 8358 5279 8359 5305
rect 8385 5279 8386 5305
rect 8358 4914 8386 5279
rect 8470 4914 8498 4919
rect 8358 4913 8498 4914
rect 8358 4887 8359 4913
rect 8385 4887 8471 4913
rect 8497 4887 8498 4913
rect 8358 4886 8498 4887
rect 8358 4881 8386 4886
rect 8470 4577 8498 4886
rect 8470 4551 8471 4577
rect 8497 4551 8498 4577
rect 8470 4521 8498 4551
rect 8470 4495 8471 4521
rect 8497 4495 8498 4521
rect 8302 4186 8386 4214
rect 7798 4103 7799 4129
rect 7825 4103 7826 4129
rect 7014 3369 7042 3374
rect 7518 3402 7546 3407
rect 6454 2561 6594 2562
rect 6454 2535 6455 2561
rect 6481 2535 6594 2561
rect 6454 2534 6594 2535
rect 6454 2505 6482 2534
rect 6454 2479 6455 2505
rect 6481 2479 6482 2505
rect 6454 2473 6482 2479
rect 6566 2506 6594 2534
rect 7518 2953 7546 3374
rect 7798 3346 7826 4103
rect 7798 3280 7826 3318
rect 8358 3793 8386 4186
rect 8358 3767 8359 3793
rect 8385 3767 8386 3793
rect 8358 3737 8386 3767
rect 8358 3711 8359 3737
rect 8385 3711 8386 3737
rect 7518 2927 7519 2953
rect 7545 2927 7546 2953
rect 6566 2473 6594 2478
rect 7014 2506 7042 2511
rect 6118 2143 6119 2169
rect 6145 2143 6146 2169
rect 6118 1778 6146 2143
rect 7014 2225 7042 2478
rect 7014 2199 7015 2225
rect 7041 2199 7042 2225
rect 7014 2169 7042 2199
rect 7014 2143 7015 2169
rect 7041 2143 7042 2169
rect 7014 2137 7042 2143
rect 7518 2170 7546 2927
rect 7518 2123 7546 2142
rect 7630 2954 7658 2959
rect 7742 2954 7770 2959
rect 7658 2953 7770 2954
rect 7658 2927 7743 2953
rect 7769 2927 7770 2953
rect 7658 2926 7770 2927
rect 6118 1745 6146 1750
rect 7462 1778 7490 1783
rect 7462 1731 7490 1750
rect 7630 1778 7658 2926
rect 7742 2921 7770 2926
rect 7966 2954 7994 2959
rect 7966 2907 7994 2926
rect 8246 2954 8274 2959
rect 8078 2561 8106 2567
rect 8078 2535 8079 2561
rect 8105 2535 8106 2561
rect 8078 2170 8106 2535
rect 8246 2562 8274 2926
rect 8246 2496 8274 2534
rect 8358 2506 8386 3711
rect 7854 1778 7882 1783
rect 7630 1777 7882 1778
rect 7630 1751 7631 1777
rect 7657 1751 7855 1777
rect 7881 1751 7882 1777
rect 7630 1750 7882 1751
rect 7630 1745 7658 1750
rect 7854 1745 7882 1750
rect 8078 1722 8106 2142
rect 8358 2225 8386 2478
rect 8470 4129 8498 4495
rect 8470 4103 8471 4129
rect 8497 4103 8498 4129
rect 8470 4074 8498 4103
rect 9534 4913 9562 5670
rect 9814 6089 9842 6510
rect 10990 6873 11018 6903
rect 10990 6847 10991 6873
rect 11017 6847 11018 6873
rect 10430 6481 10458 6487
rect 10430 6455 10431 6481
rect 10457 6455 10458 6481
rect 10430 6425 10458 6455
rect 10430 6399 10431 6425
rect 10457 6399 10458 6425
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9814 6063 9815 6089
rect 9841 6063 9842 6089
rect 9814 5698 9842 6063
rect 9814 5665 9842 5670
rect 10430 5922 10458 6399
rect 10430 5697 10458 5894
rect 10430 5671 10431 5697
rect 10457 5671 10458 5697
rect 10430 5641 10458 5671
rect 10430 5615 10431 5641
rect 10457 5615 10458 5641
rect 10430 5609 10458 5615
rect 10990 6145 11018 6847
rect 10990 6119 10991 6145
rect 11017 6119 11018 6145
rect 10990 6089 11018 6119
rect 10990 6063 10991 6089
rect 11017 6063 11018 6089
rect 10990 5922 11018 6063
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 10990 5361 11018 5894
rect 10990 5335 10991 5361
rect 11017 5335 11018 5361
rect 9534 4887 9535 4913
rect 9561 4887 9562 4913
rect 9534 4129 9562 4887
rect 10038 5305 10066 5311
rect 10038 5279 10039 5305
rect 10065 5279 10066 5305
rect 10038 4802 10066 5279
rect 10990 5305 11018 5335
rect 10990 5279 10991 5305
rect 11017 5279 11018 5305
rect 10990 5273 11018 5279
rect 11102 6538 11130 7239
rect 11998 7265 12026 7518
rect 11998 7239 11999 7265
rect 12025 7239 12026 7265
rect 11998 7209 12026 7239
rect 11998 7183 11999 7209
rect 12025 7183 12026 7209
rect 11102 6481 11130 6510
rect 11102 6455 11103 6481
rect 11129 6455 11130 6481
rect 11102 6090 11130 6455
rect 11270 6873 11298 6879
rect 11270 6847 11271 6873
rect 11297 6847 11298 6873
rect 11270 6762 11298 6847
rect 11270 6090 11298 6734
rect 11102 6089 11298 6090
rect 11102 6063 11271 6089
rect 11297 6063 11298 6089
rect 11102 6062 11298 6063
rect 11102 5697 11130 6062
rect 11270 6057 11298 6062
rect 11998 6538 12026 7183
rect 11998 6481 12026 6510
rect 11998 6455 11999 6481
rect 12025 6455 12026 6481
rect 11998 6425 12026 6455
rect 12278 8049 12306 8807
rect 12278 8023 12279 8049
rect 12305 8023 12306 8049
rect 12278 7265 12306 8023
rect 12278 7239 12279 7265
rect 12305 7239 12306 7265
rect 12278 6762 12306 7239
rect 12838 8441 12866 8447
rect 12838 8415 12839 8441
rect 12865 8415 12866 8441
rect 12838 7657 12866 8415
rect 12838 7631 12839 7657
rect 12865 7631 12866 7657
rect 12278 6481 12306 6734
rect 12278 6455 12279 6481
rect 12305 6455 12306 6481
rect 12278 6449 12306 6455
rect 12446 6929 12474 6935
rect 12446 6903 12447 6929
rect 12473 6903 12474 6929
rect 12446 6873 12474 6903
rect 12446 6847 12447 6873
rect 12473 6847 12474 6873
rect 12446 6538 12474 6847
rect 11998 6399 11999 6425
rect 12025 6399 12026 6425
rect 11102 5671 11103 5697
rect 11129 5671 11130 5697
rect 10430 4913 10458 4919
rect 10430 4887 10431 4913
rect 10457 4887 10458 4913
rect 10430 4858 10458 4887
rect 11102 4913 11130 5671
rect 11998 5922 12026 6399
rect 12446 6145 12474 6510
rect 12446 6119 12447 6145
rect 12473 6119 12474 6145
rect 12446 6089 12474 6119
rect 12446 6063 12447 6089
rect 12473 6063 12474 6089
rect 12446 6057 12474 6063
rect 12838 6873 12866 7631
rect 13342 8049 13370 9199
rect 13398 9282 13426 9982
rect 13510 10010 13538 10015
rect 13510 9963 13538 9982
rect 13398 8833 13426 9254
rect 13510 9338 13538 9343
rect 13566 9338 13594 10094
rect 13538 9310 13594 9338
rect 13510 9225 13538 9310
rect 13510 9199 13511 9225
rect 13537 9199 13538 9225
rect 13510 9193 13538 9199
rect 13398 8807 13399 8833
rect 13425 8807 13426 8833
rect 13398 8777 13426 8807
rect 13398 8751 13399 8777
rect 13425 8751 13426 8777
rect 13398 8442 13426 8751
rect 13510 8442 13538 8447
rect 13398 8441 13538 8442
rect 13398 8415 13399 8441
rect 13425 8415 13511 8441
rect 13537 8415 13538 8441
rect 13398 8414 13538 8415
rect 13398 8409 13426 8414
rect 13342 8023 13343 8049
rect 13369 8023 13370 8049
rect 13342 7993 13370 8023
rect 13342 7967 13343 7993
rect 13369 7967 13370 7993
rect 13342 7266 13370 7967
rect 13398 7658 13426 7663
rect 13510 7658 13538 8414
rect 13398 7657 13538 7658
rect 13398 7631 13399 7657
rect 13425 7631 13511 7657
rect 13537 7631 13538 7657
rect 13398 7630 13538 7631
rect 13398 7625 13426 7630
rect 13398 7266 13426 7271
rect 13342 7265 13426 7266
rect 13342 7239 13399 7265
rect 13425 7239 13426 7265
rect 13342 7238 13426 7239
rect 12838 6847 12839 6873
rect 12865 6847 12866 6873
rect 12838 6762 12866 6847
rect 12838 6089 12866 6734
rect 13398 7209 13426 7238
rect 13398 7183 13399 7209
rect 13425 7183 13426 7209
rect 13398 6538 13426 7183
rect 13398 6481 13426 6510
rect 13398 6455 13399 6481
rect 13425 6455 13426 6481
rect 13398 6425 13426 6455
rect 13398 6399 13399 6425
rect 13425 6399 13426 6425
rect 13398 6393 13426 6399
rect 12838 6063 12839 6089
rect 12865 6063 12866 6089
rect 12838 6057 12866 6063
rect 13398 6090 13426 6095
rect 13510 6090 13538 7630
rect 13398 6089 13538 6090
rect 13398 6063 13399 6089
rect 13425 6063 13511 6089
rect 13537 6063 13538 6089
rect 13398 6062 13538 6063
rect 11998 5697 12026 5894
rect 12278 5698 12306 5703
rect 11998 5671 11999 5697
rect 12025 5671 12026 5697
rect 11998 5641 12026 5671
rect 11998 5615 11999 5641
rect 12025 5615 12026 5641
rect 11998 5609 12026 5615
rect 12222 5697 12306 5698
rect 12222 5671 12279 5697
rect 12305 5671 12306 5697
rect 12222 5670 12306 5671
rect 11102 4887 11103 4913
rect 11129 4887 11130 4913
rect 10430 4857 10794 4858
rect 10430 4831 10431 4857
rect 10457 4831 10794 4857
rect 10430 4830 10794 4831
rect 10038 4774 10122 4802
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10094 4634 10122 4774
rect 10038 4606 10122 4634
rect 10038 4521 10066 4606
rect 10038 4495 10039 4521
rect 10065 4495 10066 4521
rect 10038 4214 10066 4495
rect 9534 4103 9535 4129
rect 9561 4103 9562 4129
rect 9534 4097 9562 4103
rect 9814 4186 10066 4214
rect 8750 4074 8778 4079
rect 8470 4073 8778 4074
rect 8470 4047 8751 4073
rect 8777 4047 8778 4073
rect 8470 4046 8778 4047
rect 8470 2562 8498 4046
rect 8750 4041 8778 4046
rect 9814 3737 9842 4186
rect 10038 4074 10066 4186
rect 10038 4041 10066 4046
rect 10430 4129 10458 4830
rect 10766 4577 10794 4830
rect 10766 4551 10767 4577
rect 10793 4551 10794 4577
rect 10766 4521 10794 4551
rect 10766 4495 10767 4521
rect 10793 4495 10794 4521
rect 10766 4489 10794 4495
rect 10430 4103 10431 4129
rect 10457 4103 10458 4129
rect 10430 4073 10458 4103
rect 10430 4047 10431 4073
rect 10457 4047 10458 4073
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9814 3711 9815 3737
rect 9841 3711 9842 3737
rect 9814 3705 9842 3711
rect 10374 3738 10402 3743
rect 10430 3738 10458 4047
rect 11102 4129 11130 4887
rect 11382 5305 11410 5311
rect 11382 5279 11383 5305
rect 11409 5279 11410 5305
rect 11382 4521 11410 5279
rect 11382 4495 11383 4521
rect 11409 4495 11410 4521
rect 11382 4214 11410 4495
rect 11998 4914 12026 4919
rect 11998 4857 12026 4886
rect 11998 4831 11999 4857
rect 12025 4831 12026 4857
rect 11998 4521 12026 4831
rect 11998 4495 11999 4521
rect 12025 4495 12026 4521
rect 11998 4214 12026 4495
rect 11382 4186 11578 4214
rect 11102 4103 11103 4129
rect 11129 4103 11130 4129
rect 11102 4074 11130 4103
rect 11102 4041 11130 4046
rect 11550 4074 11578 4186
rect 11550 4041 11578 4046
rect 11718 4186 12026 4214
rect 10486 3738 10514 3743
rect 10374 3737 10514 3738
rect 10374 3711 10375 3737
rect 10401 3711 10487 3737
rect 10513 3711 10514 3737
rect 10374 3710 10514 3711
rect 10374 3705 10402 3710
rect 8470 2450 8498 2534
rect 8806 3345 8834 3351
rect 8806 3319 8807 3345
rect 8833 3319 8834 3345
rect 8806 3289 8834 3319
rect 8806 3263 8807 3289
rect 8833 3263 8834 3289
rect 8806 2506 8834 3263
rect 8806 2473 8834 2478
rect 9254 3346 9282 3351
rect 9254 2954 9282 3318
rect 9758 3346 9786 3351
rect 9926 3346 9954 3351
rect 9758 3345 9954 3346
rect 9758 3319 9759 3345
rect 9785 3319 9927 3345
rect 9953 3319 9954 3345
rect 9758 3318 9954 3319
rect 9310 2954 9338 2959
rect 9254 2926 9310 2954
rect 9254 2561 9282 2926
rect 9310 2888 9338 2926
rect 9758 2954 9786 3318
rect 9926 3313 9954 3318
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9982 2954 10010 2959
rect 9758 2953 10010 2954
rect 9758 2927 9759 2953
rect 9785 2927 9983 2953
rect 10009 2927 10010 2953
rect 9758 2926 10010 2927
rect 9254 2535 9255 2561
rect 9281 2535 9282 2561
rect 8470 2417 8498 2422
rect 8358 2199 8359 2225
rect 8385 2199 8386 2225
rect 8358 2169 8386 2199
rect 8358 2143 8359 2169
rect 8385 2143 8386 2169
rect 8358 2137 8386 2143
rect 9254 2169 9282 2535
rect 9254 2143 9255 2169
rect 9281 2143 9282 2169
rect 9254 2137 9282 2143
rect 9590 2450 9618 2455
rect 9590 2114 9618 2422
rect 9758 2450 9786 2926
rect 9982 2921 10010 2926
rect 9758 2417 9786 2422
rect 10430 2561 10458 3710
rect 10486 3705 10514 3710
rect 11102 3738 11130 3743
rect 11102 3346 11130 3710
rect 11550 3738 11578 3743
rect 11550 3691 11578 3710
rect 10430 2535 10431 2561
rect 10457 2535 10458 2561
rect 10430 2506 10458 2535
rect 11046 3345 11130 3346
rect 11046 3319 11103 3345
rect 11129 3319 11130 3345
rect 11046 3318 11130 3319
rect 11046 2954 11074 3318
rect 11102 3313 11130 3318
rect 11382 3346 11410 3351
rect 11494 3346 11522 3351
rect 11382 3345 11522 3346
rect 11382 3319 11383 3345
rect 11409 3319 11495 3345
rect 11521 3319 11522 3345
rect 11382 3318 11522 3319
rect 11046 2561 11074 2926
rect 11046 2535 11047 2561
rect 11073 2535 11074 2561
rect 11046 2529 11074 2535
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10430 2225 10458 2478
rect 10430 2199 10431 2225
rect 10457 2199 10458 2225
rect 10430 2170 10458 2199
rect 10430 2123 10458 2142
rect 10878 2282 10906 2287
rect 10878 2169 10906 2254
rect 10878 2143 10879 2169
rect 10905 2143 10906 2169
rect 8078 1689 8106 1694
rect 8302 1778 8330 1783
rect 8302 400 8330 1750
rect 9422 1778 9450 1783
rect 9422 1731 9450 1750
rect 9590 1778 9618 2086
rect 9814 1778 9842 1783
rect 9590 1777 9842 1778
rect 9590 1751 9591 1777
rect 9617 1751 9815 1777
rect 9841 1751 9842 1777
rect 9590 1750 9842 1751
rect 9590 1745 9618 1750
rect 9814 1745 9842 1750
rect 10878 1778 10906 2143
rect 11158 2169 11186 2175
rect 11158 2143 11159 2169
rect 11185 2143 11186 2169
rect 11158 2114 11186 2143
rect 11158 2081 11186 2086
rect 11382 2169 11410 3318
rect 11494 3290 11522 3318
rect 11494 3257 11522 3262
rect 11718 3009 11746 4186
rect 11774 4129 11802 4186
rect 11774 4103 11775 4129
rect 11801 4103 11802 4129
rect 11774 4073 11802 4103
rect 11774 4047 11775 4073
rect 11801 4047 11802 4073
rect 11774 4041 11802 4047
rect 12222 4074 12250 5670
rect 12278 5665 12306 5670
rect 13398 5697 13426 6062
rect 13510 6057 13538 6062
rect 13398 5671 13399 5697
rect 13425 5671 13426 5697
rect 13398 5641 13426 5671
rect 13398 5615 13399 5641
rect 13425 5615 13426 5641
rect 13398 5609 13426 5615
rect 12278 5361 12306 5367
rect 12278 5335 12279 5361
rect 12305 5335 12306 5361
rect 12278 5305 12306 5335
rect 12278 5279 12279 5305
rect 12305 5279 12306 5305
rect 12278 4914 12306 5279
rect 13118 5305 13146 5311
rect 13118 5279 13119 5305
rect 13145 5279 13146 5305
rect 12278 4577 12306 4886
rect 12278 4551 12279 4577
rect 12305 4551 12306 4577
rect 12278 4214 12306 4551
rect 12558 5026 12586 5031
rect 12558 4913 12586 4998
rect 12558 4887 12559 4913
rect 12585 4887 12586 4913
rect 12278 4186 12474 4214
rect 12222 4041 12250 4046
rect 12446 3793 12474 4186
rect 12446 3767 12447 3793
rect 12473 3767 12474 3793
rect 12446 3737 12474 3767
rect 12446 3711 12447 3737
rect 12473 3711 12474 3737
rect 12446 3402 12474 3711
rect 12558 4129 12586 4887
rect 13118 5026 13146 5279
rect 13118 4521 13146 4998
rect 13118 4495 13119 4521
rect 13145 4495 13146 4521
rect 13118 4489 13146 4495
rect 13398 4914 13426 4919
rect 13398 4857 13426 4886
rect 13398 4831 13399 4857
rect 13425 4831 13426 4857
rect 13398 4214 13426 4831
rect 13342 4186 13426 4214
rect 12558 4103 12559 4129
rect 12585 4103 12586 4129
rect 12558 3738 12586 4103
rect 13230 4129 13258 4135
rect 13230 4103 13231 4129
rect 13257 4103 13258 4129
rect 13230 4073 13258 4103
rect 13230 4047 13231 4073
rect 13257 4047 13258 4073
rect 12558 3705 12586 3710
rect 13118 3738 13146 3743
rect 12446 3369 12474 3374
rect 12558 3402 12586 3407
rect 11718 2983 11719 3009
rect 11745 2983 11746 3009
rect 11662 2954 11690 2959
rect 11718 2954 11746 2983
rect 11662 2953 11746 2954
rect 11662 2927 11663 2953
rect 11689 2927 11746 2953
rect 11662 2926 11746 2927
rect 12558 3345 12586 3374
rect 13118 3402 13146 3710
rect 12558 3319 12559 3345
rect 12585 3319 12586 3345
rect 11662 2561 11690 2926
rect 11662 2535 11663 2561
rect 11689 2535 11690 2561
rect 11662 2506 11690 2535
rect 12558 2561 12586 3319
rect 12726 3345 12754 3351
rect 12726 3319 12727 3345
rect 12753 3319 12754 3345
rect 12726 3290 12754 3319
rect 12726 3257 12754 3262
rect 12950 3345 12978 3351
rect 12950 3319 12951 3345
rect 12977 3319 12978 3345
rect 12950 3290 12978 3319
rect 12950 3257 12978 3262
rect 13118 2953 13146 3374
rect 13118 2927 13119 2953
rect 13145 2927 13146 2953
rect 13118 2921 13146 2927
rect 13230 3346 13258 4047
rect 13230 2954 13258 3318
rect 13286 3737 13314 3743
rect 13286 3711 13287 3737
rect 13313 3711 13314 3737
rect 13286 3626 13314 3711
rect 13342 3626 13370 4158
rect 13566 3737 13594 3743
rect 13566 3711 13567 3737
rect 13593 3711 13594 3737
rect 13566 3626 13594 3711
rect 13286 3598 13594 3626
rect 13286 3290 13314 3598
rect 13286 3257 13314 3262
rect 13230 2921 13258 2926
rect 13454 2954 13482 2959
rect 13454 2562 13482 2926
rect 12558 2535 12559 2561
rect 12585 2535 12586 2561
rect 11774 2506 11802 2511
rect 11662 2505 11802 2506
rect 11662 2479 11775 2505
rect 11801 2479 11802 2505
rect 11662 2478 11802 2479
rect 11382 2143 11383 2169
rect 11409 2143 11410 2169
rect 11382 2114 11410 2143
rect 11382 2081 11410 2086
rect 11606 2282 11634 2287
rect 10878 1712 10906 1750
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 11606 400 11634 2254
rect 11662 2170 11690 2478
rect 11774 2473 11802 2478
rect 12558 2282 12586 2535
rect 13398 2561 13482 2562
rect 13398 2535 13455 2561
rect 13481 2535 13482 2561
rect 13398 2534 13482 2535
rect 13398 2505 13426 2534
rect 13454 2529 13482 2534
rect 13398 2479 13399 2505
rect 13425 2479 13426 2505
rect 13398 2473 13426 2479
rect 12558 2249 12586 2254
rect 13622 2450 13650 10206
rect 13678 10122 13706 29600
rect 16142 27734 16170 29600
rect 18494 28770 18522 28775
rect 17598 27846 17730 27851
rect 17626 27818 17650 27846
rect 17678 27818 17702 27846
rect 17598 27813 17730 27818
rect 16030 27706 16170 27734
rect 15302 22890 15330 22895
rect 15470 22890 15498 22895
rect 15302 22889 15498 22890
rect 15302 22863 15303 22889
rect 15329 22863 15471 22889
rect 15497 22863 15498 22889
rect 15302 22862 15498 22863
rect 15302 22857 15330 22862
rect 15470 22610 15498 22862
rect 15582 22890 15610 22895
rect 15582 22843 15610 22862
rect 15862 22890 15890 22895
rect 15862 22843 15890 22862
rect 15974 22889 16002 22895
rect 15974 22863 15975 22889
rect 16001 22863 16002 22889
rect 15974 22666 16002 22863
rect 15974 22633 16002 22638
rect 15582 22610 15610 22615
rect 15470 22582 15582 22610
rect 15582 22563 15610 22582
rect 15750 22610 15778 22615
rect 15750 22563 15778 22582
rect 15862 22553 15890 22559
rect 15862 22527 15863 22553
rect 15889 22527 15890 22553
rect 15862 21826 15890 22527
rect 15862 21793 15890 21798
rect 16030 21266 16058 27706
rect 17598 27062 17730 27067
rect 17626 27034 17650 27062
rect 17678 27034 17702 27062
rect 17598 27029 17730 27034
rect 17598 26278 17730 26283
rect 17626 26250 17650 26278
rect 17678 26250 17702 26278
rect 17598 26245 17730 26250
rect 18102 25690 18130 25695
rect 17598 25494 17730 25499
rect 17626 25466 17650 25494
rect 17678 25466 17702 25494
rect 17598 25461 17730 25466
rect 17542 25298 17570 25303
rect 16982 24906 17010 24911
rect 16814 24514 16842 24519
rect 16198 23730 16226 23735
rect 16198 23338 16226 23702
rect 16478 23730 16506 23735
rect 16478 23683 16506 23702
rect 16590 23730 16618 23735
rect 16758 23730 16786 23735
rect 16814 23730 16842 24486
rect 16982 24458 17010 24878
rect 17150 24514 17178 24519
rect 17150 24467 17178 24486
rect 17318 24514 17346 24519
rect 16590 23729 16842 23730
rect 16590 23703 16591 23729
rect 16617 23703 16759 23729
rect 16785 23703 16842 23729
rect 16590 23702 16842 23703
rect 16926 24457 17010 24458
rect 16926 24431 16983 24457
rect 17009 24431 17010 24457
rect 16926 24430 17010 24431
rect 16142 23337 16226 23338
rect 16142 23311 16199 23337
rect 16225 23311 16226 23337
rect 16142 23310 16226 23311
rect 16142 22890 16170 23310
rect 16198 23305 16226 23310
rect 16310 23338 16338 23343
rect 16478 23338 16506 23343
rect 16590 23338 16618 23702
rect 16758 23697 16786 23702
rect 16310 23337 16618 23338
rect 16310 23311 16311 23337
rect 16337 23311 16479 23337
rect 16505 23311 16618 23337
rect 16310 23310 16618 23311
rect 16310 23305 16338 23310
rect 16142 22609 16170 22862
rect 16142 22583 16143 22609
rect 16169 22583 16170 22609
rect 16142 22162 16170 22583
rect 16198 22945 16226 22951
rect 16198 22919 16199 22945
rect 16225 22919 16226 22945
rect 16198 22666 16226 22919
rect 16198 22554 16226 22638
rect 16422 22946 16450 23310
rect 16478 23305 16506 23310
rect 16534 22946 16562 22951
rect 16422 22945 16562 22946
rect 16422 22919 16423 22945
rect 16449 22919 16535 22945
rect 16561 22919 16562 22945
rect 16422 22918 16562 22919
rect 16422 22610 16450 22918
rect 16422 22577 16450 22582
rect 16310 22554 16338 22559
rect 16198 22526 16310 22554
rect 16310 22507 16338 22526
rect 16478 22554 16506 22559
rect 16478 22507 16506 22526
rect 16142 22129 16170 22134
rect 16422 22162 16450 22167
rect 16422 22115 16450 22134
rect 16534 22162 16562 22918
rect 16702 22946 16730 22951
rect 16702 22899 16730 22918
rect 16870 22946 16898 22951
rect 16870 22609 16898 22918
rect 16870 22583 16871 22609
rect 16897 22583 16898 22609
rect 16870 22577 16898 22583
rect 16702 22162 16730 22167
rect 16534 22161 16730 22162
rect 16534 22135 16535 22161
rect 16561 22135 16703 22161
rect 16729 22135 16730 22161
rect 16534 22134 16730 22135
rect 16534 22129 16562 22134
rect 16702 22129 16730 22134
rect 16870 22162 16898 22167
rect 16870 21882 16898 22134
rect 16870 21769 16898 21854
rect 16870 21743 16871 21769
rect 16897 21743 16898 21769
rect 16870 21737 16898 21743
rect 16926 21826 16954 24430
rect 16982 24425 17010 24430
rect 17262 24178 17290 24183
rect 17038 24122 17066 24127
rect 17038 23730 17066 24094
rect 17206 24122 17234 24127
rect 17206 24075 17234 24094
rect 17038 23664 17066 23702
rect 17150 23730 17178 23735
rect 17262 23730 17290 24150
rect 17150 23729 17290 23730
rect 17150 23703 17151 23729
rect 17177 23703 17263 23729
rect 17289 23703 17290 23729
rect 17150 23702 17290 23703
rect 17150 23697 17178 23702
rect 17262 23697 17290 23702
rect 17206 23506 17234 23511
rect 17206 23338 17234 23478
rect 17038 23337 17234 23338
rect 17038 23311 17207 23337
rect 17233 23311 17234 23337
rect 17038 23310 17234 23311
rect 17038 22946 17066 23310
rect 17206 23305 17234 23310
rect 17318 23394 17346 24486
rect 17542 24514 17570 25270
rect 17822 25242 17850 25247
rect 17822 24962 17850 25214
rect 18102 25241 18130 25662
rect 18326 25298 18354 25303
rect 18102 25215 18103 25241
rect 18129 25215 18130 25241
rect 17990 24962 18018 24967
rect 17822 24961 18018 24962
rect 17822 24935 17823 24961
rect 17849 24935 17991 24961
rect 18017 24935 18018 24961
rect 17822 24934 18018 24935
rect 17710 24906 17738 24911
rect 17710 24859 17738 24878
rect 17598 24710 17730 24715
rect 17626 24682 17650 24710
rect 17678 24682 17702 24710
rect 17598 24677 17730 24682
rect 17710 24514 17738 24519
rect 17542 24513 17682 24514
rect 17542 24487 17543 24513
rect 17569 24487 17682 24513
rect 17542 24486 17682 24487
rect 17542 24481 17570 24486
rect 17430 24178 17458 24183
rect 17430 24131 17458 24150
rect 17654 24178 17682 24486
rect 17710 24467 17738 24486
rect 17710 24178 17738 24183
rect 17654 24177 17738 24178
rect 17654 24151 17711 24177
rect 17737 24151 17738 24177
rect 17654 24150 17738 24151
rect 17654 24122 17682 24150
rect 17710 24145 17738 24150
rect 17822 24178 17850 24934
rect 17990 24929 18018 24934
rect 18102 24906 18130 25215
rect 18214 25242 18242 25247
rect 18214 25195 18242 25214
rect 18130 24878 18186 24906
rect 18102 24873 18130 24878
rect 17822 24112 17850 24150
rect 17878 24514 17906 24519
rect 17654 24089 17682 24094
rect 17598 23926 17730 23931
rect 17626 23898 17650 23926
rect 17678 23898 17702 23926
rect 17598 23893 17730 23898
rect 17598 23729 17626 23735
rect 17598 23703 17599 23729
rect 17625 23703 17626 23729
rect 17598 23506 17626 23703
rect 17710 23730 17738 23735
rect 17878 23730 17906 24486
rect 18102 24457 18130 24463
rect 18102 24431 18103 24457
rect 18129 24431 18130 24457
rect 17990 24178 18018 24183
rect 17990 24131 18018 24150
rect 18102 23786 18130 24431
rect 18158 24178 18186 24878
rect 18326 24905 18354 25270
rect 18494 25298 18522 28742
rect 18550 25690 18578 25695
rect 18550 25643 18578 25662
rect 18494 25265 18522 25270
rect 18326 24879 18327 24905
rect 18353 24879 18354 24905
rect 18326 24873 18354 24879
rect 18382 25242 18410 25247
rect 18382 24962 18410 25214
rect 18550 24962 18578 24967
rect 18382 24961 18578 24962
rect 18382 24935 18383 24961
rect 18409 24935 18551 24961
rect 18577 24935 18578 24961
rect 18382 24934 18578 24935
rect 18270 24514 18298 24519
rect 18270 24467 18298 24486
rect 18158 24145 18186 24150
rect 18382 24178 18410 24934
rect 18550 24929 18578 24934
rect 18438 24514 18466 24519
rect 18438 24467 18466 24486
rect 18550 24178 18578 24183
rect 18382 24177 18578 24178
rect 18382 24151 18383 24177
rect 18409 24151 18551 24177
rect 18577 24151 18578 24177
rect 18382 24150 18578 24151
rect 18326 24121 18354 24127
rect 18326 24095 18327 24121
rect 18353 24095 18354 24121
rect 18326 23786 18354 24095
rect 18102 23758 18354 23786
rect 17710 23729 17906 23730
rect 17710 23703 17711 23729
rect 17737 23703 17879 23729
rect 17905 23703 17906 23729
rect 17710 23702 17906 23703
rect 17710 23697 17738 23702
rect 17878 23697 17906 23702
rect 18158 23729 18186 23758
rect 18158 23703 18159 23729
rect 18185 23703 18186 23729
rect 17990 23674 18018 23679
rect 17710 23506 17738 23511
rect 17542 23478 17710 23506
rect 17430 23394 17458 23399
rect 17318 23393 17458 23394
rect 17318 23367 17431 23393
rect 17457 23367 17458 23393
rect 17318 23366 17458 23367
rect 17318 23337 17346 23366
rect 17430 23361 17458 23366
rect 17318 23311 17319 23337
rect 17345 23311 17346 23337
rect 17038 22880 17066 22918
rect 17150 22946 17178 22951
rect 17318 22946 17346 23311
rect 17542 22946 17570 23478
rect 17710 23393 17738 23478
rect 17990 23394 18018 23646
rect 17710 23367 17711 23393
rect 17737 23367 17738 23393
rect 17710 23361 17738 23367
rect 17878 23393 18018 23394
rect 17878 23367 17991 23393
rect 18017 23367 18018 23393
rect 17878 23366 18018 23367
rect 17878 23337 17906 23366
rect 17990 23361 18018 23366
rect 17878 23311 17879 23337
rect 17905 23311 17906 23337
rect 17598 23142 17730 23147
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17598 23109 17730 23114
rect 17150 22945 17346 22946
rect 17150 22919 17151 22945
rect 17177 22919 17319 22945
rect 17345 22919 17346 22945
rect 17150 22918 17346 22919
rect 17150 22610 17178 22918
rect 17318 22913 17346 22918
rect 17486 22945 17570 22946
rect 17486 22919 17543 22945
rect 17569 22919 17570 22945
rect 17486 22918 17570 22919
rect 17038 22582 17150 22610
rect 17038 22553 17066 22582
rect 17038 22527 17039 22553
rect 17065 22527 17066 22553
rect 17038 22521 17066 22527
rect 16982 22162 17010 22167
rect 16982 22115 17010 22134
rect 16926 21378 16954 21798
rect 17038 21770 17066 21775
rect 17094 21770 17122 22582
rect 17150 22544 17178 22582
rect 17430 22610 17458 22615
rect 17150 22162 17178 22167
rect 17318 22162 17346 22167
rect 17150 22161 17346 22162
rect 17150 22135 17151 22161
rect 17177 22135 17319 22161
rect 17345 22135 17346 22161
rect 17150 22134 17346 22135
rect 17430 22162 17458 22582
rect 17486 22553 17514 22918
rect 17542 22913 17570 22918
rect 17710 22946 17738 22951
rect 17878 22946 17906 23311
rect 18158 22946 18186 23703
rect 18214 23674 18242 23679
rect 18214 23627 18242 23646
rect 18326 23506 18354 23758
rect 18326 23337 18354 23478
rect 18326 23311 18327 23337
rect 18353 23311 18354 23337
rect 18326 23305 18354 23311
rect 18382 23729 18410 24150
rect 18550 24145 18578 24150
rect 18382 23703 18383 23729
rect 18409 23703 18410 23729
rect 18382 23674 18410 23703
rect 18382 23394 18410 23646
rect 18550 23394 18578 23399
rect 18382 23393 18578 23394
rect 18382 23367 18383 23393
rect 18409 23367 18551 23393
rect 18577 23367 18578 23393
rect 18382 23366 18578 23367
rect 17710 22945 17906 22946
rect 17710 22919 17711 22945
rect 17737 22919 17879 22945
rect 17905 22919 17906 22945
rect 17710 22918 17906 22919
rect 17710 22609 17738 22918
rect 17878 22913 17906 22918
rect 17990 22945 18186 22946
rect 17990 22919 18159 22945
rect 18185 22919 18186 22945
rect 17990 22918 18186 22919
rect 17710 22583 17711 22609
rect 17737 22583 17738 22609
rect 17710 22577 17738 22583
rect 17486 22527 17487 22553
rect 17513 22527 17514 22553
rect 17486 22521 17514 22527
rect 17542 22554 17570 22559
rect 17542 22274 17570 22526
rect 17598 22358 17730 22363
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17598 22325 17730 22330
rect 17542 22246 17626 22274
rect 17486 22162 17514 22167
rect 17430 22161 17514 22162
rect 17430 22135 17487 22161
rect 17513 22135 17514 22161
rect 17430 22134 17514 22135
rect 17150 22129 17178 22134
rect 17150 21770 17178 21775
rect 17038 21769 17178 21770
rect 17038 21743 17039 21769
rect 17065 21743 17151 21769
rect 17177 21743 17178 21769
rect 17038 21742 17178 21743
rect 17038 21737 17066 21742
rect 16982 21378 17010 21383
rect 16926 21377 17010 21378
rect 16926 21351 16983 21377
rect 17009 21351 17010 21377
rect 16926 21350 17010 21351
rect 16030 21233 16058 21238
rect 16982 21042 17010 21350
rect 17150 21378 17178 21742
rect 17318 21770 17346 22134
rect 17486 22129 17514 22134
rect 17318 21737 17346 21742
rect 17486 21882 17514 21887
rect 17486 21769 17514 21854
rect 17486 21743 17487 21769
rect 17513 21743 17514 21769
rect 17262 21378 17290 21383
rect 17150 21377 17290 21378
rect 17150 21351 17151 21377
rect 17177 21351 17263 21377
rect 17289 21351 17290 21377
rect 17150 21350 17290 21351
rect 17486 21378 17514 21743
rect 17598 21770 17626 22246
rect 17710 22106 17738 22111
rect 17710 22105 17794 22106
rect 17710 22079 17711 22105
rect 17737 22079 17794 22105
rect 17710 22078 17794 22079
rect 17710 22073 17738 22078
rect 17598 21723 17626 21742
rect 17710 21770 17738 21775
rect 17710 21723 17738 21742
rect 17598 21574 17730 21579
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17598 21541 17730 21546
rect 17542 21378 17570 21383
rect 17486 21377 17570 21378
rect 17486 21351 17543 21377
rect 17569 21351 17570 21377
rect 17486 21350 17570 21351
rect 17150 21345 17178 21350
rect 17262 21345 17290 21350
rect 17542 21345 17570 21350
rect 17710 21378 17738 21383
rect 17766 21378 17794 22078
rect 17822 22105 17850 22111
rect 17822 22079 17823 22105
rect 17849 22079 17850 22105
rect 17822 21882 17850 22079
rect 17822 21849 17850 21854
rect 17990 21602 18018 22918
rect 18158 22913 18186 22918
rect 18270 22946 18298 22951
rect 18382 22946 18410 23366
rect 18550 23361 18578 23366
rect 18270 22945 18410 22946
rect 18270 22919 18271 22945
rect 18297 22919 18383 22945
rect 18409 22919 18410 22945
rect 18270 22918 18410 22919
rect 18270 22913 18298 22918
rect 18102 22610 18130 22615
rect 18046 22553 18074 22559
rect 18046 22527 18047 22553
rect 18073 22527 18074 22553
rect 18046 21882 18074 22527
rect 18046 21769 18074 21854
rect 18046 21743 18047 21769
rect 18073 21743 18074 21769
rect 18046 21737 18074 21743
rect 18102 21770 18130 22582
rect 18270 22610 18298 22615
rect 18270 22563 18298 22582
rect 18158 22161 18186 22167
rect 18158 22135 18159 22161
rect 18185 22135 18186 22161
rect 18158 21882 18186 22135
rect 18270 22162 18298 22167
rect 18382 22162 18410 22918
rect 18270 22161 18410 22162
rect 18270 22135 18271 22161
rect 18297 22135 18383 22161
rect 18409 22135 18410 22161
rect 18270 22134 18410 22135
rect 18270 22129 18298 22134
rect 18158 21849 18186 21854
rect 18158 21770 18186 21775
rect 18326 21770 18354 21775
rect 18102 21769 18354 21770
rect 18102 21743 18159 21769
rect 18185 21743 18327 21769
rect 18353 21743 18354 21769
rect 18102 21742 18354 21743
rect 18158 21737 18186 21742
rect 17990 21574 18130 21602
rect 17710 21377 17794 21378
rect 17710 21351 17711 21377
rect 17737 21351 17794 21377
rect 17710 21350 17794 21351
rect 17710 21345 17738 21350
rect 17766 21098 17794 21350
rect 17878 21377 17906 21383
rect 17878 21351 17879 21377
rect 17905 21351 17906 21377
rect 17878 21098 17906 21351
rect 18102 21377 18130 21574
rect 18102 21351 18103 21377
rect 18129 21351 18130 21377
rect 18102 21345 18130 21351
rect 18214 21321 18242 21327
rect 18214 21295 18215 21321
rect 18241 21295 18242 21321
rect 17990 21266 18018 21271
rect 17934 21098 17962 21103
rect 17766 21070 17934 21098
rect 16982 21009 17010 21014
rect 17654 21042 17682 21047
rect 17654 20995 17682 21014
rect 17766 21041 17794 21070
rect 17766 21015 17767 21041
rect 17793 21015 17794 21041
rect 17766 21009 17794 21015
rect 17934 21041 17962 21070
rect 17934 21015 17935 21041
rect 17961 21015 17962 21041
rect 17934 21009 17962 21015
rect 17598 20790 17730 20795
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17598 20757 17730 20762
rect 14630 20258 14658 20263
rect 14574 20202 14602 20207
rect 14574 20155 14602 20174
rect 14574 19418 14602 19423
rect 14630 19418 14658 20230
rect 15246 20257 15274 20263
rect 15246 20231 15247 20257
rect 15273 20231 15274 20257
rect 15078 20202 15106 20207
rect 15078 19809 15106 20174
rect 15078 19783 15079 19809
rect 15105 19783 15106 19809
rect 14574 19417 14882 19418
rect 14574 19391 14575 19417
rect 14601 19391 14882 19417
rect 14574 19390 14882 19391
rect 14574 19385 14602 19390
rect 14854 19025 14882 19390
rect 14854 18999 14855 19025
rect 14881 18999 14882 19025
rect 14574 18633 14602 18639
rect 14574 18607 14575 18633
rect 14601 18607 14602 18633
rect 14574 17849 14602 18607
rect 14574 17823 14575 17849
rect 14601 17823 14602 17849
rect 14574 17458 14602 17823
rect 14854 18241 14882 18999
rect 15078 18298 15106 19783
rect 15078 18265 15106 18270
rect 15246 20201 15274 20231
rect 15246 20175 15247 20201
rect 15273 20175 15274 20201
rect 15246 19810 15274 20175
rect 17598 20006 17730 20011
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17598 19973 17730 19978
rect 15470 19810 15498 19815
rect 15246 19809 15498 19810
rect 15246 19783 15247 19809
rect 15273 19783 15471 19809
rect 15497 19783 15498 19809
rect 15246 19782 15498 19783
rect 15246 18690 15274 19782
rect 15470 19777 15498 19782
rect 15470 19473 15498 19479
rect 15470 19447 15471 19473
rect 15497 19447 15498 19473
rect 15470 19417 15498 19447
rect 15470 19391 15471 19417
rect 15497 19391 15498 19417
rect 15470 19026 15498 19391
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 15918 19026 15946 19031
rect 15470 19025 15946 19026
rect 15470 18999 15919 19025
rect 15945 18999 15946 19025
rect 15470 18998 15946 18999
rect 15246 18633 15274 18662
rect 15246 18607 15247 18633
rect 15273 18607 15274 18633
rect 14854 18215 14855 18241
rect 14881 18215 14882 18241
rect 14798 17458 14826 17463
rect 14574 17457 14826 17458
rect 14574 17431 14799 17457
rect 14825 17431 14826 17457
rect 14574 17430 14826 17431
rect 14574 17066 14602 17430
rect 14798 17425 14826 17430
rect 14854 17458 14882 18215
rect 14574 17000 14602 17038
rect 14798 16674 14826 16679
rect 14854 16674 14882 17430
rect 14798 16673 14882 16674
rect 14798 16647 14799 16673
rect 14825 16647 14882 16673
rect 14798 16646 14882 16647
rect 15246 17905 15274 18607
rect 15918 18969 15946 18998
rect 16254 19026 16282 19031
rect 16254 18979 16282 18998
rect 16814 19026 16842 19031
rect 16926 19026 16954 19031
rect 16814 19025 16954 19026
rect 16814 18999 16815 19025
rect 16841 18999 16927 19025
rect 16953 18999 16954 19025
rect 16814 18998 16954 18999
rect 15918 18943 15919 18969
rect 15945 18943 15946 18969
rect 15918 18242 15946 18943
rect 16814 18690 16842 18998
rect 16926 18993 16954 18998
rect 16814 18657 16842 18662
rect 17990 18689 18018 21238
rect 18214 21098 18242 21295
rect 18326 21322 18354 21742
rect 18382 21770 18410 22134
rect 18550 22553 18578 22559
rect 18550 22527 18551 22553
rect 18577 22527 18578 22553
rect 18550 21882 18578 22527
rect 18550 21825 18578 21854
rect 18550 21799 18551 21825
rect 18577 21799 18578 21825
rect 18550 21793 18578 21799
rect 18382 21737 18410 21742
rect 18382 21322 18410 21327
rect 18326 21294 18382 21322
rect 18102 21042 18130 21047
rect 18102 20593 18130 21014
rect 18214 21042 18242 21070
rect 18382 21042 18410 21294
rect 18214 21041 18466 21042
rect 18214 21015 18215 21041
rect 18241 21015 18383 21041
rect 18409 21015 18466 21041
rect 18214 21014 18466 21015
rect 18214 21009 18242 21014
rect 18382 21009 18410 21014
rect 18438 20874 18466 21014
rect 18494 20986 18522 20991
rect 18494 20939 18522 20958
rect 18438 20846 18522 20874
rect 18102 20567 18103 20593
rect 18129 20567 18130 20593
rect 18102 20561 18130 20567
rect 18270 20594 18298 20599
rect 18438 20594 18466 20599
rect 18270 20593 18438 20594
rect 18270 20567 18271 20593
rect 18297 20567 18438 20593
rect 18270 20566 18438 20567
rect 18270 20561 18298 20566
rect 18438 20547 18466 20566
rect 18102 19810 18130 19815
rect 18102 19763 18130 19782
rect 18270 19810 18298 19815
rect 18270 19763 18298 19782
rect 18494 19810 18522 20846
rect 18494 19777 18522 19782
rect 18382 19754 18410 19759
rect 18382 19707 18410 19726
rect 17990 18663 17991 18689
rect 18017 18663 18018 18689
rect 17990 18633 18018 18663
rect 17990 18607 17991 18633
rect 18017 18607 18018 18633
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 15918 18185 15946 18214
rect 16254 18298 16282 18303
rect 16254 18241 16282 18270
rect 16814 18298 16842 18303
rect 16254 18215 16255 18241
rect 16281 18215 16282 18241
rect 16254 18209 16282 18215
rect 16758 18242 16786 18247
rect 16758 18195 16786 18214
rect 15918 18159 15919 18185
rect 15945 18159 15946 18185
rect 15918 18153 15946 18159
rect 15246 17879 15247 17905
rect 15273 17879 15274 17905
rect 15246 17849 15274 17879
rect 15246 17823 15247 17849
rect 15273 17823 15274 17849
rect 15246 17458 15274 17823
rect 16814 17849 16842 18270
rect 16926 18242 16954 18247
rect 16926 18195 16954 18214
rect 17262 18242 17290 18247
rect 16814 17823 16815 17849
rect 16841 17823 16842 17849
rect 15470 17458 15498 17463
rect 15246 17457 15498 17458
rect 15246 17431 15247 17457
rect 15273 17431 15471 17457
rect 15497 17431 15498 17457
rect 15246 17430 15498 17431
rect 15246 17121 15274 17430
rect 15470 17425 15498 17430
rect 16254 17458 16282 17463
rect 16254 17411 16282 17430
rect 15246 17095 15247 17121
rect 15273 17095 15274 17121
rect 15246 17065 15274 17095
rect 15246 17039 15247 17065
rect 15273 17039 15274 17065
rect 15246 16674 15274 17039
rect 16814 17065 16842 17823
rect 16814 17039 16815 17065
rect 16841 17039 16842 17065
rect 15470 16674 15498 16679
rect 15246 16673 15498 16674
rect 15246 16647 15247 16673
rect 15273 16647 15471 16673
rect 15497 16647 15498 16673
rect 15246 16646 15498 16647
rect 14294 16281 14322 16287
rect 14294 16255 14295 16281
rect 14321 16255 14322 16281
rect 14294 15890 14322 16255
rect 14294 15498 14322 15862
rect 14798 15890 14826 16646
rect 15246 16337 15274 16646
rect 15470 16641 15498 16646
rect 16254 16673 16282 16679
rect 16254 16647 16255 16673
rect 16281 16647 16282 16673
rect 15246 16311 15247 16337
rect 15273 16311 15274 16337
rect 15246 16281 15274 16311
rect 15246 16255 15247 16281
rect 15273 16255 15274 16281
rect 15246 15974 15274 16255
rect 15246 15946 15330 15974
rect 14798 15843 14826 15862
rect 15190 15890 15218 15895
rect 14294 15451 14322 15470
rect 15190 15554 15218 15862
rect 15190 15497 15218 15526
rect 15190 15471 15191 15497
rect 15217 15471 15218 15497
rect 14798 15105 14826 15111
rect 14798 15079 14799 15105
rect 14825 15079 14826 15105
rect 14294 14713 14322 14719
rect 14294 14687 14295 14713
rect 14321 14687 14322 14713
rect 14294 13929 14322 14687
rect 14294 13903 14295 13929
rect 14321 13903 14322 13929
rect 14294 13145 14322 13903
rect 14294 13119 14295 13145
rect 14321 13119 14322 13145
rect 14294 12754 14322 13119
rect 14798 14322 14826 15079
rect 14798 13537 14826 14294
rect 14798 13511 14799 13537
rect 14825 13511 14826 13537
rect 14798 12754 14826 13511
rect 14294 12753 14826 12754
rect 14294 12727 14799 12753
rect 14825 12727 14826 12753
rect 14294 12726 14826 12727
rect 14294 12362 14322 12726
rect 14798 12721 14826 12726
rect 15190 14266 15218 15471
rect 14294 12315 14322 12334
rect 13678 10089 13706 10094
rect 14574 11970 14602 11975
rect 14574 11577 14602 11942
rect 15078 11970 15106 11975
rect 15078 11923 15106 11942
rect 14574 11551 14575 11577
rect 14601 11551 14602 11577
rect 14294 9226 14322 9231
rect 14294 8890 14322 9198
rect 14294 8441 14322 8862
rect 14574 8834 14602 11551
rect 15134 11578 15162 11583
rect 15134 11531 15162 11550
rect 15190 10094 15218 14238
rect 15246 15889 15274 15946
rect 15246 15863 15247 15889
rect 15273 15863 15274 15889
rect 15246 15106 15274 15863
rect 15302 15890 15330 15946
rect 15470 15890 15498 15895
rect 15302 15889 15498 15890
rect 15302 15863 15471 15889
rect 15497 15863 15498 15889
rect 15302 15862 15498 15863
rect 15470 15857 15498 15862
rect 16254 15889 16282 16647
rect 16814 16282 16842 17039
rect 16254 15863 16255 15889
rect 16281 15863 16282 15889
rect 15302 15554 15330 15559
rect 15302 15507 15330 15526
rect 16254 15498 16282 15863
rect 16758 16281 16842 16282
rect 16758 16255 16815 16281
rect 16841 16255 16842 16281
rect 16758 16254 16842 16255
rect 16758 15498 16786 16254
rect 16814 16249 16842 16254
rect 17262 17850 17290 18214
rect 17486 17850 17514 17855
rect 17262 17849 17514 17850
rect 17262 17823 17263 17849
rect 17289 17823 17487 17849
rect 17513 17823 17514 17849
rect 17262 17822 17514 17823
rect 17262 17457 17290 17822
rect 17486 17817 17514 17822
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17262 17431 17263 17457
rect 17289 17431 17290 17457
rect 17262 17401 17290 17431
rect 17262 17375 17263 17401
rect 17289 17375 17290 17401
rect 17262 17066 17290 17375
rect 17486 17066 17514 17071
rect 17262 17065 17514 17066
rect 17262 17039 17263 17065
rect 17289 17039 17487 17065
rect 17513 17039 17514 17065
rect 17262 17038 17514 17039
rect 17262 16673 17290 17038
rect 17486 17033 17514 17038
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17262 16647 17263 16673
rect 17289 16647 17290 16673
rect 17262 16617 17290 16647
rect 17262 16591 17263 16617
rect 17289 16591 17290 16617
rect 17262 16282 17290 16591
rect 17486 16282 17514 16287
rect 17262 16281 17514 16282
rect 17262 16255 17263 16281
rect 17289 16255 17487 16281
rect 17513 16255 17514 16281
rect 17262 16254 17514 16255
rect 17262 15974 17290 16254
rect 17486 16249 17514 16254
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17990 15974 18018 18607
rect 17206 15946 17290 15974
rect 17878 15946 18018 15974
rect 16814 15890 16842 15895
rect 16926 15890 16954 15895
rect 16842 15889 16954 15890
rect 16842 15863 16927 15889
rect 16953 15863 16954 15889
rect 16842 15862 16954 15863
rect 16814 15843 16842 15862
rect 16926 15857 16954 15862
rect 17206 15890 17234 15946
rect 17234 15862 17290 15890
rect 17206 15857 17234 15862
rect 16814 15498 16842 15503
rect 16254 15497 16842 15498
rect 16254 15471 16815 15497
rect 16841 15471 16842 15497
rect 16254 15470 16842 15471
rect 15470 15106 15498 15111
rect 15246 15105 15498 15106
rect 15246 15079 15247 15105
rect 15273 15079 15471 15105
rect 15497 15079 15498 15105
rect 15246 15078 15498 15079
rect 15246 14769 15274 15078
rect 15470 15073 15498 15078
rect 15246 14743 15247 14769
rect 15273 14743 15274 14769
rect 15246 14713 15274 14743
rect 15246 14687 15247 14713
rect 15273 14687 15274 14713
rect 15246 14322 15274 14687
rect 15470 14322 15498 14327
rect 15246 14321 15498 14322
rect 15246 14295 15247 14321
rect 15273 14295 15471 14321
rect 15497 14295 15498 14321
rect 15246 14294 15498 14295
rect 15246 13985 15274 14294
rect 15470 14289 15498 14294
rect 15246 13959 15247 13985
rect 15273 13959 15274 13985
rect 15246 13929 15274 13959
rect 15246 13903 15247 13929
rect 15273 13903 15274 13929
rect 15246 13538 15274 13903
rect 15470 13538 15498 13543
rect 15246 13537 15470 13538
rect 15246 13511 15247 13537
rect 15273 13511 15470 13537
rect 15246 13510 15470 13511
rect 15246 13201 15274 13510
rect 15470 13472 15498 13510
rect 15246 13175 15247 13201
rect 15273 13175 15274 13201
rect 15246 13145 15274 13175
rect 15246 13119 15247 13145
rect 15273 13119 15274 13145
rect 15246 12754 15274 13119
rect 15470 12754 15498 12759
rect 15246 12753 15498 12754
rect 15246 12727 15247 12753
rect 15273 12727 15471 12753
rect 15497 12727 15498 12753
rect 15246 12726 15498 12727
rect 15246 12417 15274 12726
rect 15470 12721 15498 12726
rect 16254 12753 16282 15470
rect 16814 15465 16842 15470
rect 17262 15498 17290 15862
rect 17486 15498 17514 15503
rect 17262 15497 17514 15498
rect 17262 15471 17263 15497
rect 17289 15471 17487 15497
rect 17513 15471 17514 15497
rect 17262 15470 17514 15471
rect 17262 15465 17290 15470
rect 17486 15465 17514 15470
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 16534 15105 16562 15111
rect 16534 15079 16535 15105
rect 16561 15079 16562 15105
rect 16534 14322 16562 15079
rect 17262 15105 17290 15111
rect 17262 15079 17263 15105
rect 17289 15079 17290 15105
rect 17262 15049 17290 15079
rect 17262 15023 17263 15049
rect 17289 15023 17290 15049
rect 16534 13537 16562 14294
rect 16814 14713 16842 14719
rect 16814 14687 16815 14713
rect 16841 14687 16842 14713
rect 16814 14322 16842 14687
rect 16814 13929 16842 14294
rect 16814 13903 16815 13929
rect 16841 13903 16842 13929
rect 16814 13897 16842 13903
rect 17262 14714 17290 15023
rect 17486 14714 17514 14719
rect 17262 14713 17514 14714
rect 17262 14687 17263 14713
rect 17289 14687 17487 14713
rect 17513 14687 17514 14713
rect 17262 14686 17514 14687
rect 17262 14321 17290 14686
rect 17486 14681 17514 14686
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17262 14295 17263 14321
rect 17289 14295 17290 14321
rect 17262 14265 17290 14295
rect 17262 14239 17263 14265
rect 17289 14239 17290 14265
rect 17262 13930 17290 14239
rect 17486 13930 17514 13935
rect 17262 13929 17514 13930
rect 17262 13903 17263 13929
rect 17289 13903 17487 13929
rect 17513 13903 17514 13929
rect 17262 13902 17514 13903
rect 16534 13511 16535 13537
rect 16561 13511 16562 13537
rect 16534 13505 16562 13511
rect 16814 13538 16842 13543
rect 16926 13538 16954 13543
rect 16842 13537 16954 13538
rect 16842 13511 16927 13537
rect 16953 13511 16954 13537
rect 16842 13510 16954 13511
rect 16814 13491 16842 13510
rect 16254 12727 16255 12753
rect 16281 12727 16282 12753
rect 15246 12391 15247 12417
rect 15273 12391 15274 12417
rect 15246 12361 15274 12391
rect 15246 12335 15247 12361
rect 15273 12335 15274 12361
rect 15246 11970 15274 12335
rect 15470 11970 15498 11975
rect 15246 11969 15498 11970
rect 15246 11943 15247 11969
rect 15273 11943 15471 11969
rect 15497 11943 15498 11969
rect 15246 11942 15498 11943
rect 15246 11633 15274 11942
rect 15470 11937 15498 11942
rect 16254 11970 16282 12727
rect 16814 12754 16842 12759
rect 16926 12754 16954 13510
rect 17262 13538 17290 13902
rect 17486 13897 17514 13902
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 17262 13505 17290 13510
rect 17878 13201 17906 15946
rect 17878 13175 17879 13201
rect 17905 13175 17906 13201
rect 17878 13145 17906 13175
rect 17878 13119 17879 13145
rect 17905 13119 17906 13145
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 16814 12753 16954 12754
rect 16814 12727 16815 12753
rect 16841 12727 16927 12753
rect 16953 12727 16954 12753
rect 16814 12726 16954 12727
rect 16814 12721 16842 12726
rect 16926 12721 16954 12726
rect 17878 12417 17906 13119
rect 17878 12391 17879 12417
rect 17905 12391 17906 12417
rect 17878 12361 17906 12391
rect 17878 12335 17879 12361
rect 17905 12335 17906 12361
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 16254 11937 16282 11942
rect 17486 11969 17514 11975
rect 17486 11943 17487 11969
rect 17513 11943 17514 11969
rect 15246 11607 15247 11633
rect 15273 11607 15274 11633
rect 15246 11578 15274 11607
rect 15246 11545 15274 11550
rect 15974 11185 16002 11191
rect 15974 11159 15975 11185
rect 16001 11159 16002 11185
rect 15974 11129 16002 11159
rect 15974 11103 15975 11129
rect 16001 11103 16002 11129
rect 15470 10849 15498 10855
rect 15470 10823 15471 10849
rect 15497 10823 15498 10849
rect 15470 10794 15498 10823
rect 15974 10794 16002 11103
rect 16926 11185 16954 11191
rect 16926 11159 16927 11185
rect 16953 11159 16954 11185
rect 15470 10793 16002 10794
rect 15470 10767 15471 10793
rect 15497 10767 16002 10793
rect 15470 10766 16002 10767
rect 16422 10793 16450 10799
rect 16422 10767 16423 10793
rect 16449 10767 16450 10793
rect 15470 10761 15498 10766
rect 15750 10401 15778 10766
rect 15750 10375 15751 10401
rect 15777 10375 15778 10401
rect 15750 10345 15778 10375
rect 15750 10319 15751 10345
rect 15777 10319 15778 10345
rect 15190 10066 15442 10094
rect 14742 9282 14770 9287
rect 14742 9226 14770 9254
rect 14966 9226 14994 9231
rect 14742 9225 15106 9226
rect 14742 9199 14743 9225
rect 14769 9199 14967 9225
rect 14993 9199 15106 9225
rect 14742 9198 15106 9199
rect 14742 9193 14770 9198
rect 14966 9193 14994 9198
rect 15078 9170 15106 9198
rect 15078 9142 15162 9170
rect 14574 8801 14602 8806
rect 14798 8890 14826 8895
rect 14798 8833 14826 8862
rect 14798 8807 14799 8833
rect 14825 8807 14826 8833
rect 14798 8801 14826 8807
rect 15134 8834 15162 9142
rect 15134 8801 15162 8806
rect 15246 8834 15274 8839
rect 14294 8415 14295 8441
rect 14321 8415 14322 8441
rect 14294 8050 14322 8415
rect 14294 7657 14322 8022
rect 15190 8106 15218 8111
rect 15190 8049 15218 8078
rect 15190 8023 15191 8049
rect 15217 8023 15218 8049
rect 15190 8017 15218 8023
rect 14294 7631 14295 7657
rect 14321 7631 14322 7657
rect 14294 7625 14322 7631
rect 14798 7265 14826 7271
rect 14798 7239 14799 7265
rect 14825 7239 14826 7265
rect 14014 6929 14042 6935
rect 14014 6903 14015 6929
rect 14041 6903 14042 6929
rect 14014 6873 14042 6903
rect 14014 6847 14015 6873
rect 14041 6847 14042 6873
rect 14014 6538 14042 6847
rect 14294 6873 14322 6879
rect 14294 6847 14295 6873
rect 14321 6847 14322 6873
rect 14294 6762 14322 6847
rect 14294 6729 14322 6734
rect 14798 6762 14826 7239
rect 15246 7266 15274 8806
rect 15414 8610 15442 10066
rect 15750 10010 15778 10319
rect 16422 10402 16450 10767
rect 15974 10010 16002 10015
rect 15750 10009 16002 10010
rect 15750 9983 15751 10009
rect 15777 9983 15975 10009
rect 16001 9983 16002 10009
rect 15750 9982 16002 9983
rect 15750 9977 15778 9982
rect 15974 9562 16002 9982
rect 16422 10009 16450 10374
rect 16926 10402 16954 11159
rect 17486 11185 17514 11943
rect 17766 11970 17794 11975
rect 17878 11970 17906 12335
rect 17766 11969 17906 11970
rect 17766 11943 17767 11969
rect 17793 11943 17879 11969
rect 17905 11943 17906 11969
rect 17766 11942 17906 11943
rect 17766 11937 17794 11942
rect 17878 11633 17906 11942
rect 17878 11607 17879 11633
rect 17905 11607 17906 11633
rect 17878 11577 17906 11607
rect 17878 11551 17879 11577
rect 17905 11551 17906 11577
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 17486 11159 17487 11185
rect 17513 11159 17514 11185
rect 16926 10355 16954 10374
rect 17206 10402 17234 10407
rect 16422 9983 16423 10009
rect 16449 9983 16450 10009
rect 16422 9977 16450 9983
rect 17150 10346 17178 10351
rect 15974 9529 16002 9534
rect 16254 9617 16282 9623
rect 16254 9591 16255 9617
rect 16281 9591 16282 9617
rect 16254 9562 16282 9591
rect 16254 9529 16282 9534
rect 16478 9617 16506 9623
rect 16478 9591 16479 9617
rect 16505 9591 16506 9617
rect 16478 9562 16506 9591
rect 16758 9618 16786 9623
rect 16758 9571 16786 9590
rect 17150 9618 17178 10318
rect 16478 9529 16506 9534
rect 15470 8834 15498 8839
rect 15470 8787 15498 8806
rect 15246 6929 15274 7238
rect 15246 6903 15247 6929
rect 15273 6903 15274 6929
rect 15246 6873 15274 6903
rect 15246 6847 15247 6873
rect 15273 6847 15274 6873
rect 15246 6841 15274 6847
rect 15302 8582 15442 8610
rect 14798 6729 14826 6734
rect 14014 5361 14042 6510
rect 15246 6538 15274 6543
rect 14014 5335 14015 5361
rect 14041 5335 14042 5361
rect 14014 5305 14042 5335
rect 14014 5279 14015 5305
rect 14041 5279 14042 5305
rect 14014 4914 14042 5279
rect 14574 6482 14602 6487
rect 14574 6089 14602 6454
rect 14574 6063 14575 6089
rect 14601 6063 14602 6089
rect 14574 5305 14602 6063
rect 14910 6482 14938 6487
rect 14910 5697 14938 6454
rect 15246 6481 15274 6510
rect 15246 6455 15247 6481
rect 15273 6455 15274 6481
rect 15246 6145 15274 6455
rect 15246 6119 15247 6145
rect 15273 6119 15274 6145
rect 15246 6089 15274 6119
rect 15246 6063 15247 6089
rect 15273 6063 15274 6089
rect 15246 6057 15274 6063
rect 14910 5671 14911 5697
rect 14937 5671 14938 5697
rect 14910 5665 14938 5671
rect 14574 5279 14575 5305
rect 14601 5279 14602 5305
rect 14574 5026 14602 5279
rect 14602 4998 14658 5026
rect 14574 4993 14602 4998
rect 14014 4881 14042 4886
rect 14574 4914 14602 4919
rect 14014 4577 14042 4583
rect 14014 4551 14015 4577
rect 14041 4551 14042 4577
rect 14014 4521 14042 4551
rect 14574 4522 14602 4886
rect 14014 4495 14015 4521
rect 14041 4495 14042 4521
rect 14014 3009 14042 4495
rect 14518 4521 14602 4522
rect 14518 4495 14575 4521
rect 14601 4495 14602 4521
rect 14518 4494 14602 4495
rect 14518 3738 14546 4494
rect 14574 4489 14602 4494
rect 14630 4214 14658 4998
rect 14854 4913 14882 4919
rect 14854 4887 14855 4913
rect 14881 4887 14882 4913
rect 14854 4857 14882 4887
rect 14854 4831 14855 4857
rect 14881 4831 14882 4857
rect 14854 4522 14882 4831
rect 14966 4522 14994 4527
rect 14518 3672 14546 3710
rect 14574 4186 14658 4214
rect 14742 4521 14994 4522
rect 14742 4495 14855 4521
rect 14881 4495 14967 4521
rect 14993 4495 14994 4521
rect 14742 4494 14994 4495
rect 14742 4186 14770 4494
rect 14854 4489 14882 4494
rect 14966 4489 14994 4494
rect 14014 2983 14015 3009
rect 14041 2983 14042 3009
rect 14014 2954 14042 2983
rect 14014 2907 14042 2926
rect 14350 2953 14378 2959
rect 14350 2927 14351 2953
rect 14377 2927 14378 2953
rect 13622 2226 13650 2422
rect 14350 2506 14378 2927
rect 13790 2226 13818 2231
rect 13622 2225 13818 2226
rect 13622 2199 13791 2225
rect 13817 2199 13818 2225
rect 13622 2198 13818 2199
rect 11662 1777 11690 2142
rect 12838 2169 12866 2175
rect 12838 2143 12839 2169
rect 12865 2143 12866 2169
rect 11662 1751 11663 1777
rect 11689 1751 11690 1777
rect 11662 1721 11690 1751
rect 12670 1834 12698 1839
rect 12670 1777 12698 1806
rect 12838 1834 12866 2143
rect 12838 1801 12866 1806
rect 13622 2169 13650 2198
rect 13790 2193 13818 2198
rect 14350 2226 14378 2478
rect 14350 2193 14378 2198
rect 13622 2143 13623 2169
rect 13649 2143 13650 2169
rect 12670 1751 12671 1777
rect 12697 1751 12698 1777
rect 12670 1745 12698 1751
rect 13622 1777 13650 2143
rect 14294 2169 14322 2175
rect 14294 2143 14295 2169
rect 14321 2143 14322 2169
rect 14294 2058 14322 2143
rect 14294 2025 14322 2030
rect 13622 1751 13623 1777
rect 13649 1751 13650 1777
rect 11662 1695 11663 1721
rect 11689 1695 11690 1721
rect 11662 1689 11690 1695
rect 13622 1721 13650 1751
rect 13622 1695 13623 1721
rect 13649 1695 13650 1721
rect 13622 1689 13650 1695
rect 1680 0 1736 400
rect 4984 0 5040 400
rect 8288 0 8344 400
rect 11592 0 11648 400
rect 14574 378 14602 4186
rect 14742 1777 14770 4158
rect 15302 3906 15330 8582
rect 15358 8497 15386 8503
rect 15358 8471 15359 8497
rect 15385 8471 15386 8497
rect 15358 8441 15386 8471
rect 15358 8415 15359 8441
rect 15385 8415 15386 8441
rect 15358 8106 15386 8415
rect 15358 8050 15386 8078
rect 15414 8050 15442 8055
rect 15358 8049 15442 8050
rect 15358 8023 15415 8049
rect 15441 8023 15442 8049
rect 15358 8022 15442 8023
rect 15358 7713 15386 8022
rect 15414 8017 15442 8022
rect 15694 8050 15722 8055
rect 17150 8050 17178 9590
rect 17206 9617 17234 10374
rect 17486 10402 17514 11159
rect 17766 11186 17794 11191
rect 17878 11186 17906 11551
rect 17766 11185 17906 11186
rect 17766 11159 17767 11185
rect 17793 11159 17879 11185
rect 17905 11159 17906 11185
rect 17766 11158 17906 11159
rect 17766 11153 17794 11158
rect 17878 10849 17906 11158
rect 17878 10823 17879 10849
rect 17905 10823 17906 10849
rect 17878 10793 17906 10823
rect 17878 10767 17879 10793
rect 17905 10767 17906 10793
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 17486 10355 17514 10374
rect 17766 10402 17794 10407
rect 17878 10402 17906 10767
rect 17766 10401 17906 10402
rect 17766 10375 17767 10401
rect 17793 10375 17879 10401
rect 17905 10375 17906 10401
rect 17766 10374 17906 10375
rect 17766 10369 17794 10374
rect 17878 10065 17906 10374
rect 17878 10039 17879 10065
rect 17905 10039 17906 10065
rect 17878 10010 17906 10039
rect 17878 10009 18018 10010
rect 17878 9983 17879 10009
rect 17905 9983 18018 10009
rect 17878 9982 18018 9983
rect 17878 9977 17906 9982
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 17206 9591 17207 9617
rect 17233 9591 17234 9617
rect 17206 8833 17234 9591
rect 17766 9618 17794 9623
rect 17878 9618 17906 9623
rect 17766 9617 17906 9618
rect 17766 9591 17767 9617
rect 17793 9591 17879 9617
rect 17905 9591 17906 9617
rect 17766 9590 17906 9591
rect 17766 9562 17794 9590
rect 17766 9529 17794 9534
rect 17878 9281 17906 9590
rect 17878 9255 17879 9281
rect 17905 9255 17906 9281
rect 17878 9225 17906 9255
rect 17878 9199 17879 9225
rect 17905 9199 17906 9225
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 17206 8807 17207 8833
rect 17233 8807 17234 8833
rect 17206 8801 17234 8807
rect 17766 8834 17794 8839
rect 17878 8834 17906 9199
rect 17766 8833 17906 8834
rect 17766 8807 17767 8833
rect 17793 8807 17879 8833
rect 17905 8807 17906 8833
rect 17766 8806 17906 8807
rect 17766 8801 17794 8806
rect 17878 8497 17906 8806
rect 17878 8471 17879 8497
rect 17905 8471 17906 8497
rect 17878 8441 17906 8471
rect 17878 8415 17879 8441
rect 17905 8415 17906 8441
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 17542 8106 17570 8111
rect 17206 8050 17234 8055
rect 17150 8049 17234 8050
rect 17150 8023 17207 8049
rect 17233 8023 17234 8049
rect 17150 8022 17234 8023
rect 15358 7687 15359 7713
rect 15385 7687 15386 7713
rect 15358 7657 15386 7687
rect 15358 7631 15359 7657
rect 15385 7631 15386 7657
rect 15358 6538 15386 7631
rect 15470 7266 15498 7271
rect 15470 7219 15498 7238
rect 15358 6482 15386 6510
rect 15414 6482 15442 6487
rect 15358 6481 15442 6482
rect 15358 6455 15415 6481
rect 15441 6455 15442 6481
rect 15358 6454 15442 6455
rect 15414 6449 15442 6454
rect 15694 6482 15722 8022
rect 15694 6416 15722 6454
rect 15918 7266 15946 7271
rect 15134 3878 15330 3906
rect 15470 5642 15498 5647
rect 15470 5361 15498 5614
rect 15918 5642 15946 7238
rect 16254 7265 16282 7271
rect 16254 7239 16255 7265
rect 16281 7239 16282 7265
rect 16254 7210 16282 7239
rect 16254 7144 16282 7182
rect 17150 7265 17178 7271
rect 17150 7239 17151 7265
rect 17177 7239 17178 7265
rect 17150 6482 17178 7239
rect 17150 6449 17178 6454
rect 17206 6481 17234 8022
rect 17206 6455 17207 6481
rect 17233 6455 17234 6481
rect 17206 6449 17234 6455
rect 15918 5609 15946 5614
rect 15974 5697 16002 5703
rect 15974 5671 15975 5697
rect 16001 5671 16002 5697
rect 15974 5642 16002 5671
rect 15974 5595 16002 5614
rect 16254 5697 16282 5703
rect 16254 5671 16255 5697
rect 16281 5671 16282 5697
rect 16254 5642 16282 5671
rect 16254 5576 16282 5614
rect 17150 5697 17178 5703
rect 17150 5671 17151 5697
rect 17177 5671 17178 5697
rect 15470 5335 15471 5361
rect 15497 5335 15498 5361
rect 15470 5305 15498 5335
rect 15470 5279 15471 5305
rect 15497 5279 15498 5305
rect 15134 3010 15162 3878
rect 15414 3794 15442 3799
rect 15470 3794 15498 5279
rect 15918 4914 15946 4919
rect 15918 4867 15946 4886
rect 17150 4914 17178 5671
rect 17150 4881 17178 4886
rect 17542 4522 17570 8078
rect 17766 8050 17794 8055
rect 17878 8050 17906 8415
rect 17766 8049 17906 8050
rect 17766 8023 17767 8049
rect 17793 8023 17879 8049
rect 17905 8023 17906 8049
rect 17766 8022 17906 8023
rect 17766 8017 17794 8022
rect 17878 7713 17906 8022
rect 17878 7687 17879 7713
rect 17905 7687 17906 7713
rect 17878 7657 17906 7687
rect 17878 7631 17879 7657
rect 17905 7631 17906 7657
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 17878 6929 17906 7631
rect 17878 6903 17879 6929
rect 17905 6903 17906 6929
rect 17878 6873 17906 6903
rect 17878 6847 17879 6873
rect 17905 6847 17906 6873
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17710 4914 17738 4919
rect 17878 4914 17906 6847
rect 17990 6482 18018 9982
rect 18606 9562 18634 29600
rect 18998 26474 19026 26479
rect 18662 25690 18690 25695
rect 18830 25690 18858 25695
rect 18662 25689 18858 25690
rect 18662 25663 18663 25689
rect 18689 25663 18831 25689
rect 18857 25663 18858 25689
rect 18662 25662 18858 25663
rect 18662 25242 18690 25662
rect 18830 25657 18858 25662
rect 18662 25209 18690 25214
rect 18774 25298 18802 25303
rect 18886 25298 18914 25303
rect 18774 25297 18914 25298
rect 18774 25271 18775 25297
rect 18801 25271 18887 25297
rect 18913 25271 18914 25297
rect 18774 25270 18914 25271
rect 18774 24514 18802 25270
rect 18886 25265 18914 25270
rect 18886 24514 18914 24519
rect 18802 24513 18914 24514
rect 18802 24487 18887 24513
rect 18913 24487 18914 24513
rect 18802 24486 18914 24487
rect 18774 24448 18802 24486
rect 18718 23729 18746 23735
rect 18718 23703 18719 23729
rect 18745 23703 18746 23729
rect 18718 23674 18746 23703
rect 18718 23641 18746 23646
rect 18774 22946 18802 22951
rect 18886 22946 18914 24486
rect 18998 24513 19026 26446
rect 19054 25298 19082 25303
rect 19054 25251 19082 25270
rect 18998 24487 18999 24513
rect 19025 24487 19026 24513
rect 18998 23729 19026 24487
rect 18998 23703 18999 23729
rect 19025 23703 19026 23729
rect 18942 23674 18970 23679
rect 18942 23627 18970 23646
rect 18998 23506 19026 23703
rect 18998 23473 19026 23478
rect 18774 22945 18914 22946
rect 18774 22919 18775 22945
rect 18801 22919 18887 22945
rect 18913 22919 18914 22945
rect 18774 22918 18914 22919
rect 18774 22913 18802 22918
rect 18886 22913 18914 22918
rect 19054 22889 19082 22895
rect 19054 22863 19055 22889
rect 19081 22863 19082 22889
rect 18718 22554 18746 22559
rect 18830 22554 18858 22559
rect 18718 22553 18858 22554
rect 18718 22527 18719 22553
rect 18745 22527 18831 22553
rect 18857 22527 18858 22553
rect 18718 22526 18858 22527
rect 18718 22521 18746 22526
rect 18774 22106 18802 22111
rect 18830 22106 18858 22526
rect 18886 22161 18914 22167
rect 18886 22135 18887 22161
rect 18913 22135 18914 22161
rect 18886 22106 18914 22135
rect 18774 22105 18914 22106
rect 18774 22079 18775 22105
rect 18801 22079 18914 22105
rect 18774 22078 18914 22079
rect 19054 22105 19082 22863
rect 19054 22079 19055 22105
rect 19081 22079 19082 22105
rect 18718 21770 18746 21775
rect 18774 21770 18802 22078
rect 19054 21882 19082 22079
rect 19054 21849 19082 21854
rect 18830 21770 18858 21775
rect 18746 21769 18858 21770
rect 18746 21743 18831 21769
rect 18857 21743 18858 21769
rect 18746 21742 18858 21743
rect 18718 20986 18746 21742
rect 18830 21737 18858 21742
rect 18886 21377 18914 21383
rect 18886 21351 18887 21377
rect 18913 21351 18914 21377
rect 18774 21322 18802 21327
rect 18886 21322 18914 21351
rect 18802 21294 18914 21322
rect 18998 21377 19026 21383
rect 18998 21351 18999 21377
rect 19025 21351 19026 21377
rect 18774 21275 18802 21294
rect 18774 20986 18802 20991
rect 18718 20985 18802 20986
rect 18718 20959 18775 20985
rect 18801 20959 18802 20985
rect 18718 20958 18802 20959
rect 18774 20594 18802 20958
rect 18774 20538 18802 20566
rect 18886 20985 18914 20991
rect 18886 20959 18887 20985
rect 18913 20959 18914 20985
rect 18886 20538 18914 20959
rect 18998 20986 19026 21351
rect 18998 20593 19026 20958
rect 18998 20567 18999 20593
rect 19025 20567 19026 20593
rect 18942 20538 18970 20543
rect 18774 20537 18970 20538
rect 18774 20511 18775 20537
rect 18801 20511 18943 20537
rect 18969 20511 18970 20537
rect 18774 20510 18970 20511
rect 18774 20505 18802 20510
rect 18718 20202 18746 20207
rect 18886 20202 18914 20207
rect 18718 20201 18914 20202
rect 18718 20175 18719 20201
rect 18745 20175 18887 20201
rect 18913 20175 18914 20201
rect 18718 20174 18914 20175
rect 18718 19810 18746 20174
rect 18886 20169 18914 20174
rect 18718 19362 18746 19782
rect 18774 19753 18802 19759
rect 18774 19727 18775 19753
rect 18801 19727 18802 19753
rect 18774 19474 18802 19727
rect 18942 19753 18970 20510
rect 18942 19727 18943 19753
rect 18969 19727 18970 19753
rect 18942 19474 18970 19727
rect 18998 19586 19026 20567
rect 18998 19553 19026 19558
rect 19054 20201 19082 20207
rect 19054 20175 19055 20201
rect 19081 20175 19082 20201
rect 19054 19754 19082 20175
rect 18774 19473 18970 19474
rect 18774 19447 18775 19473
rect 18801 19447 18970 19473
rect 18774 19446 18970 19447
rect 18774 19441 18802 19446
rect 18942 19417 18970 19446
rect 18942 19391 18943 19417
rect 18969 19391 18970 19417
rect 18718 19334 18858 19362
rect 18774 18634 18802 18639
rect 18606 9529 18634 9534
rect 18718 18633 18802 18634
rect 18718 18607 18775 18633
rect 18801 18607 18802 18633
rect 18718 18606 18802 18607
rect 18718 10346 18746 18606
rect 18774 18601 18802 18606
rect 18774 17066 18802 17071
rect 18830 17066 18858 19334
rect 18886 17066 18914 17071
rect 18774 17065 18914 17066
rect 18774 17039 18775 17065
rect 18801 17039 18887 17065
rect 18913 17039 18914 17065
rect 18774 17038 18914 17039
rect 18774 17033 18802 17038
rect 18886 17033 18914 17038
rect 18774 16674 18802 16679
rect 18886 16674 18914 16679
rect 18942 16674 18970 19391
rect 19054 19417 19082 19726
rect 19054 19391 19055 19417
rect 19081 19391 19082 19417
rect 19054 17290 19082 19391
rect 19054 17257 19082 17262
rect 18774 16673 18970 16674
rect 18774 16647 18775 16673
rect 18801 16647 18887 16673
rect 18913 16647 18970 16673
rect 18774 16646 18970 16647
rect 19054 17065 19082 17071
rect 19054 17039 19055 17065
rect 19081 17039 19082 17065
rect 18774 16641 18802 16646
rect 18886 16641 18914 16646
rect 19054 16617 19082 17039
rect 19054 16591 19055 16617
rect 19081 16591 19082 16617
rect 19054 14994 19082 16591
rect 19054 14961 19082 14966
rect 19054 13145 19082 13151
rect 19054 13119 19055 13145
rect 19081 13119 19082 13145
rect 19054 12698 19082 13119
rect 19054 12361 19082 12670
rect 19054 12335 19055 12361
rect 19081 12335 19082 12361
rect 19054 11577 19082 12335
rect 19054 11551 19055 11577
rect 19081 11551 19082 11577
rect 19054 10794 19082 11551
rect 18718 7658 18746 10318
rect 18774 10793 19082 10794
rect 18774 10767 19055 10793
rect 19081 10767 19082 10793
rect 18774 10766 19082 10767
rect 18774 10402 18802 10766
rect 19054 10761 19082 10766
rect 18774 10009 18802 10374
rect 18774 9983 18775 10009
rect 18801 9983 18802 10009
rect 18774 9225 18802 9983
rect 18774 9199 18775 9225
rect 18801 9199 18802 9225
rect 18774 8441 18802 9199
rect 18774 8415 18775 8441
rect 18801 8415 18802 8441
rect 18774 8409 18802 8415
rect 18774 7658 18802 7663
rect 18718 7657 18802 7658
rect 18718 7631 18775 7657
rect 18801 7631 18802 7657
rect 18718 7630 18802 7631
rect 18774 6873 18802 7630
rect 18774 6847 18775 6873
rect 18801 6847 18802 6873
rect 17990 6481 18186 6482
rect 17990 6455 17991 6481
rect 18017 6455 18186 6481
rect 17990 6454 18186 6455
rect 17990 6449 18018 6454
rect 18102 6145 18130 6454
rect 18158 6425 18186 6454
rect 18158 6399 18159 6425
rect 18185 6399 18186 6425
rect 18158 6393 18186 6399
rect 18102 6119 18103 6145
rect 18129 6119 18130 6145
rect 18102 6089 18130 6119
rect 18102 6063 18103 6089
rect 18129 6063 18130 6089
rect 18102 5361 18130 6063
rect 18102 5335 18103 5361
rect 18129 5335 18130 5361
rect 18102 5306 18130 5335
rect 18774 6089 18802 6847
rect 18774 6063 18775 6089
rect 18801 6063 18802 6089
rect 18102 5305 18466 5306
rect 18102 5279 18103 5305
rect 18129 5279 18466 5305
rect 18102 5278 18466 5279
rect 18102 5273 18130 5278
rect 17934 4914 17962 4919
rect 17710 4913 17962 4914
rect 17710 4887 17711 4913
rect 17737 4887 17935 4913
rect 17961 4887 17962 4913
rect 17710 4886 17962 4887
rect 17710 4881 17738 4886
rect 17934 4578 17962 4886
rect 18382 4913 18410 4919
rect 18382 4887 18383 4913
rect 18409 4887 18410 4913
rect 17990 4578 18018 4583
rect 17934 4577 18018 4578
rect 17934 4551 17991 4577
rect 18017 4551 18018 4577
rect 17934 4550 18018 4551
rect 17542 4489 17570 4494
rect 17990 4521 18018 4550
rect 17990 4495 17991 4521
rect 18017 4495 18018 4521
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 16478 4242 16506 4247
rect 15414 3793 15498 3794
rect 15414 3767 15415 3793
rect 15441 3767 15498 3793
rect 15414 3766 15498 3767
rect 16254 4130 16282 4135
rect 16478 4130 16506 4214
rect 17990 4242 18018 4495
rect 16254 4129 16506 4130
rect 16254 4103 16255 4129
rect 16281 4103 16479 4129
rect 16505 4103 16506 4129
rect 16254 4102 16506 4103
rect 15358 3738 15386 3743
rect 15414 3738 15442 3766
rect 15358 3737 15442 3738
rect 15358 3711 15359 3737
rect 15385 3711 15442 3737
rect 15358 3710 15442 3711
rect 15246 3010 15274 3015
rect 15134 3009 15274 3010
rect 15134 2983 15247 3009
rect 15273 2983 15274 3009
rect 15134 2982 15274 2983
rect 15134 2953 15162 2982
rect 15246 2977 15274 2982
rect 15134 2927 15135 2953
rect 15161 2927 15162 2953
rect 15134 2921 15162 2927
rect 15358 2954 15386 3710
rect 16254 3346 16282 4102
rect 16478 4097 16506 4102
rect 16758 4129 16786 4135
rect 16758 4103 16759 4129
rect 16785 4103 16786 4129
rect 16758 3458 16786 4103
rect 17710 4130 17738 4135
rect 17878 4130 17906 4135
rect 17710 4129 17878 4130
rect 17710 4103 17711 4129
rect 17737 4103 17878 4129
rect 17710 4102 17878 4103
rect 17710 4097 17738 4102
rect 17878 3793 17906 4102
rect 17878 3767 17879 3793
rect 17905 3767 17906 3793
rect 17878 3737 17906 3767
rect 17878 3711 17879 3737
rect 17905 3711 17906 3737
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 16758 3425 16786 3430
rect 17486 3458 17514 3463
rect 16366 3346 16394 3351
rect 16254 3345 16394 3346
rect 16254 3319 16255 3345
rect 16281 3319 16367 3345
rect 16393 3319 16394 3345
rect 16254 3318 16394 3319
rect 16254 3313 16282 3318
rect 16366 3313 16394 3318
rect 16926 3345 16954 3351
rect 16926 3319 16927 3345
rect 16953 3319 16954 3345
rect 14798 2561 14826 2567
rect 14798 2535 14799 2561
rect 14825 2535 14826 2561
rect 14798 2506 14826 2535
rect 14798 2473 14826 2478
rect 15246 2561 15274 2567
rect 15246 2535 15247 2561
rect 15273 2535 15274 2561
rect 15246 2450 15274 2535
rect 15246 2417 15274 2422
rect 15246 2226 15274 2231
rect 15358 2226 15386 2926
rect 15470 2561 15498 2567
rect 15470 2535 15471 2561
rect 15497 2535 15498 2561
rect 15470 2450 15498 2535
rect 16926 2562 16954 3319
rect 16926 2529 16954 2534
rect 17486 2561 17514 3430
rect 17710 3346 17738 3351
rect 17822 3346 17850 3351
rect 17878 3346 17906 3711
rect 17710 3345 17906 3346
rect 17710 3319 17711 3345
rect 17737 3319 17823 3345
rect 17849 3319 17906 3345
rect 17710 3318 17906 3319
rect 17710 3313 17738 3318
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17486 2535 17487 2561
rect 17513 2535 17514 2561
rect 17486 2529 17514 2535
rect 17766 2562 17794 2567
rect 17822 2562 17850 3318
rect 17990 3009 18018 4214
rect 18382 4522 18410 4887
rect 18382 4129 18410 4494
rect 18382 4103 18383 4129
rect 18409 4103 18410 4129
rect 18382 4097 18410 4103
rect 18438 4130 18466 5278
rect 18774 5305 18802 6063
rect 18774 5279 18775 5305
rect 18801 5279 18802 5305
rect 18774 5273 18802 5279
rect 18774 4522 18802 4527
rect 18774 4214 18802 4494
rect 18774 4186 18858 4214
rect 18438 4097 18466 4102
rect 17990 2983 17991 3009
rect 18017 2983 18018 3009
rect 17990 2953 18018 2983
rect 17990 2927 17991 2953
rect 18017 2927 18018 2953
rect 17990 2921 18018 2927
rect 18214 4074 18242 4079
rect 17878 2562 17906 2567
rect 17766 2561 17906 2562
rect 17766 2535 17767 2561
rect 17793 2535 17879 2561
rect 17905 2535 17906 2561
rect 17766 2534 17906 2535
rect 17766 2529 17794 2534
rect 15470 2417 15498 2422
rect 15246 2225 15386 2226
rect 15246 2199 15247 2225
rect 15273 2199 15386 2225
rect 15246 2198 15386 2199
rect 17878 2225 17906 2534
rect 17878 2199 17879 2225
rect 17905 2199 17906 2225
rect 15246 2169 15274 2198
rect 15246 2143 15247 2169
rect 15273 2143 15274 2169
rect 15246 2137 15274 2143
rect 17878 2169 17906 2199
rect 17878 2143 17879 2169
rect 17905 2143 17906 2169
rect 17878 2137 17906 2143
rect 14742 1751 14743 1777
rect 14769 1751 14770 1777
rect 14742 1721 14770 1751
rect 15526 2058 15554 2063
rect 15526 1777 15554 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 15526 1751 15527 1777
rect 15553 1751 15554 1777
rect 15526 1745 15554 1751
rect 14742 1695 14743 1721
rect 14769 1695 14770 1721
rect 14742 1689 14770 1695
rect 14742 462 14938 490
rect 14742 378 14770 462
rect 14910 400 14938 462
rect 18214 400 18242 4046
rect 18830 3737 18858 4186
rect 18830 3711 18831 3737
rect 18857 3711 18858 3737
rect 18830 3705 18858 3711
rect 18382 3346 18410 3351
rect 18382 3299 18410 3318
rect 18774 3346 18802 3351
rect 18774 2953 18802 3318
rect 18774 2927 18775 2953
rect 18801 2927 18802 2953
rect 18774 2921 18802 2927
rect 18774 2562 18802 2567
rect 18774 2169 18802 2534
rect 18774 2143 18775 2169
rect 18801 2143 18802 2169
rect 18774 1218 18802 2143
rect 18774 1185 18802 1190
rect 14574 350 14770 378
rect 14896 0 14952 400
rect 18200 0 18256 400
<< via2 >>
rect 1358 26894 1386 26922
rect 1750 27902 1778 27930
rect 1694 25214 1722 25242
rect 1582 23729 1610 23730
rect 1582 23703 1583 23729
rect 1583 23703 1609 23729
rect 1609 23703 1610 23729
rect 1582 23702 1610 23703
rect 1582 17654 1610 17682
rect 2238 27845 2266 27846
rect 2238 27819 2239 27845
rect 2239 27819 2265 27845
rect 2265 27819 2266 27845
rect 2238 27818 2266 27819
rect 2290 27845 2318 27846
rect 2290 27819 2291 27845
rect 2291 27819 2317 27845
rect 2317 27819 2318 27845
rect 2290 27818 2318 27819
rect 2342 27845 2370 27846
rect 2342 27819 2343 27845
rect 2343 27819 2369 27845
rect 2369 27819 2370 27845
rect 2342 27818 2370 27819
rect 2238 27061 2266 27062
rect 2238 27035 2239 27061
rect 2239 27035 2265 27061
rect 2265 27035 2266 27061
rect 2238 27034 2266 27035
rect 2290 27061 2318 27062
rect 2290 27035 2291 27061
rect 2291 27035 2317 27061
rect 2317 27035 2318 27061
rect 2290 27034 2318 27035
rect 2342 27061 2370 27062
rect 2342 27035 2343 27061
rect 2343 27035 2369 27061
rect 2369 27035 2370 27061
rect 2342 27034 2370 27035
rect 2086 26894 2114 26922
rect 3822 26865 3850 26866
rect 3822 26839 3823 26865
rect 3823 26839 3849 26865
rect 3849 26839 3850 26865
rect 3822 26838 3850 26839
rect 4494 26865 4522 26866
rect 4494 26839 4495 26865
rect 4495 26839 4521 26865
rect 4521 26839 4522 26865
rect 4494 26838 4522 26839
rect 4494 26473 4522 26474
rect 4494 26447 4495 26473
rect 4495 26447 4521 26473
rect 4521 26447 4522 26473
rect 4494 26446 4522 26447
rect 2814 26390 2842 26418
rect 2238 26277 2266 26278
rect 2238 26251 2239 26277
rect 2239 26251 2265 26277
rect 2265 26251 2266 26277
rect 2238 26250 2266 26251
rect 2290 26277 2318 26278
rect 2290 26251 2291 26277
rect 2291 26251 2317 26277
rect 2317 26251 2318 26277
rect 2290 26250 2318 26251
rect 2342 26277 2370 26278
rect 2342 26251 2343 26277
rect 2343 26251 2369 26277
rect 2369 26251 2370 26277
rect 2342 26250 2370 26251
rect 2238 25493 2266 25494
rect 2238 25467 2239 25493
rect 2239 25467 2265 25493
rect 2265 25467 2266 25493
rect 2238 25466 2266 25467
rect 2290 25493 2318 25494
rect 2290 25467 2291 25493
rect 2291 25467 2317 25493
rect 2317 25467 2318 25493
rect 2290 25466 2318 25467
rect 2342 25493 2370 25494
rect 2342 25467 2343 25493
rect 2343 25467 2369 25493
rect 2369 25467 2370 25493
rect 2342 25466 2370 25467
rect 2478 25297 2506 25298
rect 2478 25271 2479 25297
rect 2479 25271 2505 25297
rect 2505 25271 2506 25297
rect 2478 25270 2506 25271
rect 2814 25270 2842 25298
rect 3318 26054 3346 26082
rect 3094 25214 3122 25242
rect 2238 24709 2266 24710
rect 2238 24683 2239 24709
rect 2239 24683 2265 24709
rect 2265 24683 2266 24709
rect 2238 24682 2266 24683
rect 2290 24709 2318 24710
rect 2290 24683 2291 24709
rect 2291 24683 2317 24709
rect 2317 24683 2318 24709
rect 2290 24682 2318 24683
rect 2342 24709 2370 24710
rect 2342 24683 2343 24709
rect 2343 24683 2369 24709
rect 2369 24683 2370 24709
rect 2342 24682 2370 24683
rect 1918 24206 1946 24234
rect 1806 23702 1834 23730
rect 2534 24121 2562 24122
rect 2534 24095 2535 24121
rect 2535 24095 2561 24121
rect 2561 24095 2562 24121
rect 2534 24094 2562 24095
rect 2238 23925 2266 23926
rect 2238 23899 2239 23925
rect 2239 23899 2265 23925
rect 2265 23899 2266 23925
rect 2238 23898 2266 23899
rect 2290 23925 2318 23926
rect 2290 23899 2291 23925
rect 2291 23899 2317 23925
rect 2317 23899 2318 23925
rect 2290 23898 2318 23899
rect 2342 23925 2370 23926
rect 2342 23899 2343 23925
rect 2343 23899 2369 23925
rect 2369 23899 2370 23925
rect 2342 23898 2370 23899
rect 1918 23702 1946 23730
rect 3150 23729 3178 23730
rect 3150 23703 3151 23729
rect 3151 23703 3177 23729
rect 3177 23703 3178 23729
rect 3150 23702 3178 23703
rect 3318 23702 3346 23730
rect 3542 24094 3570 24122
rect 4830 26081 4858 26082
rect 4830 26055 4831 26081
rect 4831 26055 4857 26081
rect 4857 26055 4858 26081
rect 4830 26054 4858 26055
rect 5166 26054 5194 26082
rect 5726 26473 5754 26474
rect 5726 26447 5727 26473
rect 5727 26447 5753 26473
rect 5753 26447 5754 26473
rect 5726 26446 5754 26447
rect 5726 24934 5754 24962
rect 6286 25214 6314 25242
rect 5166 24878 5194 24906
rect 3766 24121 3794 24122
rect 3766 24095 3767 24121
rect 3767 24095 3793 24121
rect 3793 24095 3794 24121
rect 3766 24094 3794 24095
rect 3990 24121 4018 24122
rect 3990 24095 3991 24121
rect 3991 24095 4017 24121
rect 4017 24095 4018 24121
rect 3990 24094 4018 24095
rect 6622 24905 6650 24906
rect 6622 24879 6623 24905
rect 6623 24879 6649 24905
rect 6649 24879 6650 24905
rect 6622 24878 6650 24879
rect 6622 24374 6650 24402
rect 7126 24486 7154 24514
rect 7518 24961 7546 24962
rect 7518 24935 7519 24961
rect 7519 24935 7545 24961
rect 7545 24935 7546 24961
rect 7518 24934 7546 24935
rect 7518 24430 7546 24458
rect 7966 24457 7994 24458
rect 7966 24431 7967 24457
rect 7967 24431 7993 24457
rect 7993 24431 7994 24457
rect 7966 24430 7994 24431
rect 7070 24374 7098 24402
rect 5838 24177 5866 24178
rect 5838 24151 5839 24177
rect 5839 24151 5865 24177
rect 5865 24151 5866 24177
rect 5838 24150 5866 24151
rect 4886 24094 4914 24122
rect 3822 23646 3850 23674
rect 5166 24121 5194 24122
rect 5166 24095 5167 24121
rect 5167 24095 5193 24121
rect 5193 24095 5194 24121
rect 5166 24094 5194 24095
rect 4886 23729 4914 23730
rect 4886 23703 4887 23729
rect 4887 23703 4913 23729
rect 4913 23703 4914 23729
rect 4886 23702 4914 23703
rect 6062 24094 6090 24122
rect 5782 23673 5810 23674
rect 5782 23647 5783 23673
rect 5783 23647 5809 23673
rect 5809 23647 5810 23673
rect 5782 23646 5810 23647
rect 2238 23141 2266 23142
rect 2238 23115 2239 23141
rect 2239 23115 2265 23141
rect 2265 23115 2266 23141
rect 2238 23114 2266 23115
rect 2290 23141 2318 23142
rect 2290 23115 2291 23141
rect 2291 23115 2317 23141
rect 2317 23115 2318 23141
rect 2290 23114 2318 23115
rect 2342 23141 2370 23142
rect 2342 23115 2343 23141
rect 2343 23115 2369 23141
rect 2369 23115 2370 23141
rect 2342 23114 2370 23115
rect 2238 22357 2266 22358
rect 2238 22331 2239 22357
rect 2239 22331 2265 22357
rect 2265 22331 2266 22357
rect 2238 22330 2266 22331
rect 2290 22357 2318 22358
rect 2290 22331 2291 22357
rect 2291 22331 2317 22357
rect 2317 22331 2318 22357
rect 2290 22330 2318 22331
rect 2342 22357 2370 22358
rect 2342 22331 2343 22357
rect 2343 22331 2369 22357
rect 2369 22331 2370 22357
rect 2342 22330 2370 22331
rect 1806 20510 1834 20538
rect 2254 21742 2282 21770
rect 3038 21769 3066 21770
rect 3038 21743 3039 21769
rect 3039 21743 3065 21769
rect 3065 21743 3066 21769
rect 3038 21742 3066 21743
rect 2238 21573 2266 21574
rect 2238 21547 2239 21573
rect 2239 21547 2265 21573
rect 2265 21547 2266 21573
rect 2238 21546 2266 21547
rect 2290 21573 2318 21574
rect 2290 21547 2291 21573
rect 2291 21547 2317 21573
rect 2317 21547 2318 21573
rect 2290 21546 2318 21547
rect 2342 21573 2370 21574
rect 2342 21547 2343 21573
rect 2343 21547 2369 21573
rect 2369 21547 2370 21573
rect 2342 21546 2370 21547
rect 2478 21321 2506 21322
rect 2478 21295 2479 21321
rect 2479 21295 2505 21321
rect 2505 21295 2506 21321
rect 2478 21294 2506 21295
rect 2238 20789 2266 20790
rect 2238 20763 2239 20789
rect 2239 20763 2265 20789
rect 2265 20763 2266 20789
rect 2238 20762 2266 20763
rect 2290 20789 2318 20790
rect 2290 20763 2291 20789
rect 2291 20763 2317 20789
rect 2317 20763 2318 20789
rect 2290 20762 2318 20763
rect 2342 20789 2370 20790
rect 2342 20763 2343 20789
rect 2343 20763 2369 20789
rect 2369 20763 2370 20789
rect 2342 20762 2370 20763
rect 3038 21294 3066 21322
rect 6342 24121 6370 24122
rect 6342 24095 6343 24121
rect 6343 24095 6369 24121
rect 6369 24095 6370 24121
rect 6342 24094 6370 24095
rect 7518 24121 7546 24122
rect 7518 24095 7519 24121
rect 7519 24095 7545 24121
rect 7545 24095 7546 24121
rect 7518 24094 7546 24095
rect 8582 24513 8610 24514
rect 8582 24487 8583 24513
rect 8583 24487 8609 24513
rect 8609 24487 8610 24513
rect 8582 24486 8610 24487
rect 8358 24430 8386 24458
rect 9918 28237 9946 28238
rect 9918 28211 9919 28237
rect 9919 28211 9945 28237
rect 9945 28211 9946 28237
rect 9918 28210 9946 28211
rect 9970 28237 9998 28238
rect 9970 28211 9971 28237
rect 9971 28211 9997 28237
rect 9997 28211 9998 28237
rect 9970 28210 9998 28211
rect 10022 28237 10050 28238
rect 10022 28211 10023 28237
rect 10023 28211 10049 28237
rect 10049 28211 10050 28237
rect 10022 28210 10050 28211
rect 9918 27453 9946 27454
rect 9918 27427 9919 27453
rect 9919 27427 9945 27453
rect 9945 27427 9946 27453
rect 9918 27426 9946 27427
rect 9970 27453 9998 27454
rect 9970 27427 9971 27453
rect 9971 27427 9997 27453
rect 9997 27427 9998 27453
rect 9970 27426 9998 27427
rect 10022 27453 10050 27454
rect 10022 27427 10023 27453
rect 10023 27427 10049 27453
rect 10049 27427 10050 27453
rect 10022 27426 10050 27427
rect 9918 26669 9946 26670
rect 9918 26643 9919 26669
rect 9919 26643 9945 26669
rect 9945 26643 9946 26669
rect 9918 26642 9946 26643
rect 9970 26669 9998 26670
rect 9970 26643 9971 26669
rect 9971 26643 9997 26669
rect 9997 26643 9998 26669
rect 9970 26642 9998 26643
rect 10022 26669 10050 26670
rect 10022 26643 10023 26669
rect 10023 26643 10049 26669
rect 10049 26643 10050 26669
rect 10022 26642 10050 26643
rect 9918 25885 9946 25886
rect 9918 25859 9919 25885
rect 9919 25859 9945 25885
rect 9945 25859 9946 25885
rect 9918 25858 9946 25859
rect 9970 25885 9998 25886
rect 9970 25859 9971 25885
rect 9971 25859 9997 25885
rect 9997 25859 9998 25885
rect 9970 25858 9998 25859
rect 10022 25885 10050 25886
rect 10022 25859 10023 25885
rect 10023 25859 10049 25885
rect 10049 25859 10050 25885
rect 10022 25858 10050 25859
rect 9918 25101 9946 25102
rect 9918 25075 9919 25101
rect 9919 25075 9945 25101
rect 9945 25075 9946 25101
rect 9918 25074 9946 25075
rect 9970 25101 9998 25102
rect 9970 25075 9971 25101
rect 9971 25075 9997 25101
rect 9997 25075 9998 25101
rect 9970 25074 9998 25075
rect 10022 25101 10050 25102
rect 10022 25075 10023 25101
rect 10023 25075 10049 25101
rect 10049 25075 10050 25101
rect 10022 25074 10050 25075
rect 8750 24430 8778 24458
rect 9142 24486 9170 24514
rect 8022 24094 8050 24122
rect 2238 20005 2266 20006
rect 2238 19979 2239 20005
rect 2239 19979 2265 20005
rect 2265 19979 2266 20005
rect 2238 19978 2266 19979
rect 2290 20005 2318 20006
rect 2290 19979 2291 20005
rect 2291 19979 2317 20005
rect 2317 19979 2318 20005
rect 2290 19978 2318 19979
rect 2342 20005 2370 20006
rect 2342 19979 2343 20005
rect 2343 19979 2369 20005
rect 2369 19979 2370 20005
rect 2342 19978 2370 19979
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2478 18241 2506 18242
rect 2478 18215 2479 18241
rect 2479 18215 2505 18241
rect 2505 18215 2506 18241
rect 2478 18214 2506 18215
rect 3038 18214 3066 18242
rect 1862 17878 1890 17906
rect 3038 17849 3066 17850
rect 3038 17823 3039 17849
rect 3039 17823 3065 17849
rect 3065 17823 3066 17849
rect 3038 17822 3066 17823
rect 4214 21769 4242 21770
rect 4214 21743 4215 21769
rect 4215 21743 4241 21769
rect 4241 21743 4242 21769
rect 4214 21742 4242 21743
rect 8414 23702 8442 23730
rect 8582 24374 8610 24402
rect 9918 24317 9946 24318
rect 9918 24291 9919 24317
rect 9919 24291 9945 24317
rect 9945 24291 9946 24317
rect 9918 24290 9946 24291
rect 9970 24317 9998 24318
rect 9970 24291 9971 24317
rect 9971 24291 9997 24317
rect 9997 24291 9998 24317
rect 9970 24290 9998 24291
rect 10022 24317 10050 24318
rect 10022 24291 10023 24317
rect 10023 24291 10049 24317
rect 10049 24291 10050 24317
rect 10022 24290 10050 24291
rect 8582 23254 8610 23282
rect 9142 23310 9170 23338
rect 9422 23729 9450 23730
rect 9422 23703 9423 23729
rect 9423 23703 9449 23729
rect 9449 23703 9450 23729
rect 9422 23702 9450 23703
rect 9086 23254 9114 23282
rect 6062 21014 6090 21042
rect 7126 21014 7154 21042
rect 8022 22526 8050 22554
rect 8358 22553 8386 22554
rect 8358 22527 8359 22553
rect 8359 22527 8385 22553
rect 8385 22527 8386 22553
rect 8358 22526 8386 22527
rect 7518 21014 7546 21042
rect 3822 19025 3850 19026
rect 3822 18999 3823 19025
rect 3823 18999 3849 19025
rect 3849 18999 3850 19025
rect 3822 18998 3850 18999
rect 5278 19025 5306 19026
rect 5278 18999 5279 19025
rect 5279 18999 5305 19025
rect 5305 18999 5306 19025
rect 5278 18998 5306 18999
rect 8582 21014 8610 21042
rect 3374 17878 3402 17906
rect 4438 17849 4466 17850
rect 4438 17823 4439 17849
rect 4439 17823 4465 17849
rect 4465 17823 4466 17849
rect 4438 17822 4466 17823
rect 1862 17654 1890 17682
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2086 16814 2114 16842
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 1694 13118 1722 13146
rect 910 9422 938 9450
rect 1582 9254 1610 9282
rect 1582 8049 1610 8050
rect 1582 8023 1583 8049
rect 1583 8023 1609 8049
rect 1609 8023 1610 8049
rect 1582 8022 1610 8023
rect 1582 7265 1610 7266
rect 1582 7239 1583 7265
rect 1583 7239 1609 7265
rect 1609 7239 1610 7265
rect 1582 7238 1610 7239
rect 1862 11577 1890 11578
rect 1862 11551 1863 11577
rect 1863 11551 1889 11577
rect 1889 11551 1890 11577
rect 1862 11550 1890 11551
rect 1918 9254 1946 9282
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2534 14294 2562 14322
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2534 12361 2562 12362
rect 2534 12335 2535 12361
rect 2535 12335 2561 12361
rect 2561 12335 2562 12361
rect 2534 12334 2562 12335
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2086 8470 2114 8498
rect 1918 8022 1946 8050
rect 1918 7630 1946 7658
rect 2478 8414 2506 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2142 7657 2170 7658
rect 2142 7631 2143 7657
rect 2143 7631 2169 7657
rect 2169 7631 2170 7657
rect 2142 7630 2170 7631
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 2086 7238 2114 7266
rect 8582 19809 8610 19810
rect 8582 19783 8583 19809
rect 8583 19783 8609 19809
rect 8609 19783 8610 19809
rect 8582 19782 8610 19783
rect 6398 17849 6426 17850
rect 6398 17823 6399 17849
rect 6399 17823 6425 17849
rect 6425 17823 6426 17849
rect 6398 17822 6426 17823
rect 7574 18241 7602 18242
rect 7574 18215 7575 18241
rect 7575 18215 7601 18241
rect 7601 18215 7602 18241
rect 7574 18214 7602 18215
rect 7182 17849 7210 17850
rect 7182 17823 7183 17849
rect 7183 17823 7209 17849
rect 7209 17823 7210 17849
rect 7182 17822 7210 17823
rect 9142 19782 9170 19810
rect 9142 19417 9170 19418
rect 9142 19391 9143 19417
rect 9143 19391 9169 19417
rect 9169 19391 9170 19417
rect 9142 19390 9170 19391
rect 9478 22526 9506 22554
rect 9478 22161 9506 22162
rect 9478 22135 9479 22161
rect 9479 22135 9505 22161
rect 9505 22135 9506 22161
rect 9478 22134 9506 22135
rect 9918 23533 9946 23534
rect 9918 23507 9919 23533
rect 9919 23507 9945 23533
rect 9945 23507 9946 23533
rect 9918 23506 9946 23507
rect 9970 23533 9998 23534
rect 9970 23507 9971 23533
rect 9971 23507 9997 23533
rect 9997 23507 9998 23533
rect 9970 23506 9998 23507
rect 10022 23533 10050 23534
rect 10022 23507 10023 23533
rect 10023 23507 10049 23533
rect 10049 23507 10050 23533
rect 10022 23506 10050 23507
rect 10598 23337 10626 23338
rect 10598 23311 10599 23337
rect 10599 23311 10625 23337
rect 10625 23311 10626 23337
rect 10598 23310 10626 23311
rect 10374 23254 10402 23282
rect 9918 22749 9946 22750
rect 9918 22723 9919 22749
rect 9919 22723 9945 22749
rect 9945 22723 9946 22749
rect 9918 22722 9946 22723
rect 9970 22749 9998 22750
rect 9970 22723 9971 22749
rect 9971 22723 9997 22749
rect 9997 22723 9998 22749
rect 9970 22722 9998 22723
rect 10022 22749 10050 22750
rect 10022 22723 10023 22749
rect 10023 22723 10049 22749
rect 10049 22723 10050 22749
rect 10022 22722 10050 22723
rect 9814 22134 9842 22162
rect 10598 22918 10626 22946
rect 9918 21965 9946 21966
rect 9918 21939 9919 21965
rect 9919 21939 9945 21965
rect 9945 21939 9946 21965
rect 9918 21938 9946 21939
rect 9970 21965 9998 21966
rect 9970 21939 9971 21965
rect 9971 21939 9997 21965
rect 9997 21939 9998 21965
rect 9970 21938 9998 21939
rect 10022 21965 10050 21966
rect 10022 21939 10023 21965
rect 10023 21939 10049 21965
rect 10049 21939 10050 21965
rect 10022 21938 10050 21939
rect 9814 21854 9842 21882
rect 10038 21854 10066 21882
rect 10374 21742 10402 21770
rect 10598 21769 10626 21770
rect 10598 21743 10599 21769
rect 10599 21743 10625 21769
rect 10625 21743 10626 21769
rect 10598 21742 10626 21743
rect 9918 21181 9946 21182
rect 9918 21155 9919 21181
rect 9919 21155 9945 21181
rect 9945 21155 9946 21181
rect 9918 21154 9946 21155
rect 9970 21181 9998 21182
rect 9970 21155 9971 21181
rect 9971 21155 9997 21181
rect 9997 21155 9998 21181
rect 9970 21154 9998 21155
rect 10022 21181 10050 21182
rect 10022 21155 10023 21181
rect 10023 21155 10049 21181
rect 10049 21155 10050 21181
rect 10022 21154 10050 21155
rect 9534 21014 9562 21042
rect 9918 20397 9946 20398
rect 9918 20371 9919 20397
rect 9919 20371 9945 20397
rect 9945 20371 9946 20397
rect 9918 20370 9946 20371
rect 9970 20397 9998 20398
rect 9970 20371 9971 20397
rect 9971 20371 9997 20397
rect 9997 20371 9998 20397
rect 9970 20370 9998 20371
rect 10022 20397 10050 20398
rect 10022 20371 10023 20397
rect 10023 20371 10049 20397
rect 10049 20371 10050 20397
rect 10022 20370 10050 20371
rect 9918 19613 9946 19614
rect 9918 19587 9919 19613
rect 9919 19587 9945 19613
rect 9945 19587 9946 19613
rect 9918 19586 9946 19587
rect 9970 19613 9998 19614
rect 9970 19587 9971 19613
rect 9971 19587 9997 19613
rect 9997 19587 9998 19613
rect 9970 19586 9998 19587
rect 10022 19613 10050 19614
rect 10022 19587 10023 19613
rect 10023 19587 10049 19613
rect 10049 19587 10050 19613
rect 10022 19586 10050 19587
rect 8750 18241 8778 18242
rect 8750 18215 8751 18241
rect 8751 18215 8777 18241
rect 8777 18215 8778 18241
rect 8750 18214 8778 18215
rect 10598 19417 10626 19418
rect 10598 19391 10599 19417
rect 10599 19391 10625 19417
rect 10625 19391 10626 19417
rect 10598 19390 10626 19391
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 8974 18241 9002 18242
rect 8974 18215 8975 18241
rect 8975 18215 9001 18241
rect 9001 18215 9002 18241
rect 8974 18214 9002 18215
rect 9310 18214 9338 18242
rect 7126 15974 7154 16002
rect 4382 14321 4410 14322
rect 4382 14295 4383 14321
rect 4383 14295 4409 14321
rect 4409 14295 4410 14321
rect 4382 14294 4410 14295
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 10598 17849 10626 17850
rect 10598 17823 10599 17849
rect 10599 17823 10625 17849
rect 10625 17823 10626 17849
rect 10598 17822 10626 17823
rect 8414 15974 8442 16002
rect 5894 14294 5922 14322
rect 3766 12361 3794 12362
rect 3766 12335 3767 12361
rect 3767 12335 3793 12361
rect 3793 12335 3794 12361
rect 3766 12334 3794 12335
rect 3990 12361 4018 12362
rect 3990 12335 3991 12361
rect 3991 12335 4017 12361
rect 4017 12335 4018 12361
rect 3990 12334 4018 12335
rect 4158 12334 4186 12362
rect 4102 11969 4130 11970
rect 4102 11943 4103 11969
rect 4103 11943 4129 11969
rect 4129 11943 4130 11969
rect 4102 11942 4130 11943
rect 4214 11942 4242 11970
rect 3318 11577 3346 11578
rect 3318 11551 3319 11577
rect 3319 11551 3345 11577
rect 3345 11551 3346 11577
rect 3318 11550 3346 11551
rect 3374 11102 3402 11130
rect 4102 11158 4130 11186
rect 4214 11102 4242 11130
rect 5054 11185 5082 11186
rect 5054 11159 5055 11185
rect 5055 11159 5081 11185
rect 5081 11159 5082 11185
rect 5054 11158 5082 11159
rect 4662 11102 4690 11130
rect 3038 10009 3066 10010
rect 3038 9983 3039 10009
rect 3039 9983 3065 10009
rect 3065 9983 3066 10009
rect 3038 9982 3066 9983
rect 6342 12334 6370 12362
rect 6174 11774 6202 11802
rect 5278 11185 5306 11186
rect 5278 11159 5279 11185
rect 5279 11159 5305 11185
rect 5305 11159 5306 11185
rect 5278 11158 5306 11159
rect 5222 11102 5250 11130
rect 3766 10009 3794 10010
rect 3766 9983 3767 10009
rect 3767 9983 3793 10009
rect 3793 9983 3794 10009
rect 3766 9982 3794 9983
rect 3318 9534 3346 9562
rect 3318 9254 3346 9282
rect 3766 9254 3794 9282
rect 2814 8441 2842 8442
rect 2814 8415 2815 8441
rect 2815 8415 2841 8441
rect 2841 8415 2842 8441
rect 2814 8414 2842 8415
rect 3038 8414 3066 8442
rect 3654 8441 3682 8442
rect 3654 8415 3655 8441
rect 3655 8415 3681 8441
rect 3681 8415 3682 8441
rect 3654 8414 3682 8415
rect 3598 8358 3626 8386
rect 5110 9254 5138 9282
rect 8414 12278 8442 12306
rect 8806 14238 8834 14266
rect 8806 13454 8834 13482
rect 7574 11774 7602 11802
rect 7798 11774 7826 11802
rect 6342 9534 6370 9562
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 8974 14238 9002 14266
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9534 13929 9562 13930
rect 9534 13903 9535 13929
rect 9535 13903 9561 13929
rect 9561 13903 9562 13929
rect 9534 13902 9562 13903
rect 8862 13510 8890 13538
rect 8974 13454 9002 13482
rect 10374 13510 10402 13538
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 8862 12278 8890 12306
rect 10822 13537 10850 13538
rect 10822 13511 10823 13537
rect 10823 13511 10849 13537
rect 10849 13511 10850 13537
rect 10822 13510 10850 13511
rect 10934 15470 10962 15498
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10318 12361 10346 12362
rect 10318 12335 10319 12361
rect 10319 12335 10345 12361
rect 10345 12335 10346 12361
rect 10318 12334 10346 12335
rect 8750 11774 8778 11802
rect 4998 8358 5026 8386
rect 3598 7657 3626 7658
rect 3598 7631 3599 7657
rect 3599 7631 3625 7657
rect 3625 7631 3626 7657
rect 3598 7630 3626 7631
rect 4998 7574 5026 7602
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 966 5726 994 5754
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 3990 6734 4018 6762
rect 6342 7574 6370 7602
rect 5558 6734 5586 6762
rect 2422 5697 2450 5698
rect 2422 5671 2423 5697
rect 2423 5671 2449 5697
rect 2449 5671 2450 5697
rect 2422 5670 2450 5671
rect 1582 5166 1610 5194
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2030 4494 2058 4522
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 3374 5697 3402 5698
rect 3374 5671 3375 5697
rect 3375 5671 3401 5697
rect 3401 5671 3402 5697
rect 3374 5670 3402 5671
rect 5558 6089 5586 6090
rect 5558 6063 5559 6089
rect 5559 6063 5585 6089
rect 5585 6063 5586 6089
rect 5558 6062 5586 6063
rect 2870 5166 2898 5194
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10934 12334 10962 12362
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 7518 7265 7546 7266
rect 7518 7239 7519 7265
rect 7519 7239 7545 7265
rect 7545 7239 7546 7265
rect 7518 7238 7546 7239
rect 8974 9617 9002 9618
rect 8974 9591 8975 9617
rect 8975 9591 9001 9617
rect 9001 9591 9002 9617
rect 8974 9590 9002 9591
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10318 10094 10346 10122
rect 9254 9590 9282 9618
rect 9086 9225 9114 9226
rect 9086 9199 9087 9225
rect 9087 9199 9113 9225
rect 9113 9199 9114 9225
rect 9086 9198 9114 9199
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9534 9254 9562 9282
rect 10822 10401 10850 10402
rect 10822 10375 10823 10401
rect 10823 10375 10849 10401
rect 10849 10375 10850 10401
rect 10822 10374 10850 10375
rect 10822 10094 10850 10122
rect 11102 22945 11130 22946
rect 11102 22919 11103 22945
rect 11103 22919 11129 22945
rect 11129 22919 11130 22945
rect 11102 22918 11130 22919
rect 12278 22918 12306 22946
rect 11382 22134 11410 22162
rect 11382 21854 11410 21882
rect 11270 21798 11298 21826
rect 11102 21742 11130 21770
rect 11102 20678 11130 20706
rect 11494 21825 11522 21826
rect 11494 21799 11495 21825
rect 11495 21799 11521 21825
rect 11521 21799 11522 21825
rect 11494 21798 11522 21799
rect 12838 22161 12866 22162
rect 12838 22135 12839 22161
rect 12839 22135 12865 22161
rect 12865 22135 12866 22161
rect 12838 22134 12866 22135
rect 12950 22161 12978 22162
rect 12950 22135 12951 22161
rect 12951 22135 12977 22161
rect 12977 22135 12978 22161
rect 12950 22134 12978 22135
rect 11550 21014 11578 21042
rect 11494 19809 11522 19810
rect 11494 19783 11495 19809
rect 11495 19783 11521 19809
rect 11521 19783 11522 19809
rect 11494 19782 11522 19783
rect 12558 20958 12586 20986
rect 12558 20678 12586 20706
rect 12558 20230 12586 20258
rect 11102 17822 11130 17850
rect 12726 21014 12754 21042
rect 13286 21014 13314 21042
rect 13118 20985 13146 20986
rect 13118 20959 13119 20985
rect 13119 20959 13145 20985
rect 13145 20959 13146 20985
rect 13118 20958 13146 20959
rect 13062 20230 13090 20258
rect 13118 20174 13146 20202
rect 13510 21014 13538 21042
rect 12726 19809 12754 19810
rect 12726 19783 12727 19809
rect 12727 19783 12753 19809
rect 12753 19783 12754 19809
rect 12726 19782 12754 19783
rect 12950 19809 12978 19810
rect 12950 19783 12951 19809
rect 12951 19783 12977 19809
rect 12977 19783 12978 19809
rect 12950 19782 12978 19783
rect 13566 19782 13594 19810
rect 11102 17457 11130 17458
rect 11102 17431 11103 17457
rect 11103 17431 11129 17457
rect 11129 17431 11130 17457
rect 11102 17430 11130 17431
rect 11270 16673 11298 16674
rect 11270 16647 11271 16673
rect 11271 16647 11297 16673
rect 11297 16647 11298 16673
rect 11270 16646 11298 16647
rect 12558 17457 12586 17458
rect 12558 17431 12559 17457
rect 12559 17431 12585 17457
rect 12585 17431 12586 17457
rect 12558 17430 12586 17431
rect 11494 16673 11522 16674
rect 11494 16647 11495 16673
rect 11495 16647 11521 16673
rect 11521 16647 11522 16673
rect 11494 16646 11522 16647
rect 11326 15918 11354 15946
rect 12782 18998 12810 19026
rect 12726 15918 12754 15946
rect 11718 14238 11746 14266
rect 11494 13929 11522 13930
rect 11494 13903 11495 13929
rect 11495 13903 11521 13929
rect 11521 13903 11522 13929
rect 11494 13902 11522 13903
rect 13118 17430 13146 17458
rect 13118 17065 13146 17066
rect 13118 17039 13119 17065
rect 13119 17039 13145 17065
rect 13145 17039 13146 17065
rect 13118 17038 13146 17039
rect 12950 15918 12978 15946
rect 13454 15918 13482 15946
rect 12782 13006 12810 13034
rect 13398 14265 13426 14266
rect 13398 14239 13399 14265
rect 13399 14239 13425 14265
rect 13425 14239 13426 14265
rect 13398 14238 13426 14239
rect 11494 11577 11522 11578
rect 11494 11551 11495 11577
rect 11495 11551 11521 11577
rect 11521 11551 11522 11577
rect 11494 11550 11522 11551
rect 12278 10766 12306 10794
rect 12838 12361 12866 12362
rect 12838 12335 12839 12361
rect 12839 12335 12865 12361
rect 12865 12335 12866 12361
rect 12838 12334 12866 12335
rect 13398 11577 13426 11578
rect 13398 11551 13399 11577
rect 13399 11551 13425 11577
rect 13425 11551 13426 11577
rect 13398 11550 13426 11551
rect 12838 10793 12866 10794
rect 12838 10767 12839 10793
rect 12839 10767 12865 10793
rect 12865 10767 12866 10793
rect 12838 10766 12866 10767
rect 12278 10401 12306 10402
rect 12278 10375 12279 10401
rect 12279 10375 12305 10401
rect 12305 10375 12306 10401
rect 12278 10374 12306 10375
rect 11046 9982 11074 10010
rect 13566 10094 13594 10122
rect 10318 9225 10346 9226
rect 10318 9199 10319 9225
rect 10319 9199 10345 9225
rect 10345 9199 10346 9225
rect 10318 9198 10346 9199
rect 10990 9254 11018 9282
rect 12558 9617 12586 9618
rect 12558 9591 12559 9617
rect 12559 9591 12585 9617
rect 12585 9591 12586 9617
rect 12558 9590 12586 9591
rect 13398 10009 13426 10010
rect 13398 9983 13399 10009
rect 13399 9983 13425 10009
rect 13425 9983 13426 10009
rect 13398 9982 13426 9983
rect 12838 9590 12866 9618
rect 11270 9281 11298 9282
rect 11270 9255 11271 9281
rect 11271 9255 11297 9281
rect 11297 9255 11298 9281
rect 11270 9254 11298 9255
rect 10598 8806 10626 8834
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 11102 8833 11130 8834
rect 11102 8807 11103 8833
rect 11103 8807 11129 8833
rect 11129 8807 11130 8833
rect 11102 8806 11130 8807
rect 12838 9225 12866 9226
rect 12838 9199 12839 9225
rect 12839 9199 12865 9225
rect 12865 9199 12866 9225
rect 12838 9198 12866 9199
rect 13342 9310 13370 9338
rect 10598 8441 10626 8442
rect 10598 8415 10599 8441
rect 10599 8415 10625 8441
rect 10625 8415 10626 8441
rect 10598 8414 10626 8415
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10598 7657 10626 7658
rect 10598 7631 10599 7657
rect 10599 7631 10625 7657
rect 10625 7631 10626 7657
rect 10598 7630 10626 7631
rect 11102 7630 11130 7658
rect 8750 7265 8778 7266
rect 8750 7239 8751 7265
rect 8751 7239 8777 7265
rect 8777 7239 8778 7265
rect 8750 7238 8778 7239
rect 8974 7265 9002 7266
rect 8974 7239 8975 7265
rect 8975 7239 9001 7265
rect 9001 7239 9002 7265
rect 8974 7238 9002 7239
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9814 6510 9842 6538
rect 6790 6089 6818 6090
rect 6790 6063 6791 6089
rect 6791 6063 6817 6089
rect 6817 6063 6818 6089
rect 6790 6062 6818 6063
rect 3542 4913 3570 4914
rect 3542 4887 3543 4913
rect 3543 4887 3569 4913
rect 3569 4887 3570 4913
rect 3542 4886 3570 4887
rect 5166 4913 5194 4914
rect 5166 4887 5167 4913
rect 5167 4887 5193 4913
rect 5193 4887 5194 4913
rect 5166 4886 5194 4887
rect 5390 4913 5418 4914
rect 5390 4887 5391 4913
rect 5391 4887 5417 4913
rect 5417 4887 5418 4913
rect 5390 4886 5418 4887
rect 3374 4521 3402 4522
rect 3374 4495 3375 4521
rect 3375 4495 3401 4521
rect 3401 4495 3402 4521
rect 3374 4494 3402 4495
rect 7014 4521 7042 4522
rect 7014 4495 7015 4521
rect 7015 4495 7041 4521
rect 7041 4495 7042 4521
rect 7014 4494 7042 4495
rect 7518 4494 7546 4522
rect 5782 4158 5810 4186
rect 4046 4102 4074 4130
rect 3822 3737 3850 3738
rect 3822 3711 3823 3737
rect 3823 3711 3849 3737
rect 3849 3711 3850 3737
rect 3822 3710 3850 3711
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 966 1806 994 1834
rect 1694 2030 1722 2058
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 4046 3737 4074 3738
rect 4046 3711 4047 3737
rect 4047 3711 4073 3737
rect 4073 3711 4074 3737
rect 4046 3710 4074 3711
rect 4494 3318 4522 3346
rect 6006 4158 6034 4186
rect 6566 4158 6594 4186
rect 6454 4129 6482 4130
rect 6454 4103 6455 4129
rect 6455 4103 6481 4129
rect 6481 4103 6482 4129
rect 6454 4102 6482 4103
rect 4998 3345 5026 3346
rect 4998 3319 4999 3345
rect 4999 3319 5025 3345
rect 5025 3319 5026 3345
rect 4998 3318 5026 3319
rect 5558 3345 5586 3346
rect 5558 3319 5559 3345
rect 5559 3319 5585 3345
rect 5585 3319 5586 3345
rect 5558 3318 5586 3319
rect 3990 2561 4018 2562
rect 3990 2535 3991 2561
rect 3991 2535 4017 2561
rect 4017 2535 4018 2561
rect 3990 2534 4018 2535
rect 4494 2169 4522 2170
rect 4494 2143 4495 2169
rect 4495 2143 4521 2169
rect 4521 2143 4522 2169
rect 4494 2142 4522 2143
rect 5558 2561 5586 2562
rect 5558 2535 5559 2561
rect 5559 2535 5585 2561
rect 5585 2535 5586 2561
rect 5558 2534 5586 2535
rect 5894 2926 5922 2954
rect 5894 2590 5922 2618
rect 4998 2142 5026 2170
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 2086 1777 2114 1778
rect 2086 1751 2087 1777
rect 2087 1751 2113 1777
rect 2113 1751 2114 1777
rect 2086 1750 2114 1751
rect 2870 1806 2898 1834
rect 3822 1777 3850 1778
rect 3822 1751 3823 1777
rect 3823 1751 3849 1777
rect 3849 1751 3850 1777
rect 3822 1750 3850 1751
rect 6286 2953 6314 2954
rect 6286 2927 6287 2953
rect 6287 2927 6313 2953
rect 6313 2927 6314 2953
rect 6286 2926 6314 2927
rect 6510 2953 6538 2954
rect 6510 2927 6511 2953
rect 6511 2927 6537 2953
rect 6537 2927 6538 2953
rect 6510 2926 6538 2927
rect 6118 2534 6146 2562
rect 7014 4102 7042 4130
rect 8974 5697 9002 5698
rect 8974 5671 8975 5697
rect 8975 5671 9001 5697
rect 9001 5671 9002 5697
rect 8974 5670 9002 5671
rect 9534 5697 9562 5698
rect 9534 5671 9535 5697
rect 9535 5671 9561 5697
rect 9561 5671 9562 5697
rect 9534 5670 9562 5671
rect 7014 3374 7042 3402
rect 7518 3374 7546 3402
rect 7798 3345 7826 3346
rect 7798 3319 7799 3345
rect 7799 3319 7825 3345
rect 7825 3319 7826 3345
rect 7798 3318 7826 3319
rect 6566 2478 6594 2506
rect 7014 2478 7042 2506
rect 7518 2169 7546 2170
rect 7518 2143 7519 2169
rect 7519 2143 7545 2169
rect 7545 2143 7546 2169
rect 7518 2142 7546 2143
rect 7630 2926 7658 2954
rect 6118 1750 6146 1778
rect 7462 1777 7490 1778
rect 7462 1751 7463 1777
rect 7463 1751 7489 1777
rect 7489 1751 7490 1777
rect 7462 1750 7490 1751
rect 7966 2953 7994 2954
rect 7966 2927 7967 2953
rect 7967 2927 7993 2953
rect 7993 2927 7994 2953
rect 7966 2926 7994 2927
rect 8246 2926 8274 2954
rect 8246 2561 8274 2562
rect 8246 2535 8247 2561
rect 8247 2535 8273 2561
rect 8273 2535 8274 2561
rect 8246 2534 8274 2535
rect 8078 2142 8106 2170
rect 8358 2478 8386 2506
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9814 5670 9842 5698
rect 10430 5894 10458 5922
rect 10990 5894 11018 5922
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 11102 6510 11130 6538
rect 11270 6734 11298 6762
rect 11998 6510 12026 6538
rect 12278 6734 12306 6762
rect 12446 6510 12474 6538
rect 13510 10009 13538 10010
rect 13510 9983 13511 10009
rect 13511 9983 13537 10009
rect 13537 9983 13538 10009
rect 13510 9982 13538 9983
rect 13398 9254 13426 9282
rect 13510 9310 13538 9338
rect 12838 6734 12866 6762
rect 13398 6510 13426 6538
rect 11998 5894 12026 5922
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 10038 4046 10066 4074
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 11998 4913 12026 4914
rect 11998 4887 11999 4913
rect 11999 4887 12025 4913
rect 12025 4887 12026 4913
rect 11998 4886 12026 4887
rect 11102 4046 11130 4074
rect 11550 4046 11578 4074
rect 8470 2561 8498 2562
rect 8470 2535 8471 2561
rect 8471 2535 8497 2561
rect 8497 2535 8498 2561
rect 8470 2534 8498 2535
rect 8806 2478 8834 2506
rect 9254 3345 9282 3346
rect 9254 3319 9255 3345
rect 9255 3319 9281 3345
rect 9281 3319 9282 3345
rect 9254 3318 9282 3319
rect 9310 2953 9338 2954
rect 9310 2927 9311 2953
rect 9311 2927 9337 2953
rect 9337 2927 9338 2953
rect 9310 2926 9338 2927
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 8470 2422 8498 2450
rect 9590 2422 9618 2450
rect 9758 2422 9786 2450
rect 11102 3710 11130 3738
rect 11550 3737 11578 3738
rect 11550 3711 11551 3737
rect 11551 3711 11577 3737
rect 11577 3711 11578 3737
rect 11550 3710 11578 3711
rect 11046 2953 11074 2954
rect 11046 2927 11047 2953
rect 11047 2927 11073 2953
rect 11073 2927 11074 2953
rect 11046 2926 11074 2927
rect 10430 2505 10458 2506
rect 10430 2479 10431 2505
rect 10431 2479 10457 2505
rect 10457 2479 10458 2505
rect 10430 2478 10458 2479
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10430 2169 10458 2170
rect 10430 2143 10431 2169
rect 10431 2143 10457 2169
rect 10457 2143 10458 2169
rect 10430 2142 10458 2143
rect 10878 2254 10906 2282
rect 9590 2086 9618 2114
rect 8078 1694 8106 1722
rect 8302 1750 8330 1778
rect 9422 1777 9450 1778
rect 9422 1751 9423 1777
rect 9423 1751 9449 1777
rect 9449 1751 9450 1777
rect 9422 1750 9450 1751
rect 11158 2086 11186 2114
rect 11494 3262 11522 3290
rect 12278 4886 12306 4914
rect 12558 4998 12586 5026
rect 12222 4046 12250 4074
rect 13118 4998 13146 5026
rect 13398 4913 13426 4914
rect 13398 4887 13399 4913
rect 13399 4887 13425 4913
rect 13425 4887 13426 4913
rect 13398 4886 13426 4887
rect 13342 4158 13370 4186
rect 12558 3710 12586 3738
rect 13118 3737 13146 3738
rect 13118 3711 13119 3737
rect 13119 3711 13145 3737
rect 13145 3711 13146 3737
rect 13118 3710 13146 3711
rect 12446 3374 12474 3402
rect 12558 3374 12586 3402
rect 13118 3374 13146 3402
rect 12726 3262 12754 3290
rect 12950 3262 12978 3290
rect 13230 3318 13258 3346
rect 13286 3262 13314 3290
rect 13230 2926 13258 2954
rect 13454 2926 13482 2954
rect 11382 2086 11410 2114
rect 11606 2254 11634 2282
rect 10878 1777 10906 1778
rect 10878 1751 10879 1777
rect 10879 1751 10905 1777
rect 10905 1751 10906 1777
rect 10878 1750 10906 1751
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 12558 2254 12586 2282
rect 18494 28742 18522 28770
rect 17598 27845 17626 27846
rect 17598 27819 17599 27845
rect 17599 27819 17625 27845
rect 17625 27819 17626 27845
rect 17598 27818 17626 27819
rect 17650 27845 17678 27846
rect 17650 27819 17651 27845
rect 17651 27819 17677 27845
rect 17677 27819 17678 27845
rect 17650 27818 17678 27819
rect 17702 27845 17730 27846
rect 17702 27819 17703 27845
rect 17703 27819 17729 27845
rect 17729 27819 17730 27845
rect 17702 27818 17730 27819
rect 15582 22889 15610 22890
rect 15582 22863 15583 22889
rect 15583 22863 15609 22889
rect 15609 22863 15610 22889
rect 15582 22862 15610 22863
rect 15862 22889 15890 22890
rect 15862 22863 15863 22889
rect 15863 22863 15889 22889
rect 15889 22863 15890 22889
rect 15862 22862 15890 22863
rect 15974 22638 16002 22666
rect 15582 22609 15610 22610
rect 15582 22583 15583 22609
rect 15583 22583 15609 22609
rect 15609 22583 15610 22609
rect 15582 22582 15610 22583
rect 15750 22609 15778 22610
rect 15750 22583 15751 22609
rect 15751 22583 15777 22609
rect 15777 22583 15778 22609
rect 15750 22582 15778 22583
rect 15862 21798 15890 21826
rect 17598 27061 17626 27062
rect 17598 27035 17599 27061
rect 17599 27035 17625 27061
rect 17625 27035 17626 27061
rect 17598 27034 17626 27035
rect 17650 27061 17678 27062
rect 17650 27035 17651 27061
rect 17651 27035 17677 27061
rect 17677 27035 17678 27061
rect 17650 27034 17678 27035
rect 17702 27061 17730 27062
rect 17702 27035 17703 27061
rect 17703 27035 17729 27061
rect 17729 27035 17730 27061
rect 17702 27034 17730 27035
rect 17598 26277 17626 26278
rect 17598 26251 17599 26277
rect 17599 26251 17625 26277
rect 17625 26251 17626 26277
rect 17598 26250 17626 26251
rect 17650 26277 17678 26278
rect 17650 26251 17651 26277
rect 17651 26251 17677 26277
rect 17677 26251 17678 26277
rect 17650 26250 17678 26251
rect 17702 26277 17730 26278
rect 17702 26251 17703 26277
rect 17703 26251 17729 26277
rect 17729 26251 17730 26277
rect 17702 26250 17730 26251
rect 18102 25662 18130 25690
rect 17598 25493 17626 25494
rect 17598 25467 17599 25493
rect 17599 25467 17625 25493
rect 17625 25467 17626 25493
rect 17598 25466 17626 25467
rect 17650 25493 17678 25494
rect 17650 25467 17651 25493
rect 17651 25467 17677 25493
rect 17677 25467 17678 25493
rect 17650 25466 17678 25467
rect 17702 25493 17730 25494
rect 17702 25467 17703 25493
rect 17703 25467 17729 25493
rect 17729 25467 17730 25493
rect 17702 25466 17730 25467
rect 17542 25270 17570 25298
rect 16982 24878 17010 24906
rect 16814 24486 16842 24514
rect 16198 23702 16226 23730
rect 16478 23729 16506 23730
rect 16478 23703 16479 23729
rect 16479 23703 16505 23729
rect 16505 23703 16506 23729
rect 16478 23702 16506 23703
rect 17150 24513 17178 24514
rect 17150 24487 17151 24513
rect 17151 24487 17177 24513
rect 17177 24487 17178 24513
rect 17150 24486 17178 24487
rect 17318 24513 17346 24514
rect 17318 24487 17319 24513
rect 17319 24487 17345 24513
rect 17345 24487 17346 24513
rect 17318 24486 17346 24487
rect 16142 22862 16170 22890
rect 16198 22638 16226 22666
rect 16422 22582 16450 22610
rect 16310 22553 16338 22554
rect 16310 22527 16311 22553
rect 16311 22527 16337 22553
rect 16337 22527 16338 22553
rect 16310 22526 16338 22527
rect 16478 22553 16506 22554
rect 16478 22527 16479 22553
rect 16479 22527 16505 22553
rect 16505 22527 16506 22553
rect 16478 22526 16506 22527
rect 16142 22134 16170 22162
rect 16422 22161 16450 22162
rect 16422 22135 16423 22161
rect 16423 22135 16449 22161
rect 16449 22135 16450 22161
rect 16422 22134 16450 22135
rect 16702 22945 16730 22946
rect 16702 22919 16703 22945
rect 16703 22919 16729 22945
rect 16729 22919 16730 22945
rect 16702 22918 16730 22919
rect 16870 22918 16898 22946
rect 16870 22134 16898 22162
rect 16870 21854 16898 21882
rect 17262 24177 17290 24178
rect 17262 24151 17263 24177
rect 17263 24151 17289 24177
rect 17289 24151 17290 24177
rect 17262 24150 17290 24151
rect 17038 24094 17066 24122
rect 17206 24121 17234 24122
rect 17206 24095 17207 24121
rect 17207 24095 17233 24121
rect 17233 24095 17234 24121
rect 17206 24094 17234 24095
rect 17038 23729 17066 23730
rect 17038 23703 17039 23729
rect 17039 23703 17065 23729
rect 17065 23703 17066 23729
rect 17038 23702 17066 23703
rect 17206 23478 17234 23506
rect 17822 25214 17850 25242
rect 18326 25270 18354 25298
rect 17710 24905 17738 24906
rect 17710 24879 17711 24905
rect 17711 24879 17737 24905
rect 17737 24879 17738 24905
rect 17710 24878 17738 24879
rect 17598 24709 17626 24710
rect 17598 24683 17599 24709
rect 17599 24683 17625 24709
rect 17625 24683 17626 24709
rect 17598 24682 17626 24683
rect 17650 24709 17678 24710
rect 17650 24683 17651 24709
rect 17651 24683 17677 24709
rect 17677 24683 17678 24709
rect 17650 24682 17678 24683
rect 17702 24709 17730 24710
rect 17702 24683 17703 24709
rect 17703 24683 17729 24709
rect 17729 24683 17730 24709
rect 17702 24682 17730 24683
rect 17430 24177 17458 24178
rect 17430 24151 17431 24177
rect 17431 24151 17457 24177
rect 17457 24151 17458 24177
rect 17430 24150 17458 24151
rect 17710 24513 17738 24514
rect 17710 24487 17711 24513
rect 17711 24487 17737 24513
rect 17737 24487 17738 24513
rect 17710 24486 17738 24487
rect 18214 25241 18242 25242
rect 18214 25215 18215 25241
rect 18215 25215 18241 25241
rect 18241 25215 18242 25241
rect 18214 25214 18242 25215
rect 18102 24878 18130 24906
rect 17822 24177 17850 24178
rect 17822 24151 17823 24177
rect 17823 24151 17849 24177
rect 17849 24151 17850 24177
rect 17822 24150 17850 24151
rect 17654 24094 17682 24122
rect 17878 24513 17906 24514
rect 17878 24487 17879 24513
rect 17879 24487 17905 24513
rect 17905 24487 17906 24513
rect 17878 24486 17906 24487
rect 17598 23925 17626 23926
rect 17598 23899 17599 23925
rect 17599 23899 17625 23925
rect 17625 23899 17626 23925
rect 17598 23898 17626 23899
rect 17650 23925 17678 23926
rect 17650 23899 17651 23925
rect 17651 23899 17677 23925
rect 17677 23899 17678 23925
rect 17650 23898 17678 23899
rect 17702 23925 17730 23926
rect 17702 23899 17703 23925
rect 17703 23899 17729 23925
rect 17729 23899 17730 23925
rect 17702 23898 17730 23899
rect 17990 24177 18018 24178
rect 17990 24151 17991 24177
rect 17991 24151 18017 24177
rect 18017 24151 18018 24177
rect 17990 24150 18018 24151
rect 18550 25689 18578 25690
rect 18550 25663 18551 25689
rect 18551 25663 18577 25689
rect 18577 25663 18578 25689
rect 18550 25662 18578 25663
rect 18494 25270 18522 25298
rect 18382 25241 18410 25242
rect 18382 25215 18383 25241
rect 18383 25215 18409 25241
rect 18409 25215 18410 25241
rect 18382 25214 18410 25215
rect 18270 24513 18298 24514
rect 18270 24487 18271 24513
rect 18271 24487 18297 24513
rect 18297 24487 18298 24513
rect 18270 24486 18298 24487
rect 18158 24150 18186 24178
rect 18438 24513 18466 24514
rect 18438 24487 18439 24513
rect 18439 24487 18465 24513
rect 18465 24487 18466 24513
rect 18438 24486 18466 24487
rect 17990 23646 18018 23674
rect 17710 23478 17738 23506
rect 17038 22945 17066 22946
rect 17038 22919 17039 22945
rect 17039 22919 17065 22945
rect 17065 22919 17066 22945
rect 17038 22918 17066 22919
rect 17598 23141 17626 23142
rect 17598 23115 17599 23141
rect 17599 23115 17625 23141
rect 17625 23115 17626 23141
rect 17598 23114 17626 23115
rect 17650 23141 17678 23142
rect 17650 23115 17651 23141
rect 17651 23115 17677 23141
rect 17677 23115 17678 23141
rect 17650 23114 17678 23115
rect 17702 23141 17730 23142
rect 17702 23115 17703 23141
rect 17703 23115 17729 23141
rect 17729 23115 17730 23141
rect 17702 23114 17730 23115
rect 17150 22609 17178 22610
rect 17150 22583 17151 22609
rect 17151 22583 17177 22609
rect 17177 22583 17178 22609
rect 17150 22582 17178 22583
rect 16982 22161 17010 22162
rect 16982 22135 16983 22161
rect 16983 22135 17009 22161
rect 17009 22135 17010 22161
rect 16982 22134 17010 22135
rect 16926 21798 16954 21826
rect 17430 22582 17458 22610
rect 18214 23673 18242 23674
rect 18214 23647 18215 23673
rect 18215 23647 18241 23673
rect 18241 23647 18242 23673
rect 18214 23646 18242 23647
rect 18326 23478 18354 23506
rect 18382 23646 18410 23674
rect 17542 22553 17570 22554
rect 17542 22527 17543 22553
rect 17543 22527 17569 22553
rect 17569 22527 17570 22553
rect 17542 22526 17570 22527
rect 17598 22357 17626 22358
rect 17598 22331 17599 22357
rect 17599 22331 17625 22357
rect 17625 22331 17626 22357
rect 17598 22330 17626 22331
rect 17650 22357 17678 22358
rect 17650 22331 17651 22357
rect 17651 22331 17677 22357
rect 17677 22331 17678 22357
rect 17650 22330 17678 22331
rect 17702 22357 17730 22358
rect 17702 22331 17703 22357
rect 17703 22331 17729 22357
rect 17729 22331 17730 22357
rect 17702 22330 17730 22331
rect 16030 21238 16058 21266
rect 17318 21742 17346 21770
rect 17486 21854 17514 21882
rect 17598 21769 17626 21770
rect 17598 21743 17599 21769
rect 17599 21743 17625 21769
rect 17625 21743 17626 21769
rect 17598 21742 17626 21743
rect 17710 21769 17738 21770
rect 17710 21743 17711 21769
rect 17711 21743 17737 21769
rect 17737 21743 17738 21769
rect 17710 21742 17738 21743
rect 17598 21573 17626 21574
rect 17598 21547 17599 21573
rect 17599 21547 17625 21573
rect 17625 21547 17626 21573
rect 17598 21546 17626 21547
rect 17650 21573 17678 21574
rect 17650 21547 17651 21573
rect 17651 21547 17677 21573
rect 17677 21547 17678 21573
rect 17650 21546 17678 21547
rect 17702 21573 17730 21574
rect 17702 21547 17703 21573
rect 17703 21547 17729 21573
rect 17729 21547 17730 21573
rect 17702 21546 17730 21547
rect 17822 21854 17850 21882
rect 18102 22609 18130 22610
rect 18102 22583 18103 22609
rect 18103 22583 18129 22609
rect 18129 22583 18130 22609
rect 18102 22582 18130 22583
rect 18046 21854 18074 21882
rect 18270 22609 18298 22610
rect 18270 22583 18271 22609
rect 18271 22583 18297 22609
rect 18297 22583 18298 22609
rect 18270 22582 18298 22583
rect 18158 21854 18186 21882
rect 17990 21238 18018 21266
rect 17934 21070 17962 21098
rect 16982 21014 17010 21042
rect 17654 21041 17682 21042
rect 17654 21015 17655 21041
rect 17655 21015 17681 21041
rect 17681 21015 17682 21041
rect 17654 21014 17682 21015
rect 17598 20789 17626 20790
rect 17598 20763 17599 20789
rect 17599 20763 17625 20789
rect 17625 20763 17626 20789
rect 17598 20762 17626 20763
rect 17650 20789 17678 20790
rect 17650 20763 17651 20789
rect 17651 20763 17677 20789
rect 17677 20763 17678 20789
rect 17650 20762 17678 20763
rect 17702 20789 17730 20790
rect 17702 20763 17703 20789
rect 17703 20763 17729 20789
rect 17729 20763 17730 20789
rect 17702 20762 17730 20763
rect 14630 20230 14658 20258
rect 14574 20201 14602 20202
rect 14574 20175 14575 20201
rect 14575 20175 14601 20201
rect 14601 20175 14602 20201
rect 14574 20174 14602 20175
rect 15078 20174 15106 20202
rect 15078 18270 15106 18298
rect 17598 20005 17626 20006
rect 17598 19979 17599 20005
rect 17599 19979 17625 20005
rect 17625 19979 17626 20005
rect 17598 19978 17626 19979
rect 17650 20005 17678 20006
rect 17650 19979 17651 20005
rect 17651 19979 17677 20005
rect 17677 19979 17678 20005
rect 17650 19978 17678 19979
rect 17702 20005 17730 20006
rect 17702 19979 17703 20005
rect 17703 19979 17729 20005
rect 17729 19979 17730 20005
rect 17702 19978 17730 19979
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 15246 18689 15274 18690
rect 15246 18663 15247 18689
rect 15247 18663 15273 18689
rect 15273 18663 15274 18689
rect 15246 18662 15274 18663
rect 14854 17430 14882 17458
rect 14574 17065 14602 17066
rect 14574 17039 14575 17065
rect 14575 17039 14601 17065
rect 14601 17039 14602 17065
rect 14574 17038 14602 17039
rect 16254 19025 16282 19026
rect 16254 18999 16255 19025
rect 16255 18999 16281 19025
rect 16281 18999 16282 19025
rect 16254 18998 16282 18999
rect 16814 18662 16842 18690
rect 18550 21854 18578 21882
rect 18382 21742 18410 21770
rect 18382 21321 18410 21322
rect 18382 21295 18383 21321
rect 18383 21295 18409 21321
rect 18409 21295 18410 21321
rect 18382 21294 18410 21295
rect 18214 21070 18242 21098
rect 18102 21014 18130 21042
rect 18494 20985 18522 20986
rect 18494 20959 18495 20985
rect 18495 20959 18521 20985
rect 18521 20959 18522 20985
rect 18494 20958 18522 20959
rect 18438 20593 18466 20594
rect 18438 20567 18439 20593
rect 18439 20567 18465 20593
rect 18465 20567 18466 20593
rect 18438 20566 18466 20567
rect 18102 19809 18130 19810
rect 18102 19783 18103 19809
rect 18103 19783 18129 19809
rect 18129 19783 18130 19809
rect 18102 19782 18130 19783
rect 18270 19809 18298 19810
rect 18270 19783 18271 19809
rect 18271 19783 18297 19809
rect 18297 19783 18298 19809
rect 18270 19782 18298 19783
rect 18494 19782 18522 19810
rect 18382 19753 18410 19754
rect 18382 19727 18383 19753
rect 18383 19727 18409 19753
rect 18409 19727 18410 19753
rect 18382 19726 18410 19727
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 15918 18241 15946 18242
rect 15918 18215 15919 18241
rect 15919 18215 15945 18241
rect 15945 18215 15946 18241
rect 15918 18214 15946 18215
rect 16254 18270 16282 18298
rect 16814 18270 16842 18298
rect 16758 18241 16786 18242
rect 16758 18215 16759 18241
rect 16759 18215 16785 18241
rect 16785 18215 16786 18241
rect 16758 18214 16786 18215
rect 16926 18241 16954 18242
rect 16926 18215 16927 18241
rect 16927 18215 16953 18241
rect 16953 18215 16954 18241
rect 16926 18214 16954 18215
rect 17262 18214 17290 18242
rect 16254 17457 16282 17458
rect 16254 17431 16255 17457
rect 16255 17431 16281 17457
rect 16281 17431 16282 17457
rect 16254 17430 16282 17431
rect 14294 15862 14322 15890
rect 14798 15889 14826 15890
rect 14798 15863 14799 15889
rect 14799 15863 14825 15889
rect 14825 15863 14826 15889
rect 14798 15862 14826 15863
rect 15190 15862 15218 15890
rect 14294 15497 14322 15498
rect 14294 15471 14295 15497
rect 14295 15471 14321 15497
rect 14321 15471 14322 15497
rect 14294 15470 14322 15471
rect 15190 15526 15218 15554
rect 14798 14321 14826 14322
rect 14798 14295 14799 14321
rect 14799 14295 14825 14321
rect 14825 14295 14826 14321
rect 14798 14294 14826 14295
rect 15190 14238 15218 14266
rect 14294 12361 14322 12362
rect 14294 12335 14295 12361
rect 14295 12335 14321 12361
rect 14321 12335 14322 12361
rect 14294 12334 14322 12335
rect 13678 10094 13706 10122
rect 14574 11942 14602 11970
rect 15078 11969 15106 11970
rect 15078 11943 15079 11969
rect 15079 11943 15105 11969
rect 15105 11943 15106 11969
rect 15078 11942 15106 11943
rect 14294 9225 14322 9226
rect 14294 9199 14295 9225
rect 14295 9199 14321 9225
rect 14321 9199 14322 9225
rect 14294 9198 14322 9199
rect 14294 8862 14322 8890
rect 15134 11577 15162 11578
rect 15134 11551 15135 11577
rect 15135 11551 15161 11577
rect 15161 11551 15162 11577
rect 15134 11550 15162 11551
rect 15302 15553 15330 15554
rect 15302 15527 15303 15553
rect 15303 15527 15329 15553
rect 15329 15527 15330 15553
rect 15302 15526 15330 15527
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 16814 15889 16842 15890
rect 16814 15863 16815 15889
rect 16815 15863 16841 15889
rect 16841 15863 16842 15889
rect 16814 15862 16842 15863
rect 17206 15862 17234 15890
rect 15470 13537 15498 13538
rect 15470 13511 15471 13537
rect 15471 13511 15497 13537
rect 15497 13511 15498 13537
rect 15470 13510 15498 13511
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 16534 14321 16562 14322
rect 16534 14295 16535 14321
rect 16535 14295 16561 14321
rect 16561 14295 16562 14321
rect 16534 14294 16562 14295
rect 16814 14294 16842 14322
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 16814 13537 16842 13538
rect 16814 13511 16815 13537
rect 16815 13511 16841 13537
rect 16841 13511 16842 13537
rect 16814 13510 16842 13511
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 17262 13510 17290 13538
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 16254 11942 16282 11970
rect 15246 11550 15274 11578
rect 14742 9254 14770 9282
rect 14574 8806 14602 8834
rect 14798 8862 14826 8890
rect 15134 8806 15162 8834
rect 15246 8833 15274 8834
rect 15246 8807 15247 8833
rect 15247 8807 15273 8833
rect 15273 8807 15274 8833
rect 15246 8806 15274 8807
rect 14294 8022 14322 8050
rect 15190 8078 15218 8106
rect 14294 6734 14322 6762
rect 16422 10374 16450 10402
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 16926 10401 16954 10402
rect 16926 10375 16927 10401
rect 16927 10375 16953 10401
rect 16953 10375 16954 10401
rect 16926 10374 16954 10375
rect 17206 10374 17234 10402
rect 17150 10318 17178 10346
rect 15974 9534 16002 9562
rect 16254 9534 16282 9562
rect 16758 9617 16786 9618
rect 16758 9591 16759 9617
rect 16759 9591 16785 9617
rect 16785 9591 16786 9617
rect 16758 9590 16786 9591
rect 17150 9590 17178 9618
rect 16478 9534 16506 9562
rect 15470 8833 15498 8834
rect 15470 8807 15471 8833
rect 15471 8807 15497 8833
rect 15497 8807 15498 8833
rect 15470 8806 15498 8807
rect 15246 7265 15274 7266
rect 15246 7239 15247 7265
rect 15247 7239 15273 7265
rect 15273 7239 15274 7265
rect 15246 7238 15274 7239
rect 14798 6734 14826 6762
rect 14014 6510 14042 6538
rect 15246 6510 15274 6538
rect 14574 6454 14602 6482
rect 14910 6454 14938 6482
rect 14574 4998 14602 5026
rect 14014 4886 14042 4914
rect 14574 4886 14602 4914
rect 14518 3737 14546 3738
rect 14518 3711 14519 3737
rect 14519 3711 14545 3737
rect 14545 3711 14546 3737
rect 14518 3710 14546 3711
rect 14014 2953 14042 2954
rect 14014 2927 14015 2953
rect 14015 2927 14041 2953
rect 14041 2927 14042 2953
rect 14014 2926 14042 2927
rect 13622 2422 13650 2450
rect 14350 2478 14378 2506
rect 11662 2142 11690 2170
rect 12670 1806 12698 1834
rect 12838 1806 12866 1834
rect 14350 2198 14378 2226
rect 14294 2030 14322 2058
rect 14742 4158 14770 4186
rect 15358 8078 15386 8106
rect 15694 8049 15722 8050
rect 15694 8023 15695 8049
rect 15695 8023 15721 8049
rect 15721 8023 15722 8049
rect 15694 8022 15722 8023
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 17486 10401 17514 10402
rect 17486 10375 17487 10401
rect 17487 10375 17513 10401
rect 17513 10375 17514 10401
rect 17486 10374 17514 10375
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 17766 9534 17794 9562
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 17542 8078 17570 8106
rect 15470 7265 15498 7266
rect 15470 7239 15471 7265
rect 15471 7239 15497 7265
rect 15497 7239 15498 7265
rect 15470 7238 15498 7239
rect 15358 6510 15386 6538
rect 15694 6481 15722 6482
rect 15694 6455 15695 6481
rect 15695 6455 15721 6481
rect 15721 6455 15722 6481
rect 15694 6454 15722 6455
rect 15918 7238 15946 7266
rect 15470 5614 15498 5642
rect 16254 7209 16282 7210
rect 16254 7183 16255 7209
rect 16255 7183 16281 7209
rect 16281 7183 16282 7209
rect 16254 7182 16282 7183
rect 17150 6454 17178 6482
rect 15918 5614 15946 5642
rect 15974 5641 16002 5642
rect 15974 5615 15975 5641
rect 15975 5615 16001 5641
rect 16001 5615 16002 5641
rect 15974 5614 16002 5615
rect 16254 5641 16282 5642
rect 16254 5615 16255 5641
rect 16255 5615 16281 5641
rect 16281 5615 16282 5641
rect 16254 5614 16282 5615
rect 15918 4913 15946 4914
rect 15918 4887 15919 4913
rect 15919 4887 15945 4913
rect 15945 4887 15946 4913
rect 15918 4886 15946 4887
rect 17150 4886 17178 4914
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 18998 26446 19026 26474
rect 18662 25214 18690 25242
rect 18774 24513 18802 24514
rect 18774 24487 18775 24513
rect 18775 24487 18801 24513
rect 18801 24487 18802 24513
rect 18774 24486 18802 24487
rect 18718 23646 18746 23674
rect 19054 25297 19082 25298
rect 19054 25271 19055 25297
rect 19055 25271 19081 25297
rect 19081 25271 19082 25297
rect 19054 25270 19082 25271
rect 18942 23673 18970 23674
rect 18942 23647 18943 23673
rect 18943 23647 18969 23673
rect 18969 23647 18970 23673
rect 18942 23646 18970 23647
rect 18998 23478 19026 23506
rect 19054 21854 19082 21882
rect 18718 21769 18746 21770
rect 18718 21743 18719 21769
rect 18719 21743 18745 21769
rect 18745 21743 18746 21769
rect 18718 21742 18746 21743
rect 18774 21321 18802 21322
rect 18774 21295 18775 21321
rect 18775 21295 18801 21321
rect 18801 21295 18802 21321
rect 18774 21294 18802 21295
rect 18774 20566 18802 20594
rect 18998 20985 19026 20986
rect 18998 20959 18999 20985
rect 18999 20959 19025 20985
rect 19025 20959 19026 20985
rect 18998 20958 19026 20959
rect 18718 19782 18746 19810
rect 18998 19558 19026 19586
rect 19054 19753 19082 19754
rect 19054 19727 19055 19753
rect 19055 19727 19081 19753
rect 19081 19727 19082 19753
rect 19054 19726 19082 19727
rect 18606 9534 18634 9562
rect 19054 17262 19082 17290
rect 19054 14966 19082 14994
rect 19054 12670 19082 12698
rect 18718 10318 18746 10346
rect 18774 10374 18802 10402
rect 17542 4494 17570 4522
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 16478 4214 16506 4242
rect 17990 4214 18018 4242
rect 17878 4129 17906 4130
rect 17878 4103 17879 4129
rect 17879 4103 17905 4129
rect 17905 4103 17906 4129
rect 17878 4102 17906 4103
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 16758 3430 16786 3458
rect 17486 3430 17514 3458
rect 15358 2926 15386 2954
rect 14798 2478 14826 2506
rect 15246 2422 15274 2450
rect 16926 2534 16954 2562
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 18382 4494 18410 4522
rect 18774 4521 18802 4522
rect 18774 4495 18775 4521
rect 18775 4495 18801 4521
rect 18801 4495 18802 4521
rect 18774 4494 18802 4495
rect 18438 4102 18466 4130
rect 18214 4046 18242 4074
rect 15470 2422 15498 2450
rect 15526 2030 15554 2058
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 18382 3345 18410 3346
rect 18382 3319 18383 3345
rect 18383 3319 18409 3345
rect 18409 3319 18410 3345
rect 18382 3318 18410 3319
rect 18774 3318 18802 3346
rect 18774 2534 18802 2562
rect 18774 1190 18802 1218
<< metal3 >>
rect 19600 28770 20000 28784
rect 18489 28742 18494 28770
rect 18522 28742 20000 28770
rect 19600 28728 20000 28742
rect 9913 28210 9918 28238
rect 9946 28210 9970 28238
rect 9998 28210 10022 28238
rect 10050 28210 10055 28238
rect 0 27930 400 27944
rect 0 27902 1750 27930
rect 1778 27902 1783 27930
rect 0 27888 400 27902
rect 2233 27818 2238 27846
rect 2266 27818 2290 27846
rect 2318 27818 2342 27846
rect 2370 27818 2375 27846
rect 17593 27818 17598 27846
rect 17626 27818 17650 27846
rect 17678 27818 17702 27846
rect 17730 27818 17735 27846
rect 9913 27426 9918 27454
rect 9946 27426 9970 27454
rect 9998 27426 10022 27454
rect 10050 27426 10055 27454
rect 2233 27034 2238 27062
rect 2266 27034 2290 27062
rect 2318 27034 2342 27062
rect 2370 27034 2375 27062
rect 17593 27034 17598 27062
rect 17626 27034 17650 27062
rect 17678 27034 17702 27062
rect 17730 27034 17735 27062
rect 1353 26894 1358 26922
rect 1386 26894 2086 26922
rect 2114 26894 2119 26922
rect 3817 26838 3822 26866
rect 3850 26838 4494 26866
rect 4522 26838 4527 26866
rect 9913 26642 9918 26670
rect 9946 26642 9970 26670
rect 9998 26642 10022 26670
rect 10050 26642 10055 26670
rect 19600 26474 20000 26488
rect 4186 26446 4494 26474
rect 4522 26446 5726 26474
rect 5754 26446 5759 26474
rect 18993 26446 18998 26474
rect 19026 26446 20000 26474
rect 4186 26418 4214 26446
rect 19600 26432 20000 26446
rect 2809 26390 2814 26418
rect 2842 26390 4214 26418
rect 2233 26250 2238 26278
rect 2266 26250 2290 26278
rect 2318 26250 2342 26278
rect 2370 26250 2375 26278
rect 17593 26250 17598 26278
rect 17626 26250 17650 26278
rect 17678 26250 17702 26278
rect 17730 26250 17735 26278
rect 3313 26054 3318 26082
rect 3346 26054 4830 26082
rect 4858 26054 5166 26082
rect 5194 26054 5199 26082
rect 9913 25858 9918 25886
rect 9946 25858 9970 25886
rect 9998 25858 10022 25886
rect 10050 25858 10055 25886
rect 18097 25662 18102 25690
rect 18130 25662 18550 25690
rect 18578 25662 18583 25690
rect 2233 25466 2238 25494
rect 2266 25466 2290 25494
rect 2318 25466 2342 25494
rect 2370 25466 2375 25494
rect 17593 25466 17598 25494
rect 17626 25466 17650 25494
rect 17678 25466 17702 25494
rect 17730 25466 17735 25494
rect 2473 25270 2478 25298
rect 2506 25270 2814 25298
rect 2842 25270 2847 25298
rect 17537 25270 17542 25298
rect 17570 25270 18326 25298
rect 18354 25270 18494 25298
rect 18522 25270 19054 25298
rect 19082 25270 19087 25298
rect 1689 25214 1694 25242
rect 1722 25214 3094 25242
rect 3122 25214 3127 25242
rect 6281 25214 6286 25242
rect 6314 25214 17822 25242
rect 17850 25214 18214 25242
rect 18242 25214 18382 25242
rect 18410 25214 18662 25242
rect 18690 25214 18695 25242
rect 9913 25074 9918 25102
rect 9946 25074 9970 25102
rect 9998 25074 10022 25102
rect 10050 25074 10055 25102
rect 5721 24934 5726 24962
rect 5754 24934 7518 24962
rect 7546 24934 7551 24962
rect 5161 24878 5166 24906
rect 5194 24878 6622 24906
rect 6650 24878 6655 24906
rect 16977 24878 16982 24906
rect 17010 24878 17710 24906
rect 17738 24878 18102 24906
rect 18130 24878 18135 24906
rect 2233 24682 2238 24710
rect 2266 24682 2290 24710
rect 2318 24682 2342 24710
rect 2370 24682 2375 24710
rect 17593 24682 17598 24710
rect 17626 24682 17650 24710
rect 17678 24682 17702 24710
rect 17730 24682 17735 24710
rect 7121 24486 7126 24514
rect 7154 24486 8582 24514
rect 8610 24486 9142 24514
rect 9170 24486 9175 24514
rect 15946 24486 16814 24514
rect 16842 24486 17150 24514
rect 17178 24486 17318 24514
rect 17346 24486 17710 24514
rect 17738 24486 17878 24514
rect 17906 24486 18270 24514
rect 18298 24486 18438 24514
rect 18466 24486 18774 24514
rect 18802 24486 18807 24514
rect 15946 24458 15974 24486
rect 7513 24430 7518 24458
rect 7546 24430 7966 24458
rect 7994 24430 8358 24458
rect 8386 24430 8391 24458
rect 8745 24430 8750 24458
rect 8778 24430 15974 24458
rect 6617 24374 6622 24402
rect 6650 24374 7070 24402
rect 7098 24374 8582 24402
rect 8610 24374 8615 24402
rect 9913 24290 9918 24318
rect 9946 24290 9970 24318
rect 9998 24290 10022 24318
rect 10050 24290 10055 24318
rect 0 24234 400 24248
rect 0 24206 1918 24234
rect 1946 24206 1951 24234
rect 0 24192 400 24206
rect 19600 24178 20000 24192
rect 5833 24150 5838 24178
rect 5866 24150 7546 24178
rect 17257 24150 17262 24178
rect 17290 24150 17430 24178
rect 17458 24150 17822 24178
rect 17850 24150 17990 24178
rect 18018 24150 18023 24178
rect 18153 24150 18158 24178
rect 18186 24150 20000 24178
rect 7518 24122 7546 24150
rect 19600 24136 20000 24150
rect 2529 24094 2534 24122
rect 2562 24094 3542 24122
rect 3570 24094 3766 24122
rect 3794 24094 3990 24122
rect 4018 24094 4023 24122
rect 4881 24094 4886 24122
rect 4914 24094 5166 24122
rect 5194 24094 6062 24122
rect 6090 24094 6342 24122
rect 6370 24094 6375 24122
rect 7513 24094 7518 24122
rect 7546 24094 8022 24122
rect 8050 24094 8055 24122
rect 17033 24094 17038 24122
rect 17066 24094 17206 24122
rect 17234 24094 17654 24122
rect 17682 24094 17687 24122
rect 2233 23898 2238 23926
rect 2266 23898 2290 23926
rect 2318 23898 2342 23926
rect 2370 23898 2375 23926
rect 17593 23898 17598 23926
rect 17626 23898 17650 23926
rect 17678 23898 17702 23926
rect 17730 23898 17735 23926
rect 1577 23702 1582 23730
rect 1610 23702 1806 23730
rect 1834 23702 1839 23730
rect 1913 23702 1918 23730
rect 1946 23702 3150 23730
rect 3178 23702 3318 23730
rect 3346 23702 4886 23730
rect 4914 23702 4919 23730
rect 8409 23702 8414 23730
rect 8442 23702 9422 23730
rect 9450 23702 9455 23730
rect 16193 23702 16198 23730
rect 16226 23702 16478 23730
rect 16506 23702 17038 23730
rect 17066 23702 17071 23730
rect 3817 23646 3822 23674
rect 3850 23646 5782 23674
rect 5810 23646 5815 23674
rect 17985 23646 17990 23674
rect 18018 23646 18214 23674
rect 18242 23646 18382 23674
rect 18410 23646 18718 23674
rect 18746 23646 18942 23674
rect 18970 23646 18975 23674
rect 9913 23506 9918 23534
rect 9946 23506 9970 23534
rect 9998 23506 10022 23534
rect 10050 23506 10055 23534
rect 17201 23478 17206 23506
rect 17234 23478 17710 23506
rect 17738 23478 18326 23506
rect 18354 23478 18998 23506
rect 19026 23478 19031 23506
rect 9137 23310 9142 23338
rect 9170 23310 10598 23338
rect 10626 23310 10631 23338
rect 8577 23254 8582 23282
rect 8610 23254 9086 23282
rect 9114 23254 10374 23282
rect 10402 23254 10407 23282
rect 2233 23114 2238 23142
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2370 23114 2375 23142
rect 17593 23114 17598 23142
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17730 23114 17735 23142
rect 10593 22918 10598 22946
rect 10626 22918 11102 22946
rect 11130 22918 12278 22946
rect 12306 22918 12311 22946
rect 16697 22918 16702 22946
rect 16730 22918 16870 22946
rect 16898 22918 17038 22946
rect 17066 22918 17071 22946
rect 15577 22862 15582 22890
rect 15610 22862 15862 22890
rect 15890 22862 16142 22890
rect 16170 22862 16175 22890
rect 9913 22722 9918 22750
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 10050 22722 10055 22750
rect 15969 22638 15974 22666
rect 16002 22638 16198 22666
rect 16226 22638 16231 22666
rect 15577 22582 15582 22610
rect 15610 22582 15750 22610
rect 15778 22582 16422 22610
rect 16450 22582 16455 22610
rect 17145 22582 17150 22610
rect 17178 22582 17430 22610
rect 17458 22582 18102 22610
rect 18130 22582 18270 22610
rect 18298 22582 18303 22610
rect 8017 22526 8022 22554
rect 8050 22526 8358 22554
rect 8386 22526 9478 22554
rect 9506 22526 9511 22554
rect 16305 22526 16310 22554
rect 16338 22526 16478 22554
rect 16506 22526 17542 22554
rect 17570 22526 17575 22554
rect 2233 22330 2238 22358
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2370 22330 2375 22358
rect 17593 22330 17598 22358
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17730 22330 17735 22358
rect 9473 22134 9478 22162
rect 9506 22134 9814 22162
rect 9842 22134 9847 22162
rect 11377 22134 11382 22162
rect 11410 22134 12838 22162
rect 12866 22134 12950 22162
rect 12978 22134 12983 22162
rect 16137 22134 16142 22162
rect 16170 22134 16422 22162
rect 16450 22134 16870 22162
rect 16898 22134 16982 22162
rect 17010 22134 17015 22162
rect 9913 21938 9918 21966
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 10050 21938 10055 21966
rect 19600 21882 20000 21896
rect 9809 21854 9814 21882
rect 9842 21854 10038 21882
rect 10066 21854 11382 21882
rect 11410 21854 11415 21882
rect 16865 21854 16870 21882
rect 16898 21854 17486 21882
rect 17514 21854 17519 21882
rect 17817 21854 17822 21882
rect 17850 21854 18046 21882
rect 18074 21854 18158 21882
rect 18186 21854 18550 21882
rect 18578 21854 19054 21882
rect 19082 21854 20000 21882
rect 19600 21840 20000 21854
rect 11265 21798 11270 21826
rect 11298 21798 11494 21826
rect 11522 21798 11527 21826
rect 15857 21798 15862 21826
rect 15890 21798 16926 21826
rect 16954 21798 16959 21826
rect 2249 21742 2254 21770
rect 2282 21742 3038 21770
rect 3066 21742 4214 21770
rect 4242 21742 4247 21770
rect 10369 21742 10374 21770
rect 10402 21742 10598 21770
rect 10626 21742 11102 21770
rect 11130 21742 11135 21770
rect 17313 21742 17318 21770
rect 17346 21742 17598 21770
rect 17626 21742 17710 21770
rect 17738 21742 18382 21770
rect 18410 21742 18718 21770
rect 18746 21742 18751 21770
rect 2233 21546 2238 21574
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2370 21546 2375 21574
rect 17593 21546 17598 21574
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17730 21546 17735 21574
rect 2473 21294 2478 21322
rect 2506 21294 3038 21322
rect 3066 21294 3071 21322
rect 18377 21294 18382 21322
rect 18410 21294 18774 21322
rect 18802 21294 18807 21322
rect 16025 21238 16030 21266
rect 16058 21238 17990 21266
rect 18018 21238 18023 21266
rect 9913 21154 9918 21182
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 10050 21154 10055 21182
rect 17929 21070 17934 21098
rect 17962 21070 18214 21098
rect 18242 21070 18247 21098
rect 6057 21014 6062 21042
rect 6090 21014 7126 21042
rect 7154 21014 7159 21042
rect 7513 21014 7518 21042
rect 7546 21014 8582 21042
rect 8610 21014 8615 21042
rect 9529 21014 9534 21042
rect 9562 21014 11550 21042
rect 11578 21014 12726 21042
rect 12754 21014 13286 21042
rect 13314 21014 13510 21042
rect 13538 21014 13543 21042
rect 16977 21014 16982 21042
rect 17010 21014 17654 21042
rect 17682 21014 18102 21042
rect 18130 21014 18135 21042
rect 12553 20958 12558 20986
rect 12586 20958 13118 20986
rect 13146 20958 13151 20986
rect 18489 20958 18494 20986
rect 18522 20958 18998 20986
rect 19026 20958 19031 20986
rect 2233 20762 2238 20790
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2370 20762 2375 20790
rect 17593 20762 17598 20790
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17730 20762 17735 20790
rect 11097 20678 11102 20706
rect 11130 20678 12558 20706
rect 12586 20678 12591 20706
rect 18433 20566 18438 20594
rect 18466 20566 18774 20594
rect 18802 20566 18807 20594
rect 0 20538 400 20552
rect 0 20510 1806 20538
rect 1834 20510 1839 20538
rect 0 20496 400 20510
rect 9913 20370 9918 20398
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 10050 20370 10055 20398
rect 12553 20230 12558 20258
rect 12586 20230 13062 20258
rect 13090 20230 14630 20258
rect 14658 20230 14663 20258
rect 13113 20174 13118 20202
rect 13146 20174 14574 20202
rect 14602 20174 15078 20202
rect 15106 20174 15111 20202
rect 2233 19978 2238 20006
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2370 19978 2375 20006
rect 17593 19978 17598 20006
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17730 19978 17735 20006
rect 8577 19782 8582 19810
rect 8610 19782 9142 19810
rect 9170 19782 9175 19810
rect 11489 19782 11494 19810
rect 11522 19782 12726 19810
rect 12754 19782 12950 19810
rect 12978 19782 13566 19810
rect 13594 19782 13599 19810
rect 18097 19782 18102 19810
rect 18130 19782 18270 19810
rect 18298 19782 18494 19810
rect 18522 19782 18718 19810
rect 18746 19782 18751 19810
rect 18377 19726 18382 19754
rect 18410 19726 19054 19754
rect 19082 19726 19087 19754
rect 9913 19586 9918 19614
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 10050 19586 10055 19614
rect 19600 19586 20000 19600
rect 18993 19558 18998 19586
rect 19026 19558 20000 19586
rect 19600 19544 20000 19558
rect 9137 19390 9142 19418
rect 9170 19390 10598 19418
rect 10626 19390 10631 19418
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 3817 18998 3822 19026
rect 3850 18998 5278 19026
rect 5306 18998 5311 19026
rect 12777 18998 12782 19026
rect 12810 18998 16254 19026
rect 16282 18998 16287 19026
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 15241 18662 15246 18690
rect 15274 18662 16814 18690
rect 16842 18662 16847 18690
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 15073 18270 15078 18298
rect 15106 18270 16254 18298
rect 16282 18270 16814 18298
rect 16842 18270 16847 18298
rect 2473 18214 2478 18242
rect 2506 18214 3038 18242
rect 3066 18214 3071 18242
rect 7569 18214 7574 18242
rect 7602 18214 8750 18242
rect 8778 18214 8974 18242
rect 9002 18214 9310 18242
rect 9338 18214 9343 18242
rect 15913 18214 15918 18242
rect 15946 18214 16758 18242
rect 16786 18214 16926 18242
rect 16954 18214 17262 18242
rect 17290 18214 17295 18242
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 1857 17878 1862 17906
rect 1890 17878 3374 17906
rect 3402 17878 3407 17906
rect 3033 17822 3038 17850
rect 3066 17822 4438 17850
rect 4466 17822 4471 17850
rect 6393 17822 6398 17850
rect 6426 17822 7182 17850
rect 7210 17822 7215 17850
rect 10593 17822 10598 17850
rect 10626 17822 11102 17850
rect 11130 17822 11135 17850
rect 1577 17654 1582 17682
rect 1610 17654 1862 17682
rect 1890 17654 1895 17682
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 11097 17430 11102 17458
rect 11130 17430 12558 17458
rect 12586 17430 13118 17458
rect 13146 17430 13151 17458
rect 14849 17430 14854 17458
rect 14882 17430 16254 17458
rect 16282 17430 16287 17458
rect 19600 17290 20000 17304
rect 19049 17262 19054 17290
rect 19082 17262 20000 17290
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 19600 17248 20000 17262
rect 13113 17038 13118 17066
rect 13146 17038 14574 17066
rect 14602 17038 14607 17066
rect 0 16842 400 16856
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 0 16814 2086 16842
rect 2114 16814 2119 16842
rect 0 16800 400 16814
rect 11265 16646 11270 16674
rect 11298 16646 11494 16674
rect 11522 16646 11527 16674
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 7121 15974 7126 16002
rect 7154 15974 8414 16002
rect 8442 15974 8447 16002
rect 11321 15918 11326 15946
rect 11354 15918 12726 15946
rect 12754 15918 12950 15946
rect 12978 15918 13454 15946
rect 13482 15918 13487 15946
rect 14289 15862 14294 15890
rect 14322 15862 14798 15890
rect 14826 15862 14831 15890
rect 15185 15862 15190 15890
rect 15218 15862 16814 15890
rect 16842 15862 17206 15890
rect 17234 15862 17239 15890
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 15185 15526 15190 15554
rect 15218 15526 15302 15554
rect 15330 15526 15335 15554
rect 10929 15470 10934 15498
rect 10962 15470 14294 15498
rect 14322 15470 14327 15498
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 19600 14994 20000 15008
rect 19049 14966 19054 14994
rect 19082 14966 20000 14994
rect 19600 14952 20000 14966
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 2529 14294 2534 14322
rect 2562 14294 4382 14322
rect 4410 14294 5894 14322
rect 5922 14294 5927 14322
rect 14793 14294 14798 14322
rect 14826 14294 16534 14322
rect 16562 14294 16814 14322
rect 16842 14294 16847 14322
rect 8801 14238 8806 14266
rect 8834 14238 8974 14266
rect 9002 14238 9007 14266
rect 11713 14238 11718 14266
rect 11746 14238 13398 14266
rect 13426 14238 15190 14266
rect 15218 14238 15223 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9529 13902 9534 13930
rect 9562 13902 11494 13930
rect 11522 13902 11527 13930
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8857 13510 8862 13538
rect 8890 13510 10374 13538
rect 10402 13510 10822 13538
rect 10850 13510 10855 13538
rect 15465 13510 15470 13538
rect 15498 13510 16814 13538
rect 16842 13510 17262 13538
rect 17290 13510 17295 13538
rect 8801 13454 8806 13482
rect 8834 13454 8974 13482
rect 9002 13454 9007 13482
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 0 13146 400 13160
rect 0 13118 1694 13146
rect 1722 13118 4214 13146
rect 0 13104 400 13118
rect 4186 13034 4214 13118
rect 4186 13006 12782 13034
rect 12810 13006 12815 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 19600 12698 20000 12712
rect 19049 12670 19054 12698
rect 19082 12670 20000 12698
rect 19600 12656 20000 12670
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 2529 12334 2534 12362
rect 2562 12334 3766 12362
rect 3794 12334 3990 12362
rect 4018 12334 4158 12362
rect 4186 12334 4191 12362
rect 6337 12334 6342 12362
rect 6370 12334 10318 12362
rect 10346 12334 10934 12362
rect 10962 12334 10967 12362
rect 12833 12334 12838 12362
rect 12866 12334 14294 12362
rect 14322 12334 14327 12362
rect 8409 12278 8414 12306
rect 8442 12278 8862 12306
rect 8890 12278 8895 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 4097 11942 4102 11970
rect 4130 11942 4214 11970
rect 4242 11942 4247 11970
rect 14569 11942 14574 11970
rect 14602 11942 15078 11970
rect 15106 11942 16254 11970
rect 16282 11942 16287 11970
rect 6169 11774 6174 11802
rect 6202 11774 7574 11802
rect 7602 11774 7798 11802
rect 7826 11774 8750 11802
rect 8778 11774 8783 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 1857 11550 1862 11578
rect 1890 11550 3318 11578
rect 3346 11550 3351 11578
rect 11489 11550 11494 11578
rect 11522 11550 13398 11578
rect 13426 11550 15134 11578
rect 15162 11550 15246 11578
rect 15274 11550 15279 11578
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 4097 11158 4102 11186
rect 4130 11158 5054 11186
rect 5082 11158 5278 11186
rect 5306 11158 5311 11186
rect 3369 11102 3374 11130
rect 3402 11102 4214 11130
rect 4242 11102 4662 11130
rect 4690 11102 5222 11130
rect 5250 11102 5255 11130
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 12273 10766 12278 10794
rect 12306 10766 12838 10794
rect 12866 10766 12871 10794
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 19600 10402 20000 10416
rect 10817 10374 10822 10402
rect 10850 10374 12278 10402
rect 12306 10374 12311 10402
rect 16417 10374 16422 10402
rect 16450 10374 16926 10402
rect 16954 10374 17206 10402
rect 17234 10374 17486 10402
rect 17514 10374 18774 10402
rect 18802 10374 18807 10402
rect 18886 10374 20000 10402
rect 18886 10346 18914 10374
rect 19600 10360 20000 10374
rect 17145 10318 17150 10346
rect 17178 10318 18718 10346
rect 18746 10318 18914 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 10313 10094 10318 10122
rect 10346 10094 10822 10122
rect 10850 10094 10855 10122
rect 13561 10094 13566 10122
rect 13594 10094 13678 10122
rect 13706 10094 13711 10122
rect 3033 9982 3038 10010
rect 3066 9982 3766 10010
rect 3794 9982 3799 10010
rect 11041 9982 11046 10010
rect 11074 9982 13398 10010
rect 13426 9982 13510 10010
rect 13538 9982 13543 10010
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 8969 9590 8974 9618
rect 9002 9590 9254 9618
rect 9282 9590 9287 9618
rect 12553 9590 12558 9618
rect 12586 9590 12838 9618
rect 12866 9590 12871 9618
rect 16753 9590 16758 9618
rect 16786 9590 17150 9618
rect 17178 9590 17183 9618
rect 3313 9534 3318 9562
rect 3346 9534 6342 9562
rect 6370 9534 6375 9562
rect 15969 9534 15974 9562
rect 16002 9534 16254 9562
rect 16282 9534 16478 9562
rect 16506 9534 17766 9562
rect 17794 9534 18606 9562
rect 18634 9534 18639 9562
rect 0 9450 400 9464
rect 0 9422 910 9450
rect 938 9422 943 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 13337 9310 13342 9338
rect 13370 9310 13510 9338
rect 13538 9310 13543 9338
rect 1577 9254 1582 9282
rect 1610 9254 1918 9282
rect 1946 9254 3318 9282
rect 3346 9254 3351 9282
rect 3761 9254 3766 9282
rect 3794 9254 5110 9282
rect 5138 9254 5143 9282
rect 9529 9254 9534 9282
rect 9562 9254 10990 9282
rect 11018 9254 11270 9282
rect 11298 9254 11303 9282
rect 13393 9254 13398 9282
rect 13426 9254 14742 9282
rect 14770 9254 14775 9282
rect 9081 9198 9086 9226
rect 9114 9198 10318 9226
rect 10346 9198 10351 9226
rect 12833 9198 12838 9226
rect 12866 9198 14294 9226
rect 14322 9198 14327 9226
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 14289 8862 14294 8890
rect 14322 8862 14798 8890
rect 14826 8862 14831 8890
rect 10593 8806 10598 8834
rect 10626 8806 11102 8834
rect 11130 8806 14574 8834
rect 14602 8806 14607 8834
rect 15129 8806 15134 8834
rect 15162 8806 15246 8834
rect 15274 8806 15470 8834
rect 15498 8806 15503 8834
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 2081 8470 2086 8498
rect 2114 8470 4214 8498
rect 4186 8442 4214 8470
rect 2473 8414 2478 8442
rect 2506 8414 2814 8442
rect 2842 8414 3038 8442
rect 3066 8414 3654 8442
rect 3682 8414 3687 8442
rect 4186 8414 10598 8442
rect 10626 8414 10631 8442
rect 3593 8358 3598 8386
rect 3626 8358 4998 8386
rect 5026 8358 5031 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 19600 8106 20000 8120
rect 15185 8078 15190 8106
rect 15218 8078 15358 8106
rect 15386 8078 15391 8106
rect 17537 8078 17542 8106
rect 17570 8078 20000 8106
rect 19600 8064 20000 8078
rect 1577 8022 1582 8050
rect 1610 8022 1918 8050
rect 1946 8022 1951 8050
rect 14289 8022 14294 8050
rect 14322 8022 15694 8050
rect 15722 8022 15727 8050
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 1913 7630 1918 7658
rect 1946 7630 2142 7658
rect 2170 7630 3598 7658
rect 3626 7630 3631 7658
rect 10593 7630 10598 7658
rect 10626 7630 11102 7658
rect 11130 7630 11135 7658
rect 4993 7574 4998 7602
rect 5026 7574 6342 7602
rect 6370 7574 6375 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 1577 7238 1582 7266
rect 1610 7238 2086 7266
rect 2114 7238 2119 7266
rect 7513 7238 7518 7266
rect 7546 7238 8750 7266
rect 8778 7238 8974 7266
rect 9002 7238 9007 7266
rect 15241 7238 15246 7266
rect 15274 7238 15470 7266
rect 15498 7238 15918 7266
rect 15946 7210 15974 7266
rect 15946 7182 16254 7210
rect 16282 7182 16287 7210
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 3985 6734 3990 6762
rect 4018 6734 5558 6762
rect 5586 6734 5591 6762
rect 11265 6734 11270 6762
rect 11298 6734 12278 6762
rect 12306 6734 12838 6762
rect 12866 6734 14294 6762
rect 14322 6734 14798 6762
rect 14826 6734 14831 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9809 6510 9814 6538
rect 9842 6510 11102 6538
rect 11130 6510 11135 6538
rect 11993 6510 11998 6538
rect 12026 6510 12446 6538
rect 12474 6510 13398 6538
rect 13426 6510 14014 6538
rect 14042 6510 15246 6538
rect 15274 6510 15358 6538
rect 15386 6510 15391 6538
rect 14569 6454 14574 6482
rect 14602 6454 14910 6482
rect 14938 6454 15694 6482
rect 15722 6454 17150 6482
rect 17178 6454 17183 6482
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 5553 6062 5558 6090
rect 5586 6062 6790 6090
rect 6818 6062 6823 6090
rect 10425 5894 10430 5922
rect 10458 5894 10990 5922
rect 11018 5894 11998 5922
rect 12026 5894 12031 5922
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 19600 5810 20000 5824
rect 17817 5782 17822 5810
rect 17850 5782 20000 5810
rect 19600 5768 20000 5782
rect 0 5754 400 5768
rect 0 5726 966 5754
rect 994 5726 999 5754
rect 0 5712 400 5726
rect 2417 5670 2422 5698
rect 2450 5670 3374 5698
rect 3402 5670 3407 5698
rect 8969 5670 8974 5698
rect 9002 5670 9534 5698
rect 9562 5670 9814 5698
rect 9842 5670 9847 5698
rect 15465 5614 15470 5642
rect 15498 5614 15918 5642
rect 15946 5614 15974 5642
rect 16002 5614 16254 5642
rect 16282 5614 16287 5642
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 1577 5166 1582 5194
rect 1610 5166 2870 5194
rect 2898 5166 2903 5194
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 12553 4998 12558 5026
rect 12586 4998 13118 5026
rect 13146 4998 14574 5026
rect 14602 4998 14607 5026
rect 3537 4886 3542 4914
rect 3570 4886 5166 4914
rect 5194 4886 5390 4914
rect 5418 4886 5423 4914
rect 11993 4886 11998 4914
rect 12026 4886 12278 4914
rect 12306 4886 12311 4914
rect 13393 4886 13398 4914
rect 13426 4886 14014 4914
rect 14042 4886 14047 4914
rect 14569 4886 14574 4914
rect 14602 4886 15918 4914
rect 15946 4886 17150 4914
rect 17178 4886 17183 4914
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2025 4494 2030 4522
rect 2058 4494 3374 4522
rect 3402 4494 3407 4522
rect 7009 4494 7014 4522
rect 7042 4494 7518 4522
rect 7546 4494 7551 4522
rect 17537 4494 17542 4522
rect 17570 4494 18382 4522
rect 18410 4494 18774 4522
rect 18802 4494 18807 4522
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 16473 4214 16478 4242
rect 16506 4214 17990 4242
rect 18018 4214 18023 4242
rect 5777 4158 5782 4186
rect 5810 4158 6006 4186
rect 6034 4158 6566 4186
rect 6594 4158 6599 4186
rect 13337 4158 13342 4186
rect 13370 4158 14742 4186
rect 14770 4158 14775 4186
rect 5782 4130 5810 4158
rect 4041 4102 4046 4130
rect 4074 4102 5810 4130
rect 6449 4102 6454 4130
rect 6482 4102 7014 4130
rect 7042 4102 7047 4130
rect 17873 4102 17878 4130
rect 17906 4102 18438 4130
rect 18466 4102 18471 4130
rect 10033 4046 10038 4074
rect 10066 4046 11102 4074
rect 11130 4046 11550 4074
rect 11578 4046 12222 4074
rect 12250 4046 18214 4074
rect 18242 4046 18247 4074
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 3817 3710 3822 3738
rect 3850 3710 4046 3738
rect 4074 3710 4079 3738
rect 11097 3710 11102 3738
rect 11130 3710 11550 3738
rect 11578 3710 12558 3738
rect 12586 3710 12591 3738
rect 13113 3710 13118 3738
rect 13146 3710 14518 3738
rect 14546 3710 14551 3738
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 19600 3514 20000 3528
rect 17766 3486 20000 3514
rect 17766 3458 17794 3486
rect 19600 3472 20000 3486
rect 16753 3430 16758 3458
rect 16786 3430 17486 3458
rect 17514 3430 17794 3458
rect 7009 3374 7014 3402
rect 7042 3374 7518 3402
rect 7546 3374 7551 3402
rect 12441 3374 12446 3402
rect 12474 3374 12479 3402
rect 12553 3374 12558 3402
rect 12586 3374 13118 3402
rect 13146 3374 13151 3402
rect 12446 3346 12474 3374
rect 4489 3318 4494 3346
rect 4522 3318 4998 3346
rect 5026 3318 5558 3346
rect 5586 3318 5591 3346
rect 7793 3318 7798 3346
rect 7826 3318 9254 3346
rect 9282 3318 9287 3346
rect 12446 3318 13230 3346
rect 13258 3318 13263 3346
rect 17817 3318 17822 3346
rect 17850 3318 18382 3346
rect 18410 3318 18774 3346
rect 18802 3318 18807 3346
rect 11489 3262 11494 3290
rect 11522 3262 12726 3290
rect 12754 3262 12950 3290
rect 12978 3262 13286 3290
rect 13314 3262 13319 3290
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 5889 2926 5894 2954
rect 5922 2926 6286 2954
rect 6314 2926 6510 2954
rect 6538 2926 7630 2954
rect 7658 2926 7966 2954
rect 7994 2926 8246 2954
rect 8274 2926 8279 2954
rect 9305 2926 9310 2954
rect 9338 2926 11046 2954
rect 11074 2926 11079 2954
rect 13225 2926 13230 2954
rect 13258 2926 13454 2954
rect 13482 2926 14014 2954
rect 14042 2926 15358 2954
rect 15386 2926 15391 2954
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 4186 2590 5894 2618
rect 5922 2590 5927 2618
rect 4186 2562 4214 2590
rect 3985 2534 3990 2562
rect 4018 2534 4214 2562
rect 5553 2534 5558 2562
rect 5586 2534 6118 2562
rect 6146 2534 6151 2562
rect 8241 2534 8246 2562
rect 8274 2534 8470 2562
rect 8498 2534 8503 2562
rect 16921 2534 16926 2562
rect 16954 2534 18774 2562
rect 18802 2534 18807 2562
rect 6561 2478 6566 2506
rect 6594 2478 7014 2506
rect 7042 2478 8358 2506
rect 8386 2478 8806 2506
rect 8834 2478 10430 2506
rect 10458 2478 10463 2506
rect 14345 2478 14350 2506
rect 14378 2478 14798 2506
rect 14826 2478 14831 2506
rect 8465 2422 8470 2450
rect 8498 2422 9590 2450
rect 9618 2422 9758 2450
rect 9786 2422 9791 2450
rect 13617 2422 13622 2450
rect 13650 2422 15246 2450
rect 15274 2422 15470 2450
rect 15498 2422 15503 2450
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 10873 2254 10878 2282
rect 10906 2254 11606 2282
rect 11634 2254 12558 2282
rect 12586 2254 12591 2282
rect 4186 2198 14350 2226
rect 14378 2198 14383 2226
rect 4186 2170 4214 2198
rect 462 2142 4214 2170
rect 4489 2142 4494 2170
rect 4522 2142 4998 2170
rect 5026 2142 5031 2170
rect 7513 2142 7518 2170
rect 7546 2142 8078 2170
rect 8106 2142 8111 2170
rect 10425 2142 10430 2170
rect 10458 2142 11662 2170
rect 11690 2142 11695 2170
rect 0 2058 400 2072
rect 462 2058 490 2142
rect 9585 2086 9590 2114
rect 9618 2086 11158 2114
rect 11186 2086 11382 2114
rect 11410 2086 11415 2114
rect 0 2030 490 2058
rect 1689 2030 1694 2058
rect 1722 2030 14294 2058
rect 14322 2030 15526 2058
rect 15554 2030 15559 2058
rect 0 2016 400 2030
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 961 1806 966 1834
rect 994 1806 2870 1834
rect 2898 1806 12670 1834
rect 12698 1806 12838 1834
rect 12866 1806 12871 1834
rect 2081 1750 2086 1778
rect 2114 1750 3822 1778
rect 3850 1750 3855 1778
rect 6113 1750 6118 1778
rect 6146 1750 7462 1778
rect 7490 1750 8302 1778
rect 8330 1750 8335 1778
rect 9417 1750 9422 1778
rect 9450 1750 10878 1778
rect 10906 1750 10911 1778
rect 9422 1722 9450 1750
rect 8073 1694 8078 1722
rect 8106 1694 9450 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
rect 19600 1218 20000 1232
rect 18769 1190 18774 1218
rect 18802 1190 20000 1218
rect 19600 1176 20000 1190
<< via3 >>
rect 9918 28210 9946 28238
rect 9970 28210 9998 28238
rect 10022 28210 10050 28238
rect 2238 27818 2266 27846
rect 2290 27818 2318 27846
rect 2342 27818 2370 27846
rect 17598 27818 17626 27846
rect 17650 27818 17678 27846
rect 17702 27818 17730 27846
rect 9918 27426 9946 27454
rect 9970 27426 9998 27454
rect 10022 27426 10050 27454
rect 2238 27034 2266 27062
rect 2290 27034 2318 27062
rect 2342 27034 2370 27062
rect 17598 27034 17626 27062
rect 17650 27034 17678 27062
rect 17702 27034 17730 27062
rect 9918 26642 9946 26670
rect 9970 26642 9998 26670
rect 10022 26642 10050 26670
rect 2238 26250 2266 26278
rect 2290 26250 2318 26278
rect 2342 26250 2370 26278
rect 17598 26250 17626 26278
rect 17650 26250 17678 26278
rect 17702 26250 17730 26278
rect 9918 25858 9946 25886
rect 9970 25858 9998 25886
rect 10022 25858 10050 25886
rect 2238 25466 2266 25494
rect 2290 25466 2318 25494
rect 2342 25466 2370 25494
rect 17598 25466 17626 25494
rect 17650 25466 17678 25494
rect 17702 25466 17730 25494
rect 9918 25074 9946 25102
rect 9970 25074 9998 25102
rect 10022 25074 10050 25102
rect 2238 24682 2266 24710
rect 2290 24682 2318 24710
rect 2342 24682 2370 24710
rect 17598 24682 17626 24710
rect 17650 24682 17678 24710
rect 17702 24682 17730 24710
rect 9918 24290 9946 24318
rect 9970 24290 9998 24318
rect 10022 24290 10050 24318
rect 2238 23898 2266 23926
rect 2290 23898 2318 23926
rect 2342 23898 2370 23926
rect 17598 23898 17626 23926
rect 17650 23898 17678 23926
rect 17702 23898 17730 23926
rect 9918 23506 9946 23534
rect 9970 23506 9998 23534
rect 10022 23506 10050 23534
rect 2238 23114 2266 23142
rect 2290 23114 2318 23142
rect 2342 23114 2370 23142
rect 17598 23114 17626 23142
rect 17650 23114 17678 23142
rect 17702 23114 17730 23142
rect 9918 22722 9946 22750
rect 9970 22722 9998 22750
rect 10022 22722 10050 22750
rect 2238 22330 2266 22358
rect 2290 22330 2318 22358
rect 2342 22330 2370 22358
rect 17598 22330 17626 22358
rect 17650 22330 17678 22358
rect 17702 22330 17730 22358
rect 9918 21938 9946 21966
rect 9970 21938 9998 21966
rect 10022 21938 10050 21966
rect 2238 21546 2266 21574
rect 2290 21546 2318 21574
rect 2342 21546 2370 21574
rect 17598 21546 17626 21574
rect 17650 21546 17678 21574
rect 17702 21546 17730 21574
rect 9918 21154 9946 21182
rect 9970 21154 9998 21182
rect 10022 21154 10050 21182
rect 2238 20762 2266 20790
rect 2290 20762 2318 20790
rect 2342 20762 2370 20790
rect 17598 20762 17626 20790
rect 17650 20762 17678 20790
rect 17702 20762 17730 20790
rect 9918 20370 9946 20398
rect 9970 20370 9998 20398
rect 10022 20370 10050 20398
rect 2238 19978 2266 20006
rect 2290 19978 2318 20006
rect 2342 19978 2370 20006
rect 17598 19978 17626 20006
rect 17650 19978 17678 20006
rect 17702 19978 17730 20006
rect 9918 19586 9946 19614
rect 9970 19586 9998 19614
rect 10022 19586 10050 19614
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 17822 5782 17850 5810
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 17822 3318 17850 3346
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 27846 2384 28254
rect 2224 27818 2238 27846
rect 2266 27818 2290 27846
rect 2318 27818 2342 27846
rect 2370 27818 2384 27846
rect 2224 27062 2384 27818
rect 2224 27034 2238 27062
rect 2266 27034 2290 27062
rect 2318 27034 2342 27062
rect 2370 27034 2384 27062
rect 2224 26278 2384 27034
rect 2224 26250 2238 26278
rect 2266 26250 2290 26278
rect 2318 26250 2342 26278
rect 2370 26250 2384 26278
rect 2224 25494 2384 26250
rect 2224 25466 2238 25494
rect 2266 25466 2290 25494
rect 2318 25466 2342 25494
rect 2370 25466 2384 25494
rect 2224 24710 2384 25466
rect 2224 24682 2238 24710
rect 2266 24682 2290 24710
rect 2318 24682 2342 24710
rect 2370 24682 2384 24710
rect 2224 23926 2384 24682
rect 2224 23898 2238 23926
rect 2266 23898 2290 23926
rect 2318 23898 2342 23926
rect 2370 23898 2384 23926
rect 2224 23142 2384 23898
rect 2224 23114 2238 23142
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2370 23114 2384 23142
rect 2224 22358 2384 23114
rect 2224 22330 2238 22358
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2370 22330 2384 22358
rect 2224 21574 2384 22330
rect 2224 21546 2238 21574
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2370 21546 2384 21574
rect 2224 20790 2384 21546
rect 2224 20762 2238 20790
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2370 20762 2384 20790
rect 2224 20006 2384 20762
rect 2224 19978 2238 20006
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2370 19978 2384 20006
rect 2224 19222 2384 19978
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 28238 10064 28254
rect 9904 28210 9918 28238
rect 9946 28210 9970 28238
rect 9998 28210 10022 28238
rect 10050 28210 10064 28238
rect 9904 27454 10064 28210
rect 9904 27426 9918 27454
rect 9946 27426 9970 27454
rect 9998 27426 10022 27454
rect 10050 27426 10064 27454
rect 9904 26670 10064 27426
rect 9904 26642 9918 26670
rect 9946 26642 9970 26670
rect 9998 26642 10022 26670
rect 10050 26642 10064 26670
rect 9904 25886 10064 26642
rect 9904 25858 9918 25886
rect 9946 25858 9970 25886
rect 9998 25858 10022 25886
rect 10050 25858 10064 25886
rect 9904 25102 10064 25858
rect 9904 25074 9918 25102
rect 9946 25074 9970 25102
rect 9998 25074 10022 25102
rect 10050 25074 10064 25102
rect 9904 24318 10064 25074
rect 9904 24290 9918 24318
rect 9946 24290 9970 24318
rect 9998 24290 10022 24318
rect 10050 24290 10064 24318
rect 9904 23534 10064 24290
rect 9904 23506 9918 23534
rect 9946 23506 9970 23534
rect 9998 23506 10022 23534
rect 10050 23506 10064 23534
rect 9904 22750 10064 23506
rect 9904 22722 9918 22750
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 10050 22722 10064 22750
rect 9904 21966 10064 22722
rect 9904 21938 9918 21966
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 10050 21938 10064 21966
rect 9904 21182 10064 21938
rect 9904 21154 9918 21182
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 10050 21154 10064 21182
rect 9904 20398 10064 21154
rect 9904 20370 9918 20398
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 10050 20370 10064 20398
rect 9904 19614 10064 20370
rect 9904 19586 9918 19614
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 10050 19586 10064 19614
rect 9904 18830 10064 19586
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 27846 17744 28254
rect 17584 27818 17598 27846
rect 17626 27818 17650 27846
rect 17678 27818 17702 27846
rect 17730 27818 17744 27846
rect 17584 27062 17744 27818
rect 17584 27034 17598 27062
rect 17626 27034 17650 27062
rect 17678 27034 17702 27062
rect 17730 27034 17744 27062
rect 17584 26278 17744 27034
rect 17584 26250 17598 26278
rect 17626 26250 17650 26278
rect 17678 26250 17702 26278
rect 17730 26250 17744 26278
rect 17584 25494 17744 26250
rect 17584 25466 17598 25494
rect 17626 25466 17650 25494
rect 17678 25466 17702 25494
rect 17730 25466 17744 25494
rect 17584 24710 17744 25466
rect 17584 24682 17598 24710
rect 17626 24682 17650 24710
rect 17678 24682 17702 24710
rect 17730 24682 17744 24710
rect 17584 23926 17744 24682
rect 17584 23898 17598 23926
rect 17626 23898 17650 23926
rect 17678 23898 17702 23926
rect 17730 23898 17744 23926
rect 17584 23142 17744 23898
rect 17584 23114 17598 23142
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17730 23114 17744 23142
rect 17584 22358 17744 23114
rect 17584 22330 17598 22358
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17730 22330 17744 22358
rect 17584 21574 17744 22330
rect 17584 21546 17598 21574
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17730 21546 17744 21574
rect 17584 20790 17744 21546
rect 17584 20762 17598 20790
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17730 20762 17744 20790
rect 17584 20006 17744 20762
rect 17584 19978 17598 20006
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17730 19978 17744 20006
rect 17584 19222 17744 19978
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17822 5810 17850 5815
rect 17822 3346 17850 5782
rect 17822 3313 17850 3318
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2184 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62
timestamp 1667941163
transform 1 0 4144 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1667941163
transform 1 0 6664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 8456 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142
timestamp 1667941163
transform 1 0 8624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 10416 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 10584 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_202
timestamp 1667941163
transform 1 0 11984 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1667941163
transform 1 0 12544 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_237
timestamp 1667941163
transform 1 0 13944 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1667941163
transform 1 0 14504 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_272
timestamp 1667941163
transform 1 0 15904 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 16464 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1667941163
transform 1 0 18256 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_317
timestamp 1667941163
transform 1 0 18424 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_325 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 18872 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 19096 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1667941163
transform 1 0 784 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_27 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2184 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_43
timestamp 1667941163
transform 1 0 3080 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_45
timestamp 1667941163
transform 1 0 3192 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_89
timestamp 1667941163
transform 1 0 5656 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_115
timestamp 1667941163
transform 1 0 7112 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 8568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_144
timestamp 1667941163
transform 1 0 8736 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_176
timestamp 1667941163
transform 1 0 10528 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_202
timestamp 1667941163
transform 1 0 11984 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_210
timestamp 1667941163
transform 1 0 12432 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 12544 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1667941163
transform 1 0 12712 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_240
timestamp 1667941163
transform 1 0 14112 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_266
timestamp 1667941163
transform 1 0 15568 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_282
timestamp 1667941163
transform 1 0 16464 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_286
timestamp 1667941163
transform 1 0 16688 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_302
timestamp 1667941163
transform 1 0 17584 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_330
timestamp 1667941163
transform 1 0 19152 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_27
timestamp 1667941163
transform 1 0 2184 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_53
timestamp 1667941163
transform 1 0 3640 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_79
timestamp 1667941163
transform 1 0 5096 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_108
timestamp 1667941163
transform 1 0 6720 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_124
timestamp 1667941163
transform 1 0 7616 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_150
timestamp 1667941163
transform 1 0 9072 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 10528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1667941163
transform 1 0 10696 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_204
timestamp 1667941163
transform 1 0 12096 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_230
timestamp 1667941163
transform 1 0 13552 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_246
timestamp 1667941163
transform 1 0 14448 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1667941163
transform 1 0 14672 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_275
timestamp 1667941163
transform 1 0 16072 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_291
timestamp 1667941163
transform 1 0 16968 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_293
timestamp 1667941163
transform 1 0 17080 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1667941163
transform 1 0 18480 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_321
timestamp 1667941163
transform 1 0 18648 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_329
timestamp 1667941163
transform 1 0 19096 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_27
timestamp 1667941163
transform 1 0 2184 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_43
timestamp 1667941163
transform 1 0 3080 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_45
timestamp 1667941163
transform 1 0 3192 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_89
timestamp 1667941163
transform 1 0 5656 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_115
timestamp 1667941163
transform 1 0 7112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 8568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_144
timestamp 1667941163
transform 1 0 8736 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_152
timestamp 1667941163
transform 1 0 9184 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_177
timestamp 1667941163
transform 1 0 10584 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_203
timestamp 1667941163
transform 1 0 12040 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_211
timestamp 1667941163
transform 1 0 12488 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1667941163
transform 1 0 12712 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_240
timestamp 1667941163
transform 1 0 14112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_266
timestamp 1667941163
transform 1 0 15568 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1667941163
transform 1 0 16464 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_286
timestamp 1667941163
transform 1 0 16688 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_302
timestamp 1667941163
transform 1 0 17584 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_330
timestamp 1667941163
transform 1 0 19152 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_27
timestamp 1667941163
transform 1 0 2184 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_53
timestamp 1667941163
transform 1 0 3640 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_79
timestamp 1667941163
transform 1 0 5096 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_108
timestamp 1667941163
transform 1 0 6720 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_124
timestamp 1667941163
transform 1 0 7616 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_150
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 10528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1667941163
transform 1 0 10696 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_204
timestamp 1667941163
transform 1 0 12096 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_230
timestamp 1667941163
transform 1 0 13552 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1667941163
transform 1 0 14448 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_250
timestamp 1667941163
transform 1 0 14672 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_266
timestamp 1667941163
transform 1 0 15568 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_292
timestamp 1667941163
transform 1 0 17024 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1667941163
transform 1 0 18480 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_321
timestamp 1667941163
transform 1 0 18648 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_329
timestamp 1667941163
transform 1 0 19096 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_27
timestamp 1667941163
transform 1 0 2184 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_43
timestamp 1667941163
transform 1 0 3080 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_45
timestamp 1667941163
transform 1 0 3192 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_89
timestamp 1667941163
transform 1 0 5656 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_115
timestamp 1667941163
transform 1 0 7112 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 8568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_144
timestamp 1667941163
transform 1 0 8736 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_160
timestamp 1667941163
transform 1 0 9632 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_186
timestamp 1667941163
transform 1 0 11088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1667941163
transform 1 0 12544 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1667941163
transform 1 0 12712 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_240
timestamp 1667941163
transform 1 0 14112 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_266
timestamp 1667941163
transform 1 0 15568 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1667941163
transform 1 0 16464 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_286
timestamp 1667941163
transform 1 0 16688 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_302
timestamp 1667941163
transform 1 0 17584 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_330
timestamp 1667941163
transform 1 0 19152 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_27
timestamp 1667941163
transform 1 0 2184 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_53
timestamp 1667941163
transform 1 0 3640 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_79
timestamp 1667941163
transform 1 0 5096 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 6552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_108
timestamp 1667941163
transform 1 0 6720 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_124
timestamp 1667941163
transform 1 0 7616 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_150
timestamp 1667941163
transform 1 0 9072 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 10528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_179
timestamp 1667941163
transform 1 0 10696 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_204
timestamp 1667941163
transform 1 0 12096 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_230
timestamp 1667941163
transform 1 0 13552 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_246
timestamp 1667941163
transform 1 0 14448 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_250
timestamp 1667941163
transform 1 0 14672 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_266
timestamp 1667941163
transform 1 0 15568 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_292
timestamp 1667941163
transform 1 0 17024 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1667941163
transform 1 0 18480 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_321
timestamp 1667941163
transform 1 0 18648 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_329
timestamp 1667941163
transform 1 0 19096 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_2
timestamp 1667941163
transform 1 0 784 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_10
timestamp 1667941163
transform 1 0 1232 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_36
timestamp 1667941163
transform 1 0 2688 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_62
timestamp 1667941163
transform 1 0 4144 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 4592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1667941163
transform 1 0 4760 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_89
timestamp 1667941163
transform 1 0 5656 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_115
timestamp 1667941163
transform 1 0 7112 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 8568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_144
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1667941163
transform 1 0 9632 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_186
timestamp 1667941163
transform 1 0 11088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1667941163
transform 1 0 12544 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_215
timestamp 1667941163
transform 1 0 12712 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_240
timestamp 1667941163
transform 1 0 14112 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_266
timestamp 1667941163
transform 1 0 15568 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_282
timestamp 1667941163
transform 1 0 16464 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_286
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_302
timestamp 1667941163
transform 1 0 17584 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_330
timestamp 1667941163
transform 1 0 19152 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_2
timestamp 1667941163
transform 1 0 784 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1667941163
transform 1 0 2744 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_62
timestamp 1667941163
transform 1 0 4144 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_70
timestamp 1667941163
transform 1 0 4592 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_95
timestamp 1667941163
transform 1 0 5992 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1667941163
transform 1 0 6440 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 6552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_108
timestamp 1667941163
transform 1 0 6720 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_124
timestamp 1667941163
transform 1 0 7616 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_150
timestamp 1667941163
transform 1 0 9072 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 10528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_179
timestamp 1667941163
transform 1 0 10696 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_204
timestamp 1667941163
transform 1 0 12096 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_230
timestamp 1667941163
transform 1 0 13552 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_246
timestamp 1667941163
transform 1 0 14448 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1667941163
transform 1 0 14672 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_275
timestamp 1667941163
transform 1 0 16072 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_291
timestamp 1667941163
transform 1 0 16968 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_293
timestamp 1667941163
transform 1 0 17080 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1667941163
transform 1 0 18480 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_321
timestamp 1667941163
transform 1 0 18648 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_329
timestamp 1667941163
transform 1 0 19096 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_2
timestamp 1667941163
transform 1 0 784 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_10
timestamp 1667941163
transform 1 0 1232 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_36
timestamp 1667941163
transform 1 0 2688 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_62
timestamp 1667941163
transform 1 0 4144 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 4592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_73
timestamp 1667941163
transform 1 0 4760 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_98
timestamp 1667941163
transform 1 0 6160 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_114
timestamp 1667941163
transform 1 0 7056 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_116
timestamp 1667941163
transform 1 0 7168 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 8568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_144
timestamp 1667941163
transform 1 0 8736 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_160
timestamp 1667941163
transform 1 0 9632 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_186
timestamp 1667941163
transform 1 0 11088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1667941163
transform 1 0 12544 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1667941163
transform 1 0 12712 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_240
timestamp 1667941163
transform 1 0 14112 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_266
timestamp 1667941163
transform 1 0 15568 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_282
timestamp 1667941163
transform 1 0 16464 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_286
timestamp 1667941163
transform 1 0 16688 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_302
timestamp 1667941163
transform 1 0 17584 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_330
timestamp 1667941163
transform 1 0 19152 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1667941163
transform 1 0 784 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 2576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1667941163
transform 1 0 2744 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_62
timestamp 1667941163
transform 1 0 4144 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_70
timestamp 1667941163
transform 1 0 4592 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_95
timestamp 1667941163
transform 1 0 5992 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_103
timestamp 1667941163
transform 1 0 6440 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 6552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_108
timestamp 1667941163
transform 1 0 6720 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_124
timestamp 1667941163
transform 1 0 7616 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_150
timestamp 1667941163
transform 1 0 9072 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 10528 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1667941163
transform 1 0 10696 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_204
timestamp 1667941163
transform 1 0 12096 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_230
timestamp 1667941163
transform 1 0 13552 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_246
timestamp 1667941163
transform 1 0 14448 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1667941163
transform 1 0 14672 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_275
timestamp 1667941163
transform 1 0 16072 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_301
timestamp 1667941163
transform 1 0 17528 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_317
timestamp 1667941163
transform 1 0 18424 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_321
timestamp 1667941163
transform 1 0 18648 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_329
timestamp 1667941163
transform 1 0 19096 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_2
timestamp 1667941163
transform 1 0 784 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_10
timestamp 1667941163
transform 1 0 1232 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_36
timestamp 1667941163
transform 1 0 2688 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_44
timestamp 1667941163
transform 1 0 3136 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 4592 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_73
timestamp 1667941163
transform 1 0 4760 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_98
timestamp 1667941163
transform 1 0 6160 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_124
timestamp 1667941163
transform 1 0 7616 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_140
timestamp 1667941163
transform 1 0 8512 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_144
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_160
timestamp 1667941163
transform 1 0 9632 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_186
timestamp 1667941163
transform 1 0 11088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1667941163
transform 1 0 12544 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1667941163
transform 1 0 12712 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_240
timestamp 1667941163
transform 1 0 14112 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_266
timestamp 1667941163
transform 1 0 15568 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1667941163
transform 1 0 16464 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_286
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_302
timestamp 1667941163
transform 1 0 17584 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_330
timestamp 1667941163
transform 1 0 19152 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_2
timestamp 1667941163
transform 1 0 784 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 2576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_37
timestamp 1667941163
transform 1 0 2744 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_69
timestamp 1667941163
transform 1 0 4536 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_95
timestamp 1667941163
transform 1 0 5992 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_103
timestamp 1667941163
transform 1 0 6440 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 6552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_108
timestamp 1667941163
transform 1 0 6720 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_133
timestamp 1667941163
transform 1 0 8120 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_149
timestamp 1667941163
transform 1 0 9016 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_151
timestamp 1667941163
transform 1 0 9128 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 10528 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1667941163
transform 1 0 10696 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_204
timestamp 1667941163
transform 1 0 12096 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_230
timestamp 1667941163
transform 1 0 13552 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_246
timestamp 1667941163
transform 1 0 14448 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1667941163
transform 1 0 14672 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_275
timestamp 1667941163
transform 1 0 16072 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_291
timestamp 1667941163
transform 1 0 16968 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_293
timestamp 1667941163
transform 1 0 17080 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1667941163
transform 1 0 18480 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_321
timestamp 1667941163
transform 1 0 18648 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_329
timestamp 1667941163
transform 1 0 19096 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1667941163
transform 1 0 784 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_18
timestamp 1667941163
transform 1 0 1680 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_44
timestamp 1667941163
transform 1 0 3136 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 4592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1667941163
transform 1 0 4760 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_98
timestamp 1667941163
transform 1 0 6160 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_124
timestamp 1667941163
transform 1 0 7616 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_140
timestamp 1667941163
transform 1 0 8512 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_144
timestamp 1667941163
transform 1 0 8736 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_160
timestamp 1667941163
transform 1 0 9632 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_186
timestamp 1667941163
transform 1 0 11088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 12544 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1667941163
transform 1 0 12712 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_240
timestamp 1667941163
transform 1 0 14112 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_266
timestamp 1667941163
transform 1 0 15568 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_282
timestamp 1667941163
transform 1 0 16464 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_286
timestamp 1667941163
transform 1 0 16688 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_302
timestamp 1667941163
transform 1 0 17584 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_330
timestamp 1667941163
transform 1 0 19152 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1667941163
transform 1 0 784 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 2576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_37
timestamp 1667941163
transform 1 0 2744 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_69
timestamp 1667941163
transform 1 0 4536 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_95
timestamp 1667941163
transform 1 0 5992 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_103
timestamp 1667941163
transform 1 0 6440 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 6552 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_108
timestamp 1667941163
transform 1 0 6720 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_133
timestamp 1667941163
transform 1 0 8120 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_159
timestamp 1667941163
transform 1 0 9576 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_175
timestamp 1667941163
transform 1 0 10472 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1667941163
transform 1 0 10696 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_204
timestamp 1667941163
transform 1 0 12096 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_230
timestamp 1667941163
transform 1 0 13552 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_246
timestamp 1667941163
transform 1 0 14448 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1667941163
transform 1 0 14672 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_275
timestamp 1667941163
transform 1 0 16072 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_301
timestamp 1667941163
transform 1 0 17528 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_317
timestamp 1667941163
transform 1 0 18424 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_321
timestamp 1667941163
transform 1 0 18648 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_329
timestamp 1667941163
transform 1 0 19096 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_2
timestamp 1667941163
transform 1 0 784 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_18
timestamp 1667941163
transform 1 0 1680 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_44
timestamp 1667941163
transform 1 0 3136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 4592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_73
timestamp 1667941163
transform 1 0 4760 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_98
timestamp 1667941163
transform 1 0 6160 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_124
timestamp 1667941163
transform 1 0 7616 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_140
timestamp 1667941163
transform 1 0 8512 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_144
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 10136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_195
timestamp 1667941163
transform 1 0 11592 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_211
timestamp 1667941163
transform 1 0 12488 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_215
timestamp 1667941163
transform 1 0 12712 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_240
timestamp 1667941163
transform 1 0 14112 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_266
timestamp 1667941163
transform 1 0 15568 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_282
timestamp 1667941163
transform 1 0 16464 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_286
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_302
timestamp 1667941163
transform 1 0 17584 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_330
timestamp 1667941163
transform 1 0 19152 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_2
timestamp 1667941163
transform 1 0 784 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1667941163
transform 1 0 2576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_37
timestamp 1667941163
transform 1 0 2744 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_41
timestamp 1667941163
transform 1 0 2968 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_66
timestamp 1667941163
transform 1 0 4368 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_70
timestamp 1667941163
transform 1 0 4592 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_95
timestamp 1667941163
transform 1 0 5992 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_103
timestamp 1667941163
transform 1 0 6440 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1667941163
transform 1 0 6552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1667941163
transform 1 0 6720 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_133
timestamp 1667941163
transform 1 0 8120 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_159
timestamp 1667941163
transform 1 0 9576 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_175
timestamp 1667941163
transform 1 0 10472 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_179
timestamp 1667941163
transform 1 0 10696 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_204
timestamp 1667941163
transform 1 0 12096 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_230
timestamp 1667941163
transform 1 0 13552 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_246
timestamp 1667941163
transform 1 0 14448 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1667941163
transform 1 0 14672 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_275
timestamp 1667941163
transform 1 0 16072 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_291
timestamp 1667941163
transform 1 0 16968 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_293
timestamp 1667941163
transform 1 0 17080 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1667941163
transform 1 0 18480 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_321
timestamp 1667941163
transform 1 0 18648 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_329
timestamp 1667941163
transform 1 0 19096 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_2
timestamp 1667941163
transform 1 0 784 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_10
timestamp 1667941163
transform 1 0 1232 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_14
timestamp 1667941163
transform 1 0 1456 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_40
timestamp 1667941163
transform 1 0 2912 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1667941163
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1667941163
transform 1 0 4592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_73
timestamp 1667941163
transform 1 0 4760 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_98
timestamp 1667941163
transform 1 0 6160 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_124
timestamp 1667941163
transform 1 0 7616 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_140
timestamp 1667941163
transform 1 0 8512 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1667941163
transform 1 0 8736 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 10136 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_195
timestamp 1667941163
transform 1 0 11592 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_211
timestamp 1667941163
transform 1 0 12488 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1667941163
transform 1 0 12712 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_240
timestamp 1667941163
transform 1 0 14112 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_266
timestamp 1667941163
transform 1 0 15568 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_282
timestamp 1667941163
transform 1 0 16464 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_286
timestamp 1667941163
transform 1 0 16688 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_302
timestamp 1667941163
transform 1 0 17584 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_330
timestamp 1667941163
transform 1 0 19152 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_2
timestamp 1667941163
transform 1 0 784 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1667941163
transform 1 0 2576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_37
timestamp 1667941163
transform 1 0 2744 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_41
timestamp 1667941163
transform 1 0 2968 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_66
timestamp 1667941163
transform 1 0 4368 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_94
timestamp 1667941163
transform 1 0 5936 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_102
timestamp 1667941163
transform 1 0 6384 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_108
timestamp 1667941163
transform 1 0 6720 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_133
timestamp 1667941163
transform 1 0 8120 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_159
timestamp 1667941163
transform 1 0 9576 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_175
timestamp 1667941163
transform 1 0 10472 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1667941163
transform 1 0 10696 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_204
timestamp 1667941163
transform 1 0 12096 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_230
timestamp 1667941163
transform 1 0 13552 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_246
timestamp 1667941163
transform 1 0 14448 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1667941163
transform 1 0 14672 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_275
timestamp 1667941163
transform 1 0 16072 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_291
timestamp 1667941163
transform 1 0 16968 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_293
timestamp 1667941163
transform 1 0 17080 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1667941163
transform 1 0 18480 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_321
timestamp 1667941163
transform 1 0 18648 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_329
timestamp 1667941163
transform 1 0 19096 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_2
timestamp 1667941163
transform 1 0 784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_10
timestamp 1667941163
transform 1 0 1232 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_14
timestamp 1667941163
transform 1 0 1456 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_40
timestamp 1667941163
transform 1 0 2912 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1667941163
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1667941163
transform 1 0 4592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_73
timestamp 1667941163
transform 1 0 4760 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_98
timestamp 1667941163
transform 1 0 6160 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_124
timestamp 1667941163
transform 1 0 7616 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_140
timestamp 1667941163
transform 1 0 8512 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_144
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 10136 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_195
timestamp 1667941163
transform 1 0 11592 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_211
timestamp 1667941163
transform 1 0 12488 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_215
timestamp 1667941163
transform 1 0 12712 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_240
timestamp 1667941163
transform 1 0 14112 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_266
timestamp 1667941163
transform 1 0 15568 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_282
timestamp 1667941163
transform 1 0 16464 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_286
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_302
timestamp 1667941163
transform 1 0 17584 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_330
timestamp 1667941163
transform 1 0 19152 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_2
timestamp 1667941163
transform 1 0 784 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1667941163
transform 1 0 2576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_37
timestamp 1667941163
transform 1 0 2744 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_41
timestamp 1667941163
transform 1 0 2968 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_66
timestamp 1667941163
transform 1 0 4368 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_94
timestamp 1667941163
transform 1 0 5936 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_102
timestamp 1667941163
transform 1 0 6384 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_108
timestamp 1667941163
transform 1 0 6720 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_133
timestamp 1667941163
transform 1 0 8120 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_159
timestamp 1667941163
transform 1 0 9576 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_175
timestamp 1667941163
transform 1 0 10472 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1667941163
transform 1 0 10696 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_204
timestamp 1667941163
transform 1 0 12096 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_230
timestamp 1667941163
transform 1 0 13552 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_246
timestamp 1667941163
transform 1 0 14448 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_250
timestamp 1667941163
transform 1 0 14672 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_266
timestamp 1667941163
transform 1 0 15568 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_292
timestamp 1667941163
transform 1 0 17024 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1667941163
transform 1 0 18480 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_321
timestamp 1667941163
transform 1 0 18648 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_329
timestamp 1667941163
transform 1 0 19096 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_2
timestamp 1667941163
transform 1 0 784 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_18
timestamp 1667941163
transform 1 0 1680 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_44
timestamp 1667941163
transform 1 0 3136 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1667941163
transform 1 0 4592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_73
timestamp 1667941163
transform 1 0 4760 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_98
timestamp 1667941163
transform 1 0 6160 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_124
timestamp 1667941163
transform 1 0 7616 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_140
timestamp 1667941163
transform 1 0 8512 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_144
timestamp 1667941163
transform 1 0 8736 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 10136 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_195
timestamp 1667941163
transform 1 0 11592 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_211
timestamp 1667941163
transform 1 0 12488 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1667941163
transform 1 0 12712 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_240
timestamp 1667941163
transform 1 0 14112 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_256
timestamp 1667941163
transform 1 0 15008 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_258
timestamp 1667941163
transform 1 0 15120 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1667941163
transform 1 0 16520 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_286
timestamp 1667941163
transform 1 0 16688 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_302
timestamp 1667941163
transform 1 0 17584 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_330
timestamp 1667941163
transform 1 0 19152 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_2
timestamp 1667941163
transform 1 0 784 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1667941163
transform 1 0 2576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_37
timestamp 1667941163
transform 1 0 2744 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_41
timestamp 1667941163
transform 1 0 2968 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_43
timestamp 1667941163
transform 1 0 3080 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_68
timestamp 1667941163
transform 1 0 4480 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_94
timestamp 1667941163
transform 1 0 5936 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_102
timestamp 1667941163
transform 1 0 6384 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_108
timestamp 1667941163
transform 1 0 6720 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_133
timestamp 1667941163
transform 1 0 8120 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_159
timestamp 1667941163
transform 1 0 9576 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_175
timestamp 1667941163
transform 1 0 10472 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1667941163
transform 1 0 10696 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_204
timestamp 1667941163
transform 1 0 12096 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_230
timestamp 1667941163
transform 1 0 13552 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_246
timestamp 1667941163
transform 1 0 14448 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_250
timestamp 1667941163
transform 1 0 14672 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_266
timestamp 1667941163
transform 1 0 15568 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_292
timestamp 1667941163
transform 1 0 17024 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1667941163
transform 1 0 18480 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_321
timestamp 1667941163
transform 1 0 18648 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_329
timestamp 1667941163
transform 1 0 19096 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_2
timestamp 1667941163
transform 1 0 784 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_18
timestamp 1667941163
transform 1 0 1680 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_44
timestamp 1667941163
transform 1 0 3136 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1667941163
transform 1 0 4592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_73
timestamp 1667941163
transform 1 0 4760 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_98
timestamp 1667941163
transform 1 0 6160 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_130
timestamp 1667941163
transform 1 0 7952 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_138
timestamp 1667941163
transform 1 0 8400 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_144
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 10136 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_195
timestamp 1667941163
transform 1 0 11592 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_211
timestamp 1667941163
transform 1 0 12488 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_215
timestamp 1667941163
transform 1 0 12712 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_240
timestamp 1667941163
transform 1 0 14112 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_256
timestamp 1667941163
transform 1 0 15008 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_258
timestamp 1667941163
transform 1 0 15120 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1667941163
transform 1 0 16520 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_286
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_302
timestamp 1667941163
transform 1 0 17584 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_330
timestamp 1667941163
transform 1 0 19152 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_2
timestamp 1667941163
transform 1 0 784 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1667941163
transform 1 0 2576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_37
timestamp 1667941163
transform 1 0 2744 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_41
timestamp 1667941163
transform 1 0 2968 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_67
timestamp 1667941163
transform 1 0 4424 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_93
timestamp 1667941163
transform 1 0 5880 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1667941163
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1667941163
transform 1 0 6552 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_108
timestamp 1667941163
transform 1 0 6720 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_133
timestamp 1667941163
transform 1 0 8120 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_159
timestamp 1667941163
transform 1 0 9576 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_175
timestamp 1667941163
transform 1 0 10472 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_179
timestamp 1667941163
transform 1 0 10696 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_204
timestamp 1667941163
transform 1 0 12096 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_230
timestamp 1667941163
transform 1 0 13552 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_246
timestamp 1667941163
transform 1 0 14448 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_250
timestamp 1667941163
transform 1 0 14672 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_266
timestamp 1667941163
transform 1 0 15568 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_292
timestamp 1667941163
transform 1 0 17024 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1667941163
transform 1 0 18480 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_321
timestamp 1667941163
transform 1 0 18648 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_329
timestamp 1667941163
transform 1 0 19096 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_2
timestamp 1667941163
transform 1 0 784 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_18
timestamp 1667941163
transform 1 0 1680 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_44
timestamp 1667941163
transform 1 0 3136 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1667941163
transform 1 0 4592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_73
timestamp 1667941163
transform 1 0 4760 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_77
timestamp 1667941163
transform 1 0 4984 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_79
timestamp 1667941163
transform 1 0 5096 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_104
timestamp 1667941163
transform 1 0 6496 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_130
timestamp 1667941163
transform 1 0 7952 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_138
timestamp 1667941163
transform 1 0 8400 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_144
timestamp 1667941163
transform 1 0 8736 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 10136 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_195
timestamp 1667941163
transform 1 0 11592 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_211
timestamp 1667941163
transform 1 0 12488 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_215
timestamp 1667941163
transform 1 0 12712 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_240
timestamp 1667941163
transform 1 0 14112 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_266
timestamp 1667941163
transform 1 0 15568 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_282
timestamp 1667941163
transform 1 0 16464 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_286
timestamp 1667941163
transform 1 0 16688 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_302
timestamp 1667941163
transform 1 0 17584 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_330
timestamp 1667941163
transform 1 0 19152 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_2
timestamp 1667941163
transform 1 0 784 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1667941163
transform 1 0 2576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_37
timestamp 1667941163
transform 1 0 2744 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_53
timestamp 1667941163
transform 1 0 3640 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_79
timestamp 1667941163
transform 1 0 5096 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1667941163
transform 1 0 6552 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_108
timestamp 1667941163
transform 1 0 6720 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_133
timestamp 1667941163
transform 1 0 8120 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_159
timestamp 1667941163
transform 1 0 9576 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_175
timestamp 1667941163
transform 1 0 10472 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_179
timestamp 1667941163
transform 1 0 10696 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_204
timestamp 1667941163
transform 1 0 12096 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_230
timestamp 1667941163
transform 1 0 13552 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_246
timestamp 1667941163
transform 1 0 14448 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1667941163
transform 1 0 14672 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_275
timestamp 1667941163
transform 1 0 16072 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_291
timestamp 1667941163
transform 1 0 16968 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_293
timestamp 1667941163
transform 1 0 17080 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1667941163
transform 1 0 18480 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_321
timestamp 1667941163
transform 1 0 18648 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_329
timestamp 1667941163
transform 1 0 19096 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_2
timestamp 1667941163
transform 1 0 784 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_18
timestamp 1667941163
transform 1 0 1680 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_44
timestamp 1667941163
transform 1 0 3136 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1667941163
transform 1 0 4592 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_73
timestamp 1667941163
transform 1 0 4760 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_77
timestamp 1667941163
transform 1 0 4984 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_79
timestamp 1667941163
transform 1 0 5096 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_104
timestamp 1667941163
transform 1 0 6496 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_130
timestamp 1667941163
transform 1 0 7952 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_138
timestamp 1667941163
transform 1 0 8400 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_144
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 10136 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_195
timestamp 1667941163
transform 1 0 11592 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_211
timestamp 1667941163
transform 1 0 12488 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_215
timestamp 1667941163
transform 1 0 12712 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_240
timestamp 1667941163
transform 1 0 14112 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_266
timestamp 1667941163
transform 1 0 15568 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_282
timestamp 1667941163
transform 1 0 16464 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_286
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_302
timestamp 1667941163
transform 1 0 17584 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_330
timestamp 1667941163
transform 1 0 19152 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_2
timestamp 1667941163
transform 1 0 784 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1667941163
transform 1 0 2576 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_37
timestamp 1667941163
transform 1 0 2744 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_53
timestamp 1667941163
transform 1 0 3640 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_79
timestamp 1667941163
transform 1 0 5096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1667941163
transform 1 0 6552 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_108
timestamp 1667941163
transform 1 0 6720 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_133
timestamp 1667941163
transform 1 0 8120 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_159
timestamp 1667941163
transform 1 0 9576 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_175
timestamp 1667941163
transform 1 0 10472 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_179
timestamp 1667941163
transform 1 0 10696 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_204
timestamp 1667941163
transform 1 0 12096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_230
timestamp 1667941163
transform 1 0 13552 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_246
timestamp 1667941163
transform 1 0 14448 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_250
timestamp 1667941163
transform 1 0 14672 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_275
timestamp 1667941163
transform 1 0 16072 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_301
timestamp 1667941163
transform 1 0 17528 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_317
timestamp 1667941163
transform 1 0 18424 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_321
timestamp 1667941163
transform 1 0 18648 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_329
timestamp 1667941163
transform 1 0 19096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_2
timestamp 1667941163
transform 1 0 784 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_18
timestamp 1667941163
transform 1 0 1680 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_44
timestamp 1667941163
transform 1 0 3136 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1667941163
transform 1 0 4592 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_73
timestamp 1667941163
transform 1 0 4760 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_77
timestamp 1667941163
transform 1 0 4984 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_79
timestamp 1667941163
transform 1 0 5096 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_104
timestamp 1667941163
transform 1 0 6496 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_130
timestamp 1667941163
transform 1 0 7952 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_138
timestamp 1667941163
transform 1 0 8400 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_144
timestamp 1667941163
transform 1 0 8736 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 10136 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_195
timestamp 1667941163
transform 1 0 11592 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_211
timestamp 1667941163
transform 1 0 12488 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1667941163
transform 1 0 12712 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_240
timestamp 1667941163
transform 1 0 14112 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_266
timestamp 1667941163
transform 1 0 15568 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_282
timestamp 1667941163
transform 1 0 16464 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_286
timestamp 1667941163
transform 1 0 16688 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_302
timestamp 1667941163
transform 1 0 17584 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_330
timestamp 1667941163
transform 1 0 19152 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_2
timestamp 1667941163
transform 1 0 784 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1667941163
transform 1 0 2576 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_37
timestamp 1667941163
transform 1 0 2744 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_53
timestamp 1667941163
transform 1 0 3640 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_79
timestamp 1667941163
transform 1 0 5096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1667941163
transform 1 0 6552 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_108
timestamp 1667941163
transform 1 0 6720 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_133
timestamp 1667941163
transform 1 0 8120 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_159
timestamp 1667941163
transform 1 0 9576 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_175
timestamp 1667941163
transform 1 0 10472 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_179
timestamp 1667941163
transform 1 0 10696 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_204
timestamp 1667941163
transform 1 0 12096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_230
timestamp 1667941163
transform 1 0 13552 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_246
timestamp 1667941163
transform 1 0 14448 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_250
timestamp 1667941163
transform 1 0 14672 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_275
timestamp 1667941163
transform 1 0 16072 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_301
timestamp 1667941163
transform 1 0 17528 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_317
timestamp 1667941163
transform 1 0 18424 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_321
timestamp 1667941163
transform 1 0 18648 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_329
timestamp 1667941163
transform 1 0 19096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_2
timestamp 1667941163
transform 1 0 784 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_18
timestamp 1667941163
transform 1 0 1680 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_44
timestamp 1667941163
transform 1 0 3136 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1667941163
transform 1 0 4592 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_73
timestamp 1667941163
transform 1 0 4760 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_77
timestamp 1667941163
transform 1 0 4984 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_79
timestamp 1667941163
transform 1 0 5096 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_104
timestamp 1667941163
transform 1 0 6496 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_130
timestamp 1667941163
transform 1 0 7952 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_138
timestamp 1667941163
transform 1 0 8400 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_144
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 10136 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_195
timestamp 1667941163
transform 1 0 11592 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_211
timestamp 1667941163
transform 1 0 12488 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1667941163
transform 1 0 12712 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_240
timestamp 1667941163
transform 1 0 14112 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_266
timestamp 1667941163
transform 1 0 15568 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_282
timestamp 1667941163
transform 1 0 16464 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_286
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_311
timestamp 1667941163
transform 1 0 18088 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_327
timestamp 1667941163
transform 1 0 18984 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_2
timestamp 1667941163
transform 1 0 784 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1667941163
transform 1 0 2576 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_37
timestamp 1667941163
transform 1 0 2744 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_53
timestamp 1667941163
transform 1 0 3640 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_79
timestamp 1667941163
transform 1 0 5096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1667941163
transform 1 0 6552 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_108
timestamp 1667941163
transform 1 0 6720 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_133
timestamp 1667941163
transform 1 0 8120 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_159
timestamp 1667941163
transform 1 0 9576 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_175
timestamp 1667941163
transform 1 0 10472 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_179
timestamp 1667941163
transform 1 0 10696 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_204
timestamp 1667941163
transform 1 0 12096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_230
timestamp 1667941163
transform 1 0 13552 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_246
timestamp 1667941163
transform 1 0 14448 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1667941163
transform 1 0 14672 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_275
timestamp 1667941163
transform 1 0 16072 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_301
timestamp 1667941163
transform 1 0 17528 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1667941163
transform 1 0 18424 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_321
timestamp 1667941163
transform 1 0 18648 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_329
timestamp 1667941163
transform 1 0 19096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_2
timestamp 1667941163
transform 1 0 784 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_18
timestamp 1667941163
transform 1 0 1680 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_44
timestamp 1667941163
transform 1 0 3136 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1667941163
transform 1 0 4592 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_73
timestamp 1667941163
transform 1 0 4760 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_77
timestamp 1667941163
transform 1 0 4984 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_79
timestamp 1667941163
transform 1 0 5096 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_104
timestamp 1667941163
transform 1 0 6496 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_130
timestamp 1667941163
transform 1 0 7952 0 -1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_138
timestamp 1667941163
transform 1 0 8400 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_144
timestamp 1667941163
transform 1 0 8736 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 10136 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_195
timestamp 1667941163
transform 1 0 11592 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_211
timestamp 1667941163
transform 1 0 12488 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1667941163
transform 1 0 12712 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_240
timestamp 1667941163
transform 1 0 14112 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_266
timestamp 1667941163
transform 1 0 15568 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_282
timestamp 1667941163
transform 1 0 16464 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1667941163
transform 1 0 16688 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_311
timestamp 1667941163
transform 1 0 18088 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_327
timestamp 1667941163
transform 1 0 18984 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_2
timestamp 1667941163
transform 1 0 784 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1667941163
transform 1 0 2576 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_37
timestamp 1667941163
transform 1 0 2744 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_53
timestamp 1667941163
transform 1 0 3640 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_79
timestamp 1667941163
transform 1 0 5096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1667941163
transform 1 0 6552 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_108
timestamp 1667941163
transform 1 0 6720 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_133
timestamp 1667941163
transform 1 0 8120 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_159
timestamp 1667941163
transform 1 0 9576 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_175
timestamp 1667941163
transform 1 0 10472 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_179
timestamp 1667941163
transform 1 0 10696 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_204
timestamp 1667941163
transform 1 0 12096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_230
timestamp 1667941163
transform 1 0 13552 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_246
timestamp 1667941163
transform 1 0 14448 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1667941163
transform 1 0 14672 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_275
timestamp 1667941163
transform 1 0 16072 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_301
timestamp 1667941163
transform 1 0 17528 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1667941163
transform 1 0 18424 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_321
timestamp 1667941163
transform 1 0 18648 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_329
timestamp 1667941163
transform 1 0 19096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_2
timestamp 1667941163
transform 1 0 784 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_18
timestamp 1667941163
transform 1 0 1680 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_44
timestamp 1667941163
transform 1 0 3136 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1667941163
transform 1 0 4592 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_73
timestamp 1667941163
transform 1 0 4760 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_77
timestamp 1667941163
transform 1 0 4984 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_79
timestamp 1667941163
transform 1 0 5096 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_104
timestamp 1667941163
transform 1 0 6496 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_130
timestamp 1667941163
transform 1 0 7952 0 -1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_138
timestamp 1667941163
transform 1 0 8400 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_144
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 10136 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_195
timestamp 1667941163
transform 1 0 11592 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_211
timestamp 1667941163
transform 1 0 12488 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1667941163
transform 1 0 12712 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_240
timestamp 1667941163
transform 1 0 14112 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_266
timestamp 1667941163
transform 1 0 15568 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1667941163
transform 1 0 16464 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_286
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_311
timestamp 1667941163
transform 1 0 18088 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_327
timestamp 1667941163
transform 1 0 18984 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_2
timestamp 1667941163
transform 1 0 784 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1667941163
transform 1 0 2576 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_37
timestamp 1667941163
transform 1 0 2744 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_53
timestamp 1667941163
transform 1 0 3640 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_79
timestamp 1667941163
transform 1 0 5096 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1667941163
transform 1 0 6552 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_108
timestamp 1667941163
transform 1 0 6720 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_133
timestamp 1667941163
transform 1 0 8120 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_159
timestamp 1667941163
transform 1 0 9576 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_175
timestamp 1667941163
transform 1 0 10472 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_179
timestamp 1667941163
transform 1 0 10696 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_204
timestamp 1667941163
transform 1 0 12096 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_230
timestamp 1667941163
transform 1 0 13552 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_246
timestamp 1667941163
transform 1 0 14448 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_250
timestamp 1667941163
transform 1 0 14672 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_275
timestamp 1667941163
transform 1 0 16072 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_301
timestamp 1667941163
transform 1 0 17528 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_317
timestamp 1667941163
transform 1 0 18424 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_321
timestamp 1667941163
transform 1 0 18648 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_329
timestamp 1667941163
transform 1 0 19096 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_2
timestamp 1667941163
transform 1 0 784 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_18
timestamp 1667941163
transform 1 0 1680 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_44
timestamp 1667941163
transform 1 0 3136 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1667941163
transform 1 0 4592 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_73
timestamp 1667941163
transform 1 0 4760 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_77
timestamp 1667941163
transform 1 0 4984 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_79
timestamp 1667941163
transform 1 0 5096 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_104
timestamp 1667941163
transform 1 0 6496 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_130
timestamp 1667941163
transform 1 0 7952 0 -1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_138
timestamp 1667941163
transform 1 0 8400 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1667941163
transform 1 0 8736 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 10136 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_195
timestamp 1667941163
transform 1 0 11592 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_211
timestamp 1667941163
transform 1 0 12488 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_215
timestamp 1667941163
transform 1 0 12712 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_240
timestamp 1667941163
transform 1 0 14112 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_266
timestamp 1667941163
transform 1 0 15568 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1667941163
transform 1 0 16464 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1667941163
transform 1 0 16688 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_311
timestamp 1667941163
transform 1 0 18088 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_327
timestamp 1667941163
transform 1 0 18984 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_2
timestamp 1667941163
transform 1 0 784 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1667941163
transform 1 0 2576 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_37
timestamp 1667941163
transform 1 0 2744 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_53
timestamp 1667941163
transform 1 0 3640 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_79
timestamp 1667941163
transform 1 0 5096 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1667941163
transform 1 0 6552 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1667941163
transform 1 0 6720 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_133
timestamp 1667941163
transform 1 0 8120 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_159
timestamp 1667941163
transform 1 0 9576 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_175
timestamp 1667941163
transform 1 0 10472 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1667941163
transform 1 0 10696 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_204
timestamp 1667941163
transform 1 0 12096 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_230
timestamp 1667941163
transform 1 0 13552 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_246
timestamp 1667941163
transform 1 0 14448 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1667941163
transform 1 0 14672 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_275
timestamp 1667941163
transform 1 0 16072 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_301
timestamp 1667941163
transform 1 0 17528 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_317
timestamp 1667941163
transform 1 0 18424 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1667941163
transform 1 0 18648 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_330
timestamp 1667941163
transform 1 0 19152 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_2
timestamp 1667941163
transform 1 0 784 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_18
timestamp 1667941163
transform 1 0 1680 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_44
timestamp 1667941163
transform 1 0 3136 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1667941163
transform 1 0 4592 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_73
timestamp 1667941163
transform 1 0 4760 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_77
timestamp 1667941163
transform 1 0 4984 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_79
timestamp 1667941163
transform 1 0 5096 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_104
timestamp 1667941163
transform 1 0 6496 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_130
timestamp 1667941163
transform 1 0 7952 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_138
timestamp 1667941163
transform 1 0 8400 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1667941163
transform 1 0 8736 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 10136 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_195
timestamp 1667941163
transform 1 0 11592 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_211
timestamp 1667941163
transform 1 0 12488 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1667941163
transform 1 0 12712 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_240
timestamp 1667941163
transform 1 0 14112 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_266
timestamp 1667941163
transform 1 0 15568 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_282
timestamp 1667941163
transform 1 0 16464 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1667941163
transform 1 0 16688 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_311
timestamp 1667941163
transform 1 0 18088 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_319
timestamp 1667941163
transform 1 0 18536 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_321
timestamp 1667941163
transform 1 0 18648 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_330
timestamp 1667941163
transform 1 0 19152 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_2
timestamp 1667941163
transform 1 0 784 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1667941163
transform 1 0 2576 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_37
timestamp 1667941163
transform 1 0 2744 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_53
timestamp 1667941163
transform 1 0 3640 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_79
timestamp 1667941163
transform 1 0 5096 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1667941163
transform 1 0 6552 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_108
timestamp 1667941163
transform 1 0 6720 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_133
timestamp 1667941163
transform 1 0 8120 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_159
timestamp 1667941163
transform 1 0 9576 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_175
timestamp 1667941163
transform 1 0 10472 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1667941163
transform 1 0 10696 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_204
timestamp 1667941163
transform 1 0 12096 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_230
timestamp 1667941163
transform 1 0 13552 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_246
timestamp 1667941163
transform 1 0 14448 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1667941163
transform 1 0 14672 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_275
timestamp 1667941163
transform 1 0 16072 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_301
timestamp 1667941163
transform 1 0 17528 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_317
timestamp 1667941163
transform 1 0 18424 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_321
timestamp 1667941163
transform 1 0 18648 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_329
timestamp 1667941163
transform 1 0 19096 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_2
timestamp 1667941163
transform 1 0 784 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_18
timestamp 1667941163
transform 1 0 1680 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_44
timestamp 1667941163
transform 1 0 3136 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1667941163
transform 1 0 4592 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_73
timestamp 1667941163
transform 1 0 4760 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_77
timestamp 1667941163
transform 1 0 4984 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_79
timestamp 1667941163
transform 1 0 5096 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_104
timestamp 1667941163
transform 1 0 6496 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_130
timestamp 1667941163
transform 1 0 7952 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_138
timestamp 1667941163
transform 1 0 8400 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1667941163
transform 1 0 8736 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 10136 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_195
timestamp 1667941163
transform 1 0 11592 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_211
timestamp 1667941163
transform 1 0 12488 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1667941163
transform 1 0 12712 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_240
timestamp 1667941163
transform 1 0 14112 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_266
timestamp 1667941163
transform 1 0 15568 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_282
timestamp 1667941163
transform 1 0 16464 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1667941163
transform 1 0 16688 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_311
timestamp 1667941163
transform 1 0 18088 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_327
timestamp 1667941163
transform 1 0 18984 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_2
timestamp 1667941163
transform 1 0 784 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1667941163
transform 1 0 2576 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_37
timestamp 1667941163
transform 1 0 2744 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_53
timestamp 1667941163
transform 1 0 3640 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_79
timestamp 1667941163
transform 1 0 5096 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1667941163
transform 1 0 6552 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_108
timestamp 1667941163
transform 1 0 6720 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_133
timestamp 1667941163
transform 1 0 8120 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_159
timestamp 1667941163
transform 1 0 9576 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_175
timestamp 1667941163
transform 1 0 10472 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1667941163
transform 1 0 10696 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_204
timestamp 1667941163
transform 1 0 12096 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_230
timestamp 1667941163
transform 1 0 13552 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_246
timestamp 1667941163
transform 1 0 14448 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_250
timestamp 1667941163
transform 1 0 14672 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_275
timestamp 1667941163
transform 1 0 16072 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_301
timestamp 1667941163
transform 1 0 17528 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1667941163
transform 1 0 18424 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_321
timestamp 1667941163
transform 1 0 18648 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_329
timestamp 1667941163
transform 1 0 19096 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_2
timestamp 1667941163
transform 1 0 784 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_18
timestamp 1667941163
transform 1 0 1680 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_44
timestamp 1667941163
transform 1 0 3136 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1667941163
transform 1 0 4592 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_73
timestamp 1667941163
transform 1 0 4760 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_77
timestamp 1667941163
transform 1 0 4984 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_79
timestamp 1667941163
transform 1 0 5096 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_104
timestamp 1667941163
transform 1 0 6496 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_130
timestamp 1667941163
transform 1 0 7952 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_138
timestamp 1667941163
transform 1 0 8400 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1667941163
transform 1 0 8736 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 10136 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_195
timestamp 1667941163
transform 1 0 11592 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_211
timestamp 1667941163
transform 1 0 12488 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_215
timestamp 1667941163
transform 1 0 12712 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_240
timestamp 1667941163
transform 1 0 14112 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_266
timestamp 1667941163
transform 1 0 15568 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_282
timestamp 1667941163
transform 1 0 16464 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_286
timestamp 1667941163
transform 1 0 16688 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_302
timestamp 1667941163
transform 1 0 17584 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_330
timestamp 1667941163
transform 1 0 19152 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_2
timestamp 1667941163
transform 1 0 784 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1667941163
transform 1 0 2576 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_37
timestamp 1667941163
transform 1 0 2744 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_53
timestamp 1667941163
transform 1 0 3640 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_79
timestamp 1667941163
transform 1 0 5096 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1667941163
transform 1 0 6552 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_108
timestamp 1667941163
transform 1 0 6720 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_133
timestamp 1667941163
transform 1 0 8120 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_159
timestamp 1667941163
transform 1 0 9576 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_175
timestamp 1667941163
transform 1 0 10472 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1667941163
transform 1 0 10696 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_204
timestamp 1667941163
transform 1 0 12096 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_230
timestamp 1667941163
transform 1 0 13552 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_246
timestamp 1667941163
transform 1 0 14448 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_250
timestamp 1667941163
transform 1 0 14672 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_275
timestamp 1667941163
transform 1 0 16072 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_301
timestamp 1667941163
transform 1 0 17528 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_317
timestamp 1667941163
transform 1 0 18424 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_321
timestamp 1667941163
transform 1 0 18648 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_329
timestamp 1667941163
transform 1 0 19096 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_2
timestamp 1667941163
transform 1 0 784 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_18
timestamp 1667941163
transform 1 0 1680 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_44
timestamp 1667941163
transform 1 0 3136 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1667941163
transform 1 0 4592 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_73
timestamp 1667941163
transform 1 0 4760 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_77
timestamp 1667941163
transform 1 0 4984 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_79
timestamp 1667941163
transform 1 0 5096 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_104
timestamp 1667941163
transform 1 0 6496 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_130
timestamp 1667941163
transform 1 0 7952 0 -1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_138
timestamp 1667941163
transform 1 0 8400 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1667941163
transform 1 0 8736 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 10136 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_195
timestamp 1667941163
transform 1 0 11592 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_211
timestamp 1667941163
transform 1 0 12488 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_215
timestamp 1667941163
transform 1 0 12712 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_240
timestamp 1667941163
transform 1 0 14112 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_266
timestamp 1667941163
transform 1 0 15568 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_282
timestamp 1667941163
transform 1 0 16464 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_286
timestamp 1667941163
transform 1 0 16688 0 -1 19600
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_318
timestamp 1667941163
transform 1 0 18480 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_330
timestamp 1667941163
transform 1 0 19152 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_2
timestamp 1667941163
transform 1 0 784 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1667941163
transform 1 0 2576 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_37
timestamp 1667941163
transform 1 0 2744 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_53
timestamp 1667941163
transform 1 0 3640 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_79
timestamp 1667941163
transform 1 0 5096 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1667941163
transform 1 0 6552 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_108
timestamp 1667941163
transform 1 0 6720 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_133
timestamp 1667941163
transform 1 0 8120 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_159
timestamp 1667941163
transform 1 0 9576 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_175
timestamp 1667941163
transform 1 0 10472 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1667941163
transform 1 0 10696 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_204
timestamp 1667941163
transform 1 0 12096 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_230
timestamp 1667941163
transform 1 0 13552 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_246
timestamp 1667941163
transform 1 0 14448 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_250
timestamp 1667941163
transform 1 0 14672 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_275
timestamp 1667941163
transform 1 0 16072 0 1 19600
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_307
timestamp 1667941163
transform 1 0 17864 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_309
timestamp 1667941163
transform 1 0 17976 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1667941163
transform 1 0 18480 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_321
timestamp 1667941163
transform 1 0 18648 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_330
timestamp 1667941163
transform 1 0 19152 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_2
timestamp 1667941163
transform 1 0 784 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_18
timestamp 1667941163
transform 1 0 1680 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_44
timestamp 1667941163
transform 1 0 3136 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1667941163
transform 1 0 4592 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_73
timestamp 1667941163
transform 1 0 4760 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_89
timestamp 1667941163
transform 1 0 5656 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_114
timestamp 1667941163
transform 1 0 7056 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_140
timestamp 1667941163
transform 1 0 8512 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_144
timestamp 1667941163
transform 1 0 8736 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 10136 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_195
timestamp 1667941163
transform 1 0 11592 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_211
timestamp 1667941163
transform 1 0 12488 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1667941163
transform 1 0 12712 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_240
timestamp 1667941163
transform 1 0 14112 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_266
timestamp 1667941163
transform 1 0 15568 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_282
timestamp 1667941163
transform 1 0 16464 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_286
timestamp 1667941163
transform 1 0 16688 0 -1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_318
timestamp 1667941163
transform 1 0 18480 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_330
timestamp 1667941163
transform 1 0 19152 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_2
timestamp 1667941163
transform 1 0 784 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1667941163
transform 1 0 2576 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_37
timestamp 1667941163
transform 1 0 2744 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_53
timestamp 1667941163
transform 1 0 3640 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_79
timestamp 1667941163
transform 1 0 5096 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1667941163
transform 1 0 6552 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_108
timestamp 1667941163
transform 1 0 6720 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_133
timestamp 1667941163
transform 1 0 8120 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_159
timestamp 1667941163
transform 1 0 9576 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_175
timestamp 1667941163
transform 1 0 10472 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1667941163
transform 1 0 10696 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_204
timestamp 1667941163
transform 1 0 12096 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_230
timestamp 1667941163
transform 1 0 13552 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_246
timestamp 1667941163
transform 1 0 14448 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_250
timestamp 1667941163
transform 1 0 14672 0 1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_282
timestamp 1667941163
transform 1 0 16464 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_298
timestamp 1667941163
transform 1 0 17360 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_306
timestamp 1667941163
transform 1 0 17808 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1667941163
transform 1 0 18480 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_321
timestamp 1667941163
transform 1 0 18648 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_330
timestamp 1667941163
transform 1 0 19152 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_2
timestamp 1667941163
transform 1 0 784 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_18
timestamp 1667941163
transform 1 0 1680 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_44
timestamp 1667941163
transform 1 0 3136 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1667941163
transform 1 0 4592 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_73
timestamp 1667941163
transform 1 0 4760 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_89
timestamp 1667941163
transform 1 0 5656 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_114
timestamp 1667941163
transform 1 0 7056 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_140
timestamp 1667941163
transform 1 0 8512 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1667941163
transform 1 0 8736 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 10136 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_195
timestamp 1667941163
transform 1 0 11592 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_211
timestamp 1667941163
transform 1 0 12488 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1667941163
transform 1 0 12712 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_240
timestamp 1667941163
transform 1 0 14112 0 -1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_272
timestamp 1667941163
transform 1 0 15904 0 -1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_280
timestamp 1667941163
transform 1 0 16352 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_286
timestamp 1667941163
transform 1 0 16688 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_310
timestamp 1667941163
transform 1 0 18032 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_320
timestamp 1667941163
transform 1 0 18592 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_330
timestamp 1667941163
transform 1 0 19152 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_2
timestamp 1667941163
transform 1 0 784 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1667941163
transform 1 0 2576 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_37
timestamp 1667941163
transform 1 0 2744 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_53
timestamp 1667941163
transform 1 0 3640 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_79
timestamp 1667941163
transform 1 0 5096 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1667941163
transform 1 0 6552 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1667941163
transform 1 0 6720 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_133
timestamp 1667941163
transform 1 0 8120 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_159
timestamp 1667941163
transform 1 0 9576 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_175
timestamp 1667941163
transform 1 0 10472 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_179
timestamp 1667941163
transform 1 0 10696 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_204
timestamp 1667941163
transform 1 0 12096 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_230
timestamp 1667941163
transform 1 0 13552 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_246
timestamp 1667941163
transform 1 0 14448 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_250
timestamp 1667941163
transform 1 0 14672 0 1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_282
timestamp 1667941163
transform 1 0 16464 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_298
timestamp 1667941163
transform 1 0 17360 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_308
timestamp 1667941163
transform 1 0 17920 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1667941163
transform 1 0 18480 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_321
timestamp 1667941163
transform 1 0 18648 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_330
timestamp 1667941163
transform 1 0 19152 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_2
timestamp 1667941163
transform 1 0 784 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_18
timestamp 1667941163
transform 1 0 1680 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_44
timestamp 1667941163
transform 1 0 3136 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1667941163
transform 1 0 4592 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_73
timestamp 1667941163
transform 1 0 4760 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_89
timestamp 1667941163
transform 1 0 5656 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_114
timestamp 1667941163
transform 1 0 7056 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_140
timestamp 1667941163
transform 1 0 8512 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1667941163
transform 1 0 8736 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 10136 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_195
timestamp 1667941163
transform 1 0 11592 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_211
timestamp 1667941163
transform 1 0 12488 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_215
timestamp 1667941163
transform 1 0 12712 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_240
timestamp 1667941163
transform 1 0 14112 0 -1 21952
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_272
timestamp 1667941163
transform 1 0 15904 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_280
timestamp 1667941163
transform 1 0 16352 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_286
timestamp 1667941163
transform 1 0 16688 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_296
timestamp 1667941163
transform 1 0 17248 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_306
timestamp 1667941163
transform 1 0 17808 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_316
timestamp 1667941163
transform 1 0 18368 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_326
timestamp 1667941163
transform 1 0 18928 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_330
timestamp 1667941163
transform 1 0 19152 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_2
timestamp 1667941163
transform 1 0 784 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1667941163
transform 1 0 2576 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_37
timestamp 1667941163
transform 1 0 2744 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_53
timestamp 1667941163
transform 1 0 3640 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_79
timestamp 1667941163
transform 1 0 5096 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1667941163
transform 1 0 6552 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_108
timestamp 1667941163
transform 1 0 6720 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_133
timestamp 1667941163
transform 1 0 8120 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_159
timestamp 1667941163
transform 1 0 9576 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_175
timestamp 1667941163
transform 1 0 10472 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_179
timestamp 1667941163
transform 1 0 10696 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_204
timestamp 1667941163
transform 1 0 12096 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_230
timestamp 1667941163
transform 1 0 13552 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_246
timestamp 1667941163
transform 1 0 14448 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_250
timestamp 1667941163
transform 1 0 14672 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_266
timestamp 1667941163
transform 1 0 15568 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_274
timestamp 1667941163
transform 1 0 16016 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_278
timestamp 1667941163
transform 1 0 16240 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_288
timestamp 1667941163
transform 1 0 16800 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_298
timestamp 1667941163
transform 1 0 17360 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_308
timestamp 1667941163
transform 1 0 17920 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1667941163
transform 1 0 18480 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_321
timestamp 1667941163
transform 1 0 18648 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_330
timestamp 1667941163
transform 1 0 19152 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_2
timestamp 1667941163
transform 1 0 784 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_18
timestamp 1667941163
transform 1 0 1680 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_44
timestamp 1667941163
transform 1 0 3136 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1667941163
transform 1 0 4592 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_73
timestamp 1667941163
transform 1 0 4760 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_89
timestamp 1667941163
transform 1 0 5656 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_114
timestamp 1667941163
transform 1 0 7056 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_140
timestamp 1667941163
transform 1 0 8512 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1667941163
transform 1 0 8736 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 10136 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_195
timestamp 1667941163
transform 1 0 11592 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_211
timestamp 1667941163
transform 1 0 12488 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_215
timestamp 1667941163
transform 1 0 12712 0 -1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_247
timestamp 1667941163
transform 1 0 14504 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_263
timestamp 1667941163
transform 1 0 15400 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_273
timestamp 1667941163
transform 1 0 15960 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1667941163
transform 1 0 16520 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_286
timestamp 1667941163
transform 1 0 16688 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_296
timestamp 1667941163
transform 1 0 17248 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_306
timestamp 1667941163
transform 1 0 17808 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_316
timestamp 1667941163
transform 1 0 18368 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_326
timestamp 1667941163
transform 1 0 18928 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_330
timestamp 1667941163
transform 1 0 19152 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_2
timestamp 1667941163
transform 1 0 784 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1667941163
transform 1 0 2576 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_37
timestamp 1667941163
transform 1 0 2744 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_53
timestamp 1667941163
transform 1 0 3640 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_79
timestamp 1667941163
transform 1 0 5096 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1667941163
transform 1 0 6552 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_108
timestamp 1667941163
transform 1 0 6720 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_133
timestamp 1667941163
transform 1 0 8120 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_159
timestamp 1667941163
transform 1 0 9576 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_175
timestamp 1667941163
transform 1 0 10472 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_179
timestamp 1667941163
transform 1 0 10696 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_204
timestamp 1667941163
transform 1 0 12096 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_236
timestamp 1667941163
transform 1 0 13888 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_244
timestamp 1667941163
transform 1 0 14336 0 1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_250
timestamp 1667941163
transform 1 0 14672 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_258
timestamp 1667941163
transform 1 0 15120 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_268
timestamp 1667941163
transform 1 0 15680 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_278
timestamp 1667941163
transform 1 0 16240 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_288
timestamp 1667941163
transform 1 0 16800 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_298
timestamp 1667941163
transform 1 0 17360 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_308
timestamp 1667941163
transform 1 0 17920 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1667941163
transform 1 0 18480 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_321
timestamp 1667941163
transform 1 0 18648 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_330
timestamp 1667941163
transform 1 0 19152 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_2
timestamp 1667941163
transform 1 0 784 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_18
timestamp 1667941163
transform 1 0 1680 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_44
timestamp 1667941163
transform 1 0 3136 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1667941163
transform 1 0 4592 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_73
timestamp 1667941163
transform 1 0 4760 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_89
timestamp 1667941163
transform 1 0 5656 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_114
timestamp 1667941163
transform 1 0 7056 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_140
timestamp 1667941163
transform 1 0 8512 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_144
timestamp 1667941163
transform 1 0 8736 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 10136 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_195
timestamp 1667941163
transform 1 0 11592 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_211
timestamp 1667941163
transform 1 0 12488 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_215
timestamp 1667941163
transform 1 0 12712 0 -1 23520
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_247
timestamp 1667941163
transform 1 0 14504 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_263
timestamp 1667941163
transform 1 0 15400 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_271
timestamp 1667941163
transform 1 0 15848 0 -1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1667941163
transform 1 0 16520 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_286
timestamp 1667941163
transform 1 0 16688 0 -1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_290
timestamp 1667941163
transform 1 0 16912 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_292
timestamp 1667941163
transform 1 0 17024 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_301
timestamp 1667941163
transform 1 0 17528 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_311
timestamp 1667941163
transform 1 0 18088 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_321
timestamp 1667941163
transform 1 0 18648 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_329
timestamp 1667941163
transform 1 0 19096 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_2
timestamp 1667941163
transform 1 0 784 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1667941163
transform 1 0 2576 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_37
timestamp 1667941163
transform 1 0 2744 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_41
timestamp 1667941163
transform 1 0 2968 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_67
timestamp 1667941163
transform 1 0 4424 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_93
timestamp 1667941163
transform 1 0 5880 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1667941163
transform 1 0 6328 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1667941163
transform 1 0 6552 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_108
timestamp 1667941163
transform 1 0 6720 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_133
timestamp 1667941163
transform 1 0 8120 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_159
timestamp 1667941163
transform 1 0 9576 0 1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_175
timestamp 1667941163
transform 1 0 10472 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 10696 0 1 23520
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1667941163
transform 1 0 14280 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1667941163
transform 1 0 14504 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_250
timestamp 1667941163
transform 1 0 14672 0 1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_266
timestamp 1667941163
transform 1 0 15568 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_274
timestamp 1667941163
transform 1 0 16016 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_278
timestamp 1667941163
transform 1 0 16240 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_288
timestamp 1667941163
transform 1 0 16800 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_298
timestamp 1667941163
transform 1 0 17360 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_308
timestamp 1667941163
transform 1 0 17920 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1667941163
transform 1 0 18480 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_321
timestamp 1667941163
transform 1 0 18648 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_330
timestamp 1667941163
transform 1 0 19152 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_2
timestamp 1667941163
transform 1 0 784 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_18
timestamp 1667941163
transform 1 0 1680 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_44
timestamp 1667941163
transform 1 0 3136 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1667941163
transform 1 0 4592 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_73
timestamp 1667941163
transform 1 0 4760 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_98
timestamp 1667941163
transform 1 0 6160 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_124
timestamp 1667941163
transform 1 0 7616 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_140
timestamp 1667941163
transform 1 0 8512 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_144
timestamp 1667941163
transform 1 0 8736 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_169
timestamp 1667941163
transform 1 0 10136 0 -1 24304
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_201
timestamp 1667941163
transform 1 0 11928 0 -1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_209
timestamp 1667941163
transform 1 0 12376 0 -1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1667941163
transform 1 0 12712 0 -1 24304
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1667941163
transform 1 0 16296 0 -1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1667941163
transform 1 0 16520 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_286
timestamp 1667941163
transform 1 0 16688 0 -1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_290
timestamp 1667941163
transform 1 0 16912 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_292
timestamp 1667941163
transform 1 0 17024 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_301
timestamp 1667941163
transform 1 0 17528 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_311
timestamp 1667941163
transform 1 0 18088 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_321
timestamp 1667941163
transform 1 0 18648 0 -1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_329
timestamp 1667941163
transform 1 0 19096 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_2
timestamp 1667941163
transform 1 0 784 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1667941163
transform 1 0 2576 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_37
timestamp 1667941163
transform 1 0 2744 0 1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_41
timestamp 1667941163
transform 1 0 2968 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_66
timestamp 1667941163
transform 1 0 4368 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_68
timestamp 1667941163
transform 1 0 4480 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_93
timestamp 1667941163
transform 1 0 5880 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1667941163
transform 1 0 6328 0 1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1667941163
transform 1 0 6552 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_108
timestamp 1667941163
transform 1 0 6720 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_133
timestamp 1667941163
transform 1 0 8120 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_159
timestamp 1667941163
transform 1 0 9576 0 1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_175
timestamp 1667941163
transform 1 0 10472 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1667941163
transform 1 0 10696 0 1 24304
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1667941163
transform 1 0 14280 0 1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1667941163
transform 1 0 14504 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_250
timestamp 1667941163
transform 1 0 14672 0 1 24304
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_282
timestamp 1667941163
transform 1 0 16464 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_298
timestamp 1667941163
transform 1 0 17360 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_308
timestamp 1667941163
transform 1 0 17920 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1667941163
transform 1 0 18480 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_321
timestamp 1667941163
transform 1 0 18648 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_330
timestamp 1667941163
transform 1 0 19152 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_2
timestamp 1667941163
transform 1 0 784 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_10
timestamp 1667941163
transform 1 0 1232 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_14
timestamp 1667941163
transform 1 0 1456 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_40
timestamp 1667941163
transform 1 0 2912 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1667941163
transform 1 0 4368 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1667941163
transform 1 0 4592 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_73
timestamp 1667941163
transform 1 0 4760 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_98
timestamp 1667941163
transform 1 0 6160 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_124
timestamp 1667941163
transform 1 0 7616 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_140
timestamp 1667941163
transform 1 0 8512 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1667941163
transform 1 0 8736 0 -1 25088
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1667941163
transform 1 0 12320 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1667941163
transform 1 0 12544 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1667941163
transform 1 0 12712 0 -1 25088
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1667941163
transform 1 0 16296 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1667941163
transform 1 0 16520 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_286
timestamp 1667941163
transform 1 0 16688 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_302
timestamp 1667941163
transform 1 0 17584 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_311
timestamp 1667941163
transform 1 0 18088 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_321
timestamp 1667941163
transform 1 0 18648 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_329
timestamp 1667941163
transform 1 0 19096 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_2
timestamp 1667941163
transform 1 0 784 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1667941163
transform 1 0 2576 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_37
timestamp 1667941163
transform 1 0 2744 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_41
timestamp 1667941163
transform 1 0 2968 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_66
timestamp 1667941163
transform 1 0 4368 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_68
timestamp 1667941163
transform 1 0 4480 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_93
timestamp 1667941163
transform 1 0 5880 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1667941163
transform 1 0 6328 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1667941163
transform 1 0 6552 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_108
timestamp 1667941163
transform 1 0 6720 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_133
timestamp 1667941163
transform 1 0 8120 0 1 25088
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_165
timestamp 1667941163
transform 1 0 9912 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_173
timestamp 1667941163
transform 1 0 10360 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1667941163
transform 1 0 10696 0 1 25088
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1667941163
transform 1 0 14280 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1667941163
transform 1 0 14504 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_250
timestamp 1667941163
transform 1 0 14672 0 1 25088
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_282
timestamp 1667941163
transform 1 0 16464 0 1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_298
timestamp 1667941163
transform 1 0 17360 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_306
timestamp 1667941163
transform 1 0 17808 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1667941163
transform 1 0 18480 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_321
timestamp 1667941163
transform 1 0 18648 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_330
timestamp 1667941163
transform 1 0 19152 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_2
timestamp 1667941163
transform 1 0 784 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_10
timestamp 1667941163
transform 1 0 1232 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_14
timestamp 1667941163
transform 1 0 1456 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_40
timestamp 1667941163
transform 1 0 2912 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1667941163
transform 1 0 4368 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1667941163
transform 1 0 4592 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_73
timestamp 1667941163
transform 1 0 4760 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_98
timestamp 1667941163
transform 1 0 6160 0 -1 25872
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_130
timestamp 1667941163
transform 1 0 7952 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_138
timestamp 1667941163
transform 1 0 8400 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1667941163
transform 1 0 8736 0 -1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1667941163
transform 1 0 12320 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1667941163
transform 1 0 12544 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1667941163
transform 1 0 12712 0 -1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1667941163
transform 1 0 16296 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1667941163
transform 1 0 16520 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_286
timestamp 1667941163
transform 1 0 16688 0 -1 25872
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_326
timestamp 1667941163
transform 1 0 18928 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_330
timestamp 1667941163
transform 1 0 19152 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1667941163
transform 1 0 784 0 1 25872
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1667941163
transform 1 0 2576 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_37
timestamp 1667941163
transform 1 0 2744 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_41
timestamp 1667941163
transform 1 0 2968 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_66
timestamp 1667941163
transform 1 0 4368 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_92
timestamp 1667941163
transform 1 0 5824 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_100
timestamp 1667941163
transform 1 0 6272 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_104
timestamp 1667941163
transform 1 0 6496 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1667941163
transform 1 0 6720 0 1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1667941163
transform 1 0 10304 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1667941163
transform 1 0 10528 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1667941163
transform 1 0 10696 0 1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1667941163
transform 1 0 14280 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1667941163
transform 1 0 14504 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1667941163
transform 1 0 14672 0 1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1667941163
transform 1 0 18256 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1667941163
transform 1 0 18480 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_321
timestamp 1667941163
transform 1 0 18648 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_329
timestamp 1667941163
transform 1 0 19096 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_2
timestamp 1667941163
transform 1 0 784 0 -1 26656
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_34
timestamp 1667941163
transform 1 0 2576 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_42
timestamp 1667941163
transform 1 0 3024 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1667941163
transform 1 0 4592 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_73
timestamp 1667941163
transform 1 0 4760 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_98
timestamp 1667941163
transform 1 0 6160 0 -1 26656
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_130
timestamp 1667941163
transform 1 0 7952 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_138
timestamp 1667941163
transform 1 0 8400 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1667941163
transform 1 0 8736 0 -1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1667941163
transform 1 0 12320 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1667941163
transform 1 0 12544 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1667941163
transform 1 0 12712 0 -1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1667941163
transform 1 0 16296 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1667941163
transform 1 0 16520 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_286
timestamp 1667941163
transform 1 0 16688 0 -1 26656
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_318
timestamp 1667941163
transform 1 0 18480 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_326
timestamp 1667941163
transform 1 0 18928 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_330
timestamp 1667941163
transform 1 0 19152 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1667941163
transform 1 0 784 0 1 26656
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1667941163
transform 1 0 2576 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_37
timestamp 1667941163
transform 1 0 2744 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_45
timestamp 1667941163
transform 1 0 3192 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_71
timestamp 1667941163
transform 1 0 4648 0 1 26656
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_103
timestamp 1667941163
transform 1 0 6440 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1667941163
transform 1 0 6552 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1667941163
transform 1 0 6720 0 1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1667941163
transform 1 0 10304 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1667941163
transform 1 0 10528 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1667941163
transform 1 0 10696 0 1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1667941163
transform 1 0 14280 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1667941163
transform 1 0 14504 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1667941163
transform 1 0 14672 0 1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 18256 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1667941163
transform 1 0 18480 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_321
timestamp 1667941163
transform 1 0 18648 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_329
timestamp 1667941163
transform 1 0 19096 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1667941163
transform 1 0 784 0 -1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1667941163
transform 1 0 4368 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1667941163
transform 1 0 4592 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1667941163
transform 1 0 4760 0 -1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1667941163
transform 1 0 8344 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1667941163
transform 1 0 8568 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1667941163
transform 1 0 8736 0 -1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1667941163
transform 1 0 12320 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1667941163
transform 1 0 12544 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1667941163
transform 1 0 12712 0 -1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1667941163
transform 1 0 16296 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1667941163
transform 1 0 16520 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_286
timestamp 1667941163
transform 1 0 16688 0 -1 27440
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_318
timestamp 1667941163
transform 1 0 18480 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_326
timestamp 1667941163
transform 1 0 18928 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_330
timestamp 1667941163
transform 1 0 19152 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1667941163
transform 1 0 784 0 1 27440
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1667941163
transform 1 0 2576 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1667941163
transform 1 0 2744 0 1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1667941163
transform 1 0 6328 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1667941163
transform 1 0 6552 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1667941163
transform 1 0 6720 0 1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1667941163
transform 1 0 10304 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1667941163
transform 1 0 10528 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1667941163
transform 1 0 10696 0 1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1667941163
transform 1 0 14280 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1667941163
transform 1 0 14504 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1667941163
transform 1 0 14672 0 1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1667941163
transform 1 0 18256 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1667941163
transform 1 0 18480 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_321
timestamp 1667941163
transform 1 0 18648 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_329
timestamp 1667941163
transform 1 0 19096 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_2
timestamp 1667941163
transform 1 0 784 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_34
timestamp 1667941163
transform 1 0 2576 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_37
timestamp 1667941163
transform 1 0 2744 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_69
timestamp 1667941163
transform 1 0 4536 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_72
timestamp 1667941163
transform 1 0 4704 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_104
timestamp 1667941163
transform 1 0 6496 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_107
timestamp 1667941163
transform 1 0 6664 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1667941163
transform 1 0 8456 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_142
timestamp 1667941163
transform 1 0 8624 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_174
timestamp 1667941163
transform 1 0 10416 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_177
timestamp 1667941163
transform 1 0 10584 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1667941163
transform 1 0 12376 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_212
timestamp 1667941163
transform 1 0 12544 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_244
timestamp 1667941163
transform 1 0 14336 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_247
timestamp 1667941163
transform 1 0 14504 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_279
timestamp 1667941163
transform 1 0 16296 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_282
timestamp 1667941163
transform 1 0 16464 0 -1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_314
timestamp 1667941163
transform 1 0 18256 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_317
timestamp 1667941163
transform 1 0 18424 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_325
timestamp 1667941163
transform 1 0 18872 0 -1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_329
timestamp 1667941163
transform 1 0 19096 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 19320 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 19320 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 19320 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 19320 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 19320 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 19320 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 19320 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 19320 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 19320 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 19320 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 19320 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 19320 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 19320 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 19320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 19320 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 19320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 19320 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1667941163
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1667941163
transform -1 0 19320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1667941163
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1667941163
transform -1 0 19320 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1667941163
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1667941163
transform -1 0 19320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1667941163
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1667941163
transform -1 0 19320 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1667941163
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1667941163
transform -1 0 19320 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1667941163
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1667941163
transform -1 0 19320 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1667941163
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1667941163
transform -1 0 19320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1667941163
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1667941163
transform -1 0 19320 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1667941163
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1667941163
transform -1 0 19320 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1667941163
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1667941163
transform -1 0 19320 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1667941163
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1667941163
transform -1 0 19320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1667941163
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1667941163
transform -1 0 19320 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1667941163
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1667941163
transform -1 0 19320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1667941163
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1667941163
transform -1 0 19320 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1667941163
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1667941163
transform -1 0 19320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1667941163
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1667941163
transform -1 0 19320 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1667941163
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1667941163
transform -1 0 19320 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1667941163
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1667941163
transform -1 0 19320 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1667941163
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1667941163
transform -1 0 19320 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1667941163
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1667941163
transform -1 0 19320 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1667941163
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1667941163
transform -1 0 19320 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1667941163
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1667941163
transform -1 0 19320 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1667941163
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1667941163
transform -1 0 19320 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1667941163
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1667941163
transform -1 0 19320 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1667941163
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1667941163
transform -1 0 19320 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1667941163
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1667941163
transform -1 0 19320 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1667941163
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1667941163
transform -1 0 19320 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1667941163
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1667941163
transform -1 0 19320 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1667941163
transform 1 0 672 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1667941163
transform -1 0 19320 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1667941163
transform 1 0 672 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1667941163
transform -1 0 19320 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1667941163
transform 1 0 672 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1667941163
transform -1 0 19320 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1667941163
transform 1 0 672 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1667941163
transform -1 0 19320 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1667941163
transform 1 0 672 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1667941163
transform -1 0 19320 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1667941163
transform 1 0 672 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1667941163
transform -1 0 19320 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1667941163
transform 1 0 672 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1667941163
transform -1 0 19320 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1667941163
transform 1 0 672 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1667941163
transform -1 0 19320 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1667941163
transform 1 0 672 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1667941163
transform -1 0 19320 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1667941163
transform 1 0 672 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1667941163
transform -1 0 19320 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1667941163
transform 1 0 672 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1667941163
transform -1 0 19320 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1667941163
transform 1 0 672 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1667941163
transform -1 0 19320 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1667941163
transform 1 0 672 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1667941163
transform -1 0 19320 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1667941163
transform 1 0 672 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1667941163
transform -1 0 19320 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1667941163
transform 1 0 672 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1667941163
transform -1 0 19320 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1667941163
transform 1 0 672 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1667941163
transform -1 0 19320 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1667941163
transform 1 0 672 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1667941163
transform -1 0 19320 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1667941163
transform 1 0 672 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1667941163
transform -1 0 19320 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1667941163
transform 1 0 672 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1667941163
transform -1 0 19320 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1667941163
transform 1 0 672 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1667941163
transform -1 0 19320 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1667941163
transform 1 0 672 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1667941163
transform -1 0 19320 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1667941163
transform 1 0 672 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1667941163
transform -1 0 19320 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1667941163
transform 1 0 672 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1667941163
transform -1 0 19320 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1667941163
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1667941163
transform 1 0 8512 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1667941163
transform 1 0 10472 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1667941163
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1667941163
transform 1 0 14392 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1667941163
transform 1 0 16352 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1667941163
transform 1 0 18312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1667941163
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1667941163
transform 1 0 12600 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1667941163
transform 1 0 16576 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1667941163
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1667941163
transform 1 0 10584 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1667941163
transform 1 0 14560 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1667941163
transform 1 0 18536 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1667941163
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1667941163
transform 1 0 12600 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1667941163
transform 1 0 16576 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1667941163
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1667941163
transform 1 0 10584 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1667941163
transform 1 0 14560 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1667941163
transform 1 0 18536 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 8624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 12600 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 16576 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 10584 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 14560 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 18536 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 8624 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 12600 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 16576 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 10584 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 14560 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 18536 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 8624 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 12600 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 16576 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 10584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 14560 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 18536 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 4648 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 12600 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 16576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 6608 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 14560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 18536 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 4648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 12600 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 16576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 6608 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 14560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 18536 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 4648 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 12600 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 16576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 6608 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 14560 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 18536 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 4648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 12600 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 16576 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 6608 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 14560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 18536 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 4648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 12600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 16576 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 6608 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 14560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 18536 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 4648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 12600 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 16576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 6608 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 14560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 18536 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 4648 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 12600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 16576 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 6608 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 10584 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 14560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 18536 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 4648 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 12600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 16576 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 6608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 10584 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 14560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 18536 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 4648 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 12600 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 16576 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 6608 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 14560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 18536 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 4648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 12600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 16576 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 6608 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 14560 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 18536 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 4648 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 12600 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 16576 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 6608 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 10584 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 14560 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1667941163
transform 1 0 18536 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1667941163
transform 1 0 4648 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1667941163
transform 1 0 8624 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1667941163
transform 1 0 12600 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1667941163
transform 1 0 16576 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1667941163
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1667941163
transform 1 0 6608 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1667941163
transform 1 0 10584 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1667941163
transform 1 0 14560 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1667941163
transform 1 0 18536 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1667941163
transform 1 0 4648 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1667941163
transform 1 0 8624 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1667941163
transform 1 0 12600 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1667941163
transform 1 0 16576 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1667941163
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1667941163
transform 1 0 6608 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1667941163
transform 1 0 10584 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1667941163
transform 1 0 14560 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1667941163
transform 1 0 18536 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1667941163
transform 1 0 4648 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1667941163
transform 1 0 8624 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1667941163
transform 1 0 12600 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1667941163
transform 1 0 16576 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1667941163
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1667941163
transform 1 0 6608 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1667941163
transform 1 0 10584 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1667941163
transform 1 0 14560 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1667941163
transform 1 0 18536 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1667941163
transform 1 0 4648 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1667941163
transform 1 0 8624 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1667941163
transform 1 0 12600 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1667941163
transform 1 0 16576 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1667941163
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1667941163
transform 1 0 6608 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1667941163
transform 1 0 10584 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1667941163
transform 1 0 14560 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1667941163
transform 1 0 18536 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1667941163
transform 1 0 4648 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1667941163
transform 1 0 8624 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1667941163
transform 1 0 12600 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1667941163
transform 1 0 16576 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1667941163
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1667941163
transform 1 0 6608 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1667941163
transform 1 0 10584 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1667941163
transform 1 0 14560 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1667941163
transform 1 0 18536 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1667941163
transform 1 0 4648 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1667941163
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1667941163
transform 1 0 12600 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1667941163
transform 1 0 16576 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1667941163
transform 1 0 2632 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1667941163
transform 1 0 6608 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1667941163
transform 1 0 10584 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1667941163
transform 1 0 14560 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1667941163
transform 1 0 18536 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1667941163
transform 1 0 4648 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1667941163
transform 1 0 8624 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1667941163
transform 1 0 12600 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1667941163
transform 1 0 16576 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1667941163
transform 1 0 2632 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1667941163
transform 1 0 6608 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1667941163
transform 1 0 10584 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1667941163
transform 1 0 14560 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1667941163
transform 1 0 18536 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1667941163
transform 1 0 4648 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1667941163
transform 1 0 8624 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1667941163
transform 1 0 12600 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1667941163
transform 1 0 16576 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1667941163
transform 1 0 2632 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1667941163
transform 1 0 6608 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1667941163
transform 1 0 10584 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1667941163
transform 1 0 14560 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1667941163
transform 1 0 18536 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1667941163
transform 1 0 4648 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1667941163
transform 1 0 8624 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1667941163
transform 1 0 12600 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1667941163
transform 1 0 16576 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1667941163
transform 1 0 2632 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1667941163
transform 1 0 6608 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1667941163
transform 1 0 10584 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1667941163
transform 1 0 14560 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1667941163
transform 1 0 18536 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1667941163
transform 1 0 4648 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1667941163
transform 1 0 8624 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1667941163
transform 1 0 12600 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1667941163
transform 1 0 16576 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1667941163
transform 1 0 2632 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1667941163
transform 1 0 6608 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1667941163
transform 1 0 10584 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1667941163
transform 1 0 14560 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1667941163
transform 1 0 18536 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1667941163
transform 1 0 4648 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1667941163
transform 1 0 8624 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1667941163
transform 1 0 12600 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1667941163
transform 1 0 16576 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1667941163
transform 1 0 2632 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1667941163
transform 1 0 6608 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1667941163
transform 1 0 10584 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1667941163
transform 1 0 14560 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1667941163
transform 1 0 18536 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1667941163
transform 1 0 4648 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1667941163
transform 1 0 8624 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1667941163
transform 1 0 12600 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1667941163
transform 1 0 16576 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1667941163
transform 1 0 2632 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1667941163
transform 1 0 6608 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1667941163
transform 1 0 10584 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1667941163
transform 1 0 14560 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1667941163
transform 1 0 18536 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1667941163
transform 1 0 4648 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1667941163
transform 1 0 8624 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1667941163
transform 1 0 12600 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1667941163
transform 1 0 16576 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1667941163
transform 1 0 2632 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1667941163
transform 1 0 6608 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1667941163
transform 1 0 10584 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1667941163
transform 1 0 14560 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1667941163
transform 1 0 18536 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1667941163
transform 1 0 4648 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1667941163
transform 1 0 8624 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1667941163
transform 1 0 12600 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1667941163
transform 1 0 16576 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1667941163
transform 1 0 2632 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1667941163
transform 1 0 6608 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1667941163
transform 1 0 10584 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1667941163
transform 1 0 14560 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1667941163
transform 1 0 18536 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1667941163
transform 1 0 4648 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1667941163
transform 1 0 8624 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1667941163
transform 1 0 12600 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1667941163
transform 1 0 16576 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1667941163
transform 1 0 2632 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1667941163
transform 1 0 6608 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1667941163
transform 1 0 10584 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1667941163
transform 1 0 14560 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1667941163
transform 1 0 18536 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1667941163
transform 1 0 4648 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1667941163
transform 1 0 8624 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1667941163
transform 1 0 12600 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1667941163
transform 1 0 16576 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1667941163
transform 1 0 2632 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1667941163
transform 1 0 6608 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1667941163
transform 1 0 10584 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1667941163
transform 1 0 14560 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1667941163
transform 1 0 18536 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1667941163
transform 1 0 4648 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1667941163
transform 1 0 8624 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1667941163
transform 1 0 12600 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1667941163
transform 1 0 16576 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1667941163
transform 1 0 2632 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1667941163
transform 1 0 6608 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1667941163
transform 1 0 10584 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1667941163
transform 1 0 14560 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1667941163
transform 1 0 18536 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1667941163
transform 1 0 2632 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1667941163
transform 1 0 4592 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1667941163
transform 1 0 6552 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1667941163
transform 1 0 8512 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1667941163
transform 1 0 10472 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1667941163
transform 1 0 12432 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1667941163
transform 1 0 14392 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1667941163
transform 1 0 16352 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1667941163
transform 1 0 18312 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 13552 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyn2
timestamp 1667941163
transform -1 0 9072 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 14112 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyp2
timestamp 1667941163
transform -1 0 10528 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 12544 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyn2
timestamp 1667941163
transform -1 0 14112 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 13552 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyp2
timestamp 1667941163
transform -1 0 13552 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 11592 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyn2
timestamp 1667941163
transform -1 0 10584 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 13552 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyp2
timestamp 1667941163
transform -1 0 14112 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 12096 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyn2
timestamp 1667941163
transform -1 0 15568 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 14112 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyp2
timestamp 1667941163
transform -1 0 14112 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 12544 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyn2
timestamp 1667941163
transform -1 0 9072 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 14112 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyp2
timestamp 1667941163
transform -1 0 16072 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 13552 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyn2
timestamp 1667941163
transform -1 0 15568 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 12096 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyp2
timestamp 1667941163
transform -1 0 16072 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 11088 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyn2
timestamp 1667941163
transform 1 0 14728 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 16072 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyp2
timestamp 1667941163
transform 1 0 5768 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 10528 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyn2
timestamp 1667941163
transform -1 0 8568 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 12544 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyp2
timestamp 1667941163
transform -1 0 12096 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 13552 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyn2
timestamp 1667941163
transform -1 0 13552 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyp2
timestamp 1667941163
transform -1 0 15568 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 12096 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyn2
timestamp 1667941163
transform 1 0 14728 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyp2
timestamp 1667941163
transform -1 0 15568 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 11088 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyn2
timestamp 1667941163
transform -1 0 12096 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyp2
timestamp 1667941163
transform -1 0 12544 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyn2
timestamp 1667941163
transform -1 0 8568 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyp2
timestamp 1667941163
transform 1 0 16184 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 12096 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyn2
timestamp 1667941163
transform -1 0 13552 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyp2
timestamp 1667941163
transform -1 0 10528 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 10528 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyn2
timestamp 1667941163
transform -1 0 14112 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 12096 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyp2
timestamp 1667941163
transform -1 0 9072 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 11088 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyn2
timestamp 1667941163
transform -1 0 15568 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyp1
timestamp 1667941163
transform -1 0 12544 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyp2
timestamp 1667941163
transform -1 0 8568 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 12096 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyn2
timestamp 1667941163
transform -1 0 10528 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyp1
timestamp 1667941163
transform 1 0 7728 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyp2
timestamp 1667941163
transform -1 0 12040 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 10416 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 11984 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 9072 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyp1
timestamp 1667941163
transform 1 0 16184 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 8568 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 8568 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 11984 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 13552 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 13552 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyp1
timestamp 1667941163
transform 1 0 5768 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 14112 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 15568 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyn1
timestamp 1667941163
transform 1 0 14728 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyp1
timestamp 1667941163
transform 1 0 5208 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 6552 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 7112 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 8456 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyp1
timestamp 1667941163
transform 1 0 3752 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyn1
timestamp 1667941163
transform 1 0 3752 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 6552 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 7112 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyp1
timestamp 1667941163
transform 1 0 3248 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 6496 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyp1
timestamp 1667941163
transform 1 0 3248 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyn1
timestamp 1667941163
transform 1 0 3752 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyp1
timestamp 1667941163
transform 1 0 3248 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyn1
timestamp 1667941163
transform 1 0 14560 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 2912 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 5992 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 5992 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_p
timestamp 1667941163
transform -1 0 5992 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_p
timestamp 1667941163
transform -1 0 5936 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_p
timestamp 1667941163
transform -1 0 5992 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[64\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[64\].u_shunt_p
timestamp 1667941163
transform -1 0 4536 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[65\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[65\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[66\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[66\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[67\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[67\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[68\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[68\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[69\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[69\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[70\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[70\].u_shunt_p
timestamp 1667941163
transform -1 0 4424 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[71\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[71\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[72\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[72\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[73\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[73\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[74\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[74\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[75\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[75\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[76\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[76\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[77\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[77\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[78\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[78\].u_shunt_p
timestamp 1667941163
transform -1 0 5992 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[79\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[79\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[80\].u_shunt_n
timestamp 1667941163
transform -1 0 7952 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[80\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[81\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[81\].u_shunt_p
timestamp 1667941163
transform -1 0 5936 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[82\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[82\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[83\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[83\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[84\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[84\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[85\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[85\].u_shunt_p
timestamp 1667941163
transform -1 0 4536 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[86\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[86\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[87\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[87\].u_shunt_p
timestamp 1667941163
transform -1 0 4480 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[88\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[88\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[89\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[89\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[90\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[90\].u_shunt_p
timestamp 1667941163
transform -1 0 5936 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[91\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[91\].u_shunt_p
timestamp 1667941163
transform -1 0 5880 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[92\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[92\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[93\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[93\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[94\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[94\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[95\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[95\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 8512 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 7056 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 8512 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 8512 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 8512 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 6496 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 5880 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 5880 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 7056 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 7056 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 7056 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 5880 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 7056 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 8512 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 4424 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 4648 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 2912 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 2912 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 2912 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 6160 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 5824 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 7616 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 8120 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 6160 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 4368 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 2688 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 4144 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 4144 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 4144 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 2688 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 2688 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 4144 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 4144 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 13944 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g8\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g8\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 16520 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 17360 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 17360 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18088 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 16800 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 18480 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 16520 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18480 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 17920 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 17920 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18648 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 17920 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 17528 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18648 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 18704 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 17248 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 17248 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 17360 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18480 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 18704 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 18480 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 17528 0 -1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18648 0 -1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 16800 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 16352 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 16240 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 17920 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15232 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 18704 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 17808 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 17808 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 17360 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 18368 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18480 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 18704 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 17360 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 18704 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18480 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18928 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15512 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 17472 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18928 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 18032 0 -1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 18368 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18928 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18480 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 18144 0 -1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 18704 0 -1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 18704 0 -1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 18704 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 18704 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 18032 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 18704 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 18704 0 -1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_n
timestamp 1667941163
transform 1 0 18704 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_p
timestamp 1667941163
transform 1 0 18704 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15176 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15680 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15680 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17808 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18480 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15176 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18480 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17808 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18480 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 15680 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 18480 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17808 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17808 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17808 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17808 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17136 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17136 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 17808 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 15680 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn3
timestamp 1667941163
transform 1 0 15680 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 17136 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 18480 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp3
timestamp 1667941163
transform 1 0 17808 0 -1 2352
box -43 -43 1387 435
<< labels >>
flabel metal2 s 18592 29600 18648 30000 0 FreeSans 224 90 0 0 cap_series_gygyn
port 0 nsew signal bidirectional
flabel metal2 s 16128 29600 16184 30000 0 FreeSans 224 90 0 0 cap_series_gygyp
port 1 nsew signal bidirectional
flabel metal2 s 13664 29600 13720 30000 0 FreeSans 224 90 0 0 cap_series_gyn
port 2 nsew signal bidirectional
flabel metal2 s 11200 29600 11256 30000 0 FreeSans 224 90 0 0 cap_series_gyp
port 3 nsew signal bidirectional
flabel metal2 s 8736 29600 8792 30000 0 FreeSans 224 90 0 0 cap_shunt_gyn
port 4 nsew signal bidirectional
flabel metal2 s 6272 29600 6328 30000 0 FreeSans 224 90 0 0 cap_shunt_gyp
port 5 nsew signal bidirectional
flabel metal2 s 3808 29600 3864 30000 0 FreeSans 224 90 0 0 cap_shunt_n
port 6 nsew signal bidirectional
flabel metal2 s 1344 29600 1400 30000 0 FreeSans 224 90 0 0 cap_shunt_p
port 7 nsew signal bidirectional
flabel metal2 s 1680 0 1736 400 0 FreeSans 224 90 0 0 tune_series_gy[0]
port 8 nsew signal input
flabel metal2 s 4984 0 5040 400 0 FreeSans 224 90 0 0 tune_series_gy[1]
port 9 nsew signal input
flabel metal2 s 8288 0 8344 400 0 FreeSans 224 90 0 0 tune_series_gy[2]
port 10 nsew signal input
flabel metal2 s 11592 0 11648 400 0 FreeSans 224 90 0 0 tune_series_gy[3]
port 11 nsew signal input
flabel metal2 s 14896 0 14952 400 0 FreeSans 224 90 0 0 tune_series_gy[4]
port 12 nsew signal input
flabel metal2 s 18200 0 18256 400 0 FreeSans 224 90 0 0 tune_series_gy[5]
port 13 nsew signal input
flabel metal3 s 19600 1176 20000 1232 0 FreeSans 224 0 0 0 tune_series_gygy[0]
port 14 nsew signal input
flabel metal3 s 19600 3472 20000 3528 0 FreeSans 224 0 0 0 tune_series_gygy[1]
port 15 nsew signal input
flabel metal3 s 19600 5768 20000 5824 0 FreeSans 224 0 0 0 tune_series_gygy[2]
port 16 nsew signal input
flabel metal3 s 19600 8064 20000 8120 0 FreeSans 224 0 0 0 tune_series_gygy[3]
port 17 nsew signal input
flabel metal3 s 19600 10360 20000 10416 0 FreeSans 224 0 0 0 tune_series_gygy[4]
port 18 nsew signal input
flabel metal3 s 19600 12656 20000 12712 0 FreeSans 224 0 0 0 tune_series_gygy[5]
port 19 nsew signal input
flabel metal3 s 0 2016 400 2072 0 FreeSans 224 0 0 0 tune_shunt[0]
port 20 nsew signal input
flabel metal3 s 0 5712 400 5768 0 FreeSans 224 0 0 0 tune_shunt[1]
port 21 nsew signal input
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 tune_shunt[2]
port 22 nsew signal input
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 tune_shunt[3]
port 23 nsew signal input
flabel metal3 s 0 16800 400 16856 0 FreeSans 224 0 0 0 tune_shunt[4]
port 24 nsew signal input
flabel metal3 s 0 20496 400 20552 0 FreeSans 224 0 0 0 tune_shunt[5]
port 25 nsew signal input
flabel metal3 s 0 24192 400 24248 0 FreeSans 224 0 0 0 tune_shunt[6]
port 26 nsew signal input
flabel metal3 s 0 27888 400 27944 0 FreeSans 224 0 0 0 tune_shunt[7]
port 27 nsew signal input
flabel metal3 s 19600 14952 20000 15008 0 FreeSans 224 0 0 0 tune_shunt_gy[0]
port 28 nsew signal input
flabel metal3 s 19600 17248 20000 17304 0 FreeSans 224 0 0 0 tune_shunt_gy[1]
port 29 nsew signal input
flabel metal3 s 19600 19544 20000 19600 0 FreeSans 224 0 0 0 tune_shunt_gy[2]
port 30 nsew signal input
flabel metal3 s 19600 21840 20000 21896 0 FreeSans 224 0 0 0 tune_shunt_gy[3]
port 31 nsew signal input
flabel metal3 s 19600 24136 20000 24192 0 FreeSans 224 0 0 0 tune_shunt_gy[4]
port 32 nsew signal input
flabel metal3 s 19600 26432 20000 26488 0 FreeSans 224 0 0 0 tune_shunt_gy[5]
port 33 nsew signal input
flabel metal3 s 19600 28728 20000 28784 0 FreeSans 224 0 0 0 tune_shunt_gy[6]
port 34 nsew signal input
flabel metal4 s 2224 1538 2384 28254 0 FreeSans 640 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 17584 1538 17744 28254 0 FreeSans 640 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 9904 1538 10064 28254 0 FreeSans 640 90 0 0 vss
port 36 nsew ground bidirectional
rlabel metal1 9996 27832 9996 27832 0 vdd
rlabel via1 9996 28224 9996 28224 0 vss
rlabel metal2 15484 10808 15484 10808 0 cap_series_gygyn
rlabel metal2 17892 2184 17892 2184 0 cap_series_gygyp
rlabel metal2 3892 4088 3892 4088 0 cap_series_gyn
rlabel metal2 4060 3920 4060 3920 0 cap_series_gyp
rlabel metal3 15680 22596 15680 22596 0 cap_shunt_gyn
rlabel metal2 17836 25088 17836 25088 0 cap_shunt_gyp
rlabel metal2 3836 1736 3836 1736 0 cap_shunt_n
rlabel metal2 2044 2968 2044 2968 0 cap_shunt_p
rlabel metal2 1708 1211 1708 1211 0 tune_series_gy[0]
rlabel metal2 5124 1764 5124 1764 0 tune_series_gy[1]
rlabel metal3 7896 1764 7896 1764 0 tune_series_gy[2]
rlabel metal3 13832 3724 13832 3724 0 tune_series_gy[3]
rlabel metal3 12068 3724 12068 3724 0 tune_series_gy[4]
rlabel metal3 11900 4060 11900 4060 0 tune_series_gy[5]
rlabel metal2 18788 2352 18788 2352 0 tune_series_gygy[0]
rlabel metal2 17500 2996 17500 2996 0 tune_series_gygy[1]
rlabel metal3 18592 3332 18592 3332 0 tune_series_gygy[2]
rlabel metal2 18844 3962 18844 3962 0 tune_series_gygy[3]
rlabel metal3 19257 10388 19257 10388 0 tune_series_gygy[4]
rlabel metal2 19068 12516 19068 12516 0 tune_series_gygy[5]
rlabel metal3 427 2044 427 2044 0 tune_shunt[0]
rlabel metal2 2884 1792 2884 1792 0 tune_shunt[1]
rlabel metal2 924 2352 924 2352 0 tune_shunt[2]
rlabel metal2 12684 22148 12684 22148 0 tune_shunt[3]
rlabel metal2 14588 11760 14588 11760 0 tune_shunt[4]
rlabel metal2 1428 10780 1428 10780 0 tune_shunt[5]
rlabel metal2 3612 22932 3612 22932 0 tune_shunt[6]
rlabel metal2 1876 15092 1876 15092 0 tune_shunt[7]
rlabel metal3 19341 14980 19341 14980 0 tune_shunt_gy[0]
rlabel metal2 19068 18340 19068 18340 0 tune_shunt_gy[1]
rlabel metal2 19012 20076 19012 20076 0 tune_shunt_gy[2]
rlabel metal2 19068 21980 19068 21980 0 tune_shunt_gy[3]
rlabel metal2 15876 22176 15876 22176 0 tune_shunt_gy[4]
rlabel metal2 19012 25480 19012 25480 0 tune_shunt_gy[5]
rlabel metal3 15736 22876 15736 22876 0 tune_shunt_gy[6]
<< properties >>
string FIXED_BBOX 0 0 20000 30000
<< end >>
