// This is the unpowered netlist.
module caparray_s2 (cap_series_gygyn,
    cap_series_gygyp,
    cap_series_gyn,
    cap_series_gyp,
    cap_shunt_gyn,
    cap_shunt_gyp,
    cap_shunt_n,
    cap_shunt_p,
    tune_series_gy,
    tune_series_gygy,
    tune_shunt,
    tune_shunt_gy);
 inout cap_series_gygyn;
 inout cap_series_gygyp;
 inout cap_series_gyn;
 inout cap_series_gyp;
 inout cap_shunt_gyn;
 inout cap_shunt_gyp;
 inout cap_shunt_n;
 inout cap_shunt_p;
 input [7:0] tune_series_gy;
 input [7:0] tune_series_gygy;
 input [10:0] tune_shunt;
 input [4:0] tune_shunt_gy;

 wire \gen_series_gy_g1[0].d1 ;
 wire \gen_series_gy_g1[0].d2 ;
 wire \gen_series_gy_g1[10].d1 ;
 wire \gen_series_gy_g1[10].d2 ;
 wire \gen_series_gy_g1[11].d1 ;
 wire \gen_series_gy_g1[11].d2 ;
 wire \gen_series_gy_g1[12].d1 ;
 wire \gen_series_gy_g1[12].d2 ;
 wire \gen_series_gy_g1[13].d1 ;
 wire \gen_series_gy_g1[13].d2 ;
 wire \gen_series_gy_g1[14].d1 ;
 wire \gen_series_gy_g1[14].d2 ;
 wire \gen_series_gy_g1[15].d1 ;
 wire \gen_series_gy_g1[15].d2 ;
 wire \gen_series_gy_g1[16].d1 ;
 wire \gen_series_gy_g1[16].d2 ;
 wire \gen_series_gy_g1[17].d1 ;
 wire \gen_series_gy_g1[17].d2 ;
 wire \gen_series_gy_g1[18].d1 ;
 wire \gen_series_gy_g1[18].d2 ;
 wire \gen_series_gy_g1[19].d1 ;
 wire \gen_series_gy_g1[19].d2 ;
 wire \gen_series_gy_g1[1].d1 ;
 wire \gen_series_gy_g1[1].d2 ;
 wire \gen_series_gy_g1[20].d1 ;
 wire \gen_series_gy_g1[20].d2 ;
 wire \gen_series_gy_g1[21].d1 ;
 wire \gen_series_gy_g1[21].d2 ;
 wire \gen_series_gy_g1[22].d1 ;
 wire \gen_series_gy_g1[22].d2 ;
 wire \gen_series_gy_g1[23].d1 ;
 wire \gen_series_gy_g1[23].d2 ;
 wire \gen_series_gy_g1[24].d1 ;
 wire \gen_series_gy_g1[24].d2 ;
 wire \gen_series_gy_g1[25].d1 ;
 wire \gen_series_gy_g1[25].d2 ;
 wire \gen_series_gy_g1[26].d1 ;
 wire \gen_series_gy_g1[26].d2 ;
 wire \gen_series_gy_g1[27].d1 ;
 wire \gen_series_gy_g1[27].d2 ;
 wire \gen_series_gy_g1[28].d1 ;
 wire \gen_series_gy_g1[28].d2 ;
 wire \gen_series_gy_g1[29].d1 ;
 wire \gen_series_gy_g1[29].d2 ;
 wire \gen_series_gy_g1[2].d1 ;
 wire \gen_series_gy_g1[2].d2 ;
 wire \gen_series_gy_g1[30].d1 ;
 wire \gen_series_gy_g1[30].d2 ;
 wire \gen_series_gy_g1[31].d1 ;
 wire \gen_series_gy_g1[31].d2 ;
 wire \gen_series_gy_g1[3].d1 ;
 wire \gen_series_gy_g1[3].d2 ;
 wire \gen_series_gy_g1[4].d1 ;
 wire \gen_series_gy_g1[4].d2 ;
 wire \gen_series_gy_g1[5].d1 ;
 wire \gen_series_gy_g1[5].d2 ;
 wire \gen_series_gy_g1[6].d1 ;
 wire \gen_series_gy_g1[6].d2 ;
 wire \gen_series_gy_g1[7].d1 ;
 wire \gen_series_gy_g1[7].d2 ;
 wire \gen_series_gy_g1[8].d1 ;
 wire \gen_series_gy_g1[8].d2 ;
 wire \gen_series_gy_g1[9].d1 ;
 wire \gen_series_gy_g1[9].d2 ;
 wire \gen_series_gy_g2[0].d1 ;
 wire \gen_series_gy_g2[0].d2 ;
 wire \gen_series_gy_g2[10].d1 ;
 wire \gen_series_gy_g2[10].d2 ;
 wire \gen_series_gy_g2[11].d1 ;
 wire \gen_series_gy_g2[11].d2 ;
 wire \gen_series_gy_g2[12].d1 ;
 wire \gen_series_gy_g2[12].d2 ;
 wire \gen_series_gy_g2[13].d1 ;
 wire \gen_series_gy_g2[13].d2 ;
 wire \gen_series_gy_g2[14].d1 ;
 wire \gen_series_gy_g2[14].d2 ;
 wire \gen_series_gy_g2[15].d1 ;
 wire \gen_series_gy_g2[15].d2 ;
 wire \gen_series_gy_g2[1].d1 ;
 wire \gen_series_gy_g2[1].d2 ;
 wire \gen_series_gy_g2[2].d1 ;
 wire \gen_series_gy_g2[2].d2 ;
 wire \gen_series_gy_g2[3].d1 ;
 wire \gen_series_gy_g2[3].d2 ;
 wire \gen_series_gy_g2[4].d1 ;
 wire \gen_series_gy_g2[4].d2 ;
 wire \gen_series_gy_g2[5].d1 ;
 wire \gen_series_gy_g2[5].d2 ;
 wire \gen_series_gy_g2[6].d1 ;
 wire \gen_series_gy_g2[6].d2 ;
 wire \gen_series_gy_g2[7].d1 ;
 wire \gen_series_gy_g2[7].d2 ;
 wire \gen_series_gy_g2[8].d1 ;
 wire \gen_series_gy_g2[8].d2 ;
 wire \gen_series_gy_g2[9].d1 ;
 wire \gen_series_gy_g2[9].d2 ;
 wire \gen_series_gy_g3[0].d1 ;
 wire \gen_series_gy_g3[0].d2 ;
 wire \gen_series_gy_g3[0].d3 ;
 wire \gen_series_gy_g3[0].d4 ;
 wire \gen_series_gy_g3[1].d1 ;
 wire \gen_series_gy_g3[1].d2 ;
 wire \gen_series_gy_g3[1].d3 ;
 wire \gen_series_gy_g3[1].d4 ;
 wire \gen_series_gy_g3[2].d1 ;
 wire \gen_series_gy_g3[2].d2 ;
 wire \gen_series_gy_g3[2].d3 ;
 wire \gen_series_gy_g3[2].d4 ;
 wire \gen_series_gy_g3[3].d1 ;
 wire \gen_series_gy_g3[3].d2 ;
 wire \gen_series_gy_g3[3].d3 ;
 wire \gen_series_gy_g3[3].d4 ;
 wire \gen_series_gy_g3[4].d1 ;
 wire \gen_series_gy_g3[4].d2 ;
 wire \gen_series_gy_g3[4].d3 ;
 wire \gen_series_gy_g3[4].d4 ;
 wire \gen_series_gy_g3[5].d1 ;
 wire \gen_series_gy_g3[5].d2 ;
 wire \gen_series_gy_g3[5].d3 ;
 wire \gen_series_gy_g3[5].d4 ;
 wire \gen_series_gy_g3[6].d1 ;
 wire \gen_series_gy_g3[6].d2 ;
 wire \gen_series_gy_g3[6].d3 ;
 wire \gen_series_gy_g3[6].d4 ;
 wire \gen_series_gy_g3[7].d1 ;
 wire \gen_series_gy_g3[7].d2 ;
 wire \gen_series_gy_g3[7].d3 ;
 wire \gen_series_gy_g3[7].d4 ;
 wire \gen_series_gy_g4[0].d1 ;
 wire \gen_series_gy_g4[0].d2 ;
 wire \gen_series_gy_g4[0].d3 ;
 wire \gen_series_gy_g4[0].d4 ;
 wire \gen_series_gy_g4[1].d1 ;
 wire \gen_series_gy_g4[1].d2 ;
 wire \gen_series_gy_g4[1].d3 ;
 wire \gen_series_gy_g4[1].d4 ;
 wire \gen_series_gy_g4[2].d1 ;
 wire \gen_series_gy_g4[2].d2 ;
 wire \gen_series_gy_g4[2].d3 ;
 wire \gen_series_gy_g4[2].d4 ;
 wire \gen_series_gy_g4[3].d1 ;
 wire \gen_series_gy_g4[3].d2 ;
 wire \gen_series_gy_g4[3].d3 ;
 wire \gen_series_gy_g4[3].d4 ;
 wire \gen_series_gy_g5[0].d1 ;
 wire \gen_series_gy_g5[0].d2 ;
 wire \gen_series_gy_g5[1].d1 ;
 wire \gen_series_gy_g5[1].d2 ;
 wire \gen_series_gy_g6[0].d1 ;
 wire \gen_series_gy_g6[0].d2 ;
 wire \gen_shunt_g1[0].d1 ;
 wire \gen_shunt_g1[0].d2 ;
 wire \gen_shunt_g1[10].d1 ;
 wire \gen_shunt_g1[10].d2 ;
 wire \gen_shunt_g1[11].d1 ;
 wire \gen_shunt_g1[11].d2 ;
 wire \gen_shunt_g1[12].d1 ;
 wire \gen_shunt_g1[12].d2 ;
 wire \gen_shunt_g1[13].d1 ;
 wire \gen_shunt_g1[13].d2 ;
 wire \gen_shunt_g1[14].d1 ;
 wire \gen_shunt_g1[14].d2 ;
 wire \gen_shunt_g1[15].d1 ;
 wire \gen_shunt_g1[15].d2 ;
 wire \gen_shunt_g1[16].d1 ;
 wire \gen_shunt_g1[16].d2 ;
 wire \gen_shunt_g1[17].d1 ;
 wire \gen_shunt_g1[17].d2 ;
 wire \gen_shunt_g1[18].d1 ;
 wire \gen_shunt_g1[18].d2 ;
 wire \gen_shunt_g1[19].d1 ;
 wire \gen_shunt_g1[19].d2 ;
 wire \gen_shunt_g1[1].d1 ;
 wire \gen_shunt_g1[1].d2 ;
 wire \gen_shunt_g1[20].d1 ;
 wire \gen_shunt_g1[20].d2 ;
 wire \gen_shunt_g1[21].d1 ;
 wire \gen_shunt_g1[21].d2 ;
 wire \gen_shunt_g1[22].d1 ;
 wire \gen_shunt_g1[22].d2 ;
 wire \gen_shunt_g1[23].d1 ;
 wire \gen_shunt_g1[23].d2 ;
 wire \gen_shunt_g1[24].d1 ;
 wire \gen_shunt_g1[24].d2 ;
 wire \gen_shunt_g1[25].d1 ;
 wire \gen_shunt_g1[25].d2 ;
 wire \gen_shunt_g1[26].d1 ;
 wire \gen_shunt_g1[26].d2 ;
 wire \gen_shunt_g1[27].d1 ;
 wire \gen_shunt_g1[27].d2 ;
 wire \gen_shunt_g1[28].d1 ;
 wire \gen_shunt_g1[28].d2 ;
 wire \gen_shunt_g1[29].d1 ;
 wire \gen_shunt_g1[29].d2 ;
 wire \gen_shunt_g1[2].d1 ;
 wire \gen_shunt_g1[2].d2 ;
 wire \gen_shunt_g1[30].d1 ;
 wire \gen_shunt_g1[30].d2 ;
 wire \gen_shunt_g1[31].d1 ;
 wire \gen_shunt_g1[31].d2 ;
 wire \gen_shunt_g1[32].d1 ;
 wire \gen_shunt_g1[32].d2 ;
 wire \gen_shunt_g1[33].d1 ;
 wire \gen_shunt_g1[33].d2 ;
 wire \gen_shunt_g1[34].d1 ;
 wire \gen_shunt_g1[34].d2 ;
 wire \gen_shunt_g1[35].d1 ;
 wire \gen_shunt_g1[35].d2 ;
 wire \gen_shunt_g1[36].d1 ;
 wire \gen_shunt_g1[36].d2 ;
 wire \gen_shunt_g1[37].d1 ;
 wire \gen_shunt_g1[37].d2 ;
 wire \gen_shunt_g1[38].d1 ;
 wire \gen_shunt_g1[38].d2 ;
 wire \gen_shunt_g1[39].d1 ;
 wire \gen_shunt_g1[39].d2 ;
 wire \gen_shunt_g1[3].d1 ;
 wire \gen_shunt_g1[3].d2 ;
 wire \gen_shunt_g1[40].d1 ;
 wire \gen_shunt_g1[40].d2 ;
 wire \gen_shunt_g1[41].d1 ;
 wire \gen_shunt_g1[41].d2 ;
 wire \gen_shunt_g1[42].d1 ;
 wire \gen_shunt_g1[42].d2 ;
 wire \gen_shunt_g1[43].d1 ;
 wire \gen_shunt_g1[43].d2 ;
 wire \gen_shunt_g1[44].d1 ;
 wire \gen_shunt_g1[44].d2 ;
 wire \gen_shunt_g1[45].d1 ;
 wire \gen_shunt_g1[45].d2 ;
 wire \gen_shunt_g1[46].d1 ;
 wire \gen_shunt_g1[46].d2 ;
 wire \gen_shunt_g1[47].d1 ;
 wire \gen_shunt_g1[47].d2 ;
 wire \gen_shunt_g1[48].d1 ;
 wire \gen_shunt_g1[48].d2 ;
 wire \gen_shunt_g1[49].d1 ;
 wire \gen_shunt_g1[49].d2 ;
 wire \gen_shunt_g1[4].d1 ;
 wire \gen_shunt_g1[4].d2 ;
 wire \gen_shunt_g1[50].d1 ;
 wire \gen_shunt_g1[50].d2 ;
 wire \gen_shunt_g1[51].d1 ;
 wire \gen_shunt_g1[51].d2 ;
 wire \gen_shunt_g1[52].d1 ;
 wire \gen_shunt_g1[52].d2 ;
 wire \gen_shunt_g1[53].d1 ;
 wire \gen_shunt_g1[53].d2 ;
 wire \gen_shunt_g1[54].d1 ;
 wire \gen_shunt_g1[54].d2 ;
 wire \gen_shunt_g1[55].d1 ;
 wire \gen_shunt_g1[55].d2 ;
 wire \gen_shunt_g1[56].d1 ;
 wire \gen_shunt_g1[56].d2 ;
 wire \gen_shunt_g1[57].d1 ;
 wire \gen_shunt_g1[57].d2 ;
 wire \gen_shunt_g1[58].d1 ;
 wire \gen_shunt_g1[58].d2 ;
 wire \gen_shunt_g1[59].d1 ;
 wire \gen_shunt_g1[59].d2 ;
 wire \gen_shunt_g1[5].d1 ;
 wire \gen_shunt_g1[5].d2 ;
 wire \gen_shunt_g1[60].d1 ;
 wire \gen_shunt_g1[60].d2 ;
 wire \gen_shunt_g1[61].d1 ;
 wire \gen_shunt_g1[61].d2 ;
 wire \gen_shunt_g1[62].d1 ;
 wire \gen_shunt_g1[62].d2 ;
 wire \gen_shunt_g1[63].d1 ;
 wire \gen_shunt_g1[63].d2 ;
 wire \gen_shunt_g1[6].d1 ;
 wire \gen_shunt_g1[6].d2 ;
 wire \gen_shunt_g1[7].d1 ;
 wire \gen_shunt_g1[7].d2 ;
 wire \gen_shunt_g1[8].d1 ;
 wire \gen_shunt_g1[8].d2 ;
 wire \gen_shunt_g1[9].d1 ;
 wire \gen_shunt_g1[9].d2 ;
 wire \gen_shunt_g2[0].d1 ;
 wire \gen_shunt_g2[0].d2 ;
 wire \gen_shunt_g2[0].d3 ;
 wire \gen_shunt_g2[0].d4 ;
 wire \gen_shunt_g2[10].d1 ;
 wire \gen_shunt_g2[10].d2 ;
 wire \gen_shunt_g2[10].d3 ;
 wire \gen_shunt_g2[10].d4 ;
 wire \gen_shunt_g2[11].d1 ;
 wire \gen_shunt_g2[11].d2 ;
 wire \gen_shunt_g2[11].d3 ;
 wire \gen_shunt_g2[11].d4 ;
 wire \gen_shunt_g2[12].d1 ;
 wire \gen_shunt_g2[12].d2 ;
 wire \gen_shunt_g2[12].d3 ;
 wire \gen_shunt_g2[12].d4 ;
 wire \gen_shunt_g2[13].d1 ;
 wire \gen_shunt_g2[13].d2 ;
 wire \gen_shunt_g2[13].d3 ;
 wire \gen_shunt_g2[13].d4 ;
 wire \gen_shunt_g2[14].d1 ;
 wire \gen_shunt_g2[14].d2 ;
 wire \gen_shunt_g2[14].d3 ;
 wire \gen_shunt_g2[14].d4 ;
 wire \gen_shunt_g2[15].d1 ;
 wire \gen_shunt_g2[15].d2 ;
 wire \gen_shunt_g2[15].d3 ;
 wire \gen_shunt_g2[15].d4 ;
 wire \gen_shunt_g2[16].d1 ;
 wire \gen_shunt_g2[16].d2 ;
 wire \gen_shunt_g2[16].d3 ;
 wire \gen_shunt_g2[16].d4 ;
 wire \gen_shunt_g2[17].d1 ;
 wire \gen_shunt_g2[17].d2 ;
 wire \gen_shunt_g2[17].d3 ;
 wire \gen_shunt_g2[17].d4 ;
 wire \gen_shunt_g2[18].d1 ;
 wire \gen_shunt_g2[18].d2 ;
 wire \gen_shunt_g2[18].d3 ;
 wire \gen_shunt_g2[18].d4 ;
 wire \gen_shunt_g2[19].d1 ;
 wire \gen_shunt_g2[19].d2 ;
 wire \gen_shunt_g2[19].d3 ;
 wire \gen_shunt_g2[19].d4 ;
 wire \gen_shunt_g2[1].d1 ;
 wire \gen_shunt_g2[1].d2 ;
 wire \gen_shunt_g2[1].d3 ;
 wire \gen_shunt_g2[1].d4 ;
 wire \gen_shunt_g2[20].d1 ;
 wire \gen_shunt_g2[20].d2 ;
 wire \gen_shunt_g2[20].d3 ;
 wire \gen_shunt_g2[20].d4 ;
 wire \gen_shunt_g2[21].d1 ;
 wire \gen_shunt_g2[21].d2 ;
 wire \gen_shunt_g2[21].d3 ;
 wire \gen_shunt_g2[21].d4 ;
 wire \gen_shunt_g2[22].d1 ;
 wire \gen_shunt_g2[22].d2 ;
 wire \gen_shunt_g2[22].d3 ;
 wire \gen_shunt_g2[22].d4 ;
 wire \gen_shunt_g2[23].d1 ;
 wire \gen_shunt_g2[23].d2 ;
 wire \gen_shunt_g2[23].d3 ;
 wire \gen_shunt_g2[23].d4 ;
 wire \gen_shunt_g2[24].d1 ;
 wire \gen_shunt_g2[24].d2 ;
 wire \gen_shunt_g2[24].d3 ;
 wire \gen_shunt_g2[24].d4 ;
 wire \gen_shunt_g2[25].d1 ;
 wire \gen_shunt_g2[25].d2 ;
 wire \gen_shunt_g2[25].d3 ;
 wire \gen_shunt_g2[25].d4 ;
 wire \gen_shunt_g2[26].d1 ;
 wire \gen_shunt_g2[26].d2 ;
 wire \gen_shunt_g2[26].d3 ;
 wire \gen_shunt_g2[26].d4 ;
 wire \gen_shunt_g2[27].d1 ;
 wire \gen_shunt_g2[27].d2 ;
 wire \gen_shunt_g2[27].d3 ;
 wire \gen_shunt_g2[27].d4 ;
 wire \gen_shunt_g2[28].d1 ;
 wire \gen_shunt_g2[28].d2 ;
 wire \gen_shunt_g2[28].d3 ;
 wire \gen_shunt_g2[28].d4 ;
 wire \gen_shunt_g2[29].d1 ;
 wire \gen_shunt_g2[29].d2 ;
 wire \gen_shunt_g2[29].d3 ;
 wire \gen_shunt_g2[29].d4 ;
 wire \gen_shunt_g2[2].d1 ;
 wire \gen_shunt_g2[2].d2 ;
 wire \gen_shunt_g2[2].d3 ;
 wire \gen_shunt_g2[2].d4 ;
 wire \gen_shunt_g2[30].d1 ;
 wire \gen_shunt_g2[30].d2 ;
 wire \gen_shunt_g2[30].d3 ;
 wire \gen_shunt_g2[30].d4 ;
 wire \gen_shunt_g2[31].d1 ;
 wire \gen_shunt_g2[31].d2 ;
 wire \gen_shunt_g2[31].d3 ;
 wire \gen_shunt_g2[31].d4 ;
 wire \gen_shunt_g2[3].d1 ;
 wire \gen_shunt_g2[3].d2 ;
 wire \gen_shunt_g2[3].d3 ;
 wire \gen_shunt_g2[3].d4 ;
 wire \gen_shunt_g2[4].d1 ;
 wire \gen_shunt_g2[4].d2 ;
 wire \gen_shunt_g2[4].d3 ;
 wire \gen_shunt_g2[4].d4 ;
 wire \gen_shunt_g2[5].d1 ;
 wire \gen_shunt_g2[5].d2 ;
 wire \gen_shunt_g2[5].d3 ;
 wire \gen_shunt_g2[5].d4 ;
 wire \gen_shunt_g2[6].d1 ;
 wire \gen_shunt_g2[6].d2 ;
 wire \gen_shunt_g2[6].d3 ;
 wire \gen_shunt_g2[6].d4 ;
 wire \gen_shunt_g2[7].d1 ;
 wire \gen_shunt_g2[7].d2 ;
 wire \gen_shunt_g2[7].d3 ;
 wire \gen_shunt_g2[7].d4 ;
 wire \gen_shunt_g2[8].d1 ;
 wire \gen_shunt_g2[8].d2 ;
 wire \gen_shunt_g2[8].d3 ;
 wire \gen_shunt_g2[8].d4 ;
 wire \gen_shunt_g2[9].d1 ;
 wire \gen_shunt_g2[9].d2 ;
 wire \gen_shunt_g2[9].d3 ;
 wire \gen_shunt_g2[9].d4 ;
 wire \gen_shunt_g3[0].d1 ;
 wire \gen_shunt_g3[0].d2 ;
 wire \gen_shunt_g3[0].d3 ;
 wire \gen_shunt_g3[0].d4 ;
 wire \gen_shunt_g3[10].d1 ;
 wire \gen_shunt_g3[10].d2 ;
 wire \gen_shunt_g3[10].d3 ;
 wire \gen_shunt_g3[10].d4 ;
 wire \gen_shunt_g3[11].d1 ;
 wire \gen_shunt_g3[11].d2 ;
 wire \gen_shunt_g3[11].d3 ;
 wire \gen_shunt_g3[11].d4 ;
 wire \gen_shunt_g3[12].d1 ;
 wire \gen_shunt_g3[12].d2 ;
 wire \gen_shunt_g3[12].d3 ;
 wire \gen_shunt_g3[12].d4 ;
 wire \gen_shunt_g3[13].d1 ;
 wire \gen_shunt_g3[13].d2 ;
 wire \gen_shunt_g3[13].d3 ;
 wire \gen_shunt_g3[13].d4 ;
 wire \gen_shunt_g3[14].d1 ;
 wire \gen_shunt_g3[14].d2 ;
 wire \gen_shunt_g3[14].d3 ;
 wire \gen_shunt_g3[14].d4 ;
 wire \gen_shunt_g3[15].d1 ;
 wire \gen_shunt_g3[15].d2 ;
 wire \gen_shunt_g3[15].d3 ;
 wire \gen_shunt_g3[15].d4 ;
 wire \gen_shunt_g3[1].d1 ;
 wire \gen_shunt_g3[1].d2 ;
 wire \gen_shunt_g3[1].d3 ;
 wire \gen_shunt_g3[1].d4 ;
 wire \gen_shunt_g3[2].d1 ;
 wire \gen_shunt_g3[2].d2 ;
 wire \gen_shunt_g3[2].d3 ;
 wire \gen_shunt_g3[2].d4 ;
 wire \gen_shunt_g3[3].d1 ;
 wire \gen_shunt_g3[3].d2 ;
 wire \gen_shunt_g3[3].d3 ;
 wire \gen_shunt_g3[3].d4 ;
 wire \gen_shunt_g3[4].d1 ;
 wire \gen_shunt_g3[4].d2 ;
 wire \gen_shunt_g3[4].d3 ;
 wire \gen_shunt_g3[4].d4 ;
 wire \gen_shunt_g3[5].d1 ;
 wire \gen_shunt_g3[5].d2 ;
 wire \gen_shunt_g3[5].d3 ;
 wire \gen_shunt_g3[5].d4 ;
 wire \gen_shunt_g3[6].d1 ;
 wire \gen_shunt_g3[6].d2 ;
 wire \gen_shunt_g3[6].d3 ;
 wire \gen_shunt_g3[6].d4 ;
 wire \gen_shunt_g3[7].d1 ;
 wire \gen_shunt_g3[7].d2 ;
 wire \gen_shunt_g3[7].d3 ;
 wire \gen_shunt_g3[7].d4 ;
 wire \gen_shunt_g3[8].d1 ;
 wire \gen_shunt_g3[8].d2 ;
 wire \gen_shunt_g3[8].d3 ;
 wire \gen_shunt_g3[8].d4 ;
 wire \gen_shunt_g3[9].d1 ;
 wire \gen_shunt_g3[9].d2 ;
 wire \gen_shunt_g3[9].d3 ;
 wire \gen_shunt_g3[9].d4 ;
 wire \gen_shunt_g4[0].d1 ;
 wire \gen_shunt_g4[0].d2 ;
 wire \gen_shunt_g4[0].d3 ;
 wire \gen_shunt_g4[0].d4 ;
 wire \gen_shunt_g4[1].d1 ;
 wire \gen_shunt_g4[1].d2 ;
 wire \gen_shunt_g4[1].d3 ;
 wire \gen_shunt_g4[1].d4 ;
 wire \gen_shunt_g4[2].d1 ;
 wire \gen_shunt_g4[2].d2 ;
 wire \gen_shunt_g4[2].d3 ;
 wire \gen_shunt_g4[2].d4 ;
 wire \gen_shunt_g4[3].d1 ;
 wire \gen_shunt_g4[3].d2 ;
 wire \gen_shunt_g4[3].d3 ;
 wire \gen_shunt_g4[3].d4 ;
 wire \gen_shunt_g4[4].d1 ;
 wire \gen_shunt_g4[4].d2 ;
 wire \gen_shunt_g4[4].d3 ;
 wire \gen_shunt_g4[4].d4 ;
 wire \gen_shunt_g4[5].d1 ;
 wire \gen_shunt_g4[5].d2 ;
 wire \gen_shunt_g4[5].d3 ;
 wire \gen_shunt_g4[5].d4 ;
 wire \gen_shunt_g4[6].d1 ;
 wire \gen_shunt_g4[6].d2 ;
 wire \gen_shunt_g4[6].d3 ;
 wire \gen_shunt_g4[6].d4 ;
 wire \gen_shunt_g4[7].d1 ;
 wire \gen_shunt_g4[7].d2 ;
 wire \gen_shunt_g4[7].d3 ;
 wire \gen_shunt_g4[7].d4 ;
 wire \gen_shunt_g5[0].d1 ;
 wire \gen_shunt_g5[0].d2 ;
 wire \gen_shunt_g5[1].d1 ;
 wire \gen_shunt_g5[1].d2 ;
 wire \gen_shunt_g5[2].d1 ;
 wire \gen_shunt_g5[2].d2 ;
 wire \gen_shunt_g5[3].d1 ;
 wire \gen_shunt_g5[3].d2 ;
 wire \gen_shunt_g6[0].d1 ;
 wire \gen_shunt_g6[0].d2 ;
 wire \gen_shunt_g6[0].d3 ;
 wire \gen_shunt_g6[0].d4 ;
 wire \gen_shunt_g6[1].d1 ;
 wire \gen_shunt_g6[1].d2 ;
 wire \gen_shunt_g6[1].d3 ;
 wire \gen_shunt_g6[1].d4 ;
 wire \gen_shunt_g7[0].d1 ;
 wire \gen_shunt_g7[0].d2 ;
 wire \gen_shunt_gy_g1[0].d1 ;
 wire \gen_shunt_gy_g1[0].d2 ;
 wire \gen_shunt_gy_g1[0].d3 ;
 wire \gen_shunt_gy_g1[0].d4 ;
 wire \gen_shunt_gy_g1[1].d1 ;
 wire \gen_shunt_gy_g1[1].d2 ;
 wire \gen_shunt_gy_g1[1].d3 ;
 wire \gen_shunt_gy_g1[1].d4 ;
 wire \gen_shunt_gy_g1[2].d1 ;
 wire \gen_shunt_gy_g1[2].d2 ;
 wire \gen_shunt_gy_g1[2].d3 ;
 wire \gen_shunt_gy_g1[2].d4 ;
 wire \gen_shunt_gy_g1[3].d1 ;
 wire \gen_shunt_gy_g1[3].d2 ;
 wire \gen_shunt_gy_g1[3].d3 ;
 wire \gen_shunt_gy_g1[3].d4 ;
 wire \gen_shunt_gy_g1[4].d1 ;
 wire \gen_shunt_gy_g1[4].d2 ;
 wire \gen_shunt_gy_g1[4].d3 ;
 wire \gen_shunt_gy_g1[4].d4 ;
 wire \gen_shunt_gy_g1[5].d1 ;
 wire \gen_shunt_gy_g1[5].d2 ;
 wire \gen_shunt_gy_g1[5].d3 ;
 wire \gen_shunt_gy_g1[5].d4 ;
 wire \gen_shunt_gy_g1[6].d1 ;
 wire \gen_shunt_gy_g1[6].d2 ;
 wire \gen_shunt_gy_g1[6].d3 ;
 wire \gen_shunt_gy_g1[6].d4 ;
 wire \gen_shunt_gy_g1[7].d1 ;
 wire \gen_shunt_gy_g1[7].d2 ;
 wire \gen_shunt_gy_g1[7].d3 ;
 wire \gen_shunt_gy_g1[7].d4 ;
 wire \gen_shunt_gy_g2[0].d1 ;
 wire \gen_shunt_gy_g2[0].d2 ;
 wire \gen_shunt_gy_g2[0].d3 ;
 wire \gen_shunt_gy_g2[0].d4 ;
 wire \gen_shunt_gy_g2[1].d1 ;
 wire \gen_shunt_gy_g2[1].d2 ;
 wire \gen_shunt_gy_g2[1].d3 ;
 wire \gen_shunt_gy_g2[1].d4 ;
 wire \gen_shunt_gy_g2[2].d1 ;
 wire \gen_shunt_gy_g2[2].d2 ;
 wire \gen_shunt_gy_g2[2].d3 ;
 wire \gen_shunt_gy_g2[2].d4 ;
 wire \gen_shunt_gy_g2[3].d1 ;
 wire \gen_shunt_gy_g2[3].d2 ;
 wire \gen_shunt_gy_g2[3].d3 ;
 wire \gen_shunt_gy_g2[3].d4 ;
 wire \gen_shunt_gy_g3[0].d1 ;
 wire \gen_shunt_gy_g3[0].d2 ;
 wire \gen_shunt_gy_g3[1].d1 ;
 wire \gen_shunt_gy_g3[1].d2 ;
 wire \gen_shunt_gy_g4[0].d1 ;
 wire \gen_shunt_gy_g4[0].d2 ;
 wire \gen_shunt_gygy_g1[0].d1 ;
 wire \gen_shunt_gygy_g1[0].d2 ;
 wire \gen_shunt_gygy_g1[0].d3 ;
 wire \gen_shunt_gygy_g1[0].d4 ;
 wire \gen_shunt_gygy_g1[10].d1 ;
 wire \gen_shunt_gygy_g1[10].d2 ;
 wire \gen_shunt_gygy_g1[10].d3 ;
 wire \gen_shunt_gygy_g1[10].d4 ;
 wire \gen_shunt_gygy_g1[11].d1 ;
 wire \gen_shunt_gygy_g1[11].d2 ;
 wire \gen_shunt_gygy_g1[11].d3 ;
 wire \gen_shunt_gygy_g1[11].d4 ;
 wire \gen_shunt_gygy_g1[12].d1 ;
 wire \gen_shunt_gygy_g1[12].d2 ;
 wire \gen_shunt_gygy_g1[12].d3 ;
 wire \gen_shunt_gygy_g1[12].d4 ;
 wire \gen_shunt_gygy_g1[13].d1 ;
 wire \gen_shunt_gygy_g1[13].d2 ;
 wire \gen_shunt_gygy_g1[13].d3 ;
 wire \gen_shunt_gygy_g1[13].d4 ;
 wire \gen_shunt_gygy_g1[14].d1 ;
 wire \gen_shunt_gygy_g1[14].d2 ;
 wire \gen_shunt_gygy_g1[14].d3 ;
 wire \gen_shunt_gygy_g1[14].d4 ;
 wire \gen_shunt_gygy_g1[15].d1 ;
 wire \gen_shunt_gygy_g1[15].d2 ;
 wire \gen_shunt_gygy_g1[15].d3 ;
 wire \gen_shunt_gygy_g1[15].d4 ;
 wire \gen_shunt_gygy_g1[1].d1 ;
 wire \gen_shunt_gygy_g1[1].d2 ;
 wire \gen_shunt_gygy_g1[1].d3 ;
 wire \gen_shunt_gygy_g1[1].d4 ;
 wire \gen_shunt_gygy_g1[2].d1 ;
 wire \gen_shunt_gygy_g1[2].d2 ;
 wire \gen_shunt_gygy_g1[2].d3 ;
 wire \gen_shunt_gygy_g1[2].d4 ;
 wire \gen_shunt_gygy_g1[3].d1 ;
 wire \gen_shunt_gygy_g1[3].d2 ;
 wire \gen_shunt_gygy_g1[3].d3 ;
 wire \gen_shunt_gygy_g1[3].d4 ;
 wire \gen_shunt_gygy_g1[4].d1 ;
 wire \gen_shunt_gygy_g1[4].d2 ;
 wire \gen_shunt_gygy_g1[4].d3 ;
 wire \gen_shunt_gygy_g1[4].d4 ;
 wire \gen_shunt_gygy_g1[5].d1 ;
 wire \gen_shunt_gygy_g1[5].d2 ;
 wire \gen_shunt_gygy_g1[5].d3 ;
 wire \gen_shunt_gygy_g1[5].d4 ;
 wire \gen_shunt_gygy_g1[6].d1 ;
 wire \gen_shunt_gygy_g1[6].d2 ;
 wire \gen_shunt_gygy_g1[6].d3 ;
 wire \gen_shunt_gygy_g1[6].d4 ;
 wire \gen_shunt_gygy_g1[7].d1 ;
 wire \gen_shunt_gygy_g1[7].d2 ;
 wire \gen_shunt_gygy_g1[7].d3 ;
 wire \gen_shunt_gygy_g1[7].d4 ;
 wire \gen_shunt_gygy_g1[8].d1 ;
 wire \gen_shunt_gygy_g1[8].d2 ;
 wire \gen_shunt_gygy_g1[8].d3 ;
 wire \gen_shunt_gygy_g1[8].d4 ;
 wire \gen_shunt_gygy_g1[9].d1 ;
 wire \gen_shunt_gygy_g1[9].d2 ;
 wire \gen_shunt_gygy_g1[9].d3 ;
 wire \gen_shunt_gygy_g1[9].d4 ;
 wire \gen_shunt_gygy_g2[0].d1 ;
 wire \gen_shunt_gygy_g2[0].d2 ;
 wire \gen_shunt_gygy_g2[0].d3 ;
 wire \gen_shunt_gygy_g2[0].d4 ;
 wire \gen_shunt_gygy_g2[1].d1 ;
 wire \gen_shunt_gygy_g2[1].d2 ;
 wire \gen_shunt_gygy_g2[1].d3 ;
 wire \gen_shunt_gygy_g2[1].d4 ;
 wire \gen_shunt_gygy_g2[2].d1 ;
 wire \gen_shunt_gygy_g2[2].d2 ;
 wire \gen_shunt_gygy_g2[2].d3 ;
 wire \gen_shunt_gygy_g2[2].d4 ;
 wire \gen_shunt_gygy_g2[3].d1 ;
 wire \gen_shunt_gygy_g2[3].d2 ;
 wire \gen_shunt_gygy_g2[3].d3 ;
 wire \gen_shunt_gygy_g2[3].d4 ;
 wire \gen_shunt_gygy_g2[4].d1 ;
 wire \gen_shunt_gygy_g2[4].d2 ;
 wire \gen_shunt_gygy_g2[4].d3 ;
 wire \gen_shunt_gygy_g2[4].d4 ;
 wire \gen_shunt_gygy_g2[5].d1 ;
 wire \gen_shunt_gygy_g2[5].d2 ;
 wire \gen_shunt_gygy_g2[5].d3 ;
 wire \gen_shunt_gygy_g2[5].d4 ;
 wire \gen_shunt_gygy_g2[6].d1 ;
 wire \gen_shunt_gygy_g2[6].d2 ;
 wire \gen_shunt_gygy_g2[6].d3 ;
 wire \gen_shunt_gygy_g2[6].d4 ;
 wire \gen_shunt_gygy_g2[7].d1 ;
 wire \gen_shunt_gygy_g2[7].d2 ;
 wire \gen_shunt_gygy_g2[7].d3 ;
 wire \gen_shunt_gygy_g2[7].d4 ;
 wire \gen_shunt_gygy_g3[0].d1 ;
 wire \gen_shunt_gygy_g3[0].d2 ;
 wire \gen_shunt_gygy_g3[1].d1 ;
 wire \gen_shunt_gygy_g3[1].d2 ;
 wire \gen_shunt_gygy_g3[2].d1 ;
 wire \gen_shunt_gygy_g3[2].d2 ;
 wire \gen_shunt_gygy_g3[3].d1 ;
 wire \gen_shunt_gygy_g3[3].d2 ;
 wire \gen_shunt_gygy_g4[0].d1 ;
 wire \gen_shunt_gygy_g4[0].d2 ;
 wire \gen_shunt_gygy_g4[0].d3 ;
 wire \gen_shunt_gygy_g4[0].d4 ;
 wire \gen_shunt_gygy_g4[1].d1 ;
 wire \gen_shunt_gygy_g4[1].d2 ;
 wire \gen_shunt_gygy_g4[1].d3 ;
 wire \gen_shunt_gygy_g4[1].d4 ;
 wire \gen_shunt_gygy_g5[0].d1 ;
 wire \gen_shunt_gygy_g5[0].d2 ;

 gf180mcu_fd_sc_mcu7t5v0__tiel _0_ (.ZN(\gen_shunt_gy_g2[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1_ (.ZN(\gen_shunt_gy_g2[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2_ (.ZN(\gen_shunt_gy_g2[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3_ (.ZN(\gen_shunt_gy_g2[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _4_ (.ZN(\gen_shunt_gy_g2[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _5_ (.ZN(\gen_shunt_gy_g2[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _6_ (.ZN(\gen_shunt_gy_g2[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _7_ (.ZN(\gen_shunt_gy_g2[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[10].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[10].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[10].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[11].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[11].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[11].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[12].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[12].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[12].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[13].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[13].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[13].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[14].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[14].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[14].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[15].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[15].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[15].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[16].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[16].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[16].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[16].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[17].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[17].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[17].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[17].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[18].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[18].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[18].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[18].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[19].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[19].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[19].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[19].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[20].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[20].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[20].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[20].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[21].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[21].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[21].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[21].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[22].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[22].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[22].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[22].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[23].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[23].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[23].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[23].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[24].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[24].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[24].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[24].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[25].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[25].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[25].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[25].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[26].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[26].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[26].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[26].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[27].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[27].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[27].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[27].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[28].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[28].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[28].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[28].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[29].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[29].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[29].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[29].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[30].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[30].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[30].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[30].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[31].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[31].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[31].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[31].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[8].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[8].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[8].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[9].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g1[9].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[7]),
    .ZN(\gen_series_gy_g1[9].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[10].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[10].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[10].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[10].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[11].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[11].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[11].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[11].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[12].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[12].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[12].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[12].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[13].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[13].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[13].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[13].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[14].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[14].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[14].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[14].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[15].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[15].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[15].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[15].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[8].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[8].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[8].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[8].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[9].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[9].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g2[9].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[6]),
    .ZN(\gen_series_gy_g2[9].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[0].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[1].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[2].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[3].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[4].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[5].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[6].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[5]),
    .ZN(\gen_series_gy_g3[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g3[7].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[4]),
    .ZN(\gen_series_gy_g3[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[0].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[1].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[2].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyn2  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[3]),
    .ZN(\gen_series_gy_g4[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g4[3].u_series_gyp2  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[2]),
    .ZN(\gen_series_gy_g4[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[1].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g5[1].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[1]),
    .ZN(\gen_series_gy_g5[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g6[0].u_series_gyn1  (.A1(cap_series_gyn),
    .A2(cap_series_gyn),
    .B(tune_series_gy[0]),
    .ZN(\gen_series_gy_g6[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_series_gy_g6[0].u_series_gyp1  (.A1(cap_series_gyp),
    .A2(cap_series_gyp),
    .B(tune_series_gy[0]),
    .ZN(\gen_series_gy_g6[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[10].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[10].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[10].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[10].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[11].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[11].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[11].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[11].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[12].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[12].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[12].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[12].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[13].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[13].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[13].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[13].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[14].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[14].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[14].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[14].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[15].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[15].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[15].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[15].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[16].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[16].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[16].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[16].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[17].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[17].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[17].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[17].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[18].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[18].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[18].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[18].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[19].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[19].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[19].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[19].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[20].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[20].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[20].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[20].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[21].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[21].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[21].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[21].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[22].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[22].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[22].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[22].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[23].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[23].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[23].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[23].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[24].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[24].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[24].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[24].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[25].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[25].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[25].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[25].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[26].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[26].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[26].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[26].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[27].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[27].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[27].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[27].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[28].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[28].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[28].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[28].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[29].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[29].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[29].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[29].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[30].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[30].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[30].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[30].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[31].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[31].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[31].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[31].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[32].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[32].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[32].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[32].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[33].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[33].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[33].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[33].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[34].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[34].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[34].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[34].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[35].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[35].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[35].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[35].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[36].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[36].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[36].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[36].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[37].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[37].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[37].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[37].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[38].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[38].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[38].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[38].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[39].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[39].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[39].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[39].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[40].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[40].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[40].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[40].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[41].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[41].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[41].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[41].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[42].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[42].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[42].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[42].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[43].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[43].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[43].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[43].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[44].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[44].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[44].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[44].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[45].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[45].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[45].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[45].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[46].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[46].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[46].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[46].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[47].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[47].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[47].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[47].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[48].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[48].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[48].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[48].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[49].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[49].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[49].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[49].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[4].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[4].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[50].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[50].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[50].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[50].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[51].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[51].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[51].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[51].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[52].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[52].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[52].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[52].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[53].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[53].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[53].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[53].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[54].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[54].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[54].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[54].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[55].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[55].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[55].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[55].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[56].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[56].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[56].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[56].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[57].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[57].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[57].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[57].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[58].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[58].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[58].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[58].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[59].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[59].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[59].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[59].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[5].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[5].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[60].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[60].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[60].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[60].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[61].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[61].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[61].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[61].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[62].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[62].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[62].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[62].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[63].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[63].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[63].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[63].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[6].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[6].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[7].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[7].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[8].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[8].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[8].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[8].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[9].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[9].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g1[9].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[10]),
    .ZN(\gen_shunt_g1[9].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[10].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[10].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[10].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[10].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[10].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[11].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[11].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[11].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[11].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[11].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[12].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[12].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[12].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[12].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[12].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[13].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[13].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[13].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[13].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[13].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[14].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[14].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[14].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[14].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[14].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[15].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[15].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[15].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[15].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[15].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[16].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[16].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[16].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[16].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[16].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[17].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[17].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[17].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[17].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[17].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[18].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[18].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[18].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[18].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[18].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[19].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[19].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[19].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[19].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[19].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[20].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[20].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[20].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[20].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[20].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[21].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[21].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[21].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[21].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[21].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[22].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[22].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[22].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[22].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[22].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[23].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[23].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[23].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[23].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[23].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[24].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[24].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[24].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[24].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[24].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[25].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[25].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[25].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[25].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[25].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[26].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[26].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[26].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[26].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[26].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[27].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[27].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[27].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[27].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[27].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[28].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[28].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[28].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[28].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[28].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[29].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[29].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[29].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[29].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[29].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[2].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[30].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[30].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[30].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[30].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[30].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[31].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[31].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[31].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[31].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[31].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[3].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[4].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[5].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[6].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[7].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[8].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[8].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[8].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[8].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[8].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[9].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[9].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[9]),
    .ZN(\gen_shunt_g2[9].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g2[9].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[8]),
    .ZN(\gen_shunt_g2[9].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[10].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[10].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[10].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[10].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[10].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[11].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[11].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[11].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[11].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[11].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[12].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[12].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[12].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[12].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[12].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[13].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[13].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[13].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[13].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[13].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[14].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[14].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[14].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[14].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[14].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[15].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[15].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[15].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[15].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[15].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[2].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[3].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[4].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[5].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[6].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[7].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[8].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[8].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[8].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[8].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[8].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[9].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[9].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[7]),
    .ZN(\gen_shunt_g3[9].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g3[9].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[6]),
    .ZN(\gen_shunt_g3[9].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[2].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[3].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[4].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[5].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[6].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[5]),
    .ZN(\gen_shunt_g4[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g4[7].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[4]),
    .ZN(\gen_shunt_g4[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[1].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[1].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[2].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[2].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[3].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g5[3].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[3]),
    .ZN(\gen_shunt_g5[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[0].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_n1  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_n2  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_p1  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[2]),
    .ZN(\gen_shunt_g6[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g6[1].u_shunt_p2  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[1]),
    .ZN(\gen_shunt_g6[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[0].u_shunt_n  (.A1(cap_shunt_n),
    .A2(cap_shunt_n),
    .B(tune_shunt[0]),
    .ZN(\gen_shunt_g7[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_g7[0].u_shunt_p  (.A1(cap_shunt_p),
    .A2(cap_shunt_p),
    .B(tune_shunt[0]),
    .ZN(\gen_shunt_g7[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[2].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[3].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[4].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[5].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[6].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyn1  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyp1  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[4]),
    .ZN(\gen_shunt_gy_g1[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g1[7].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[3]),
    .ZN(\gen_shunt_gy_g1[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[2].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g2[3].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[2]),
    .ZN(\gen_shunt_gy_g2[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[0].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyn2  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g3[1].u_shunt_gyp2  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[1]),
    .ZN(\gen_shunt_gy_g3[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g4[0].u_shunt_n  (.A1(cap_shunt_gyn),
    .A2(cap_shunt_gyn),
    .B(tune_shunt_gy[0]),
    .ZN(\gen_shunt_gy_g4[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \gen_shunt_gy_g4[0].u_shunt_p  (.A1(cap_shunt_gyp),
    .A2(cap_shunt_gyp),
    .B(tune_shunt_gy[0]),
    .ZN(\gen_shunt_gy_g4[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[0].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[10].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[10].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[10].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[10].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[10].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[11].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[11].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[11].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[11].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[11].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[12].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[12].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[12].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[12].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[12].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[13].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[13].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[13].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[13].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[13].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[14].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[14].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[14].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[14].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[14].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[15].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[15].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[15].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[15].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[15].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[1].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[2].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[3].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[4].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[5].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[6].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[7].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[8].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[8].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[8].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[8].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[8].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[9].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[9].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[7]),
    .ZN(\gen_shunt_gygy_g1[9].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g1[9].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[6]),
    .ZN(\gen_shunt_gygy_g1[9].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[0].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[1].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[2].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[2].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[2].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[3].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[3].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[3].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[4].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[4].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[4].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[4].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[4].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[5].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[5].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[5].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[5].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[5].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[6].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[6].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[6].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[6].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[6].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[7].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[7].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[5]),
    .ZN(\gen_shunt_gygy_g2[7].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g2[7].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[4]),
    .ZN(\gen_shunt_gygy_g2[7].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[2].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[2].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[2].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[2].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[3].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[3].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g3[3].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[3]),
    .ZN(\gen_shunt_gygy_g3[3].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[0].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[0].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[0].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[1].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyn2  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[1].d4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[2]),
    .ZN(\gen_shunt_gygy_g4[1].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g4[1].u_series_gygyp2  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[1]),
    .ZN(\gen_shunt_gygy_g4[1].d3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g5[0].u_series_gygyn1  (.A1(cap_series_gygyn),
    .A2(cap_series_gygyn),
    .B(tune_series_gygy[0]),
    .ZN(\gen_shunt_gygy_g5[0].d2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \gen_shunt_gygy_g5[0].u_series_gygyp1  (.A1(cap_series_gygyp),
    .A2(cap_series_gygyp),
    .B(tune_series_gygy[0]),
    .ZN(\gen_shunt_gygy_g5[0].d1 ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_687 ();
endmodule

