VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 5tc_flat
  CLASS BLOCK ;
  FOREIGN 5tc_flat ;
  ORIGIN -0.490 -0.820 ;
  SIZE 2.920 BY 20.480 ;
END 5tc_flat
END LIBRARY

