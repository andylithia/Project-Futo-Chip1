magic
tech sky130A
magscale 1 2
timestamp 1669997259
<< dnwell >>
rect -2000 -2000 18000 18000
<< nwell >>
rect -2080 17794 18080 18080
rect -2080 -1794 -1794 17794
rect 17794 -1794 18080 17794
rect -2080 -2080 18080 -1794
<< nsubdiff >>
rect -2043 18023 18043 18043
rect -2043 17989 -1963 18023
rect 17963 17989 18043 18023
rect -2043 17969 18043 17989
rect -2043 17963 -1969 17969
rect -2043 -1963 -2023 17963
rect -1989 -1963 -1969 17963
rect -2043 -1969 -1969 -1963
rect 17969 17963 18043 17969
rect 17969 -1963 17989 17963
rect 18023 -1963 18043 17963
rect 17969 -1969 18043 -1963
rect -2043 -1989 18043 -1969
rect -2043 -2023 -1963 -1989
rect 17963 -2023 18043 -1989
rect -2043 -2043 18043 -2023
<< nsubdiffcont >>
rect -1963 17989 17963 18023
rect -2023 -1963 -1989 17963
rect 17989 -1963 18023 17963
rect -1963 -2023 17963 -1989
<< locali >>
rect -2023 17989 -1963 18023
rect 17963 17989 18023 18023
rect -2023 17963 -1989 17989
rect -2023 -1989 -1989 -1963
rect 17989 17963 18023 17989
rect 17989 -1989 18023 -1963
rect -2023 -2023 -1963 -1989
rect 17963 -2023 18023 -1989
<< end >>
