// This is the unpowered netlist.
module gyrator (nbus,
    nload,
    pbus,
    pload);
 inout nbus;
 inout nload;
 inout pbus;
 inout pload;


 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[0].fbn  (.I(nload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[0].fbp  (.I(pload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[1].fbn  (.I(nload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[1].fbp  (.I(pload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[2].fbn  (.I(nload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[2].fbp  (.I(pload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[3].fbn  (.I(nload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_FB[3].fbp  (.I(pload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[0].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[0].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[1].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[1].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[2].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[2].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[3].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[3].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[4].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[4].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[5].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[5].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[6].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[6].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[7].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[7].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[8].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[8].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[9].thrun  (.I(pbus),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_T[9].thrup  (.I(nbus),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[0].crossn  (.I(pload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[0].crossp  (.I(nload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[1].crossn  (.I(pload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[1].crossp  (.I(nload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[2].crossn  (.I(pload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[2].crossp  (.I(nload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[3].crossn  (.I(pload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[3].crossp  (.I(nload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[4].crossn  (.I(pload),
    .ZN(nload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_f.gen_X[4].crossp  (.I(nload),
    .ZN(pload));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[0].fbn  (.I(nbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[0].fbp  (.I(pbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[1].fbn  (.I(nbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[1].fbp  (.I(pbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[2].fbn  (.I(nbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[2].fbp  (.I(pbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[3].fbn  (.I(nbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_FB[3].fbp  (.I(pbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[0].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[0].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[1].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[1].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[2].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[2].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[3].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[3].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[4].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[4].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[5].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[5].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[6].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[6].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[7].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[7].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[8].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[8].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[9].thrun  (.I(nload),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_T[9].thrup  (.I(pload),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[0].crossn  (.I(pbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[0].crossp  (.I(nbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[1].crossn  (.I(pbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[1].crossp  (.I(nbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[2].crossn  (.I(pbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[2].crossp  (.I(nbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[3].crossn  (.I(pbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[3].crossp  (.I(nbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[4].crossn  (.I(pbus),
    .ZN(nbus));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_nauta_r.gen_X[4].crossp  (.I(nbus),
    .ZN(pbus));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_98 ();
endmodule

