magic
tech gf180mcuC
magscale 1 10
timestamp 1669581115
<< error_p >>
rect -34 38 -23 84
rect -118 -54 -107 -8
rect 50 -54 61 -8
<< pwell >>
rect -144 -121 144 121
<< nmos >>
rect -28 -53 28 -9
<< ndiff >>
rect -120 -8 -48 5
rect -120 -54 -107 -8
rect -61 -9 -48 -8
rect 48 -8 120 5
rect 48 -9 61 -8
rect -61 -53 -28 -9
rect 28 -53 61 -9
rect -61 -54 -48 -53
rect -120 -67 -48 -54
rect 48 -54 61 -53
rect 107 -54 120 -8
rect 48 -67 120 -54
<< ndiffc >>
rect -107 -54 -61 -8
rect 61 -54 107 -8
<< polysilicon >>
rect -36 84 36 97
rect -36 38 -23 84
rect 23 38 36 84
rect -36 25 36 38
rect -28 -9 28 25
rect -28 -97 28 -53
<< polycontact >>
rect -23 38 23 84
<< metal1 >>
rect -34 38 -23 84
rect 23 38 34 84
rect -118 -54 -107 -8
rect -61 -54 -50 -8
rect 50 -54 61 -8
rect 107 -54 118 -8
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.22 l 0.280 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
