* NGSPICE file created from gf180mcu_fd_io__asig_5p0_flat.ext - technology: gf180mcuC

.subckt gf180mcu_fd_io__asig_5p0_flat ASIG5V DVDD DVSS VDD VSS
X0 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X1 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X2 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D0 DVSS ASIG5V diode_nd2ps_06v0 pj=0.106n area=0.15n
X3 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X4 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X5 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X6 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X7 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X8 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D1 DVSS ASIG5V diode_nd2ps_06v0 pj=0.106n area=0.15n
D2 ASIG5V DVDD diode_pd2nw_06v0 pj=0.106n area=0.15n
X9 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X10 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X11 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X12 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X13 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X14 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X15 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X16 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X17 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X18 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X19 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D3 ASIG5V DVDD diode_pd2nw_06v0 pj=0.106n area=0.15n
D4 DVSS ASIG5V diode_nd2ps_06v0 pj=0.106n area=0.15n
X20 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X21 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D5 ASIG5V DVDD diode_pd2nw_06v0 pj=0.106n area=0.15n
X22 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X23 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X24 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X25 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D6 DVSS DVDD diode_nd2ps_06v0 pj=82p area=40p
X26 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X27 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X28 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X29 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D7 DVSS DVDD diode_nd2ps_06v0 pj=82p area=40p
D8 DVSS ASIG5V diode_nd2ps_06v0 pj=0.106n area=0.15n
X30 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D9 DVSS DVDD diode_nd2ps_06v0 pj=82p area=40p
X31 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D10 ASIG5V DVDD diode_pd2nw_06v0 pj=0.106n area=0.15n
X32 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
D11 DVSS DVDD diode_nd2ps_06v0 pj=82p area=40p
X33 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X34 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X35 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
C0 DVSS DVDD 1.56p
C1 VDD ASIG5V 21.9f
C2 DVSS ASIG5V 0.486p
C3 DVDD ASIG5V 0.626p
C4 DVSS VDD 51f
C5 VDD DVDD 48.2f
C6 VDD VSS 36.1f
C7 ASIG5V VSS 0.151p
C8 DVDD VSS 0.479p
C9 DVSS VSS 0.361p
.ends
