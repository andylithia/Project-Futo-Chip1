magic
tech gf180mcuC
magscale 1 5
timestamp 1669830058
<< obsm1 >>
rect 672 1538 9376 4342
<< metal2 >>
rect 1232 5600 1288 6000
rect 3696 5600 3752 6000
rect 6160 5600 6216 6000
rect 8624 5600 8680 6000
rect 1232 0 1288 400
rect 3696 0 3752 400
rect 6160 0 6216 400
rect 8624 0 8680 400
<< obsm2 >>
rect 910 5570 1202 5600
rect 1318 5570 3666 5600
rect 3782 5570 6130 5600
rect 6246 5570 8594 5600
rect 8710 5570 9362 5600
rect 910 430 9362 5570
rect 910 400 1202 430
rect 1318 400 3666 430
rect 3782 400 6130 430
rect 6246 400 8594 430
rect 8710 400 9362 430
<< metal3 >>
rect 0 4424 400 4480
rect 9600 4424 10000 4480
rect 0 1456 400 1512
rect 9600 1456 10000 1512
<< obsm3 >>
rect 430 4394 9570 4466
rect 400 1542 9600 4394
rect 430 1470 9570 1542
<< metal4 >>
rect 1670 1538 1830 4342
rect 2748 1538 2908 4342
rect 3826 1538 3986 4342
rect 4904 1538 5064 4342
rect 5982 1538 6142 4342
rect 7060 1538 7220 4342
rect 8138 1538 8298 4342
rect 9216 1538 9376 4342
<< labels >>
rlabel metal3 s 0 1456 400 1512 6 enable
port 1 nsew signal input
rlabel metal3 s 9600 4424 10000 4480 6 outn
port 2 nsew signal bidirectional
rlabel metal3 s 9600 1456 10000 1512 6 outp
port 3 nsew signal bidirectional
rlabel metal3 s 0 4424 400 4480 6 signal
port 4 nsew signal input
rlabel metal2 s 1232 0 1288 400 6 trim_n[0]
port 5 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 trim_n[1]
port 6 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 trim_n[2]
port 7 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 trim_n[3]
port 8 nsew signal input
rlabel metal2 s 1232 5600 1288 6000 6 trim_p[0]
port 9 nsew signal input
rlabel metal2 s 3696 5600 3752 6000 6 trim_p[1]
port 10 nsew signal input
rlabel metal2 s 6160 5600 6216 6000 6 trim_p[2]
port 11 nsew signal input
rlabel metal2 s 8624 5600 8680 6000 6 trim_p[3]
port 12 nsew signal input
rlabel metal4 s 1670 1538 1830 4342 6 vdd
port 13 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 4342 6 vdd
port 13 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 4342 6 vdd
port 13 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 4342 6 vdd
port 13 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 4342 6 vss
port 14 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 4342 6 vss
port 14 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 4342 6 vss
port 14 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 4342 6 vss
port 14 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 6000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 151602
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/injector/runs/22_11_30_12_40/results/signoff/injector.magic.gds
string GDS_START 34854
<< end >>

