* NGSPICE file created from gf180mcu_fd_io__bi_t.ext - technology: gf180mcuC

.subckt gf180mcu_fd_io__bi_t DVDD DVSS PAD PU SL A Y PDRV1 PDRV0 PD CS OE IE VDD VSS
X0 a_11617_50285# SL VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
D0 DVSS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN diode_nd2ps_06v0 pj=42p area=20p
X1 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_8850_42732# DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X2 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X3 a_4157_63027# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD DVDD pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X4 a_2031_61071# a_1751_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
X5 a_12966_56686# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X6 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X7 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X8 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<0> DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X9 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X10 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_y_<0> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
D1 IE VDD diode_pd2nw_06v0 pj=4p area=1p
X11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X12 PAD GF_NI_BI_T_BASE_0.pdrive_y_<0> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.111n pd=85.6u as=11.2p ps=80.6u w=40u l=0.7u  
X13 GF_NI_BI_T_BASE_0.pdrive_y_<1> DVDD GF_NI_BI_T_BASE_0.pdrive_x_<1> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X14 a_5463_64256# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_4235_64204# DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X15 GF_NI_BI_T_BASE_0.ndrive_y_<0> DVSS GF_NI_BI_T_BASE_0.ndrive_x_<0> DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X16 PAD GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.144n pd=83.6u as=10.6p ps=76.6u w=38u l=1.15u  
X17 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_11294_42688# DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X18 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X19 a_5463_64256# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X20 PU a_12527_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X21 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X22 VDD PU a_12715_59749# VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X23 DVSS a_3891_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X24 a_2591_61071# a_2311_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
X25 PAD GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.111n pd=85.6u as=11.2p ps=80.6u w=40u l=0.7u  
X26 GF_NI_BI_T_BASE_0.ndrive_x_<3> a_12354_42732# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X27 GF_NI_BI_T_BASE_0.ndrive_Y_<1> a_5346_42732# DVDD DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X28 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X29 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X30 a_1260_51889# PDRV0 VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X31 a_7790_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X32 DVSS a_11294_42688# GF_NI_BI_T_BASE_0.pdrive_y_<3> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X33 a_5575_63014# a_4157_63027# DVSS DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X34 PAD GF_NI_BI_T_BASE_0.ndrive_x_<0> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.144n pd=83.6u as=10.6p ps=76.6u w=38u l=1.15u  
X35 DVSS a_12354_42732# GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X36 a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X37 DVSS a_4157_63027# a_5575_63014# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X38 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X39 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_7790_42688# DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X40 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_6824_66100# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X41 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X42 DVSS a_7790_42688# GF_NI_BI_T_BASE_0.ndrive_y_<2> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X43 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X44 DVDD a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X45 PAD GF_NI_BI_T_BASE_0.pdrive_x_<3> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.111n pd=85.6u as=11.2p ps=80.6u w=40u l=0.7u  
X46 a_3891_66144# IE VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X47 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X48 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=1.54p ps=7.88u w=3.5u l=0.7u
X49 DVSS a_12068_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X50 GF_NI_BI_T_BASE_0.pdrive_y_<1> a_4286_42688# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X51 DVDD a_1842_42732# GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X52 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z a_9135_66144# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X53 a_1191_61071# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z DVDD DVDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X54 DVDD a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_y_<2> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X55 DVSS a_2947_62989# a_3430_64204# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X56 DVSS a_8953_50157# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X57 DVSS a_1842_42732# GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
D2 VSS OE diode_pd2nw_06v0 pj=1.92p area=0.23p
X58 GF_NI_BI_T_BASE_0.pdrive_y_<0> a_1842_42732# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X59 a_5346_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X60 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X61 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_4157_63027# DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X62 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN a_1842_42732# DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X63 DVDD a_12354_42732# GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X64 DVDD a_4286_42688# GF_NI_BI_T_BASE_0.pdrive_y_<1> DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X65 VDD CS a_6824_66100# VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X66 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X67 a_5463_64256# a_3430_64204# DVDD DVSS nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
X68 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<3> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X69 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X70 a_2031_61071# a_2311_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
X71 a_6504_51889# OE a_6504_50201# VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X72 PAD GF_NI_BI_T_BASE_0.pdrive_y_<2> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.111n pd=85.6u as=11.2p ps=80.6u w=40u l=0.7u  
X73 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<3> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X74 GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X75 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<3> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X76 a_4235_64204# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=1.41p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X77 a_6504_50201# VDD VSS VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X78 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<2> DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X79 VDD PDRV1 a_3961_50157# VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X80 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z a_12527_59749# a_12715_59749# VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X81 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X82 GF_NI_BI_T_BASE_0.pdrive_y_<0> a_1842_42732# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X83 a_3961_50157# OE VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X84 VDD OE a_9197_50157# VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X85 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X86 a_9197_50157# A VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X87 GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X88 VSS PU a_12966_56686# VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X89 a_11617_50285# SL VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X90 a_2591_61071# a_2871_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
X91 DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<3> PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.6p pd=76.6u as=0.144n ps=83.6u w=38u l=1.15u  
X92 VDD PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X93 GF_NI_BI_T_BASE_0.ndrive_Y_<1> a_5346_42732# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X94 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z a_9536_64061# VDD VDD pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
X95 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<3> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.2p pd=80.6u as=0.111n ps=85.6u w=40u l=0.7u  
X96 DVDD a_11294_42688# GF_NI_BI_T_BASE_0.pdrive_x_<3> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X97 a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS DVSS nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
D3 VSS OE diode_pd2nw_06v0 pj=1.92p area=0.23p
D4 VSS VDD diode_pd2nw_06v0 pj=1.92p area=0.23p
X98 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_4286_42688# DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X99 a_11294_42688# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_12354_42732# DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X100 GF_NI_BI_T_BASE_0.pdrive_y_<1> a_4286_42688# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X101 a_5463_64256# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_4235_64204# DVSS nfet_06v0 ad=1.17p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X102 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_5463_64256# DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X103 GF_NI_BI_T_BASE_0.pdrive_x_<3> a_11294_42688# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X104 a_1260_51889# OE a_1260_50201# VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X105 DVSS GF_NI_BI_T_BASE_0.ndrive_y_<0> PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.6p pd=76.6u as=0.144n ps=83.6u w=38u l=1.15u  
X106 DVSS a_6824_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X107 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X108 VDD a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
X109 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB a_1842_42732# DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X110 DVSS a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X111 GF_NI_BI_T_BASE_0.ndrive_y_<2> a_7790_42688# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X112 DVDD a_3891_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
D5 A VDD diode_pd2nw_06v0 pj=4p area=1p
X113 GF_NI_BI_T_BASE_0.pdrive_y_<2> a_8850_42732# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X114 a_7790_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_8850_42732# DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X115 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_4157_63027# DVDD pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X116 a_3430_64204# a_2947_62989# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X117 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_2871_53829# DVDD ppolyf_u r_width=0.8u r_length=23u
X118 DVSS a_11617_50285# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X119 a_4235_64204# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_5463_64256# DVSS nfet_06v0 ad=0.689p pd=3.17u as=1.17p ps=6.18u w=2.65u l=0.7u
X120 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X121 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X122 VSS PU a_12715_59749# VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X123 DVSS a_6504_51889# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X124 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<0> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X125 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<1> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.2p pd=80.6u as=0.111n ps=85.6u w=40u l=0.7u  
X126 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X127 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X128 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X129 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X130 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z a_12068_66100# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X131 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS VSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X132 DVDD a_8953_50157# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X133 a_11294_42688# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN a_12354_42732# DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X134 a_4286_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X135 GF_NI_BI_T_BASE_0.pdrive_y_<3> DVDD GF_NI_BI_T_BASE_0.pdrive_x_<3> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X136 DVSS a_4286_42688# GF_NI_BI_T_BASE_0.pdrive_y_<1> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X137 GF_NI_BI_T_BASE_0.pdrive_y_<2> a_8850_42732# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X138 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X139 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_3891_66144# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X140 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VDD pfet_06v0 ad=1.54p pd=7.88u as=0.91p ps=4.02u w=3.5u l=0.7u
X141 PAD GF_NI_BI_T_BASE_0.ndrive_x_<2> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.144n pd=83.6u as=10.6p ps=76.6u w=38u l=1.15u  
X142 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X143 DVDD a_12068_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X144 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X145 a_5575_63014# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X146 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X147 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z a_9135_66144# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X148 a_1191_61071# a_1191_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
D6 VSS OE diode_pd2nw_06v0 pj=1.92p area=0.23p
D7 SL VDD diode_pd2nw_06v0 pj=4p area=1p
X149 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_y_<2> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X150 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_12068_66100# VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X151 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X152 GF_NI_BI_T_BASE_0.ndrive_y_<2> DVSS GF_NI_BI_T_BASE_0.ndrive_x_<2> DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X153 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X154 GF_NI_BI_T_BASE_0.pdrive_x_<0> a_1842_42732# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X155 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X156 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_11617_50285# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X157 DVSS a_782_42688# GF_NI_BI_T_BASE_0.ndrive_x_<0> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X158 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X159 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X160 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_5346_42732# DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
D8 PU VDD diode_pd2nw_06v0 pj=4p area=1p
X161 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_4235_64204# DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X162 a_12527_59749# PD VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X163 GF_NI_BI_T_BASE_0.pdrive_y_<3> a_11294_42688# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X164 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<1> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X165 DVDD a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X166 a_4235_64204# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=1.41p ps=7.28u w=3.2u l=0.7u
X167 a_1842_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X168 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<0> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.2p pd=80.6u as=0.111n ps=85.6u w=40u l=0.7u  
X169 a_3891_66144# IE VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X170 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z PD a_12715_59749# VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X171 a_12354_42732# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X172 DVDD a_11294_42688# GF_NI_BI_T_BASE_0.pdrive_y_<3> DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X173 VDD OE a_6504_51889# VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X174 PAD GF_NI_BI_T_BASE_0.pdrive_x_<1> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.111n pd=85.6u as=11.2p ps=80.6u w=40u l=0.7u  
X175 a_6504_51889# VDD VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X176 DVSS a_12354_42732# GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X177 a_2947_62989# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS DVSS nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X178 DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<1> PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.6p pd=76.6u as=0.144n ps=83.6u w=38u l=1.15u  
D9 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN DVDD diode_pd2nw_06v0 pj=42p area=20p
X179 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_3961_50157# DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X180 GF_NI_BI_T_BASE_0.ndrive_y_<0> a_782_42688# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X181 DVDD a_6824_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X182 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD DVDD ppolyf_u r_width=2.5u r_length=2.8u
X183 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X184 DVSS a_1260_51889# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X185 a_2947_62989# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD DVDD pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X186 a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X187 a_3430_64204# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X188 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_9536_64061# DVSS nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X189 DVDD a_6504_51889# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X190 GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X191 DVDD a_4286_42688# GF_NI_BI_T_BASE_0.pdrive_x_<1> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X192 a_5575_63014# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN DVDD DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X193 a_1471_61071# a_1191_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
D10 DVSS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN diode_nd2ps_06v0 pj=42p area=20p
X194 a_1260_50201# PDRV0 VSS VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X195 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X196 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z a_9536_64061# VDD VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X197 DVSS GF_NI_BI_T_BASE_0.ndrive_y_<2> PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.6p pd=76.6u as=0.144n ps=83.6u w=38u l=1.15u  
X198 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<1> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.2p pd=80.6u as=0.111n ps=85.6u w=40u l=0.7u  
X199 GF_NI_BI_T_BASE_0.ndrive_x_<1> a_5346_42732# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X200 DVDD GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_5575_63014# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X201 GF_NI_BI_T_BASE_0.ndrive_Y_<3> a_12354_42732# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X202 DVSS a_5346_42732# GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X203 VDD a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X204 a_8953_50157# a_9197_50157# DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X205 DVDD a_11617_50285# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X206 GF_NI_BI_T_BASE_0.pdrive_y_<3> a_11294_42688# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X207 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z a_12000_56686# VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X208 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X209 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X210 PU PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
D11 VSS PDRV1 diode_pd2nw_06v0 pj=1.92p area=0.23p
X211 GF_NI_BI_T_BASE_0.ndrive_Y_<3> a_12354_42732# DVDD DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X212 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X213 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z a_12068_66100# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X214 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X215 GF_NI_BI_T_BASE_0.ndrive_x_<0> a_782_42688# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X216 DVSS a_7790_42688# GF_NI_BI_T_BASE_0.ndrive_x_<2> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X217 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X218 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X219 VDD OE a_1260_51889# VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X220 VSS CS a_6824_66100# VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X221 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X222 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_3891_66144# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X223 a_8850_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
D12 PD VDD diode_pd2nw_06v0 pj=4p area=1p
X224 VSS a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X225 PAD GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.144n pd=83.6u as=10.6p ps=76.6u w=38u l=1.15u  
X226 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<3> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.2p pd=80.6u as=0.111n ps=85.6u w=40u l=0.7u  
X227 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z a_9536_64061# VSS VSS nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
X228 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
D13 VSS PDRV0 diode_pd2nw_06v0 pj=1.92p area=0.23p
X229 a_4286_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_5346_42732# DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X230 DVDD a_1842_42732# GF_NI_BI_T_BASE_0.pdrive_y_<0> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X231 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD DVDD ppolyf_u r_width=2.5u r_length=2.8u
X232 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_1842_42732# DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X233 a_5463_64256# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X234 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X235 DVDD a_5346_42732# GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X236 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_6824_66100# DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X237 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X238 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_5463_64256# DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X239 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X240 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<2> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X241 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X242 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X243 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<1> DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X244 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X245 DVSS a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X246 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X247 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_5575_63014# DVDD pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X248 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X249 a_7790_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_8850_42732# DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
D14 CS VDD diode_pd2nw_06v0 pj=4p area=1p
X250 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<1> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X251 a_11294_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X252 GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X253 VSS PDRV1 a_5502_50201# VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X254 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_11617_50285# DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X255 GF_NI_BI_T_BASE_0.ndrive_y_<2> a_7790_42688# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X256 DVDD a_782_42688# GF_NI_BI_T_BASE_0.ndrive_y_<0> DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X257 a_12000_56686# PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X258 a_5502_50201# OE a_3961_50157# VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X259 a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X260 VSS OE a_10720_50201# VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X261 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X262 a_10720_50201# A a_9197_50157# VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X263 GF_NI_BI_T_BASE_0.ndrive_x_<2> a_7790_42688# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X264 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A PD VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X265 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X266 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<2> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.2p pd=80.6u as=0.111n ps=85.6u w=40u l=0.7u  
X267 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X268 a_1471_61071# a_1751_53829# DVDD ppolyf_u r_width=0.8u r_length=35.7u
X269 a_12527_59749# PD VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X270 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_3961_50157# DVDD DVDD pfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X271 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X272 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X273 DVDD a_1260_51889# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.9u w=6u l=0.7u
X274 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN a_782_42688# DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X275 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_2947_62989# DVSS nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X276 PAD GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.111n pd=85.6u as=11.2p ps=80.6u w=40u l=0.7u  
X277 GF_NI_BI_T_BASE_0.pdrive_x_<2> a_8850_42732# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=3.12p ps=12.5u w=12u l=0.7u
X278 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_2947_62989# a_4157_63027# DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X279 a_1191_61071# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB DVSS DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X280 DVSS a_782_42688# GF_NI_BI_T_BASE_0.ndrive_y_<0> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X281 a_4235_64204# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_5463_64256# DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
D15 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN DVDD diode_pd2nw_06v0 pj=42p area=20p
X282 GF_NI_BI_T_BASE_0.ndrive_y_<0> a_782_42688# DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X283 a_4286_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_5346_42732# DVDD pfet_06v0 ad=5.28p pd=24.9u as=3.12p ps=12.5u w=12u l=0.7u
X284 GF_NI_BI_T_BASE_0.pdrive_x_<1> a_4286_42688# DVDD DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X285 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X286 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_12068_66100# VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X287 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD DVDD ppolyf_u r_width=2.5u r_length=2.8u
X288 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_12354_42732# DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X289 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_4235_64204# DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X290 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_2947_62989# DVDD pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X291 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X292 a_4235_64204# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X293 DVDD a_7790_42688# GF_NI_BI_T_BASE_0.ndrive_y_<2> DVDD pfet_06v0 ad=3.12p pd=12.5u as=5.28p ps=24.9u w=12u l=0.7u
X294 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD DVDD ppolyf_u r_width=2.5u r_length=2.8u
X295 a_8953_50157# a_9197_50157# DVDD DVDD pfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
X296 DVSS a_5346_42732# GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS nfet_06v0 ad=2.64p pd=12.9u as=1.56p ps=6.52u w=6u l=0.7u
C0 a_1191_61071# PD 0.106f
C1 a_3891_66144# DVSS 1.41f
C2 a_12527_59749# SL 0.00318f
C3 a_12715_59749# VDD 0.74f
C4 DVSS a_3430_64204# 2.04f
C5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_7790_42688# 0.519f
C6 a_10720_50201# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 4.99e-19
C7 a_9135_66144# PD 0.0222f
C8 a_6824_66100# PD 7.47e-19
C9 OE VDD 9.92f
C10 a_9197_50157# SL 0.0108f
C11 a_4286_42688# PDRV1 0.0019f
C12 GF_NI_BI_T_BASE_0.pdrive_y_<0> DVDD 18f
C13 Y SL 0.122f
C14 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 1.11f
C15 DVSS PDRV0 2.24f
C16 a_6824_66100# a_5463_64256# 1.67e-19
C17 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.0352f
C18 A VDD 3.81f
C19 PD SL 0.00209f
C20 a_12000_56686# PD 0.0273f
C21 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_4286_42688# 0.505f
C22 a_3961_50157# DVDD 0.492f
C23 GF_NI_BI_T_BASE_0.ndrive_Y_<1> a_1842_42732# 0.00137f
C24 a_3891_66144# a_3430_64204# 0.00136f
C25 a_2947_62989# a_4235_64204# 1.21e-19
C26 a_12715_59749# a_12527_59749# 0.59f
C27 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z SL 0.586f
C28 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z a_12000_56686# 0.0273f
C29 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_8953_50157# 1.29e-20
C30 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN GF_NI_BI_T_BASE_0.ndrive_Y_<1> 3.42e-19
C31 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.ndrive_Y_<1> 3.42e-19
C32 DVDD a_12068_66100# 1.29f
C33 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.823f
C34 PAD DVDD 0.312p
C35 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 2.19f
C36 PU VDD 3.27f
C37 OE a_9197_50157# 0.182f
C38 a_12715_59749# PD 0.1f
C39 OE Y 2.47f
C40 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.858f
C41 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.00359f
C42 a_12966_56686# DVSS 0.0121f
C43 A a_9197_50157# 0.652f
C44 A Y 0.0658f
C45 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB VDD 0.135f
C46 a_12715_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 1.12f
C47 GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVSS 16.1f
C48 DVDD a_12354_42732# 5.62f
C49 a_782_42688# GF_NI_BI_T_BASE_0.ndrive_x_<0> 1.8f
C50 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<1> 30.2f
C51 a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_x_<3> 5.58e-20
C52 a_6504_51889# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 0.00882f
C53 OE a_6504_50201# 0.0328f
C54 PU a_12527_59749# 0.272f
C55 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL PDRV1 2.27e-19
C56 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN PDRV1 0.0864f
C57 a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 4.06e-20
C58 PU Y 0.228f
C59 a_10720_50201# SL 2.49e-19
C60 a_6504_51889# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 0.609f
C61 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.809f
C62 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 8.49f
C63 PU PD 0.774f
C64 a_5346_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.00353f
C65 a_1260_51889# a_1260_50201# 0.152f
C66 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.0045f
C67 a_782_42688# a_1842_42732# 1.9f
C68 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<2> 1.53e-19
C69 a_8850_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.0263f
C70 PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 1.31f
C71 GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS 9.78f
C72 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 4.77f
C73 DVSS a_2947_62989# 0.664f
C74 a_7790_42688# DVDD 5.24f
C75 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_11294_42688# 0.012f
C76 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.346f
C77 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 2.3f
C78 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 0.561f
C79 VDD GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.977f
C80 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 0.00151f
C81 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 2.47f
C82 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 0.042f
C83 PDRV0 a_1191_53829# 0.0456f
C84 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_9536_64061# 0.0665f
C85 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<2> 30.2f
C86 OE a_10720_50201# 0.0273f
C87 a_8850_42732# GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.0351f
C88 DVSS PDRV1 3.25f
C89 A a_10720_50201# 0.0273f
C90 a_2947_62989# a_3430_64204# 0.217f
C91 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 0.00225f
C92 a_12068_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.00105f
C93 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 11f
C94 a_8953_50157# DVDD 1.06f
C95 a_5346_42732# GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.0268f
C96 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_11617_50285# 0.0167f
C97 a_2947_62989# PDRV0 9.62e-20
C98 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.584f
C99 PU IE 1.65e-19
C100 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 0.00773f
C101 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_y_<0> 1.13f
C102 DVSS GF_NI_BI_T_BASE_0.pdrive_y_<2> 2.51f
C103 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_4157_63027# 0.332f
C104 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PD 0.00202f
C105 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN a_11617_50285# 8.15e-19
C106 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z CS 0.054f
C107 DVSS a_11294_42688# 4.63f
C108 a_2031_61071# a_2591_61071# 0.0346f
C109 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL SL 3.57e-19
C110 PDRV0 PDRV1 6.88f
C111 a_5463_64256# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 2.1f
C112 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN a_2311_53829# 1.01e-19
C113 GF_NI_BI_T_BASE_0.ndrive_x_<0> DVDD 7.91f
C114 a_3961_50157# VDD 1.2f
C115 GF_NI_BI_T_BASE_0.pdrive_x_<0> a_4286_42688# 5.58e-20
C116 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB 0.615f
C117 a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.025f
C118 a_12068_66100# VDD 0.537f
C119 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB a_4286_42688# 0.0268f
C120 PAD VDD 1.41f
C121 DVSS a_1191_61071# 1.08f
C122 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.227f
C123 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.00109f
C124 DVSS GF_NI_BI_T_BASE_0.ndrive_y_<0> 12.2f
C125 a_9135_66144# DVSS 1.55f
C126 a_6824_66100# DVSS 1.43f
C127 a_1751_53829# a_1191_53829# 0.0346f
C128 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB a_1191_61071# 1.1f
C129 DVDD a_1842_42732# 4f
C130 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL A 5.38e-19
C131 a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB 0.027f
C132 DVDD GF_NI_BI_T_BASE_0.ndrive_y_<2> 11.7f
C133 DVSS SL 3.47f
C134 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A a_9536_64061# 0.152f
C135 DVSS a_12000_56686# 0.0149f
C136 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN DVDD 1.76f
C137 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB DVDD 1.3f
C138 a_1191_61071# a_3430_64204# 5.42e-20
C139 a_5346_42732# PAD 0.29f
C140 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.613f
C141 PAD a_9197_50157# 0.00324f
C142 a_1191_53829# PDRV1 0.0312f
C143 a_12068_66100# Y 8.4e-19
C144 a_6824_66100# a_3430_64204# 0.00135f
C145 a_1191_61071# PDRV0 0.195f
C146 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB DVDD 1.31f
C147 GF_NI_BI_T_BASE_0.pdrive_y_<1> a_4286_42688# 2.81f
C148 DVDD GF_NI_BI_T_BASE_0.ndrive_x_<3> 5.84f
C149 a_12715_59749# DVSS 0.378f
C150 a_5346_42732# GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.184f
C151 GF_NI_BI_T_BASE_0.ndrive_Y_<3> a_11294_42688# 1.27f
C152 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.361f
C153 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 9.57f
C154 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.0882f
C155 OE DVSS 3.49f
C156 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN DVDD 1.75f
C157 a_1751_53829# PDRV1 0.0095f
C158 DVDD a_1260_51889# 0.493f
C159 a_2947_62989# PDRV1 0.00291f
C160 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB a_12715_59749# 3.68e-20
C161 A DVSS 2.11f
C162 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_6504_51889# 7.24e-20
C163 DVSS GF_NI_BI_T_BASE_0.pdrive_x_<3> 5.57f
C164 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.00192f
C165 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.00332f
C166 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.862f
C167 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A CS 0.0325f
C168 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN a_4235_64204# 1.12f
C169 DVDD a_9536_64061# 0.416f
C170 PU DVSS 6.93f
C171 a_5346_42732# a_7790_42688# 0.032f
C172 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A PDRV1 0.00363f
C173 a_8953_50157# VDD 0.29f
C174 DVSS GF_NI_BI_T_BASE_0.pdrive_x_<0> 5.52f
C175 GF_NI_BI_T_BASE_0.pdrive_y_<0> a_4286_42688# 0.025f
C176 OE PDRV0 0.527f
C177 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.00656f
C178 a_12966_56686# SL 0.00398f
C179 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB PU 0.052f
C180 a_8850_42732# a_7790_42688# 1.9f
C181 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.00504f
C182 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<1> 1.53e-19
C183 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 17.3f
C184 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.0037f
C185 a_2031_61071# a_1471_61071# 0.0346f
C186 a_3891_66144# PU 3.68e-19
C187 a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.864f
C188 PU a_3430_64204# 0.0299f
C189 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.064f
C190 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A 0.753f
C191 DVDD a_2031_61071# 0.353f
C192 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_11294_42688# 0.492f
C193 a_1191_61071# a_2947_62989# 0.00101f
C194 DVSS GF_NI_BI_T_BASE_0.ndrive_x_<2> 11f
C195 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z a_1191_61071# 0.427f
C196 a_8953_50157# a_9197_50157# 0.589f
C197 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<3> 1.53e-19
C198 PU PDRV0 1.15f
C199 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.ndrive_y_<0> 10f
C200 a_4157_63027# DVDD 1.44f
C201 a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 8.53e-19
C202 CS DVDD 1.36f
C203 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.584f
C204 GF_NI_BI_T_BASE_0.pdrive_x_<1> a_4286_42688# 0.864f
C205 a_1191_61071# PDRV1 0.0921f
C206 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z SL 1.61e-19
C207 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB DVDD 0.584f
C208 GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVDD 17.8f
C209 GF_NI_BI_T_BASE_0.pdrive_y_<1> DVSS 2.58f
C210 OE a_1191_53829# 3.29e-19
C211 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 1.53e-19
C212 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.pdrive_x_<3> 4.4e-19
C213 DVSS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 33.9f
C214 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_9536_64061# 6.92e-19
C215 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_9536_64061# 0.52f
C216 a_5575_63014# a_4157_63027# 0.194f
C217 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD 3.54f
C218 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_3961_50157# 4.94e-20
C219 a_3961_50157# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.594f
C220 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.00192f
C221 a_12966_56686# PU 0.0273f
C222 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 1.62e-21
C223 a_6504_51889# DVDD 0.493f
C224 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB VDD 0.137f
C225 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN VDD 0.292f
C226 a_12715_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 3.11e-20
C227 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A DVDD 0.84f
C228 a_9536_64061# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 1.02f
C229 DVDD a_2591_61071# 0.373f
C230 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A SL 5.29e-20
C231 DVSS GF_NI_BI_T_BASE_0.pdrive_y_<3> 2.52f
C232 OE a_1751_53829# 5.33e-19
C233 a_3430_64204# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.064f
C234 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL PAD 0.599f
C235 PAD GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.11f
C236 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB VDD 0.137f
C237 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_5575_63014# 0.0121f
C238 A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 9.24e-21
C239 a_5346_42732# GF_NI_BI_T_BASE_0.ndrive_y_<2> 3.7e-19
C240 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN VDD 0.415f
C241 OE PDRV1 2.66f
C242 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_12354_42732# 0.33f
C243 a_1260_51889# VDD 1.19f
C244 GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS 2.4f
C245 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.0138f
C246 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.0551f
C247 a_8850_42732# GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.29f
C248 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_4157_63027# 0.575f
C249 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_4157_63027# 0.424f
C250 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.00329f
C251 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z CS 0.0455f
C252 a_3961_50157# DVSS 0.625f
C253 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.00648f
C254 PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 0.2f
C255 PU a_2947_62989# 2.31e-19
C256 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.0744f
C257 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_9197_50157# 1.6e-19
C258 A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.00133f
C259 a_9536_64061# VDD 1.48f
C260 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.00224f
C261 DVSS a_12068_66100# 1.43f
C262 a_782_42688# DVDD 5.46f
C263 a_8850_42732# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 1.8e-19
C264 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 0.0037f
C265 a_9135_66144# a_6824_66100# 0.0136f
C266 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB DVDD 1.74f
C267 PAD DVSS 0.239p
C268 a_5502_50201# VDD 0.012f
C269 PU PDRV1 0.0348f
C270 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.29f
C271 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN a_9197_50157# 0.00159f
C272 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 1.53f
C273 DVDD a_11617_50285# 0.988f
C274 a_8850_42732# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 2.31e-19
C275 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z 0.0032f
C276 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_7790_42688# 0.325f
C277 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_7790_42688# 2.3f
C278 GF_NI_BI_T_BASE_0.pdrive_x_<3> a_11294_42688# 0.718f
C279 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.00226f
C280 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB PDRV1 1.35e-19
C281 DVSS a_12354_42732# 2.76f
C282 DVSS GF_NI_BI_T_BASE_0.pdrive_x_<1> 4.81f
C283 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.00599f
C284 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.055f
C285 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.215f
C286 a_9536_64061# Y 0.00264f
C287 a_2031_61071# VDD 0.00125f
C288 a_9536_64061# PD 0.223f
C289 a_2871_53829# PDRV1 9.06e-19
C290 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.318f
C291 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A DVDD 0.852f
C292 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.737f
C293 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_8953_50157# 4.94e-20
C294 a_4157_63027# VDD 0.363f
C295 a_8953_50157# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 4.38e-19
C296 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.0694f
C297 a_2311_53829# DVDD 0.436f
C298 CS VDD 2.83f
C299 a_1842_42732# a_4286_42688# 0.00366f
C300 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 9.39e-21
C301 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.00656f
C302 a_12715_59749# SL 0.397f
C303 a_2947_62989# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 1.13f
C304 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.00138f
C305 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB a_11294_42688# 0.0268f
C306 OE SL 2.07f
C307 DVSS a_7790_42688# 2.82f
C308 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB VDD 0.00656f
C309 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.465f
C310 A SL 8.86f
C311 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PDRV1 0.0155f
C312 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVDD 1.63f
C313 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z VDD 0.172f
C314 GF_NI_BI_T_BASE_0.ndrive_x_<2> a_11294_42688# 0.00137f
C315 DVSS GF_NI_BI_T_BASE_0.pdrive_x_<2> 4.8f
C316 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.87f
C317 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.064f
C318 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0> 7.63e-19
C319 a_6824_66100# PU 3.68e-19
C320 a_6504_51889# VDD 1.29f
C321 a_9135_66144# PU 3.68e-19
C322 GF_NI_BI_T_BASE_0.ndrive_Y_<3> PAD 5.1f
C323 DVDD a_1471_61071# 0.352f
C324 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A VDD 2.05f
C325 a_1260_50201# VDD 0.012f
C326 a_2591_61071# VDD 0.00134f
C327 PU SL 1.24f
C328 CS PD 4.8f
C329 DVSS a_8953_50157# 0.734f
C330 a_5346_42732# GF_NI_BI_T_BASE_0.ndrive_Y_<1> 1.9f
C331 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.0694f
C332 a_4157_63027# a_5463_64256# 0.447f
C333 OE A 7.47f
C334 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.299f
C335 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.056f
C336 GF_NI_BI_T_BASE_0.ndrive_Y_<3> a_12354_42732# 1.92f
C337 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_1842_42732# 0.012f
C338 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_12527_59749# 0.139f
C339 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.00154f
C340 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z PD 0.0469f
C341 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.125f
C342 a_12715_59749# PU 0.841f
C343 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.11f
C344 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.ndrive_y_<2> 6.12e-19
C345 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z a_12068_66100# 0.771f
C346 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.00151f
C347 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 0.407f
C348 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.0115f
C349 GF_NI_BI_T_BASE_0.ndrive_x_<1> PAD 5.88f
C350 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 0.051f
C351 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_5463_64256# 0.00101f
C352 GF_NI_BI_T_BASE_0.ndrive_x_<0> DVSS 17.8f
C353 a_5575_63014# DVDD 1.29f
C354 GF_NI_BI_T_BASE_0.pdrive_y_<3> a_11294_42688# 2.92f
C355 OE PU 1.85f
C356 a_3961_50157# PDRV1 0.221f
C357 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A Y 0.109f
C358 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.056f
C359 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A PD 0.361f
C360 PU A 0.0977f
C361 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.0153f
C362 a_1191_61071# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.135f
C363 a_6504_51889# a_6504_50201# 0.152f
C364 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 0.247f
C365 a_3961_50157# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 5.93e-20
C366 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.00532f
C367 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.00106f
C368 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.865f
C369 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB VDD 0.137f
C370 a_4157_63027# IE 3.48e-20
C371 PAD PDRV1 7.17e-21
C372 a_6824_66100# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 9.14e-19
C373 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.157f
C374 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 0.906f
C375 CS IE 0.00244f
C376 VDD a_11617_50285# 0.969f
C377 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.545f
C378 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.713f
C379 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 0.0989f
C380 PAD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.107f
C381 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_1260_51889# 4.94e-20
C382 DVSS a_1842_42732# 4.61f
C383 OE a_2871_53829# 5.25e-19
C384 DVSS GF_NI_BI_T_BASE_0.ndrive_y_<2> 9.63f
C385 PAD GF_NI_BI_T_BASE_0.pdrive_y_<2> 10.2f
C386 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 2.26f
C387 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB DVSS 2.65f
C388 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z IE 0.0016f
C389 a_5346_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB 0.562f
C390 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD 2.37f
C391 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD 3.13f
C392 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.981f
C393 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.545f
C394 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.0511f
C395 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_12354_42732# 1.68f
C396 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VDD 3.26f
C397 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_8850_42732# 2.43f
C398 a_9197_50157# a_11617_50285# 0.00349f
C399 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 2.57f
C400 GF_NI_BI_T_BASE_0.ndrive_Y_<1> a_4286_42688# 1.27f
C401 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_y_<0> 2.38e-19
C402 DVSS GF_NI_BI_T_BASE_0.ndrive_x_<3> 12f
C403 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.00556f
C404 a_11294_42688# a_12354_42732# 1.9f
C405 a_5575_63014# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 0.00326f
C406 a_4157_63027# a_4235_64204# 0.228f
C407 a_5575_63014# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.531f
C408 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 2.65f
C409 DVSS a_1260_51889# 0.625f
C410 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A a_12527_59749# 0.0161f
C411 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB PDRV0 0.00682f
C412 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN PDRV0 0.0114f
C413 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z VDD 0.0339f
C414 PAD GF_NI_BI_T_BASE_0.ndrive_y_<0> 5.88f
C415 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_7790_42688# 1.68f
C416 PU GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.00486f
C417 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A PD 2.43f
C418 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_x_<3> 2.34f
C419 DVSS a_9536_64061# 1.24f
C420 a_12068_66100# SL 0.0347f
C421 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.0511f
C422 a_1471_61071# VDD 8.9e-19
C423 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_4235_64204# 0.576f
C424 a_7790_42688# GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.0268f
C425 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.737f
C426 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB a_9536_64061# 0.0842f
C427 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 0.402f
C428 DVDD VDD 49.7f
C429 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2> 2.31f
C430 a_1260_51889# PDRV0 0.222f
C431 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.00389f
C432 OE a_3961_50157# 0.77f
C433 a_8953_50157# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.517f
C434 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 3.37f
C435 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_Y_<1> 1.12f
C436 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN GF_NI_BI_T_BASE_0.ndrive_Y_<1> 3.42e-19
C437 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.00382f
C438 a_9536_64061# a_3430_64204# 6.63e-20
C439 a_11294_42688# GF_NI_BI_T_BASE_0.pdrive_x_<2> 5.58e-20
C440 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.737f
C441 OE a_12068_66100# 0.00128f
C442 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_6504_51889# 4.94e-20
C443 a_6504_51889# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 9.04e-20
C444 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_4286_42688# 2.43f
C445 a_12527_59749# DVDD 0.0715f
C446 OE PAD 1.53f
C447 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 1.39e-19
C448 a_5575_63014# VDD 1.09f
C449 DVSS a_2031_61071# 0.07f
C450 A a_12068_66100# 0.00442f
C451 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 0.36f
C452 a_5346_42732# DVDD 5.24f
C453 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0> 2.35f
C454 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_1260_50201# 8.26e-20
C455 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3> 10.3f
C456 DVDD a_9197_50157# 0.492f
C457 a_4157_63027# DVSS 0.763f
C458 PAD GF_NI_BI_T_BASE_0.pdrive_x_<3> 20.2f
C459 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 7.02e-19
C460 DVDD Y 2.1f
C461 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.298f
C462 DVSS CS 4.28f
C463 GF_NI_BI_T_BASE_0.ndrive_x_<1> a_1842_42732# 0.00245f
C464 a_8850_42732# DVDD 3.93f
C465 DVDD PD 2.85f
C466 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.159f
C467 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.737f
C468 DVDD a_5463_64256# 0.355f
C469 PU a_12068_66100# 9.13e-19
C470 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 6.12e-19
C471 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 6.12e-19
C472 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.024f
C473 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB DVSS 0.298f
C474 DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<1> 10.8f
C475 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z DVDD 0.775f
C476 a_3891_66144# a_4157_63027# 5.15e-20
C477 GF_NI_BI_T_BASE_0.pdrive_x_<3> a_12354_42732# 8.77e-19
C478 PAD GF_NI_BI_T_BASE_0.pdrive_x_<0> 20.2f
C479 a_1260_51889# a_1191_53829# 1.01e-19
C480 a_4157_63027# a_3430_64204# 1.99f
C481 a_3891_66144# CS 0.0206f
C482 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS 5.6f
C483 CS a_3430_64204# 0.0168f
C484 a_6504_51889# DVSS 0.616f
C485 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_1842_42732# 0.505f
C486 PAD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.102f
C487 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A VDD 0.607f
C488 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN PDRV1 5.15e-19
C489 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z VDD 0.181f
C490 a_3891_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB 0.0223f
C491 a_5575_63014# a_5463_64256# 0.00384f
C492 DVSS a_2591_61071# 0.074f
C493 CS PDRV0 0.0377f
C494 a_6824_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.0223f
C495 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A DVSS 1.66f
C496 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.329f
C497 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.00122f
C498 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB a_3430_64204# 5.12e-19
C499 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.0482f
C500 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB 0.342f
C501 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 5.45f
C502 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.329f
C503 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.658f
C504 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_3891_66144# 0.937f
C505 OE a_7790_42688# 0.00103f
C506 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_3430_64204# 0.317f
C507 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB 0.00382f
C508 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.125f
C509 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB a_12354_42732# 0.0142f
C510 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 2.99f
C511 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_11617_50285# 0.763f
C512 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.545f
C513 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.0692f
C514 PAD GF_NI_BI_T_BASE_0.ndrive_x_<2> 7.42f
C515 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_y_<0> 10.4f
C516 DVDD IE 1.18f
C517 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.0916f
C518 a_11294_42688# GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.00245f
C519 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.00197f
C520 a_1260_51889# PDRV1 6.18e-19
C521 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z a_9536_64061# 0.0604f
C522 a_9536_64061# a_2947_62989# 7.55e-19
C523 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.0482f
C524 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A PD 0.0556f
C525 OE a_8953_50157# 2.94e-19
C526 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.835f
C527 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_1260_51889# 5.93e-20
C528 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PD 2.63f
C529 a_1260_50201# PDRV0 0.0647f
C530 a_12527_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 9.9e-19
C531 GF_NI_BI_T_BASE_0.pdrive_y_<1> PAD 10.2f
C532 DVDD a_4286_42688# 3.94f
C533 A a_8953_50157# 0.0015f
C534 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_11294_42688# 2.42f
C535 PAD GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.341f
C536 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_5463_64256# 0.894f
C537 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_5463_64256# 0.0506f
C538 GF_NI_BI_T_BASE_0.ndrive_x_<3> a_11294_42688# 0.04f
C539 a_782_42688# DVSS 2.85f
C540 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y 2.42f
C541 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB DVSS 4.89f
C542 GF_NI_BI_T_BASE_0.ndrive_y_<0> a_1842_42732# 1.29f
C543 a_7790_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.00353f
C544 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z PD 0.00118f
C545 a_5502_50201# PDRV1 0.0647f
C546 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN a_11294_42688# 2.22f
C547 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.pdrive_x_<1> 2.29f
C548 DVSS a_11617_50285# 1.54f
C549 PAD GF_NI_BI_T_BASE_0.pdrive_y_<3> 10.2f
C550 a_5502_50201# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 1.66e-19
C551 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.545f
C552 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.00714f
C553 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.372f
C554 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 5.21e-19
C555 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_12966_56686# 0.169f
C556 a_7790_42688# GF_NI_BI_T_BASE_0.ndrive_x_<2> 1.78f
C557 DVDD a_4235_64204# 6.16e-19
C558 a_4157_63027# a_2947_62989# 1.01f
C559 CS a_2947_62989# 9.64e-20
C560 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.613f
C561 GF_NI_BI_T_BASE_0.pdrive_y_<3> a_12354_42732# 0.0205f
C562 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.524f
C563 a_782_42688# PDRV0 0.0011f
C564 a_12527_59749# VDD 0.512f
C565 a_2031_61071# PDRV1 0.0032f
C566 GF_NI_BI_T_BASE_0.pdrive_y_<0> PAD 10.2f
C567 a_5346_42732# VDD 0.00255f
C568 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z IE 1.4e-19
C569 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A DVSS 2.41f
C570 a_9197_50157# VDD 1.3f
C571 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB SL 1.29e-19
C572 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 14.8f
C573 VDD Y 1.79f
C574 OE a_1842_42732# 9.09e-19
C575 a_5575_63014# a_4235_64204# 0.00124f
C576 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVDD 7f
C577 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN DVDD 2.36f
C578 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0> 4.33e-19
C579 CS PDRV1 0.0399f
C580 VDD PD 4.66f
C581 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB 1.35f
C582 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_2947_62989# 0.665f
C583 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN SL 9.91e-20
C584 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.0715f
C585 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 0.0408f
C586 a_1191_61071# a_9536_64061# 0.017f
C587 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 0.206f
C588 a_6504_50201# VDD 0.0767f
C589 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z VDD 1.49f
C590 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.0744f
C591 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 0.0247f
C592 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z 1.6f
C593 a_12527_59749# PD 0.823f
C594 OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 0.0238f
C595 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 6.85e-19
C596 a_6504_51889# PDRV1 0.0023f
C597 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z 0.633f
C598 a_1842_42732# GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.718f
C599 A GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 1.54e-19
C600 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.0715f
C601 PAD GF_NI_BI_T_BASE_0.pdrive_x_<1> 20.9f
C602 DVSS a_1471_61071# 0.0534f
C603 Y PD 1.13e-19
C604 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.pdrive_x_<3> 6.39e-19
C605 a_2591_61071# PDRV1 9.81e-19
C606 a_12527_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 0.24f
C607 a_6504_51889# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 5.93e-20
C608 OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 0.0321f
C609 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.pdrive_x_<3> 7.34e-19
C610 OE a_1260_51889# 0.769f
C611 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_4235_64204# 0.00726f
C612 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB a_1842_42732# 0.0245f
C613 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN GF_NI_BI_T_BASE_0.pdrive_x_<0> 9.2e-19
C614 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.pdrive_x_<0> 6.39e-19
C615 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_4235_64204# 0.0794f
C616 DVSS DVDD 0.361p
C617 A GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 1.16e-19
C618 a_2031_61071# a_1191_61071# 4.22e-19
C619 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z Y 7.07e-20
C620 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.pdrive_x_<3> 9.56e-19
C621 VDD IE 1.31f
C622 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 4.24e-20
C623 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z PD 0.381f
C624 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 5.97e-20
C625 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB DVDD 0.606f
C626 a_4157_63027# a_1191_61071# 0.00154f
C627 a_10720_50201# VDD 0.012f
C628 a_3891_66144# DVDD 1.29f
C629 a_6824_66100# a_4157_63027# 2.86e-20
C630 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.0127f
C631 DVDD a_3430_64204# 0.0953f
C632 OE a_5502_50201# 0.0328f
C633 a_5575_63014# DVSS 0.282f
C634 a_9135_66144# CS 0.00184f
C635 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.212f
C636 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.ndrive_y_<2> 14.7f
C637 a_1471_61071# PDRV0 0.0175f
C638 a_6824_66100# CS 0.424f
C639 PAD a_7790_42688# 0.29f
C640 a_2871_53829# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 2.39e-19
C641 a_2871_53829# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 1.01e-19
C642 DVDD PDRV0 3.3f
C643 PAD GF_NI_BI_T_BASE_0.pdrive_x_<2> 20.9f
C644 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.0313f
C645 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.0396f
C646 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_1191_61071# 0.00239f
C647 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB PDRV1 4.26e-19
C648 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.ndrive_x_<2> 3.42e-19
C649 a_10720_50201# a_9197_50157# 0.152f
C650 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.00321f
C651 IE PD 0.815f
C652 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z a_6824_66100# 3.3e-21
C653 PU a_9536_64061# 0.0212f
C654 a_782_42688# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 1.68f
C655 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 4.44f
C656 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_1191_61071# 3.14e-19
C657 PAD a_8953_50157# 0.00582f
C658 a_2591_61071# a_1191_61071# 4.05e-19
C659 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_x_<0> 1.64e-19
C660 a_2871_53829# a_1260_51889# 2.93e-19
C661 a_5346_42732# a_4286_42688# 1.9f
C662 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.926f
C663 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.ndrive_x_<2> 3.42e-19
C664 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 0.101f
C665 a_1751_53829# a_2311_53829# 0.0346f
C666 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS 1.44f
C667 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS 4.88f
C668 a_12966_56686# DVDD 0.0274f
C669 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A SL 0.704f
C670 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.07f
C671 GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVDD 12.4f
C672 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB 9.98e-19
C673 GF_NI_BI_T_BASE_0.ndrive_x_<0> PAD 5.05f
C674 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL VDD 0.671f
C675 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.0133f
C676 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN VDD 0.366f
C677 a_2311_53829# PDRV1 0.00198f
C678 GF_NI_BI_T_BASE_0.pdrive_y_<0> a_1842_42732# 2.92f
C679 DVDD a_1191_53829# 0.427f
C680 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 0.0296f
C681 a_3891_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 5.09e-19
C682 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_3430_64204# 0.505f
C683 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_3430_64204# 0.303f
C684 OE a_6504_51889# 0.732f
C685 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3> 3.33e-19
C686 a_7790_42688# GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.184f
C687 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_12715_59749# 0.0928f
C688 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 8.1e-20
C689 PU CS 0.371f
C690 OE GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A 0.00464f
C691 OE a_1260_50201# 0.0328f
C692 a_782_42688# GF_NI_BI_T_BASE_0.ndrive_y_<0> 1.89f
C693 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PDRV0 1.79e-19
C694 a_5463_64256# a_4235_64204# 1.04f
C695 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A A 0.00702f
C696 GF_NI_BI_T_BASE_0.ndrive_x_<1> DVDD 9.37f
C697 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z DVDD 2.29f
C698 a_5346_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.33f
C699 a_1751_53829# DVDD 0.433f
C700 a_5346_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 2.31f
C701 DVDD a_2947_62989# 1.95f
C702 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.981f
C703 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_9197_50157# 4.94e-20
C704 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z PU 0.0534f
C705 PAD GF_NI_BI_T_BASE_0.ndrive_y_<2> 6.37f
C706 a_1471_61071# PDRV1 0.0479f
C707 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_8850_42732# 0.012f
C708 a_8850_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 2.22f
C709 a_11617_50285# SL 0.4f
C710 DVSS VDD 31.8f
C711 DVDD PDRV1 4.98f
C712 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A PU 1.15f
C713 a_1842_42732# GF_NI_BI_T_BASE_0.pdrive_x_<1> 5.58e-20
C714 a_5575_63014# a_2947_62989# 0.063f
C715 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_6504_50201# 6.69e-20
C716 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A a_1191_61071# 0.0635f
C717 PAD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB 0.00592f
C718 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB VDD 0.6f
C719 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD 3.81f
C720 PAD GF_NI_BI_T_BASE_0.ndrive_x_<3> 6.1f
C721 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.136f
C722 a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A 0.373f
C723 a_6824_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A 0.00184f
C724 a_3891_66144# VDD 0.575f
C725 OE GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB 0.0374f
C726 VDD a_3430_64204# 0.0742f
C727 a_4157_63027# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.311f
C728 PAD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 0.228f
C729 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<2> 16.8f
C730 a_12527_59749# DVSS 0.242f
C731 a_5346_42732# DVSS 2.76f
C732 CS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.0014f
C733 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_12354_42732# 0.561f
C734 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A a_12000_56686# 0.178f
C735 OE a_11617_50285# 0.00143f
C736 GF_NI_BI_T_BASE_0.ndrive_x_<3> a_12354_42732# 1.77f
C737 DVSS a_9197_50157# 0.628f
C738 DVDD a_11294_42688# 4f
C739 a_5502_50201# a_3961_50157# 0.152f
C740 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB a_12527_59749# 2.7e-20
C741 DVSS Y 0.979f
C742 VDD PDRV0 2.4f
C743 a_8850_42732# DVSS 4.61f
C744 A a_11617_50285# 9.54e-19
C745 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.464f
C746 DVSS PD 6.47f
C747 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 7.86e-20
C748 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN a_12354_42732# 2.3f
C749 a_9135_66144# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z 0.751f
C750 a_7790_42688# GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.88f
C751 DVSS a_5463_64256# 0.759f
C752 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB PD 0.0137f
C753 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.0477f
C754 a_782_42688# GF_NI_BI_T_BASE_0.pdrive_x_<0> 8.77e-19
C755 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 0.00182f
C756 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_2947_62989# 1.98f
C757 a_1471_61071# a_1191_61071# 0.0352f
C758 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A a_12715_59749# 0.00487f
C759 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_2947_62989# 3.4f
C760 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z DVSS 1.63f
C761 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.00333f
C762 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.217f
C763 a_3891_66144# PD 7.47e-19
C764 DVDD a_1191_61071# 5.17f
C765 a_3430_64204# PD 0.0113f
C766 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.0773f
C767 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_7790_42688# 1.28e-19
C768 OE a_2311_53829# 5.25e-19
C769 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL a_4286_42688# 0.012f
C770 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN a_4286_42688# 2.22f
C771 DVDD GF_NI_BI_T_BASE_0.ndrive_y_<0> 8.54f
C772 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 4.33e-19
C773 a_12966_56686# VDD 1.11e-20
C774 a_6824_66100# DVDD 1.28f
C775 a_5463_64256# a_3430_64204# 0.396f
C776 a_9135_66144# DVDD 1.29f
C777 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PDRV1 0.0478f
C778 PD PDRV0 7.52e-20
C779 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB a_11617_50285# 0.0306f
C780 DVDD SL 3.76f
C781 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN a_7790_42688# 6.5e-19
C782 a_12000_56686# DVDD 0.0273f
C783 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.158f
C784 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.00753f
C785 a_5575_63014# a_1191_61071# 0.00522f
C786 VDD a_1191_53829# 0.00259f
C787 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A PU 1.72f
C788 DVSS IE 1.19f
C789 a_12068_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB 0.0223f
C790 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB a_8953_50157# 0.00164f
C791 DVSS a_10720_50201# 0.00289f
C792 GF_NI_BI_T_BASE_0.ndrive_x_<0> a_1842_42732# 0.0338f
C793 a_12715_59749# DVDD 0.163f
C794 a_6504_51889# a_3961_50157# 0.00675f
C795 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 0.00298f
C796 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB 0.00719f
C797 a_8953_50157# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 0.015f
C798 PAD GF_NI_BI_T_BASE_0.ndrive_Y_<1> 8f
C799 a_3891_66144# IE 0.348f
C800 a_1751_53829# VDD 0.00106f
C801 OE DVDD 7.85f
C802 DVSS a_4286_42688# 4.61f
C803 VDD a_2947_62989# 0.179f
C804 IE a_3430_64204# 5.96e-20
C805 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z VDD 0.53f
C806 PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z 3.68e-19
C807 A DVDD 4.11f
C808 a_12966_56686# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 0.0414f
C809 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 0.0866f
C810 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<3> 29.8f
C811 a_6504_51889# PAD 0.302f
C812 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A a_12068_66100# 0.441f
C813 a_2871_53829# a_2311_53829# 0.0346f
C814 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A a_1191_61071# 0.00103f
C815 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.669f
C816 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_1191_61071# 0.0024f
C817 VDD PDRV1 3.12f
C818 a_12527_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z 2e-20
C819 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB a_1842_42732# 2.43f
C820 a_6824_66100# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 8.96e-20
C821 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z a_6824_66100# 0.769f
C822 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN a_1842_42732# 2.22f
C823 a_5346_42732# GF_NI_BI_T_BASE_0.ndrive_x_<1> 1.77f
C824 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A VDD 0.157f
C825 DVSS a_4235_64204# 1.72f
C826 PU DVDD 3.58f
C827 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<0> 29.7f
C828 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN 1.47f
C829 a_782_42688# GF_NI_BI_T_BASE_0.pdrive_y_<0> 0.0205f
C830 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z PD 1.54f
C831 a_2947_62989# PD 1.33e-19
C832 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVDD 0.478f
C833 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.ndrive_y_<2> 7.22e-19
C834 a_3891_66144# a_4235_64204# 2.37e-19
C835 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_y_<2> 9.96f
C836 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB a_3961_50157# 0.0139f
C837 a_3430_64204# a_4235_64204# 0.179f
C838 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z SL 0.00491f
C839 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN 3.77f
C840 GF_NI_BI_T_BASE_0.ndrive_Y_<1> a_7790_42688# 3.7e-19
C841 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS 9.65f
C842 a_5346_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 1.68f
C843 PD PDRV1 0.032f
C844 a_2871_53829# DVDD 0.462f
C845 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A a_9197_50157# 0.0458f
C846 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.ndrive_y_<2> 6.12e-19
C847 DVDD GF_NI_BI_T_BASE_0.ndrive_x_<2> 15.3f
C848 a_8850_42732# GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.505f
C849 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN a_1260_51889# 0.594f
C850 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB a_1260_51889# 0.0139f
C851 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB PAD 0.116f
C852 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.0143f
C853 a_12715_59749# GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 4.85e-19
C854 a_8850_42732# GF_NI_BI_T_BASE_0.pdrive_y_<2> 2.81f
C855 a_1191_61071# VDD 1.57f
C856 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN 5.39f
C857 OE GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.00202f
C858 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.00748f
C859 GF_NI_BI_T_BASE_0.pdrive_y_<1> DVDD 16.8f
C860 a_9135_66144# VDD 0.565f
C861 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.0352f
C862 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.024f
C863 a_6824_66100# VDD 0.565f
C864 a_8850_42732# a_11294_42688# 0.00366f
C865 DVDD GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 50.7f
C866 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL PDRV0 0.0251f
C867 A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.00283f
C868 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB 0.00379f
C869 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A PU 0.00136f
C870 VDD SL 3.37f
C871 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PU 2.63f
C872 a_12000_56686# VDD 1.11e-20
C873 a_12527_59749# a_1191_61071# 0.00326f
C874 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB DVSS 2f
C875 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.00221f
C876 GF_NI_BI_T_BASE_0.pdrive_y_<3> DVDD 17.9f
C877 GF_NI_BI_T_BASE_0.ndrive_x_<1> a_4286_42688# 0.0416f
C878 a_5575_63014# GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN 0.719f
C879 PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z 0.203f
C880 A VSS 2.59f
C881 SL VSS 2.93f
C882 Y VSS 2.9f
C883 PD VSS 6.58f
C884 PU VSS 9.77f
C885 CS VSS 4.51f
C886 IE VSS 1.56f
C887 PDRV1 VSS 6.06f
C888 OE VSS 14.9f
C889 PDRV0 VSS 6.94f
C890 VDD VSS 0.149p
C891 DVSS VSS 0.199p
C892 PAD VSS 92.7f
C893 DVDD VSS 1.08p
C894 GF_NI_BI_T_BASE_0.ndrive_x_<3> VSS 1.04f $ **FLOATING
C895 GF_NI_BI_T_BASE_0.ndrive_Y_<3> VSS 0.773f $ **FLOATING
C896 GF_NI_BI_T_BASE_0.pdrive_y_<3> VSS 1.1f $ **FLOATING
C897 GF_NI_BI_T_BASE_0.pdrive_x_<3> VSS 1.74f $ **FLOATING
C898 a_12354_42732# VSS 1.07f $ **FLOATING
C899 a_11294_42688# VSS 1.04f $ **FLOATING
C900 GF_NI_BI_T_BASE_0.pdrive_x_<2> VSS 1.82f $ **FLOATING
C901 GF_NI_BI_T_BASE_0.pdrive_y_<2> VSS 1.15f $ **FLOATING
C902 GF_NI_BI_T_BASE_0.ndrive_y_<2> VSS 1.83f $ **FLOATING
C903 GF_NI_BI_T_BASE_0.ndrive_x_<2> VSS 2.19f $ **FLOATING
C904 a_8850_42732# VSS 1.04f $ **FLOATING
C905 a_7790_42688# VSS 1.03f $ **FLOATING
C906 GF_NI_BI_T_BASE_0.ndrive_x_<1> VSS 1.77f $ **FLOATING
C907 GF_NI_BI_T_BASE_0.ndrive_Y_<1> VSS 2.29f $ **FLOATING
C908 GF_NI_BI_T_BASE_0.pdrive_y_<1> VSS 1.15f $ **FLOATING
C909 GF_NI_BI_T_BASE_0.pdrive_x_<1> VSS 1.8f $ **FLOATING
C910 a_5346_42732# VSS 1.04f $ **FLOATING
C911 a_4286_42688# VSS 1.04f $ **FLOATING
C912 GF_NI_BI_T_BASE_0.pdrive_x_<0> VSS 1.74f $ **FLOATING
C913 GF_NI_BI_T_BASE_0.pdrive_y_<0> VSS 1.09f $ **FLOATING
C914 GF_NI_BI_T_BASE_0.ndrive_y_<0> VSS 1.15f $ **FLOATING
C915 GF_NI_BI_T_BASE_0.ndrive_x_<0> VSS 0.908f $ **FLOATING
C916 a_1842_42732# VSS 1.04f $ **FLOATING
C917 a_782_42688# VSS 1.08f $ **FLOATING
C918 a_10720_50201# VSS 0.245f $ **FLOATING
C919 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB VSS 2.91f $ **FLOATING
C920 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL VSS 4.39f $ **FLOATING
C921 a_11617_50285# VSS 1.49f $ **FLOATING
C922 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A VSS 4.9f $ **FLOATING
C923 a_9197_50157# VSS 1.03f $ **FLOATING
C924 a_8953_50157# VSS 0.327f $ **FLOATING
C925 a_6504_50201# VSS 0.236f $ **FLOATING
C926 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.ENB VSS 2.82f $ **FLOATING
C927 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.EN VSS 2.53f $ **FLOATING
C928 a_5502_50201# VSS 0.236f $ **FLOATING
C929 a_6504_51889# VSS 0.967f $ **FLOATING
C930 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.ENB VSS 2.39f $ **FLOATING
C931 a_3961_50157# VSS 0.977f $ **FLOATING
C932 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.EN VSS 4.74f $ **FLOATING
C933 a_1260_50201# VSS 0.236f $ **FLOATING
C934 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.ENB VSS 1.66f $ **FLOATING
C935 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.EN VSS 2.36f $ **FLOATING
C936 a_1260_51889# VSS 1.01f $ **FLOATING
C937 a_12966_56686# VSS 0.203f $ **FLOATING
C938 a_12000_56686# VSS 0.203f $ **FLOATING
C939 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z VSS 1.71f $ **FLOATING
C940 a_12715_59749# VSS 0.81f $ **FLOATING
C941 a_12527_59749# VSS 1.06f $ **FLOATING
C942 a_2871_53829# VSS 0.153f $ **FLOATING
C943 a_2591_61071# VSS 0.151f $ **FLOATING
C944 a_2311_53829# VSS 0.151f $ **FLOATING
C945 a_2031_61071# VSS 0.149f $ **FLOATING
C946 a_1751_53829# VSS 0.152f $ **FLOATING
C947 a_1471_61071# VSS 0.149f $ **FLOATING
C948 a_1191_53829# VSS 0.163f $ **FLOATING
C949 a_1191_61071# VSS 3.42f $ **FLOATING
C950 a_5575_63014# VSS 0.132f $ **FLOATING
C951 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS 6.37f $ **FLOATING
C952 a_9536_64061# VSS 4.02f $ **FLOATING
C953 a_4157_63027# VSS 2.67f $ **FLOATING
C954 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A VSS 2.53f $ **FLOATING
C955 a_5463_64256# VSS 0.962f $ **FLOATING
C956 a_4235_64204# VSS 0.629f $ **FLOATING
C957 a_3430_64204# VSS 2.94f $ **FLOATING
C958 a_2947_62989# VSS 1.1f $ **FLOATING
C959 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN VSS 6.08f $ **FLOATING
C960 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A VSS 3.54f $ **FLOATING
C961 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB VSS 0.148f $ **FLOATING
C962 a_12068_66100# VSS 1.49f $ **FLOATING
C963 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.Z VSS 1.91f $ **FLOATING
C964 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.ZB VSS 1.17f $ **FLOATING
C965 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z VSS 0.601f $ **FLOATING
C966 a_9135_66144# VSS 1.42f $ **FLOATING
C967 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VSS 3.51f $ **FLOATING
C968 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB VSS 0.148f $ **FLOATING
C969 a_6824_66100# VSS 1.54f $ **FLOATING
C970 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z VSS 4.07f $ **FLOATING
C971 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB VSS 0.148f $ **FLOATING
C972 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z VSS 2.94f $ **FLOATING
C973 a_3891_66144# VSS 1.47f $ **FLOATING
.ends
