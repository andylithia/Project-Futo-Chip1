magic
tech gf180mcuC
magscale 1 10
timestamp 1669692783
<< metal1 >>
rect 1344 36874 38640 36908
rect 1344 36822 5876 36874
rect 5928 36822 5980 36874
rect 6032 36822 6084 36874
rect 6136 36822 15200 36874
rect 15252 36822 15304 36874
rect 15356 36822 15408 36874
rect 15460 36822 24524 36874
rect 24576 36822 24628 36874
rect 24680 36822 24732 36874
rect 24784 36822 33848 36874
rect 33900 36822 33952 36874
rect 34004 36822 34056 36874
rect 34108 36822 38640 36874
rect 1344 36788 38640 36822
rect 1344 36090 38800 36124
rect 1344 36038 10538 36090
rect 10590 36038 10642 36090
rect 10694 36038 10746 36090
rect 10798 36038 19862 36090
rect 19914 36038 19966 36090
rect 20018 36038 20070 36090
rect 20122 36038 29186 36090
rect 29238 36038 29290 36090
rect 29342 36038 29394 36090
rect 29446 36038 38510 36090
rect 38562 36038 38614 36090
rect 38666 36038 38718 36090
rect 38770 36038 38800 36090
rect 1344 36004 38800 36038
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 1344 34522 38800 34556
rect 1344 34470 10538 34522
rect 10590 34470 10642 34522
rect 10694 34470 10746 34522
rect 10798 34470 19862 34522
rect 19914 34470 19966 34522
rect 20018 34470 20070 34522
rect 20122 34470 29186 34522
rect 29238 34470 29290 34522
rect 29342 34470 29394 34522
rect 29446 34470 38510 34522
rect 38562 34470 38614 34522
rect 38666 34470 38718 34522
rect 38770 34470 38800 34522
rect 1344 34436 38800 34470
rect 1344 33738 38640 33772
rect 1344 33686 5876 33738
rect 5928 33686 5980 33738
rect 6032 33686 6084 33738
rect 6136 33686 15200 33738
rect 15252 33686 15304 33738
rect 15356 33686 15408 33738
rect 15460 33686 24524 33738
rect 24576 33686 24628 33738
rect 24680 33686 24732 33738
rect 24784 33686 33848 33738
rect 33900 33686 33952 33738
rect 34004 33686 34056 33738
rect 34108 33686 38640 33738
rect 1344 33652 38640 33686
rect 1344 32954 38800 32988
rect 1344 32902 10538 32954
rect 10590 32902 10642 32954
rect 10694 32902 10746 32954
rect 10798 32902 19862 32954
rect 19914 32902 19966 32954
rect 20018 32902 20070 32954
rect 20122 32902 29186 32954
rect 29238 32902 29290 32954
rect 29342 32902 29394 32954
rect 29446 32902 38510 32954
rect 38562 32902 38614 32954
rect 38666 32902 38718 32954
rect 38770 32902 38800 32954
rect 1344 32868 38800 32902
rect 1344 32170 38640 32204
rect 1344 32118 5876 32170
rect 5928 32118 5980 32170
rect 6032 32118 6084 32170
rect 6136 32118 15200 32170
rect 15252 32118 15304 32170
rect 15356 32118 15408 32170
rect 15460 32118 24524 32170
rect 24576 32118 24628 32170
rect 24680 32118 24732 32170
rect 24784 32118 33848 32170
rect 33900 32118 33952 32170
rect 34004 32118 34056 32170
rect 34108 32118 38640 32170
rect 1344 32084 38640 32118
rect 1344 31386 38800 31420
rect 1344 31334 10538 31386
rect 10590 31334 10642 31386
rect 10694 31334 10746 31386
rect 10798 31334 19862 31386
rect 19914 31334 19966 31386
rect 20018 31334 20070 31386
rect 20122 31334 29186 31386
rect 29238 31334 29290 31386
rect 29342 31334 29394 31386
rect 29446 31334 38510 31386
rect 38562 31334 38614 31386
rect 38666 31334 38718 31386
rect 38770 31334 38800 31386
rect 1344 31300 38800 31334
rect 1344 30602 38640 30636
rect 1344 30550 5876 30602
rect 5928 30550 5980 30602
rect 6032 30550 6084 30602
rect 6136 30550 15200 30602
rect 15252 30550 15304 30602
rect 15356 30550 15408 30602
rect 15460 30550 24524 30602
rect 24576 30550 24628 30602
rect 24680 30550 24732 30602
rect 24784 30550 33848 30602
rect 33900 30550 33952 30602
rect 34004 30550 34056 30602
rect 34108 30550 38640 30602
rect 1344 30516 38640 30550
rect 1344 29818 38800 29852
rect 1344 29766 10538 29818
rect 10590 29766 10642 29818
rect 10694 29766 10746 29818
rect 10798 29766 19862 29818
rect 19914 29766 19966 29818
rect 20018 29766 20070 29818
rect 20122 29766 29186 29818
rect 29238 29766 29290 29818
rect 29342 29766 29394 29818
rect 29446 29766 38510 29818
rect 38562 29766 38614 29818
rect 38666 29766 38718 29818
rect 38770 29766 38800 29818
rect 1344 29732 38800 29766
rect 1344 29034 38640 29068
rect 1344 28982 5876 29034
rect 5928 28982 5980 29034
rect 6032 28982 6084 29034
rect 6136 28982 15200 29034
rect 15252 28982 15304 29034
rect 15356 28982 15408 29034
rect 15460 28982 24524 29034
rect 24576 28982 24628 29034
rect 24680 28982 24732 29034
rect 24784 28982 33848 29034
rect 33900 28982 33952 29034
rect 34004 28982 34056 29034
rect 34108 28982 38640 29034
rect 1344 28948 38640 28982
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 1344 27466 38640 27500
rect 1344 27414 5876 27466
rect 5928 27414 5980 27466
rect 6032 27414 6084 27466
rect 6136 27414 15200 27466
rect 15252 27414 15304 27466
rect 15356 27414 15408 27466
rect 15460 27414 24524 27466
rect 24576 27414 24628 27466
rect 24680 27414 24732 27466
rect 24784 27414 33848 27466
rect 33900 27414 33952 27466
rect 34004 27414 34056 27466
rect 34108 27414 38640 27466
rect 1344 27380 38640 27414
rect 1344 26682 38800 26716
rect 1344 26630 10538 26682
rect 10590 26630 10642 26682
rect 10694 26630 10746 26682
rect 10798 26630 19862 26682
rect 19914 26630 19966 26682
rect 20018 26630 20070 26682
rect 20122 26630 29186 26682
rect 29238 26630 29290 26682
rect 29342 26630 29394 26682
rect 29446 26630 38510 26682
rect 38562 26630 38614 26682
rect 38666 26630 38718 26682
rect 38770 26630 38800 26682
rect 1344 26596 38800 26630
rect 1344 25898 38640 25932
rect 1344 25846 5876 25898
rect 5928 25846 5980 25898
rect 6032 25846 6084 25898
rect 6136 25846 15200 25898
rect 15252 25846 15304 25898
rect 15356 25846 15408 25898
rect 15460 25846 24524 25898
rect 24576 25846 24628 25898
rect 24680 25846 24732 25898
rect 24784 25846 33848 25898
rect 33900 25846 33952 25898
rect 34004 25846 34056 25898
rect 34108 25846 38640 25898
rect 1344 25812 38640 25846
rect 1344 25114 38800 25148
rect 1344 25062 10538 25114
rect 10590 25062 10642 25114
rect 10694 25062 10746 25114
rect 10798 25062 19862 25114
rect 19914 25062 19966 25114
rect 20018 25062 20070 25114
rect 20122 25062 29186 25114
rect 29238 25062 29290 25114
rect 29342 25062 29394 25114
rect 29446 25062 38510 25114
rect 38562 25062 38614 25114
rect 38666 25062 38718 25114
rect 38770 25062 38800 25114
rect 1344 25028 38800 25062
rect 1344 24330 38640 24364
rect 1344 24278 5876 24330
rect 5928 24278 5980 24330
rect 6032 24278 6084 24330
rect 6136 24278 15200 24330
rect 15252 24278 15304 24330
rect 15356 24278 15408 24330
rect 15460 24278 24524 24330
rect 24576 24278 24628 24330
rect 24680 24278 24732 24330
rect 24784 24278 33848 24330
rect 33900 24278 33952 24330
rect 34004 24278 34056 24330
rect 34108 24278 38640 24330
rect 1344 24244 38640 24278
rect 1344 23546 38800 23580
rect 1344 23494 10538 23546
rect 10590 23494 10642 23546
rect 10694 23494 10746 23546
rect 10798 23494 19862 23546
rect 19914 23494 19966 23546
rect 20018 23494 20070 23546
rect 20122 23494 29186 23546
rect 29238 23494 29290 23546
rect 29342 23494 29394 23546
rect 29446 23494 38510 23546
rect 38562 23494 38614 23546
rect 38666 23494 38718 23546
rect 38770 23494 38800 23546
rect 1344 23460 38800 23494
rect 1344 22762 38640 22796
rect 1344 22710 5876 22762
rect 5928 22710 5980 22762
rect 6032 22710 6084 22762
rect 6136 22710 15200 22762
rect 15252 22710 15304 22762
rect 15356 22710 15408 22762
rect 15460 22710 24524 22762
rect 24576 22710 24628 22762
rect 24680 22710 24732 22762
rect 24784 22710 33848 22762
rect 33900 22710 33952 22762
rect 34004 22710 34056 22762
rect 34108 22710 38640 22762
rect 1344 22676 38640 22710
rect 1344 21978 38800 22012
rect 1344 21926 10538 21978
rect 10590 21926 10642 21978
rect 10694 21926 10746 21978
rect 10798 21926 19862 21978
rect 19914 21926 19966 21978
rect 20018 21926 20070 21978
rect 20122 21926 29186 21978
rect 29238 21926 29290 21978
rect 29342 21926 29394 21978
rect 29446 21926 38510 21978
rect 38562 21926 38614 21978
rect 38666 21926 38718 21978
rect 38770 21926 38800 21978
rect 1344 21892 38800 21926
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 1344 20410 38800 20444
rect 1344 20358 10538 20410
rect 10590 20358 10642 20410
rect 10694 20358 10746 20410
rect 10798 20358 19862 20410
rect 19914 20358 19966 20410
rect 20018 20358 20070 20410
rect 20122 20358 29186 20410
rect 29238 20358 29290 20410
rect 29342 20358 29394 20410
rect 29446 20358 38510 20410
rect 38562 20358 38614 20410
rect 38666 20358 38718 20410
rect 38770 20358 38800 20410
rect 1344 20324 38800 20358
rect 1344 19626 38640 19660
rect 1344 19574 5876 19626
rect 5928 19574 5980 19626
rect 6032 19574 6084 19626
rect 6136 19574 15200 19626
rect 15252 19574 15304 19626
rect 15356 19574 15408 19626
rect 15460 19574 24524 19626
rect 24576 19574 24628 19626
rect 24680 19574 24732 19626
rect 24784 19574 33848 19626
rect 33900 19574 33952 19626
rect 34004 19574 34056 19626
rect 34108 19574 38640 19626
rect 1344 19540 38640 19574
rect 1344 18842 38800 18876
rect 1344 18790 10538 18842
rect 10590 18790 10642 18842
rect 10694 18790 10746 18842
rect 10798 18790 19862 18842
rect 19914 18790 19966 18842
rect 20018 18790 20070 18842
rect 20122 18790 29186 18842
rect 29238 18790 29290 18842
rect 29342 18790 29394 18842
rect 29446 18790 38510 18842
rect 38562 18790 38614 18842
rect 38666 18790 38718 18842
rect 38770 18790 38800 18842
rect 1344 18756 38800 18790
rect 1344 18058 38640 18092
rect 1344 18006 5876 18058
rect 5928 18006 5980 18058
rect 6032 18006 6084 18058
rect 6136 18006 15200 18058
rect 15252 18006 15304 18058
rect 15356 18006 15408 18058
rect 15460 18006 24524 18058
rect 24576 18006 24628 18058
rect 24680 18006 24732 18058
rect 24784 18006 33848 18058
rect 33900 18006 33952 18058
rect 34004 18006 34056 18058
rect 34108 18006 38640 18058
rect 1344 17972 38640 18006
rect 1344 17274 38800 17308
rect 1344 17222 10538 17274
rect 10590 17222 10642 17274
rect 10694 17222 10746 17274
rect 10798 17222 19862 17274
rect 19914 17222 19966 17274
rect 20018 17222 20070 17274
rect 20122 17222 29186 17274
rect 29238 17222 29290 17274
rect 29342 17222 29394 17274
rect 29446 17222 38510 17274
rect 38562 17222 38614 17274
rect 38666 17222 38718 17274
rect 38770 17222 38800 17274
rect 1344 17188 38800 17222
rect 1344 16490 38640 16524
rect 1344 16438 5876 16490
rect 5928 16438 5980 16490
rect 6032 16438 6084 16490
rect 6136 16438 15200 16490
rect 15252 16438 15304 16490
rect 15356 16438 15408 16490
rect 15460 16438 24524 16490
rect 24576 16438 24628 16490
rect 24680 16438 24732 16490
rect 24784 16438 33848 16490
rect 33900 16438 33952 16490
rect 34004 16438 34056 16490
rect 34108 16438 38640 16490
rect 1344 16404 38640 16438
rect 1344 15706 38800 15740
rect 1344 15654 10538 15706
rect 10590 15654 10642 15706
rect 10694 15654 10746 15706
rect 10798 15654 19862 15706
rect 19914 15654 19966 15706
rect 20018 15654 20070 15706
rect 20122 15654 29186 15706
rect 29238 15654 29290 15706
rect 29342 15654 29394 15706
rect 29446 15654 38510 15706
rect 38562 15654 38614 15706
rect 38666 15654 38718 15706
rect 38770 15654 38800 15706
rect 1344 15620 38800 15654
rect 1344 14922 38640 14956
rect 1344 14870 5876 14922
rect 5928 14870 5980 14922
rect 6032 14870 6084 14922
rect 6136 14870 15200 14922
rect 15252 14870 15304 14922
rect 15356 14870 15408 14922
rect 15460 14870 24524 14922
rect 24576 14870 24628 14922
rect 24680 14870 24732 14922
rect 24784 14870 33848 14922
rect 33900 14870 33952 14922
rect 34004 14870 34056 14922
rect 34108 14870 38640 14922
rect 1344 14836 38640 14870
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 1344 13354 38640 13388
rect 1344 13302 5876 13354
rect 5928 13302 5980 13354
rect 6032 13302 6084 13354
rect 6136 13302 15200 13354
rect 15252 13302 15304 13354
rect 15356 13302 15408 13354
rect 15460 13302 24524 13354
rect 24576 13302 24628 13354
rect 24680 13302 24732 13354
rect 24784 13302 33848 13354
rect 33900 13302 33952 13354
rect 34004 13302 34056 13354
rect 34108 13302 38640 13354
rect 1344 13268 38640 13302
rect 1344 12570 38800 12604
rect 1344 12518 10538 12570
rect 10590 12518 10642 12570
rect 10694 12518 10746 12570
rect 10798 12518 19862 12570
rect 19914 12518 19966 12570
rect 20018 12518 20070 12570
rect 20122 12518 29186 12570
rect 29238 12518 29290 12570
rect 29342 12518 29394 12570
rect 29446 12518 38510 12570
rect 38562 12518 38614 12570
rect 38666 12518 38718 12570
rect 38770 12518 38800 12570
rect 1344 12484 38800 12518
rect 1344 11786 38640 11820
rect 1344 11734 5876 11786
rect 5928 11734 5980 11786
rect 6032 11734 6084 11786
rect 6136 11734 15200 11786
rect 15252 11734 15304 11786
rect 15356 11734 15408 11786
rect 15460 11734 24524 11786
rect 24576 11734 24628 11786
rect 24680 11734 24732 11786
rect 24784 11734 33848 11786
rect 33900 11734 33952 11786
rect 34004 11734 34056 11786
rect 34108 11734 38640 11786
rect 1344 11700 38640 11734
rect 1344 11002 38800 11036
rect 1344 10950 10538 11002
rect 10590 10950 10642 11002
rect 10694 10950 10746 11002
rect 10798 10950 19862 11002
rect 19914 10950 19966 11002
rect 20018 10950 20070 11002
rect 20122 10950 29186 11002
rect 29238 10950 29290 11002
rect 29342 10950 29394 11002
rect 29446 10950 38510 11002
rect 38562 10950 38614 11002
rect 38666 10950 38718 11002
rect 38770 10950 38800 11002
rect 1344 10916 38800 10950
rect 1344 10218 38640 10252
rect 1344 10166 5876 10218
rect 5928 10166 5980 10218
rect 6032 10166 6084 10218
rect 6136 10166 15200 10218
rect 15252 10166 15304 10218
rect 15356 10166 15408 10218
rect 15460 10166 24524 10218
rect 24576 10166 24628 10218
rect 24680 10166 24732 10218
rect 24784 10166 33848 10218
rect 33900 10166 33952 10218
rect 34004 10166 34056 10218
rect 34108 10166 38640 10218
rect 1344 10132 38640 10166
rect 1344 9434 38800 9468
rect 1344 9382 10538 9434
rect 10590 9382 10642 9434
rect 10694 9382 10746 9434
rect 10798 9382 19862 9434
rect 19914 9382 19966 9434
rect 20018 9382 20070 9434
rect 20122 9382 29186 9434
rect 29238 9382 29290 9434
rect 29342 9382 29394 9434
rect 29446 9382 38510 9434
rect 38562 9382 38614 9434
rect 38666 9382 38718 9434
rect 38770 9382 38800 9434
rect 1344 9348 38800 9382
rect 24222 8930 24274 8942
rect 24222 8866 24274 8878
rect 24670 8930 24722 8942
rect 24670 8866 24722 8878
rect 25678 8930 25730 8942
rect 25678 8866 25730 8878
rect 26126 8930 26178 8942
rect 26126 8866 26178 8878
rect 26574 8930 26626 8942
rect 26574 8866 26626 8878
rect 26910 8930 26962 8942
rect 26910 8866 26962 8878
rect 1344 8650 38640 8684
rect 1344 8598 5876 8650
rect 5928 8598 5980 8650
rect 6032 8598 6084 8650
rect 6136 8598 15200 8650
rect 15252 8598 15304 8650
rect 15356 8598 15408 8650
rect 15460 8598 24524 8650
rect 24576 8598 24628 8650
rect 24680 8598 24732 8650
rect 24784 8598 33848 8650
rect 33900 8598 33952 8650
rect 34004 8598 34056 8650
rect 34108 8598 38640 8650
rect 1344 8564 38640 8598
rect 23214 8034 23266 8046
rect 23214 7970 23266 7982
rect 23886 8034 23938 8046
rect 23886 7970 23938 7982
rect 24446 8034 24498 8046
rect 24446 7970 24498 7982
rect 24782 8034 24834 8046
rect 24782 7970 24834 7982
rect 25342 8034 25394 8046
rect 25342 7970 25394 7982
rect 26014 8034 26066 8046
rect 26014 7970 26066 7982
rect 26574 8034 26626 8046
rect 26574 7970 26626 7982
rect 26910 8034 26962 8046
rect 26910 7970 26962 7982
rect 27358 8034 27410 8046
rect 27358 7970 27410 7982
rect 27918 8034 27970 8046
rect 27918 7970 27970 7982
rect 28254 8034 28306 8046
rect 28254 7970 28306 7982
rect 28702 8034 28754 8046
rect 28702 7970 28754 7982
rect 1344 7866 38800 7900
rect 1344 7814 10538 7866
rect 10590 7814 10642 7866
rect 10694 7814 10746 7866
rect 10798 7814 19862 7866
rect 19914 7814 19966 7866
rect 20018 7814 20070 7866
rect 20122 7814 29186 7866
rect 29238 7814 29290 7866
rect 29342 7814 29394 7866
rect 29446 7814 38510 7866
rect 38562 7814 38614 7866
rect 38666 7814 38718 7866
rect 38770 7814 38800 7866
rect 1344 7780 38800 7814
rect 28702 7474 28754 7486
rect 28702 7410 28754 7422
rect 29150 7474 29202 7486
rect 29150 7410 29202 7422
rect 22430 7362 22482 7374
rect 22430 7298 22482 7310
rect 22766 7362 22818 7374
rect 22766 7298 22818 7310
rect 23214 7362 23266 7374
rect 23214 7298 23266 7310
rect 23886 7362 23938 7374
rect 23886 7298 23938 7310
rect 24558 7362 24610 7374
rect 24558 7298 24610 7310
rect 25566 7362 25618 7374
rect 25566 7298 25618 7310
rect 26014 7362 26066 7374
rect 26014 7298 26066 7310
rect 26462 7362 26514 7374
rect 26462 7298 26514 7310
rect 26910 7362 26962 7374
rect 26910 7298 26962 7310
rect 27358 7362 27410 7374
rect 27358 7298 27410 7310
rect 27806 7362 27858 7374
rect 27806 7298 27858 7310
rect 29710 7362 29762 7374
rect 29710 7298 29762 7310
rect 30046 7362 30098 7374
rect 30046 7298 30098 7310
rect 28590 7250 28642 7262
rect 29026 7198 29038 7250
rect 29090 7247 29102 7250
rect 29698 7247 29710 7250
rect 29090 7201 29710 7247
rect 29090 7198 29102 7201
rect 29698 7198 29710 7201
rect 29762 7198 29774 7250
rect 28590 7186 28642 7198
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 21858 6862 21870 6914
rect 21922 6911 21934 6914
rect 22418 6911 22430 6914
rect 21922 6865 22430 6911
rect 21922 6862 21934 6865
rect 22418 6862 22430 6865
rect 22482 6862 22494 6914
rect 27470 6802 27522 6814
rect 27470 6738 27522 6750
rect 28814 6802 28866 6814
rect 28814 6738 28866 6750
rect 22878 6690 22930 6702
rect 22878 6626 22930 6638
rect 23550 6690 23602 6702
rect 23550 6626 23602 6638
rect 24894 6690 24946 6702
rect 24894 6626 24946 6638
rect 25566 6690 25618 6702
rect 25566 6626 25618 6638
rect 24222 6578 24274 6590
rect 24222 6514 24274 6526
rect 26238 6578 26290 6590
rect 26238 6514 26290 6526
rect 26910 6578 26962 6590
rect 26910 6514 26962 6526
rect 28254 6578 28306 6590
rect 28254 6514 28306 6526
rect 29598 6578 29650 6590
rect 29598 6514 29650 6526
rect 29710 6578 29762 6590
rect 29710 6514 29762 6526
rect 30158 6578 30210 6590
rect 30158 6514 30210 6526
rect 21870 6466 21922 6478
rect 21870 6402 21922 6414
rect 22318 6466 22370 6478
rect 22318 6402 22370 6414
rect 22990 6466 23042 6478
rect 22990 6402 23042 6414
rect 23662 6466 23714 6478
rect 23662 6402 23714 6414
rect 24334 6466 24386 6478
rect 24334 6402 24386 6414
rect 25006 6466 25058 6478
rect 25006 6402 25058 6414
rect 25678 6466 25730 6478
rect 25678 6402 25730 6414
rect 26350 6466 26402 6478
rect 26350 6402 26402 6414
rect 27022 6466 27074 6478
rect 27022 6402 27074 6414
rect 28366 6466 28418 6478
rect 28366 6402 28418 6414
rect 30606 6466 30658 6478
rect 30606 6402 30658 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 31502 6466 31554 6478
rect 31502 6402 31554 6414
rect 31950 6466 32002 6478
rect 31950 6402 32002 6414
rect 1344 6298 38800 6332
rect 1344 6246 10538 6298
rect 10590 6246 10642 6298
rect 10694 6246 10746 6298
rect 10798 6246 19862 6298
rect 19914 6246 19966 6298
rect 20018 6246 20070 6298
rect 20122 6246 29186 6298
rect 29238 6246 29290 6298
rect 29342 6246 29394 6298
rect 29446 6246 38510 6298
rect 38562 6246 38614 6298
rect 38666 6246 38718 6298
rect 38770 6246 38800 6298
rect 1344 6212 38800 6246
rect 25790 6130 25842 6142
rect 25790 6066 25842 6078
rect 26462 6130 26514 6142
rect 26462 6066 26514 6078
rect 27134 6130 27186 6142
rect 27134 6066 27186 6078
rect 27806 6130 27858 6142
rect 27806 6066 27858 6078
rect 28478 6130 28530 6142
rect 28478 6066 28530 6078
rect 29822 6130 29874 6142
rect 29822 6066 29874 6078
rect 30942 6130 30994 6142
rect 30942 6066 30994 6078
rect 31390 6130 31442 6142
rect 31390 6066 31442 6078
rect 31838 6130 31890 6142
rect 31838 6066 31890 6078
rect 27694 6018 27746 6030
rect 27694 5954 27746 5966
rect 29038 6018 29090 6030
rect 29038 5954 29090 5966
rect 29150 6018 29202 6030
rect 29150 5954 29202 5966
rect 30382 6018 30434 6030
rect 30382 5954 30434 5966
rect 21982 5906 22034 5918
rect 21982 5842 22034 5854
rect 22654 5906 22706 5918
rect 22654 5842 22706 5854
rect 23326 5906 23378 5918
rect 23326 5842 23378 5854
rect 23998 5906 24050 5918
rect 23998 5842 24050 5854
rect 24670 5906 24722 5918
rect 24670 5842 24722 5854
rect 25678 5906 25730 5918
rect 25678 5842 25730 5854
rect 26350 5906 26402 5918
rect 26350 5842 26402 5854
rect 27022 5906 27074 5918
rect 27022 5842 27074 5854
rect 28366 5906 28418 5918
rect 28366 5842 28418 5854
rect 29710 5906 29762 5918
rect 29710 5842 29762 5854
rect 20526 5794 20578 5806
rect 20526 5730 20578 5742
rect 20974 5794 21026 5806
rect 20974 5730 21026 5742
rect 21422 5794 21474 5806
rect 21422 5730 21474 5742
rect 32286 5794 32338 5806
rect 32286 5730 32338 5742
rect 32734 5794 32786 5806
rect 32734 5730 32786 5742
rect 33518 5794 33570 5806
rect 33518 5730 33570 5742
rect 22094 5682 22146 5694
rect 20962 5630 20974 5682
rect 21026 5679 21038 5682
rect 21746 5679 21758 5682
rect 21026 5633 21758 5679
rect 21026 5630 21038 5633
rect 21746 5630 21758 5633
rect 21810 5630 21822 5682
rect 22094 5618 22146 5630
rect 22766 5682 22818 5694
rect 22766 5618 22818 5630
rect 23438 5682 23490 5694
rect 23438 5618 23490 5630
rect 24110 5682 24162 5694
rect 24110 5618 24162 5630
rect 24782 5682 24834 5694
rect 24782 5618 24834 5630
rect 30494 5682 30546 5694
rect 30494 5618 30546 5630
rect 1344 5514 38640 5548
rect 1344 5462 5876 5514
rect 5928 5462 5980 5514
rect 6032 5462 6084 5514
rect 6136 5462 15200 5514
rect 15252 5462 15304 5514
rect 15356 5462 15408 5514
rect 15460 5462 24524 5514
rect 24576 5462 24628 5514
rect 24680 5462 24732 5514
rect 24784 5462 33848 5514
rect 33900 5462 33952 5514
rect 34004 5462 34056 5514
rect 34108 5462 38640 5514
rect 1344 5428 38640 5462
rect 21870 5346 21922 5358
rect 21870 5282 21922 5294
rect 23214 5346 23266 5358
rect 23214 5282 23266 5294
rect 23886 5346 23938 5358
rect 23886 5282 23938 5294
rect 24558 5346 24610 5358
rect 24558 5282 24610 5294
rect 25230 5346 25282 5358
rect 25230 5282 25282 5294
rect 26574 5346 26626 5358
rect 26574 5282 26626 5294
rect 27246 5346 27298 5358
rect 27246 5282 27298 5294
rect 27918 5346 27970 5358
rect 27918 5282 27970 5294
rect 28590 5346 28642 5358
rect 28590 5282 28642 5294
rect 29710 5346 29762 5358
rect 29710 5282 29762 5294
rect 30382 5346 30434 5358
rect 30382 5282 30434 5294
rect 19630 5234 19682 5246
rect 19630 5170 19682 5182
rect 20414 5234 20466 5246
rect 20414 5170 20466 5182
rect 20862 5234 20914 5246
rect 20862 5170 20914 5182
rect 21758 5122 21810 5134
rect 21758 5058 21810 5070
rect 23102 5122 23154 5134
rect 23102 5058 23154 5070
rect 23774 5122 23826 5134
rect 23774 5058 23826 5070
rect 25118 5122 25170 5134
rect 25118 5058 25170 5070
rect 25790 5122 25842 5134
rect 25790 5058 25842 5070
rect 25902 5122 25954 5134
rect 25902 5058 25954 5070
rect 26462 5122 26514 5134
rect 26462 5058 26514 5070
rect 27806 5122 27858 5134
rect 27806 5058 27858 5070
rect 28478 5122 28530 5134
rect 28478 5058 28530 5070
rect 29598 5122 29650 5134
rect 29598 5058 29650 5070
rect 30270 5122 30322 5134
rect 30270 5058 30322 5070
rect 30942 5122 30994 5134
rect 30942 5058 30994 5070
rect 22430 5010 22482 5022
rect 22430 4946 22482 4958
rect 24446 5010 24498 5022
rect 24446 4946 24498 4958
rect 27134 5010 27186 5022
rect 27134 4946 27186 4958
rect 31054 5010 31106 5022
rect 31054 4946 31106 4958
rect 31614 5010 31666 5022
rect 31614 4946 31666 4958
rect 31726 5010 31778 5022
rect 31726 4946 31778 4958
rect 33518 5010 33570 5022
rect 33518 4946 33570 4958
rect 19070 4898 19122 4910
rect 19070 4834 19122 4846
rect 19966 4898 20018 4910
rect 19966 4834 20018 4846
rect 22542 4898 22594 4910
rect 22542 4834 22594 4846
rect 32174 4898 32226 4910
rect 32174 4834 32226 4846
rect 32622 4898 32674 4910
rect 32622 4834 32674 4846
rect 33070 4898 33122 4910
rect 33070 4834 33122 4846
rect 33966 4898 34018 4910
rect 33966 4834 34018 4846
rect 34414 4898 34466 4910
rect 34414 4834 34466 4846
rect 1344 4730 38800 4764
rect 1344 4678 10538 4730
rect 10590 4678 10642 4730
rect 10694 4678 10746 4730
rect 10798 4678 19862 4730
rect 19914 4678 19966 4730
rect 20018 4678 20070 4730
rect 20122 4678 29186 4730
rect 29238 4678 29290 4730
rect 29342 4678 29394 4730
rect 29446 4678 38510 4730
rect 38562 4678 38614 4730
rect 38666 4678 38718 4730
rect 38770 4678 38800 4730
rect 1344 4644 38800 4678
rect 18846 4562 18898 4574
rect 18846 4498 18898 4510
rect 19182 4562 19234 4574
rect 19182 4498 19234 4510
rect 23662 4562 23714 4574
rect 23662 4498 23714 4510
rect 24334 4562 24386 4574
rect 24334 4498 24386 4510
rect 24782 4562 24834 4574
rect 24782 4498 24834 4510
rect 25790 4562 25842 4574
rect 25790 4498 25842 4510
rect 27806 4562 27858 4574
rect 27806 4498 27858 4510
rect 28478 4562 28530 4574
rect 28478 4498 28530 4510
rect 29150 4562 29202 4574
rect 29150 4498 29202 4510
rect 29822 4562 29874 4574
rect 29822 4498 29874 4510
rect 31166 4562 31218 4574
rect 31166 4498 31218 4510
rect 31838 4562 31890 4574
rect 31838 4498 31890 4510
rect 34862 4562 34914 4574
rect 34862 4498 34914 4510
rect 20862 4450 20914 4462
rect 20862 4386 20914 4398
rect 21534 4450 21586 4462
rect 21534 4386 21586 4398
rect 22206 4450 22258 4462
rect 22206 4386 22258 4398
rect 26350 4450 26402 4462
rect 26350 4386 26402 4398
rect 26462 4450 26514 4462
rect 26462 4386 26514 4398
rect 27022 4450 27074 4462
rect 27022 4386 27074 4398
rect 30382 4450 30434 4462
rect 30382 4386 30434 4398
rect 30494 4450 30546 4462
rect 30494 4386 30546 4398
rect 31054 4450 31106 4462
rect 31054 4386 31106 4398
rect 31726 4450 31778 4462
rect 31726 4386 31778 4398
rect 20190 4338 20242 4350
rect 20190 4274 20242 4286
rect 22878 4338 22930 4350
rect 22878 4274 22930 4286
rect 23550 4338 23602 4350
rect 23550 4274 23602 4286
rect 24222 4338 24274 4350
rect 24222 4274 24274 4286
rect 25678 4338 25730 4350
rect 25678 4274 25730 4286
rect 27694 4338 27746 4350
rect 27694 4274 27746 4286
rect 28366 4338 28418 4350
rect 28366 4274 28418 4286
rect 29038 4338 29090 4350
rect 29038 4274 29090 4286
rect 29710 4338 29762 4350
rect 29710 4274 29762 4286
rect 32398 4338 32450 4350
rect 32398 4274 32450 4286
rect 19630 4226 19682 4238
rect 19630 4162 19682 4174
rect 33518 4226 33570 4238
rect 33518 4162 33570 4174
rect 33966 4226 34018 4238
rect 33966 4162 34018 4174
rect 34414 4226 34466 4238
rect 34414 4162 34466 4174
rect 20302 4114 20354 4126
rect 20302 4050 20354 4062
rect 20974 4114 21026 4126
rect 20974 4050 21026 4062
rect 21646 4114 21698 4126
rect 21646 4050 21698 4062
rect 22318 4114 22370 4126
rect 22318 4050 22370 4062
rect 22990 4114 23042 4126
rect 22990 4050 23042 4062
rect 27134 4114 27186 4126
rect 27134 4050 27186 4062
rect 32510 4114 32562 4126
rect 32510 4050 32562 4062
rect 1344 3946 38640 3980
rect 1344 3894 5876 3946
rect 5928 3894 5980 3946
rect 6032 3894 6084 3946
rect 6136 3894 15200 3946
rect 15252 3894 15304 3946
rect 15356 3894 15408 3946
rect 15460 3894 24524 3946
rect 24576 3894 24628 3946
rect 24680 3894 24732 3946
rect 24784 3894 33848 3946
rect 33900 3894 33952 3946
rect 34004 3894 34056 3946
rect 34108 3894 38640 3946
rect 1344 3860 38640 3894
rect 16606 3778 16658 3790
rect 16606 3714 16658 3726
rect 19294 3778 19346 3790
rect 19294 3714 19346 3726
rect 19966 3778 20018 3790
rect 19966 3714 20018 3726
rect 24222 3778 24274 3790
rect 24222 3714 24274 3726
rect 25454 3778 25506 3790
rect 25454 3714 25506 3726
rect 26126 3778 26178 3790
rect 26126 3714 26178 3726
rect 26798 3778 26850 3790
rect 26798 3714 26850 3726
rect 27358 3778 27410 3790
rect 27358 3714 27410 3726
rect 29262 3778 29314 3790
rect 29262 3714 29314 3726
rect 29934 3778 29986 3790
rect 29934 3714 29986 3726
rect 30606 3778 30658 3790
rect 30606 3714 30658 3726
rect 31390 3778 31442 3790
rect 31390 3714 31442 3726
rect 20638 3666 20690 3678
rect 20638 3602 20690 3614
rect 21646 3666 21698 3678
rect 21646 3602 21698 3614
rect 22318 3666 22370 3678
rect 22318 3602 22370 3614
rect 22990 3666 23042 3678
rect 22990 3602 23042 3614
rect 23662 3666 23714 3678
rect 23662 3602 23714 3614
rect 28030 3666 28082 3678
rect 28030 3602 28082 3614
rect 34414 3666 34466 3678
rect 34414 3602 34466 3614
rect 34862 3666 34914 3678
rect 34862 3602 34914 3614
rect 35310 3666 35362 3678
rect 35310 3602 35362 3614
rect 17726 3554 17778 3566
rect 17726 3490 17778 3502
rect 18174 3554 18226 3566
rect 18174 3490 18226 3502
rect 18622 3554 18674 3566
rect 18622 3490 18674 3502
rect 19182 3554 19234 3566
rect 19182 3490 19234 3502
rect 19854 3554 19906 3566
rect 19854 3490 19906 3502
rect 20526 3554 20578 3566
rect 20526 3490 20578 3502
rect 21534 3554 21586 3566
rect 21534 3490 21586 3502
rect 22206 3554 22258 3566
rect 22206 3490 22258 3502
rect 22878 3554 22930 3566
rect 22878 3490 22930 3502
rect 23550 3554 23602 3566
rect 23550 3490 23602 3502
rect 24334 3554 24386 3566
rect 24334 3490 24386 3502
rect 25342 3554 25394 3566
rect 25342 3490 25394 3502
rect 26014 3554 26066 3566
rect 26014 3490 26066 3502
rect 26686 3554 26738 3566
rect 26686 3490 26738 3502
rect 27470 3554 27522 3566
rect 27470 3490 27522 3502
rect 28142 3554 28194 3566
rect 28142 3490 28194 3502
rect 29374 3554 29426 3566
rect 29374 3490 29426 3502
rect 30046 3554 30098 3566
rect 30046 3490 30098 3502
rect 30718 3554 30770 3566
rect 30718 3490 30770 3502
rect 31278 3554 31330 3566
rect 31278 3490 31330 3502
rect 31950 3554 32002 3566
rect 31950 3490 32002 3502
rect 16046 3442 16098 3454
rect 16046 3378 16098 3390
rect 16494 3442 16546 3454
rect 16494 3378 16546 3390
rect 32062 3442 32114 3454
rect 32062 3378 32114 3390
rect 33182 3442 33234 3454
rect 33182 3378 33234 3390
rect 33294 3442 33346 3454
rect 33294 3378 33346 3390
rect 33854 3442 33906 3454
rect 33854 3378 33906 3390
rect 33966 3442 34018 3454
rect 33966 3378 34018 3390
rect 35758 3442 35810 3454
rect 35758 3378 35810 3390
rect 1344 3162 38800 3196
rect 1344 3110 10538 3162
rect 10590 3110 10642 3162
rect 10694 3110 10746 3162
rect 10798 3110 19862 3162
rect 19914 3110 19966 3162
rect 20018 3110 20070 3162
rect 20122 3110 29186 3162
rect 29238 3110 29290 3162
rect 29342 3110 29394 3162
rect 29446 3110 38510 3162
rect 38562 3110 38614 3162
rect 38666 3110 38718 3162
rect 38770 3110 38800 3162
rect 1344 3076 38800 3110
<< via1 >>
rect 5876 36822 5928 36874
rect 5980 36822 6032 36874
rect 6084 36822 6136 36874
rect 15200 36822 15252 36874
rect 15304 36822 15356 36874
rect 15408 36822 15460 36874
rect 24524 36822 24576 36874
rect 24628 36822 24680 36874
rect 24732 36822 24784 36874
rect 33848 36822 33900 36874
rect 33952 36822 34004 36874
rect 34056 36822 34108 36874
rect 10538 36038 10590 36090
rect 10642 36038 10694 36090
rect 10746 36038 10798 36090
rect 19862 36038 19914 36090
rect 19966 36038 20018 36090
rect 20070 36038 20122 36090
rect 29186 36038 29238 36090
rect 29290 36038 29342 36090
rect 29394 36038 29446 36090
rect 38510 36038 38562 36090
rect 38614 36038 38666 36090
rect 38718 36038 38770 36090
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 10538 34470 10590 34522
rect 10642 34470 10694 34522
rect 10746 34470 10798 34522
rect 19862 34470 19914 34522
rect 19966 34470 20018 34522
rect 20070 34470 20122 34522
rect 29186 34470 29238 34522
rect 29290 34470 29342 34522
rect 29394 34470 29446 34522
rect 38510 34470 38562 34522
rect 38614 34470 38666 34522
rect 38718 34470 38770 34522
rect 5876 33686 5928 33738
rect 5980 33686 6032 33738
rect 6084 33686 6136 33738
rect 15200 33686 15252 33738
rect 15304 33686 15356 33738
rect 15408 33686 15460 33738
rect 24524 33686 24576 33738
rect 24628 33686 24680 33738
rect 24732 33686 24784 33738
rect 33848 33686 33900 33738
rect 33952 33686 34004 33738
rect 34056 33686 34108 33738
rect 10538 32902 10590 32954
rect 10642 32902 10694 32954
rect 10746 32902 10798 32954
rect 19862 32902 19914 32954
rect 19966 32902 20018 32954
rect 20070 32902 20122 32954
rect 29186 32902 29238 32954
rect 29290 32902 29342 32954
rect 29394 32902 29446 32954
rect 38510 32902 38562 32954
rect 38614 32902 38666 32954
rect 38718 32902 38770 32954
rect 5876 32118 5928 32170
rect 5980 32118 6032 32170
rect 6084 32118 6136 32170
rect 15200 32118 15252 32170
rect 15304 32118 15356 32170
rect 15408 32118 15460 32170
rect 24524 32118 24576 32170
rect 24628 32118 24680 32170
rect 24732 32118 24784 32170
rect 33848 32118 33900 32170
rect 33952 32118 34004 32170
rect 34056 32118 34108 32170
rect 10538 31334 10590 31386
rect 10642 31334 10694 31386
rect 10746 31334 10798 31386
rect 19862 31334 19914 31386
rect 19966 31334 20018 31386
rect 20070 31334 20122 31386
rect 29186 31334 29238 31386
rect 29290 31334 29342 31386
rect 29394 31334 29446 31386
rect 38510 31334 38562 31386
rect 38614 31334 38666 31386
rect 38718 31334 38770 31386
rect 5876 30550 5928 30602
rect 5980 30550 6032 30602
rect 6084 30550 6136 30602
rect 15200 30550 15252 30602
rect 15304 30550 15356 30602
rect 15408 30550 15460 30602
rect 24524 30550 24576 30602
rect 24628 30550 24680 30602
rect 24732 30550 24784 30602
rect 33848 30550 33900 30602
rect 33952 30550 34004 30602
rect 34056 30550 34108 30602
rect 10538 29766 10590 29818
rect 10642 29766 10694 29818
rect 10746 29766 10798 29818
rect 19862 29766 19914 29818
rect 19966 29766 20018 29818
rect 20070 29766 20122 29818
rect 29186 29766 29238 29818
rect 29290 29766 29342 29818
rect 29394 29766 29446 29818
rect 38510 29766 38562 29818
rect 38614 29766 38666 29818
rect 38718 29766 38770 29818
rect 5876 28982 5928 29034
rect 5980 28982 6032 29034
rect 6084 28982 6136 29034
rect 15200 28982 15252 29034
rect 15304 28982 15356 29034
rect 15408 28982 15460 29034
rect 24524 28982 24576 29034
rect 24628 28982 24680 29034
rect 24732 28982 24784 29034
rect 33848 28982 33900 29034
rect 33952 28982 34004 29034
rect 34056 28982 34108 29034
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 5876 27414 5928 27466
rect 5980 27414 6032 27466
rect 6084 27414 6136 27466
rect 15200 27414 15252 27466
rect 15304 27414 15356 27466
rect 15408 27414 15460 27466
rect 24524 27414 24576 27466
rect 24628 27414 24680 27466
rect 24732 27414 24784 27466
rect 33848 27414 33900 27466
rect 33952 27414 34004 27466
rect 34056 27414 34108 27466
rect 10538 26630 10590 26682
rect 10642 26630 10694 26682
rect 10746 26630 10798 26682
rect 19862 26630 19914 26682
rect 19966 26630 20018 26682
rect 20070 26630 20122 26682
rect 29186 26630 29238 26682
rect 29290 26630 29342 26682
rect 29394 26630 29446 26682
rect 38510 26630 38562 26682
rect 38614 26630 38666 26682
rect 38718 26630 38770 26682
rect 5876 25846 5928 25898
rect 5980 25846 6032 25898
rect 6084 25846 6136 25898
rect 15200 25846 15252 25898
rect 15304 25846 15356 25898
rect 15408 25846 15460 25898
rect 24524 25846 24576 25898
rect 24628 25846 24680 25898
rect 24732 25846 24784 25898
rect 33848 25846 33900 25898
rect 33952 25846 34004 25898
rect 34056 25846 34108 25898
rect 10538 25062 10590 25114
rect 10642 25062 10694 25114
rect 10746 25062 10798 25114
rect 19862 25062 19914 25114
rect 19966 25062 20018 25114
rect 20070 25062 20122 25114
rect 29186 25062 29238 25114
rect 29290 25062 29342 25114
rect 29394 25062 29446 25114
rect 38510 25062 38562 25114
rect 38614 25062 38666 25114
rect 38718 25062 38770 25114
rect 5876 24278 5928 24330
rect 5980 24278 6032 24330
rect 6084 24278 6136 24330
rect 15200 24278 15252 24330
rect 15304 24278 15356 24330
rect 15408 24278 15460 24330
rect 24524 24278 24576 24330
rect 24628 24278 24680 24330
rect 24732 24278 24784 24330
rect 33848 24278 33900 24330
rect 33952 24278 34004 24330
rect 34056 24278 34108 24330
rect 10538 23494 10590 23546
rect 10642 23494 10694 23546
rect 10746 23494 10798 23546
rect 19862 23494 19914 23546
rect 19966 23494 20018 23546
rect 20070 23494 20122 23546
rect 29186 23494 29238 23546
rect 29290 23494 29342 23546
rect 29394 23494 29446 23546
rect 38510 23494 38562 23546
rect 38614 23494 38666 23546
rect 38718 23494 38770 23546
rect 5876 22710 5928 22762
rect 5980 22710 6032 22762
rect 6084 22710 6136 22762
rect 15200 22710 15252 22762
rect 15304 22710 15356 22762
rect 15408 22710 15460 22762
rect 24524 22710 24576 22762
rect 24628 22710 24680 22762
rect 24732 22710 24784 22762
rect 33848 22710 33900 22762
rect 33952 22710 34004 22762
rect 34056 22710 34108 22762
rect 10538 21926 10590 21978
rect 10642 21926 10694 21978
rect 10746 21926 10798 21978
rect 19862 21926 19914 21978
rect 19966 21926 20018 21978
rect 20070 21926 20122 21978
rect 29186 21926 29238 21978
rect 29290 21926 29342 21978
rect 29394 21926 29446 21978
rect 38510 21926 38562 21978
rect 38614 21926 38666 21978
rect 38718 21926 38770 21978
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 10538 20358 10590 20410
rect 10642 20358 10694 20410
rect 10746 20358 10798 20410
rect 19862 20358 19914 20410
rect 19966 20358 20018 20410
rect 20070 20358 20122 20410
rect 29186 20358 29238 20410
rect 29290 20358 29342 20410
rect 29394 20358 29446 20410
rect 38510 20358 38562 20410
rect 38614 20358 38666 20410
rect 38718 20358 38770 20410
rect 5876 19574 5928 19626
rect 5980 19574 6032 19626
rect 6084 19574 6136 19626
rect 15200 19574 15252 19626
rect 15304 19574 15356 19626
rect 15408 19574 15460 19626
rect 24524 19574 24576 19626
rect 24628 19574 24680 19626
rect 24732 19574 24784 19626
rect 33848 19574 33900 19626
rect 33952 19574 34004 19626
rect 34056 19574 34108 19626
rect 10538 18790 10590 18842
rect 10642 18790 10694 18842
rect 10746 18790 10798 18842
rect 19862 18790 19914 18842
rect 19966 18790 20018 18842
rect 20070 18790 20122 18842
rect 29186 18790 29238 18842
rect 29290 18790 29342 18842
rect 29394 18790 29446 18842
rect 38510 18790 38562 18842
rect 38614 18790 38666 18842
rect 38718 18790 38770 18842
rect 5876 18006 5928 18058
rect 5980 18006 6032 18058
rect 6084 18006 6136 18058
rect 15200 18006 15252 18058
rect 15304 18006 15356 18058
rect 15408 18006 15460 18058
rect 24524 18006 24576 18058
rect 24628 18006 24680 18058
rect 24732 18006 24784 18058
rect 33848 18006 33900 18058
rect 33952 18006 34004 18058
rect 34056 18006 34108 18058
rect 10538 17222 10590 17274
rect 10642 17222 10694 17274
rect 10746 17222 10798 17274
rect 19862 17222 19914 17274
rect 19966 17222 20018 17274
rect 20070 17222 20122 17274
rect 29186 17222 29238 17274
rect 29290 17222 29342 17274
rect 29394 17222 29446 17274
rect 38510 17222 38562 17274
rect 38614 17222 38666 17274
rect 38718 17222 38770 17274
rect 5876 16438 5928 16490
rect 5980 16438 6032 16490
rect 6084 16438 6136 16490
rect 15200 16438 15252 16490
rect 15304 16438 15356 16490
rect 15408 16438 15460 16490
rect 24524 16438 24576 16490
rect 24628 16438 24680 16490
rect 24732 16438 24784 16490
rect 33848 16438 33900 16490
rect 33952 16438 34004 16490
rect 34056 16438 34108 16490
rect 10538 15654 10590 15706
rect 10642 15654 10694 15706
rect 10746 15654 10798 15706
rect 19862 15654 19914 15706
rect 19966 15654 20018 15706
rect 20070 15654 20122 15706
rect 29186 15654 29238 15706
rect 29290 15654 29342 15706
rect 29394 15654 29446 15706
rect 38510 15654 38562 15706
rect 38614 15654 38666 15706
rect 38718 15654 38770 15706
rect 5876 14870 5928 14922
rect 5980 14870 6032 14922
rect 6084 14870 6136 14922
rect 15200 14870 15252 14922
rect 15304 14870 15356 14922
rect 15408 14870 15460 14922
rect 24524 14870 24576 14922
rect 24628 14870 24680 14922
rect 24732 14870 24784 14922
rect 33848 14870 33900 14922
rect 33952 14870 34004 14922
rect 34056 14870 34108 14922
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 5876 13302 5928 13354
rect 5980 13302 6032 13354
rect 6084 13302 6136 13354
rect 15200 13302 15252 13354
rect 15304 13302 15356 13354
rect 15408 13302 15460 13354
rect 24524 13302 24576 13354
rect 24628 13302 24680 13354
rect 24732 13302 24784 13354
rect 33848 13302 33900 13354
rect 33952 13302 34004 13354
rect 34056 13302 34108 13354
rect 10538 12518 10590 12570
rect 10642 12518 10694 12570
rect 10746 12518 10798 12570
rect 19862 12518 19914 12570
rect 19966 12518 20018 12570
rect 20070 12518 20122 12570
rect 29186 12518 29238 12570
rect 29290 12518 29342 12570
rect 29394 12518 29446 12570
rect 38510 12518 38562 12570
rect 38614 12518 38666 12570
rect 38718 12518 38770 12570
rect 5876 11734 5928 11786
rect 5980 11734 6032 11786
rect 6084 11734 6136 11786
rect 15200 11734 15252 11786
rect 15304 11734 15356 11786
rect 15408 11734 15460 11786
rect 24524 11734 24576 11786
rect 24628 11734 24680 11786
rect 24732 11734 24784 11786
rect 33848 11734 33900 11786
rect 33952 11734 34004 11786
rect 34056 11734 34108 11786
rect 10538 10950 10590 11002
rect 10642 10950 10694 11002
rect 10746 10950 10798 11002
rect 19862 10950 19914 11002
rect 19966 10950 20018 11002
rect 20070 10950 20122 11002
rect 29186 10950 29238 11002
rect 29290 10950 29342 11002
rect 29394 10950 29446 11002
rect 38510 10950 38562 11002
rect 38614 10950 38666 11002
rect 38718 10950 38770 11002
rect 5876 10166 5928 10218
rect 5980 10166 6032 10218
rect 6084 10166 6136 10218
rect 15200 10166 15252 10218
rect 15304 10166 15356 10218
rect 15408 10166 15460 10218
rect 24524 10166 24576 10218
rect 24628 10166 24680 10218
rect 24732 10166 24784 10218
rect 33848 10166 33900 10218
rect 33952 10166 34004 10218
rect 34056 10166 34108 10218
rect 10538 9382 10590 9434
rect 10642 9382 10694 9434
rect 10746 9382 10798 9434
rect 19862 9382 19914 9434
rect 19966 9382 20018 9434
rect 20070 9382 20122 9434
rect 29186 9382 29238 9434
rect 29290 9382 29342 9434
rect 29394 9382 29446 9434
rect 38510 9382 38562 9434
rect 38614 9382 38666 9434
rect 38718 9382 38770 9434
rect 24222 8878 24274 8930
rect 24670 8878 24722 8930
rect 25678 8878 25730 8930
rect 26126 8878 26178 8930
rect 26574 8878 26626 8930
rect 26910 8878 26962 8930
rect 5876 8598 5928 8650
rect 5980 8598 6032 8650
rect 6084 8598 6136 8650
rect 15200 8598 15252 8650
rect 15304 8598 15356 8650
rect 15408 8598 15460 8650
rect 24524 8598 24576 8650
rect 24628 8598 24680 8650
rect 24732 8598 24784 8650
rect 33848 8598 33900 8650
rect 33952 8598 34004 8650
rect 34056 8598 34108 8650
rect 23214 7982 23266 8034
rect 23886 7982 23938 8034
rect 24446 7982 24498 8034
rect 24782 7982 24834 8034
rect 25342 7982 25394 8034
rect 26014 7982 26066 8034
rect 26574 7982 26626 8034
rect 26910 7982 26962 8034
rect 27358 7982 27410 8034
rect 27918 7982 27970 8034
rect 28254 7982 28306 8034
rect 28702 7982 28754 8034
rect 10538 7814 10590 7866
rect 10642 7814 10694 7866
rect 10746 7814 10798 7866
rect 19862 7814 19914 7866
rect 19966 7814 20018 7866
rect 20070 7814 20122 7866
rect 29186 7814 29238 7866
rect 29290 7814 29342 7866
rect 29394 7814 29446 7866
rect 38510 7814 38562 7866
rect 38614 7814 38666 7866
rect 38718 7814 38770 7866
rect 28702 7422 28754 7474
rect 29150 7422 29202 7474
rect 22430 7310 22482 7362
rect 22766 7310 22818 7362
rect 23214 7310 23266 7362
rect 23886 7310 23938 7362
rect 24558 7310 24610 7362
rect 25566 7310 25618 7362
rect 26014 7310 26066 7362
rect 26462 7310 26514 7362
rect 26910 7310 26962 7362
rect 27358 7310 27410 7362
rect 27806 7310 27858 7362
rect 29710 7310 29762 7362
rect 30046 7310 30098 7362
rect 28590 7198 28642 7250
rect 29038 7198 29090 7250
rect 29710 7198 29762 7250
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 21870 6862 21922 6914
rect 22430 6862 22482 6914
rect 27470 6750 27522 6802
rect 28814 6750 28866 6802
rect 22878 6638 22930 6690
rect 23550 6638 23602 6690
rect 24894 6638 24946 6690
rect 25566 6638 25618 6690
rect 24222 6526 24274 6578
rect 26238 6526 26290 6578
rect 26910 6526 26962 6578
rect 28254 6526 28306 6578
rect 29598 6526 29650 6578
rect 29710 6526 29762 6578
rect 30158 6526 30210 6578
rect 21870 6414 21922 6466
rect 22318 6414 22370 6466
rect 22990 6414 23042 6466
rect 23662 6414 23714 6466
rect 24334 6414 24386 6466
rect 25006 6414 25058 6466
rect 25678 6414 25730 6466
rect 26350 6414 26402 6466
rect 27022 6414 27074 6466
rect 28366 6414 28418 6466
rect 30606 6414 30658 6466
rect 31054 6414 31106 6466
rect 31502 6414 31554 6466
rect 31950 6414 32002 6466
rect 10538 6246 10590 6298
rect 10642 6246 10694 6298
rect 10746 6246 10798 6298
rect 19862 6246 19914 6298
rect 19966 6246 20018 6298
rect 20070 6246 20122 6298
rect 29186 6246 29238 6298
rect 29290 6246 29342 6298
rect 29394 6246 29446 6298
rect 38510 6246 38562 6298
rect 38614 6246 38666 6298
rect 38718 6246 38770 6298
rect 25790 6078 25842 6130
rect 26462 6078 26514 6130
rect 27134 6078 27186 6130
rect 27806 6078 27858 6130
rect 28478 6078 28530 6130
rect 29822 6078 29874 6130
rect 30942 6078 30994 6130
rect 31390 6078 31442 6130
rect 31838 6078 31890 6130
rect 27694 5966 27746 6018
rect 29038 5966 29090 6018
rect 29150 5966 29202 6018
rect 30382 5966 30434 6018
rect 21982 5854 22034 5906
rect 22654 5854 22706 5906
rect 23326 5854 23378 5906
rect 23998 5854 24050 5906
rect 24670 5854 24722 5906
rect 25678 5854 25730 5906
rect 26350 5854 26402 5906
rect 27022 5854 27074 5906
rect 28366 5854 28418 5906
rect 29710 5854 29762 5906
rect 20526 5742 20578 5794
rect 20974 5742 21026 5794
rect 21422 5742 21474 5794
rect 32286 5742 32338 5794
rect 32734 5742 32786 5794
rect 33518 5742 33570 5794
rect 20974 5630 21026 5682
rect 21758 5630 21810 5682
rect 22094 5630 22146 5682
rect 22766 5630 22818 5682
rect 23438 5630 23490 5682
rect 24110 5630 24162 5682
rect 24782 5630 24834 5682
rect 30494 5630 30546 5682
rect 5876 5462 5928 5514
rect 5980 5462 6032 5514
rect 6084 5462 6136 5514
rect 15200 5462 15252 5514
rect 15304 5462 15356 5514
rect 15408 5462 15460 5514
rect 24524 5462 24576 5514
rect 24628 5462 24680 5514
rect 24732 5462 24784 5514
rect 33848 5462 33900 5514
rect 33952 5462 34004 5514
rect 34056 5462 34108 5514
rect 21870 5294 21922 5346
rect 23214 5294 23266 5346
rect 23886 5294 23938 5346
rect 24558 5294 24610 5346
rect 25230 5294 25282 5346
rect 26574 5294 26626 5346
rect 27246 5294 27298 5346
rect 27918 5294 27970 5346
rect 28590 5294 28642 5346
rect 29710 5294 29762 5346
rect 30382 5294 30434 5346
rect 19630 5182 19682 5234
rect 20414 5182 20466 5234
rect 20862 5182 20914 5234
rect 21758 5070 21810 5122
rect 23102 5070 23154 5122
rect 23774 5070 23826 5122
rect 25118 5070 25170 5122
rect 25790 5070 25842 5122
rect 25902 5070 25954 5122
rect 26462 5070 26514 5122
rect 27806 5070 27858 5122
rect 28478 5070 28530 5122
rect 29598 5070 29650 5122
rect 30270 5070 30322 5122
rect 30942 5070 30994 5122
rect 22430 4958 22482 5010
rect 24446 4958 24498 5010
rect 27134 4958 27186 5010
rect 31054 4958 31106 5010
rect 31614 4958 31666 5010
rect 31726 4958 31778 5010
rect 33518 4958 33570 5010
rect 19070 4846 19122 4898
rect 19966 4846 20018 4898
rect 22542 4846 22594 4898
rect 32174 4846 32226 4898
rect 32622 4846 32674 4898
rect 33070 4846 33122 4898
rect 33966 4846 34018 4898
rect 34414 4846 34466 4898
rect 10538 4678 10590 4730
rect 10642 4678 10694 4730
rect 10746 4678 10798 4730
rect 19862 4678 19914 4730
rect 19966 4678 20018 4730
rect 20070 4678 20122 4730
rect 29186 4678 29238 4730
rect 29290 4678 29342 4730
rect 29394 4678 29446 4730
rect 38510 4678 38562 4730
rect 38614 4678 38666 4730
rect 38718 4678 38770 4730
rect 18846 4510 18898 4562
rect 19182 4510 19234 4562
rect 23662 4510 23714 4562
rect 24334 4510 24386 4562
rect 24782 4510 24834 4562
rect 25790 4510 25842 4562
rect 27806 4510 27858 4562
rect 28478 4510 28530 4562
rect 29150 4510 29202 4562
rect 29822 4510 29874 4562
rect 31166 4510 31218 4562
rect 31838 4510 31890 4562
rect 34862 4510 34914 4562
rect 20862 4398 20914 4450
rect 21534 4398 21586 4450
rect 22206 4398 22258 4450
rect 26350 4398 26402 4450
rect 26462 4398 26514 4450
rect 27022 4398 27074 4450
rect 30382 4398 30434 4450
rect 30494 4398 30546 4450
rect 31054 4398 31106 4450
rect 31726 4398 31778 4450
rect 20190 4286 20242 4338
rect 22878 4286 22930 4338
rect 23550 4286 23602 4338
rect 24222 4286 24274 4338
rect 25678 4286 25730 4338
rect 27694 4286 27746 4338
rect 28366 4286 28418 4338
rect 29038 4286 29090 4338
rect 29710 4286 29762 4338
rect 32398 4286 32450 4338
rect 19630 4174 19682 4226
rect 33518 4174 33570 4226
rect 33966 4174 34018 4226
rect 34414 4174 34466 4226
rect 20302 4062 20354 4114
rect 20974 4062 21026 4114
rect 21646 4062 21698 4114
rect 22318 4062 22370 4114
rect 22990 4062 23042 4114
rect 27134 4062 27186 4114
rect 32510 4062 32562 4114
rect 5876 3894 5928 3946
rect 5980 3894 6032 3946
rect 6084 3894 6136 3946
rect 15200 3894 15252 3946
rect 15304 3894 15356 3946
rect 15408 3894 15460 3946
rect 24524 3894 24576 3946
rect 24628 3894 24680 3946
rect 24732 3894 24784 3946
rect 33848 3894 33900 3946
rect 33952 3894 34004 3946
rect 34056 3894 34108 3946
rect 16606 3726 16658 3778
rect 19294 3726 19346 3778
rect 19966 3726 20018 3778
rect 24222 3726 24274 3778
rect 25454 3726 25506 3778
rect 26126 3726 26178 3778
rect 26798 3726 26850 3778
rect 27358 3726 27410 3778
rect 29262 3726 29314 3778
rect 29934 3726 29986 3778
rect 30606 3726 30658 3778
rect 31390 3726 31442 3778
rect 20638 3614 20690 3666
rect 21646 3614 21698 3666
rect 22318 3614 22370 3666
rect 22990 3614 23042 3666
rect 23662 3614 23714 3666
rect 28030 3614 28082 3666
rect 34414 3614 34466 3666
rect 34862 3614 34914 3666
rect 35310 3614 35362 3666
rect 17726 3502 17778 3554
rect 18174 3502 18226 3554
rect 18622 3502 18674 3554
rect 19182 3502 19234 3554
rect 19854 3502 19906 3554
rect 20526 3502 20578 3554
rect 21534 3502 21586 3554
rect 22206 3502 22258 3554
rect 22878 3502 22930 3554
rect 23550 3502 23602 3554
rect 24334 3502 24386 3554
rect 25342 3502 25394 3554
rect 26014 3502 26066 3554
rect 26686 3502 26738 3554
rect 27470 3502 27522 3554
rect 28142 3502 28194 3554
rect 29374 3502 29426 3554
rect 30046 3502 30098 3554
rect 30718 3502 30770 3554
rect 31278 3502 31330 3554
rect 31950 3502 32002 3554
rect 16046 3390 16098 3442
rect 16494 3390 16546 3442
rect 32062 3390 32114 3442
rect 33182 3390 33234 3442
rect 33294 3390 33346 3442
rect 33854 3390 33906 3442
rect 33966 3390 34018 3442
rect 35758 3390 35810 3442
rect 10538 3110 10590 3162
rect 10642 3110 10694 3162
rect 10746 3110 10798 3162
rect 19862 3110 19914 3162
rect 19966 3110 20018 3162
rect 20070 3110 20122 3162
rect 29186 3110 29238 3162
rect 29290 3110 29342 3162
rect 29394 3110 29446 3162
rect 38510 3110 38562 3162
rect 38614 3110 38666 3162
rect 38718 3110 38770 3162
<< metal2 >>
rect 5874 36876 6138 36886
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 5874 36810 6138 36820
rect 15198 36876 15462 36886
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15198 36810 15462 36820
rect 24522 36876 24786 36886
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24522 36810 24786 36820
rect 33846 36876 34110 36886
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 33846 36810 34110 36820
rect 10536 36092 10800 36102
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10536 36026 10800 36036
rect 19860 36092 20124 36102
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 19860 36026 20124 36036
rect 29184 36092 29448 36102
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29184 36026 29448 36036
rect 38508 36092 38772 36102
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38508 36026 38772 36036
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 10536 34524 10800 34534
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10536 34458 10800 34468
rect 19860 34524 20124 34534
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 19860 34458 20124 34468
rect 29184 34524 29448 34534
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29184 34458 29448 34468
rect 38508 34524 38772 34534
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38508 34458 38772 34468
rect 5874 33740 6138 33750
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 5874 33674 6138 33684
rect 15198 33740 15462 33750
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15198 33674 15462 33684
rect 24522 33740 24786 33750
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24522 33674 24786 33684
rect 33846 33740 34110 33750
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 33846 33674 34110 33684
rect 10536 32956 10800 32966
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10536 32890 10800 32900
rect 19860 32956 20124 32966
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 19860 32890 20124 32900
rect 29184 32956 29448 32966
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29184 32890 29448 32900
rect 38508 32956 38772 32966
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38508 32890 38772 32900
rect 5874 32172 6138 32182
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 5874 32106 6138 32116
rect 15198 32172 15462 32182
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15198 32106 15462 32116
rect 24522 32172 24786 32182
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24522 32106 24786 32116
rect 33846 32172 34110 32182
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 33846 32106 34110 32116
rect 10536 31388 10800 31398
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10536 31322 10800 31332
rect 19860 31388 20124 31398
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 19860 31322 20124 31332
rect 29184 31388 29448 31398
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29184 31322 29448 31332
rect 38508 31388 38772 31398
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38508 31322 38772 31332
rect 5874 30604 6138 30614
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 5874 30538 6138 30548
rect 15198 30604 15462 30614
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15198 30538 15462 30548
rect 24522 30604 24786 30614
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24522 30538 24786 30548
rect 33846 30604 34110 30614
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 33846 30538 34110 30548
rect 10536 29820 10800 29830
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10536 29754 10800 29764
rect 19860 29820 20124 29830
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 19860 29754 20124 29764
rect 29184 29820 29448 29830
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29184 29754 29448 29764
rect 38508 29820 38772 29830
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38508 29754 38772 29764
rect 5874 29036 6138 29046
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 5874 28970 6138 28980
rect 15198 29036 15462 29046
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15198 28970 15462 28980
rect 24522 29036 24786 29046
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24522 28970 24786 28980
rect 33846 29036 34110 29046
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 33846 28970 34110 28980
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 5874 27468 6138 27478
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 5874 27402 6138 27412
rect 15198 27468 15462 27478
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15198 27402 15462 27412
rect 24522 27468 24786 27478
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24522 27402 24786 27412
rect 33846 27468 34110 27478
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 33846 27402 34110 27412
rect 10536 26684 10800 26694
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10536 26618 10800 26628
rect 19860 26684 20124 26694
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 19860 26618 20124 26628
rect 29184 26684 29448 26694
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29184 26618 29448 26628
rect 38508 26684 38772 26694
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38508 26618 38772 26628
rect 5874 25900 6138 25910
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 5874 25834 6138 25844
rect 15198 25900 15462 25910
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15198 25834 15462 25844
rect 24522 25900 24786 25910
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24522 25834 24786 25844
rect 33846 25900 34110 25910
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 33846 25834 34110 25844
rect 10536 25116 10800 25126
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10536 25050 10800 25060
rect 19860 25116 20124 25126
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 19860 25050 20124 25060
rect 29184 25116 29448 25126
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29184 25050 29448 25060
rect 38508 25116 38772 25126
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38508 25050 38772 25060
rect 5874 24332 6138 24342
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 5874 24266 6138 24276
rect 15198 24332 15462 24342
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15198 24266 15462 24276
rect 24522 24332 24786 24342
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24522 24266 24786 24276
rect 33846 24332 34110 24342
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 33846 24266 34110 24276
rect 10536 23548 10800 23558
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10536 23482 10800 23492
rect 19860 23548 20124 23558
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 19860 23482 20124 23492
rect 29184 23548 29448 23558
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29184 23482 29448 23492
rect 38508 23548 38772 23558
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38508 23482 38772 23492
rect 5874 22764 6138 22774
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 5874 22698 6138 22708
rect 15198 22764 15462 22774
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15198 22698 15462 22708
rect 24522 22764 24786 22774
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24522 22698 24786 22708
rect 33846 22764 34110 22774
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 33846 22698 34110 22708
rect 10536 21980 10800 21990
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10536 21914 10800 21924
rect 19860 21980 20124 21990
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 19860 21914 20124 21924
rect 29184 21980 29448 21990
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29184 21914 29448 21924
rect 38508 21980 38772 21990
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38508 21914 38772 21924
rect 5874 21196 6138 21206
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 10536 20412 10800 20422
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10536 20346 10800 20356
rect 19860 20412 20124 20422
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 19860 20346 20124 20356
rect 29184 20412 29448 20422
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29184 20346 29448 20356
rect 38508 20412 38772 20422
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38508 20346 38772 20356
rect 5874 19628 6138 19638
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 5874 19562 6138 19572
rect 15198 19628 15462 19638
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15198 19562 15462 19572
rect 24522 19628 24786 19638
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24522 19562 24786 19572
rect 33846 19628 34110 19638
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 33846 19562 34110 19572
rect 10536 18844 10800 18854
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10536 18778 10800 18788
rect 19860 18844 20124 18854
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 19860 18778 20124 18788
rect 29184 18844 29448 18854
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29184 18778 29448 18788
rect 38508 18844 38772 18854
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38508 18778 38772 18788
rect 5874 18060 6138 18070
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 5874 17994 6138 18004
rect 15198 18060 15462 18070
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15198 17994 15462 18004
rect 24522 18060 24786 18070
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24522 17994 24786 18004
rect 33846 18060 34110 18070
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 33846 17994 34110 18004
rect 10536 17276 10800 17286
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10536 17210 10800 17220
rect 19860 17276 20124 17286
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 19860 17210 20124 17220
rect 29184 17276 29448 17286
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29184 17210 29448 17220
rect 38508 17276 38772 17286
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38508 17210 38772 17220
rect 5874 16492 6138 16502
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 5874 16426 6138 16436
rect 15198 16492 15462 16502
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15198 16426 15462 16436
rect 24522 16492 24786 16502
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24522 16426 24786 16436
rect 33846 16492 34110 16502
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 33846 16426 34110 16436
rect 10536 15708 10800 15718
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10536 15642 10800 15652
rect 19860 15708 20124 15718
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 19860 15642 20124 15652
rect 29184 15708 29448 15718
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29184 15642 29448 15652
rect 38508 15708 38772 15718
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38508 15642 38772 15652
rect 5874 14924 6138 14934
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 5874 14858 6138 14868
rect 15198 14924 15462 14934
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15198 14858 15462 14868
rect 24522 14924 24786 14934
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24522 14858 24786 14868
rect 33846 14924 34110 14934
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 33846 14858 34110 14868
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 5874 13356 6138 13366
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 5874 13290 6138 13300
rect 15198 13356 15462 13366
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15198 13290 15462 13300
rect 24522 13356 24786 13366
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24522 13290 24786 13300
rect 33846 13356 34110 13366
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 33846 13290 34110 13300
rect 10536 12572 10800 12582
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10536 12506 10800 12516
rect 19860 12572 20124 12582
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 19860 12506 20124 12516
rect 29184 12572 29448 12582
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29184 12506 29448 12516
rect 38508 12572 38772 12582
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38508 12506 38772 12516
rect 5874 11788 6138 11798
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 5874 11722 6138 11732
rect 15198 11788 15462 11798
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15198 11722 15462 11732
rect 24522 11788 24786 11798
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24522 11722 24786 11732
rect 33846 11788 34110 11798
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 33846 11722 34110 11732
rect 10536 11004 10800 11014
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10536 10938 10800 10948
rect 19860 11004 20124 11014
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 19860 10938 20124 10948
rect 29184 11004 29448 11014
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29184 10938 29448 10948
rect 38508 11004 38772 11014
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38508 10938 38772 10948
rect 5874 10220 6138 10230
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 5874 10154 6138 10164
rect 15198 10220 15462 10230
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15198 10154 15462 10164
rect 24522 10220 24786 10230
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24522 10154 24786 10164
rect 33846 10220 34110 10230
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 33846 10154 34110 10164
rect 10536 9436 10800 9446
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10536 9370 10800 9380
rect 19860 9436 20124 9446
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 19860 9370 20124 9380
rect 29184 9436 29448 9446
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29184 9370 29448 9380
rect 38508 9436 38772 9446
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38508 9370 38772 9380
rect 24220 8932 24276 8942
rect 5874 8652 6138 8662
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 5874 8586 6138 8596
rect 15198 8652 15462 8662
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15198 8586 15462 8596
rect 23212 8036 23268 8046
rect 23100 7980 23212 8036
rect 10536 7868 10800 7878
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10536 7802 10800 7812
rect 19860 7868 20124 7878
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 19860 7802 20124 7812
rect 22428 7362 22484 7374
rect 22428 7310 22430 7362
rect 22482 7310 22484 7362
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 21868 6914 21924 6926
rect 21868 6862 21870 6914
rect 21922 6862 21924 6914
rect 19628 6804 19684 6814
rect 10536 6300 10800 6310
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10536 6234 10800 6244
rect 5874 5516 6138 5526
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 5874 5450 6138 5460
rect 15198 5516 15462 5526
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15198 5450 15462 5460
rect 19628 5234 19684 6748
rect 21868 6692 21924 6862
rect 22428 6914 22484 7310
rect 22428 6862 22430 6914
rect 22482 6862 22484 6914
rect 22428 6850 22484 6862
rect 22764 7364 22820 7374
rect 23100 7364 23156 7980
rect 23212 7904 23268 7980
rect 23884 8034 23940 8046
rect 23884 7982 23886 8034
rect 23938 7982 23940 8034
rect 22764 7362 23156 7364
rect 22764 7310 22766 7362
rect 22818 7310 23156 7362
rect 22764 7308 23156 7310
rect 23212 7362 23268 7374
rect 23212 7310 23214 7362
rect 23266 7310 23268 7362
rect 21756 6636 21924 6692
rect 21980 6804 22036 6814
rect 19860 6300 20124 6310
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 19860 6234 20124 6244
rect 21420 5908 21476 5918
rect 20524 5794 20580 5806
rect 20524 5742 20526 5794
rect 20578 5742 20580 5794
rect 19628 5182 19630 5234
rect 19682 5182 19684 5234
rect 19628 5170 19684 5182
rect 20412 5236 20468 5246
rect 20524 5236 20580 5742
rect 20972 5794 21028 5806
rect 20972 5742 20974 5794
rect 21026 5742 21028 5794
rect 20972 5682 21028 5742
rect 20972 5630 20974 5682
rect 21026 5630 21028 5682
rect 20412 5234 20580 5236
rect 20412 5182 20414 5234
rect 20466 5182 20580 5234
rect 20412 5180 20580 5182
rect 20860 5236 20916 5246
rect 20972 5236 21028 5630
rect 20860 5234 21028 5236
rect 20860 5182 20862 5234
rect 20914 5182 21028 5234
rect 20860 5180 21028 5182
rect 21420 5794 21476 5852
rect 21420 5742 21422 5794
rect 21474 5742 21476 5794
rect 19068 4900 19124 4910
rect 19964 4900 20020 4910
rect 20412 4900 20468 5180
rect 19068 4898 19236 4900
rect 19068 4846 19070 4898
rect 19122 4846 19236 4898
rect 19068 4844 19236 4846
rect 19068 4834 19124 4844
rect 10536 4732 10800 4742
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10536 4666 10800 4676
rect 18844 4564 18900 4574
rect 18844 4470 18900 4508
rect 19180 4564 19236 4844
rect 5874 3948 6138 3958
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 5874 3882 6138 3892
rect 15198 3948 15462 3958
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15198 3882 15462 3892
rect 16604 3780 16660 3790
rect 16604 3686 16660 3724
rect 12572 3556 12628 3566
rect 2716 3444 2772 3454
rect 2716 800 2772 3388
rect 10536 3164 10800 3174
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10536 3098 10800 3108
rect 12572 800 12628 3500
rect 17724 3556 17780 3566
rect 17724 3462 17780 3500
rect 18172 3556 18228 3566
rect 18172 3462 18228 3500
rect 18620 3556 18676 3566
rect 18620 3462 18676 3500
rect 19180 3554 19236 4508
rect 19628 4898 20468 4900
rect 19628 4846 19966 4898
rect 20018 4846 20468 4898
rect 19628 4844 20468 4846
rect 19628 4226 19684 4844
rect 19964 4834 20020 4844
rect 19860 4732 20124 4742
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 19860 4666 20124 4676
rect 20188 4564 20244 4574
rect 20188 4452 20244 4508
rect 19628 4174 19630 4226
rect 19682 4174 19684 4226
rect 19292 4116 19348 4126
rect 19292 3778 19348 4060
rect 19292 3726 19294 3778
rect 19346 3726 19348 3778
rect 19292 3714 19348 3726
rect 19180 3502 19182 3554
rect 19234 3502 19236 3554
rect 19180 3490 19236 3502
rect 19628 3556 19684 4174
rect 19964 4396 20244 4452
rect 19964 3778 20020 4396
rect 19964 3726 19966 3778
rect 20018 3726 20020 3778
rect 19964 3714 20020 3726
rect 20188 4338 20244 4396
rect 20860 4450 20916 5180
rect 20860 4398 20862 4450
rect 20914 4398 20916 4450
rect 20860 4386 20916 4398
rect 20188 4286 20190 4338
rect 20242 4286 20244 4338
rect 20188 3668 20244 4286
rect 20300 4116 20356 4126
rect 20300 4022 20356 4060
rect 20972 4114 21028 4126
rect 20972 4062 20974 4114
rect 21026 4062 21028 4114
rect 20188 3602 20244 3612
rect 20636 3668 20692 3678
rect 20636 3574 20692 3612
rect 20972 3668 21028 4062
rect 21420 4116 21476 5742
rect 21756 5682 21812 6636
rect 21868 6468 21924 6478
rect 21980 6468 22036 6748
rect 22316 6468 22372 6478
rect 21868 6466 22372 6468
rect 21868 6414 21870 6466
rect 21922 6414 22318 6466
rect 22370 6414 22372 6466
rect 21868 6412 22372 6414
rect 21868 6402 21924 6412
rect 21980 5908 22036 5918
rect 22316 5908 22372 6412
rect 22652 5908 22708 5918
rect 22764 5908 22820 7308
rect 22876 6692 22932 6702
rect 23212 6692 23268 7310
rect 23884 7362 23940 7982
rect 24220 8036 24276 8876
rect 24668 8932 24724 8942
rect 25676 8932 25732 8942
rect 24668 8930 24948 8932
rect 24668 8878 24670 8930
rect 24722 8878 24948 8930
rect 24668 8876 24948 8878
rect 24668 8866 24724 8876
rect 24522 8652 24786 8662
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24522 8586 24786 8596
rect 24220 7970 24276 7980
rect 24444 8036 24500 8046
rect 23884 7310 23886 7362
rect 23938 7310 23940 7362
rect 23548 6692 23604 6702
rect 23884 6692 23940 7310
rect 24444 7252 24500 7980
rect 24780 8036 24836 8046
rect 24892 8036 24948 8876
rect 25676 8838 25732 8876
rect 26124 8932 26180 8942
rect 26124 8838 26180 8876
rect 26572 8932 26628 8942
rect 26572 8838 26628 8876
rect 26908 8932 26964 8942
rect 26908 8838 26964 8876
rect 33846 8652 34110 8662
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 33846 8586 34110 8596
rect 24780 8034 24948 8036
rect 24780 7982 24782 8034
rect 24834 7982 24948 8034
rect 24780 7980 24948 7982
rect 24780 7970 24836 7980
rect 24556 7362 24612 7374
rect 24556 7310 24558 7362
rect 24610 7310 24612 7362
rect 24556 7252 24612 7310
rect 22876 6690 23940 6692
rect 22876 6638 22878 6690
rect 22930 6638 23550 6690
rect 23602 6638 23940 6690
rect 22876 6636 23940 6638
rect 22876 6626 22932 6636
rect 23548 6626 23604 6636
rect 22988 6468 23044 6478
rect 22988 6374 23044 6412
rect 23660 6468 23716 6478
rect 23324 5908 23380 5918
rect 22316 5906 23380 5908
rect 22316 5854 22654 5906
rect 22706 5854 23326 5906
rect 23378 5854 23380 5906
rect 22316 5852 23380 5854
rect 21980 5814 22036 5852
rect 22652 5842 22708 5852
rect 21756 5630 21758 5682
rect 21810 5630 21812 5682
rect 21756 5124 21812 5630
rect 22092 5682 22148 5694
rect 22092 5630 22094 5682
rect 22146 5630 22148 5682
rect 21868 5348 21924 5358
rect 22092 5348 22148 5630
rect 22764 5684 22820 5694
rect 22764 5590 22820 5628
rect 23212 5684 23268 5694
rect 21868 5346 22148 5348
rect 21868 5294 21870 5346
rect 21922 5294 22148 5346
rect 21868 5292 22148 5294
rect 21868 5282 21924 5292
rect 21420 4050 21476 4060
rect 21532 5122 21812 5124
rect 21532 5070 21758 5122
rect 21810 5070 21812 5122
rect 21532 5068 21812 5070
rect 21532 4452 21588 5068
rect 21756 5058 21812 5068
rect 22092 5012 22148 5292
rect 23212 5346 23268 5628
rect 23212 5294 23214 5346
rect 23266 5294 23268 5346
rect 23212 5282 23268 5294
rect 23100 5124 23156 5134
rect 23324 5124 23380 5852
rect 23436 5684 23492 5694
rect 23660 5684 23716 6412
rect 23884 5908 23940 6636
rect 24332 7196 24612 7252
rect 24220 6580 24276 6590
rect 24332 6580 24388 7196
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 24892 6692 24948 7980
rect 25340 8036 25396 8046
rect 25340 7942 25396 7980
rect 26012 8034 26068 8046
rect 26572 8036 26628 8046
rect 26012 7982 26014 8034
rect 26066 7982 26068 8034
rect 25564 7364 25620 7374
rect 25564 6692 25620 7308
rect 26012 7364 26068 7982
rect 26012 7270 26068 7308
rect 26460 8034 26628 8036
rect 26460 7982 26574 8034
rect 26626 7982 26628 8034
rect 26460 7980 26628 7982
rect 26460 7362 26516 7980
rect 26572 7970 26628 7980
rect 26908 8034 26964 8046
rect 26908 7982 26910 8034
rect 26962 7982 26964 8034
rect 26460 7310 26462 7362
rect 26514 7310 26516 7362
rect 24892 6690 25620 6692
rect 24892 6638 24894 6690
rect 24946 6638 25566 6690
rect 25618 6638 25620 6690
rect 24892 6636 25620 6638
rect 24892 6626 24948 6636
rect 24220 6578 24388 6580
rect 24220 6526 24222 6578
rect 24274 6526 24388 6578
rect 24220 6524 24388 6526
rect 24220 6514 24276 6524
rect 24332 6466 24388 6524
rect 24332 6414 24334 6466
rect 24386 6414 24388 6466
rect 23996 5908 24052 5918
rect 23884 5906 24052 5908
rect 23884 5854 23998 5906
rect 24050 5854 24052 5906
rect 23884 5852 24052 5854
rect 23492 5628 23716 5684
rect 23436 5590 23492 5628
rect 23100 5122 23492 5124
rect 23100 5070 23102 5122
rect 23154 5070 23492 5122
rect 23100 5068 23492 5070
rect 23100 5058 23156 5068
rect 22428 5012 22484 5022
rect 22092 5010 22596 5012
rect 22092 4958 22430 5010
rect 22482 4958 22596 5010
rect 22092 4956 22596 4958
rect 22428 4946 22484 4956
rect 22540 4898 22596 4956
rect 22540 4846 22542 4898
rect 22594 4846 22596 4898
rect 20972 3602 21028 3612
rect 19628 3490 19684 3500
rect 19852 3556 19908 3566
rect 19852 3462 19908 3500
rect 20524 3556 20580 3566
rect 20524 3462 20580 3500
rect 21532 3556 21588 4396
rect 22204 4452 22260 4462
rect 21644 4114 21700 4126
rect 21644 4062 21646 4114
rect 21698 4062 21700 4114
rect 21644 3668 21700 4062
rect 21644 3574 21700 3612
rect 16044 3444 16100 3454
rect 16044 3350 16100 3388
rect 16492 3444 16548 3454
rect 21532 3424 21588 3500
rect 22204 3556 22260 4396
rect 22540 4340 22596 4846
rect 22876 4340 22932 4350
rect 23436 4340 23492 5068
rect 23660 4562 23716 5628
rect 23884 5348 23940 5358
rect 23996 5348 24052 5852
rect 24108 5684 24164 5694
rect 24332 5684 24388 6414
rect 25004 6468 25060 6478
rect 25004 6374 25060 6412
rect 24668 5906 24724 5918
rect 24668 5854 24670 5906
rect 24722 5854 24724 5906
rect 24668 5684 24724 5854
rect 24164 5628 24724 5684
rect 24780 5684 24836 5694
rect 24780 5682 24948 5684
rect 24780 5630 24782 5682
rect 24834 5630 24948 5682
rect 24780 5628 24948 5630
rect 24108 5590 24164 5628
rect 23884 5346 24052 5348
rect 23884 5294 23886 5346
rect 23938 5294 24052 5346
rect 23884 5292 24052 5294
rect 23772 5124 23828 5134
rect 23884 5124 23940 5292
rect 23772 5122 23940 5124
rect 23772 5070 23774 5122
rect 23826 5070 23940 5122
rect 23772 5068 23940 5070
rect 23772 5058 23828 5068
rect 23996 5012 24052 5292
rect 23996 4946 24052 4956
rect 24332 5348 24388 5628
rect 24780 5618 24836 5628
rect 24522 5516 24786 5526
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24522 5450 24786 5460
rect 24556 5348 24612 5358
rect 24892 5348 24948 5628
rect 25228 5348 25284 6636
rect 25564 6626 25620 6636
rect 26236 6804 26292 6814
rect 26236 6578 26292 6748
rect 26460 6804 26516 7310
rect 26460 6738 26516 6748
rect 26908 7364 26964 7982
rect 27356 8036 27412 8046
rect 27916 8036 27972 8046
rect 27356 7364 27412 7980
rect 26964 7362 27412 7364
rect 26964 7310 27358 7362
rect 27410 7310 27412 7362
rect 26964 7308 27412 7310
rect 26236 6526 26238 6578
rect 26290 6526 26292 6578
rect 25676 6468 25732 6478
rect 25676 6374 25732 6412
rect 25788 6132 25844 6142
rect 25788 6038 25844 6076
rect 24332 5346 24612 5348
rect 24332 5294 24558 5346
rect 24610 5294 24612 5346
rect 24332 5292 24612 5294
rect 24332 5124 24388 5292
rect 24556 5282 24612 5292
rect 24780 5346 25284 5348
rect 24780 5294 25230 5346
rect 25282 5294 25284 5346
rect 24780 5292 25284 5294
rect 23660 4510 23662 4562
rect 23714 4510 23716 4562
rect 23660 4498 23716 4510
rect 24332 4562 24388 5068
rect 24332 4510 24334 4562
rect 24386 4510 24388 4562
rect 24332 4498 24388 4510
rect 24444 5010 24500 5022
rect 24444 4958 24446 5010
rect 24498 4958 24500 5010
rect 23548 4340 23604 4350
rect 22540 4338 23044 4340
rect 22540 4286 22878 4338
rect 22930 4286 23044 4338
rect 22540 4284 23044 4286
rect 22876 4274 22932 4284
rect 22316 4114 22372 4126
rect 22316 4062 22318 4114
rect 22370 4062 22372 4114
rect 22316 3668 22372 4062
rect 22316 3574 22372 3612
rect 22988 4114 23044 4284
rect 22988 4062 22990 4114
rect 23042 4062 23044 4114
rect 22988 3668 23044 4062
rect 22988 3574 23044 3612
rect 23436 4284 23548 4340
rect 22204 3424 22260 3500
rect 22876 3556 22932 3566
rect 22876 3462 22932 3500
rect 16492 3350 16548 3388
rect 19860 3164 20124 3174
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 19860 3098 20124 3108
rect 22428 924 22820 980
rect 22428 800 22484 924
rect 2688 0 2800 800
rect 7616 0 7728 800
rect 12544 0 12656 800
rect 17472 0 17584 800
rect 22400 0 22512 800
rect 22764 756 22820 924
rect 23436 756 23492 4284
rect 23548 4208 23604 4284
rect 24220 4340 24276 4350
rect 24444 4340 24500 4958
rect 24276 4284 24500 4340
rect 24780 5012 24836 5292
rect 25228 5282 25284 5292
rect 25676 5906 25732 5918
rect 25676 5854 25678 5906
rect 25730 5854 25732 5906
rect 25116 5124 25172 5134
rect 25116 5030 25172 5068
rect 25676 5124 25732 5854
rect 25788 5124 25844 5134
rect 25900 5124 25956 5134
rect 25732 5122 25956 5124
rect 25732 5070 25790 5122
rect 25842 5070 25902 5122
rect 25954 5070 25956 5122
rect 25732 5068 25956 5070
rect 25676 5058 25732 5068
rect 24780 4562 24836 4956
rect 25788 4564 25844 5068
rect 25900 5058 25956 5068
rect 26236 4564 26292 6526
rect 26908 6578 26964 7308
rect 27356 7298 27412 7308
rect 27804 8034 27972 8036
rect 27804 7982 27918 8034
rect 27970 7982 27972 8034
rect 27804 7980 27972 7982
rect 27804 7362 27860 7980
rect 27916 7970 27972 7980
rect 28252 8036 28308 8046
rect 28252 7942 28308 7980
rect 28700 8036 28756 8046
rect 28700 7942 28756 7980
rect 29184 7868 29448 7878
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29184 7802 29448 7812
rect 38508 7868 38772 7878
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38508 7802 38772 7812
rect 28700 7476 28756 7486
rect 29148 7476 29204 7486
rect 27804 7310 27806 7362
rect 27858 7310 27860 7362
rect 27468 6804 27524 6814
rect 27804 6804 27860 7310
rect 27524 6748 27860 6804
rect 28588 7474 29204 7476
rect 28588 7422 28702 7474
rect 28754 7422 29150 7474
rect 29202 7422 29204 7474
rect 28588 7420 29204 7422
rect 28588 7250 28644 7420
rect 28700 7410 28756 7420
rect 29148 7410 29204 7420
rect 29708 7362 29764 7374
rect 29708 7310 29710 7362
rect 29762 7310 29764 7362
rect 28588 7198 28590 7250
rect 28642 7198 28644 7250
rect 27468 6710 27524 6748
rect 26908 6526 26910 6578
rect 26962 6526 26964 6578
rect 26348 6466 26404 6478
rect 26348 6414 26350 6466
rect 26402 6414 26404 6466
rect 26348 6132 26404 6414
rect 26348 6066 26404 6076
rect 26460 6468 26516 6478
rect 26460 6130 26516 6412
rect 26460 6078 26462 6130
rect 26514 6078 26516 6130
rect 26348 5906 26404 5918
rect 26348 5854 26350 5906
rect 26402 5854 26404 5906
rect 26348 5124 26404 5854
rect 26460 5348 26516 6078
rect 26908 5908 26964 6526
rect 27020 6468 27076 6478
rect 27020 6132 27076 6412
rect 27132 6132 27188 6142
rect 27020 6130 27188 6132
rect 27020 6078 27134 6130
rect 27186 6078 27188 6130
rect 27020 6076 27188 6078
rect 27020 5908 27076 5918
rect 26908 5906 27076 5908
rect 26908 5854 27022 5906
rect 27074 5854 27076 5906
rect 26908 5852 27076 5854
rect 26572 5348 26628 5358
rect 26460 5346 26628 5348
rect 26460 5294 26574 5346
rect 26626 5294 26628 5346
rect 26460 5292 26628 5294
rect 26572 5282 26628 5292
rect 26460 5124 26516 5134
rect 26348 5122 26964 5124
rect 26348 5070 26462 5122
rect 26514 5070 26964 5122
rect 26348 5068 26964 5070
rect 26460 5058 26516 5068
rect 26908 5012 26964 5068
rect 27020 5012 27076 5852
rect 27132 5348 27188 6076
rect 27692 6018 27748 6748
rect 28252 6578 28308 6590
rect 28252 6526 28254 6578
rect 28306 6526 28308 6578
rect 27692 5966 27694 6018
rect 27746 5966 27748 6018
rect 27244 5348 27300 5358
rect 27132 5346 27300 5348
rect 27132 5294 27246 5346
rect 27298 5294 27300 5346
rect 27132 5292 27300 5294
rect 27132 5012 27188 5022
rect 26908 5010 27188 5012
rect 26908 4958 27134 5010
rect 27186 4958 27188 5010
rect 26908 4956 27188 4958
rect 27132 4900 27188 4956
rect 27132 4834 27188 4844
rect 24780 4510 24782 4562
rect 24834 4510 24836 4562
rect 24220 4246 24276 4284
rect 24780 4116 24836 4510
rect 25452 4562 26292 4564
rect 25452 4510 25790 4562
rect 25842 4510 26292 4562
rect 25452 4508 26292 4510
rect 24332 4060 24836 4116
rect 25340 4340 25396 4350
rect 24220 3780 24276 3790
rect 24332 3780 24388 4060
rect 24522 3948 24786 3958
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24522 3882 24786 3892
rect 24220 3778 24388 3780
rect 24220 3726 24222 3778
rect 24274 3726 24388 3778
rect 24220 3724 24388 3726
rect 24220 3714 24276 3724
rect 23660 3668 23716 3678
rect 23660 3574 23716 3612
rect 24332 3668 24388 3724
rect 23548 3556 23604 3566
rect 23548 3462 23604 3500
rect 24332 3554 24388 3612
rect 24332 3502 24334 3554
rect 24386 3502 24388 3554
rect 24332 3490 24388 3502
rect 25340 3556 25396 4284
rect 25452 3778 25508 4508
rect 25788 4498 25844 4508
rect 25676 4340 25732 4350
rect 25676 4246 25732 4284
rect 25452 3726 25454 3778
rect 25506 3726 25508 3778
rect 25452 3714 25508 3726
rect 26124 3778 26180 4508
rect 26236 4452 26292 4508
rect 27244 4564 27300 5292
rect 27692 5124 27748 5966
rect 27804 6132 27860 6142
rect 27804 5348 27860 6076
rect 28252 6132 28308 6526
rect 28588 6580 28644 7198
rect 29036 7250 29092 7262
rect 29036 7198 29038 7250
rect 29090 7198 29092 7250
rect 28812 6804 28868 6814
rect 28812 6710 28868 6748
rect 28364 6468 28420 6478
rect 28364 6374 28420 6412
rect 28476 6132 28532 6142
rect 28588 6132 28644 6524
rect 28308 6130 28644 6132
rect 28308 6078 28478 6130
rect 28530 6078 28644 6130
rect 28308 6076 28644 6078
rect 28252 6066 28308 6076
rect 28476 6066 28532 6076
rect 28364 5906 28420 5918
rect 28364 5854 28366 5906
rect 28418 5854 28420 5906
rect 27916 5348 27972 5358
rect 27804 5346 27972 5348
rect 27804 5294 27918 5346
rect 27970 5294 27972 5346
rect 27804 5292 27972 5294
rect 27916 5282 27972 5292
rect 27804 5124 27860 5134
rect 28364 5124 28420 5854
rect 28588 5346 28644 6076
rect 29036 6468 29092 7198
rect 29708 7250 29764 7310
rect 29708 7198 29710 7250
rect 29762 7198 29764 7250
rect 29708 7186 29764 7198
rect 30044 7362 30100 7374
rect 30044 7310 30046 7362
rect 30098 7310 30100 7362
rect 30044 6804 30100 7310
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 30044 6738 30100 6748
rect 30940 6692 30996 6702
rect 30996 6636 31892 6692
rect 29596 6580 29652 6590
rect 29708 6580 29764 6590
rect 29652 6578 29764 6580
rect 29652 6526 29710 6578
rect 29762 6526 29764 6578
rect 29652 6524 29764 6526
rect 29596 6486 29652 6524
rect 29036 6020 29092 6412
rect 29184 6300 29448 6310
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29184 6234 29448 6244
rect 29708 6132 29764 6524
rect 30156 6580 30212 6590
rect 30212 6524 30436 6580
rect 30156 6486 30212 6524
rect 30380 6468 30436 6524
rect 30604 6468 30660 6478
rect 30380 6466 30660 6468
rect 30380 6414 30606 6466
rect 30658 6414 30660 6466
rect 30380 6412 30660 6414
rect 29820 6132 29876 6142
rect 29708 6130 29876 6132
rect 29708 6078 29822 6130
rect 29874 6078 29876 6130
rect 29708 6076 29876 6078
rect 29820 6066 29876 6076
rect 29148 6020 29204 6030
rect 29036 6018 29764 6020
rect 29036 5966 29038 6018
rect 29090 5966 29150 6018
rect 29202 5966 29764 6018
rect 29036 5964 29764 5966
rect 29036 5954 29092 5964
rect 29148 5954 29204 5964
rect 28588 5294 28590 5346
rect 28642 5294 28644 5346
rect 28588 5282 28644 5294
rect 29708 5906 29764 5964
rect 29708 5854 29710 5906
rect 29762 5854 29764 5906
rect 29708 5346 29764 5854
rect 29708 5294 29710 5346
rect 29762 5294 29764 5346
rect 29708 5236 29764 5294
rect 30380 6018 30436 6412
rect 30604 6402 30660 6412
rect 30940 6130 30996 6636
rect 30940 6078 30942 6130
rect 30994 6078 30996 6130
rect 30940 6066 30996 6078
rect 31052 6466 31108 6478
rect 31052 6414 31054 6466
rect 31106 6414 31108 6466
rect 30380 5966 30382 6018
rect 30434 5966 30436 6018
rect 30380 5346 30436 5966
rect 30380 5294 30382 5346
rect 30434 5294 30436 5346
rect 29708 5180 30324 5236
rect 28476 5124 28532 5134
rect 27692 5122 28532 5124
rect 27692 5070 27806 5122
rect 27858 5070 28478 5122
rect 28530 5070 28532 5122
rect 27692 5068 28532 5070
rect 27804 5058 27860 5068
rect 28476 5058 28532 5068
rect 29596 5124 29652 5134
rect 29708 5124 29764 5180
rect 29596 5122 29764 5124
rect 29596 5070 29598 5122
rect 29650 5070 29764 5122
rect 29596 5068 29764 5070
rect 30268 5122 30324 5180
rect 30268 5070 30270 5122
rect 30322 5070 30324 5122
rect 29596 5058 29652 5068
rect 29820 5012 29876 5022
rect 27244 4498 27300 4508
rect 27692 4900 27748 4910
rect 26348 4452 26404 4462
rect 26460 4452 26516 4462
rect 27020 4452 27076 4462
rect 26236 4450 27076 4452
rect 26236 4398 26350 4450
rect 26402 4398 26462 4450
rect 26514 4398 27022 4450
rect 27074 4398 27076 4450
rect 26236 4396 27076 4398
rect 26348 4386 26404 4396
rect 26460 4386 26516 4396
rect 26124 3726 26126 3778
rect 26178 3726 26180 3778
rect 26124 3714 26180 3726
rect 26796 3778 26852 4396
rect 27020 4340 27076 4396
rect 27020 4284 27412 4340
rect 27132 4116 27188 4126
rect 27132 4022 27188 4060
rect 26796 3726 26798 3778
rect 26850 3726 26852 3778
rect 26796 3714 26852 3726
rect 27244 3780 27300 3790
rect 25340 3424 25396 3500
rect 26012 3556 26068 3566
rect 26012 3462 26068 3500
rect 26684 3556 26740 3566
rect 26684 3462 26740 3500
rect 27244 1876 27300 3724
rect 27356 3778 27412 4284
rect 27356 3726 27358 3778
rect 27410 3726 27412 3778
rect 27356 3556 27412 3726
rect 27692 4338 27748 4844
rect 29184 4732 29448 4742
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29184 4666 29448 4676
rect 27804 4564 27860 4574
rect 27804 4470 27860 4508
rect 28476 4564 28532 4574
rect 28476 4470 28532 4508
rect 29148 4564 29204 4574
rect 29148 4470 29204 4508
rect 29820 4564 29876 4956
rect 29260 4452 29316 4462
rect 27692 4286 27694 4338
rect 27746 4286 27748 4338
rect 27692 4116 27748 4286
rect 27692 3668 27748 4060
rect 28364 4338 28420 4350
rect 28364 4286 28366 4338
rect 28418 4286 28420 4338
rect 27692 3602 27748 3612
rect 28028 3668 28084 3678
rect 28028 3574 28084 3612
rect 28364 3668 28420 4286
rect 28364 3602 28420 3612
rect 29036 4340 29092 4350
rect 27468 3556 27524 3566
rect 27356 3500 27468 3556
rect 27468 3424 27524 3500
rect 28140 3556 28196 3566
rect 28140 3462 28196 3500
rect 29036 3556 29092 4284
rect 29260 3778 29316 4396
rect 29708 4340 29764 4350
rect 29708 4246 29764 4284
rect 29260 3726 29262 3778
rect 29314 3726 29316 3778
rect 29260 3714 29316 3726
rect 29820 3780 29876 4508
rect 30268 4452 30324 5070
rect 30380 5012 30436 5294
rect 30380 4946 30436 4956
rect 30492 5682 30548 5694
rect 30492 5630 30494 5682
rect 30546 5630 30548 5682
rect 30492 5124 30548 5630
rect 31052 5236 31108 6414
rect 31388 6130 31444 6636
rect 31388 6078 31390 6130
rect 31442 6078 31444 6130
rect 31388 6066 31444 6078
rect 31500 6466 31556 6478
rect 31500 6414 31502 6466
rect 31554 6414 31556 6466
rect 30940 5180 31220 5236
rect 30940 5124 30996 5180
rect 30492 5122 30996 5124
rect 30492 5070 30942 5122
rect 30994 5070 30996 5122
rect 30492 5068 30996 5070
rect 30380 4452 30436 4462
rect 30492 4452 30548 5068
rect 30940 5058 30996 5068
rect 30268 4450 30548 4452
rect 30268 4398 30382 4450
rect 30434 4398 30494 4450
rect 30546 4398 30548 4450
rect 30268 4396 30548 4398
rect 30380 4386 30436 4396
rect 30492 4386 30548 4396
rect 31052 5012 31108 5022
rect 31052 4450 31108 4956
rect 31164 4900 31220 5180
rect 31500 5012 31556 6414
rect 31836 6130 31892 6636
rect 31836 6078 31838 6130
rect 31890 6078 31892 6130
rect 31836 5124 31892 6078
rect 31948 6466 32004 6478
rect 31948 6414 31950 6466
rect 32002 6414 32004 6466
rect 31948 5796 32004 6414
rect 38508 6300 38772 6310
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38508 6234 38772 6244
rect 32284 5796 32340 5806
rect 32732 5796 32788 5806
rect 31948 5794 32788 5796
rect 31948 5742 32286 5794
rect 32338 5742 32734 5794
rect 32786 5742 32788 5794
rect 31948 5740 32788 5742
rect 31836 5058 31892 5068
rect 31500 4946 31556 4956
rect 31612 5010 31668 5022
rect 31612 4958 31614 5010
rect 31666 4958 31668 5010
rect 31164 4564 31220 4844
rect 31612 4900 31668 4958
rect 31612 4834 31668 4844
rect 31724 5012 31780 5022
rect 31164 4562 31444 4564
rect 31164 4510 31166 4562
rect 31218 4510 31444 4562
rect 31164 4508 31444 4510
rect 31164 4498 31220 4508
rect 31052 4398 31054 4450
rect 31106 4398 31108 4450
rect 31052 4386 31108 4398
rect 29932 3780 29988 3790
rect 29820 3724 29932 3780
rect 29036 3490 29092 3500
rect 29372 3668 29428 3678
rect 29932 3648 29988 3724
rect 30604 3780 30660 3790
rect 30604 3686 30660 3724
rect 31388 3778 31444 4508
rect 31724 4450 31780 4956
rect 31836 4900 31892 4910
rect 31836 4562 31892 4844
rect 32172 4900 32228 4910
rect 32172 4806 32228 4844
rect 31836 4510 31838 4562
rect 31890 4510 31892 4562
rect 31836 4498 31892 4510
rect 31724 4398 31726 4450
rect 31778 4398 31780 4450
rect 31724 4340 31780 4398
rect 32284 4340 32340 5740
rect 32732 5730 32788 5740
rect 33516 5794 33572 5806
rect 33516 5742 33518 5794
rect 33570 5742 33572 5794
rect 33516 5012 33572 5742
rect 33846 5516 34110 5526
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 33846 5450 34110 5460
rect 33516 4918 33572 4956
rect 34412 5012 34468 5022
rect 32620 4900 32676 4910
rect 32396 4340 32452 4350
rect 31724 4284 32004 4340
rect 31388 3726 31390 3778
rect 31442 3726 31444 3778
rect 29372 3554 29428 3612
rect 29372 3502 29374 3554
rect 29426 3502 29428 3554
rect 29372 3490 29428 3502
rect 30044 3556 30100 3566
rect 30044 3462 30100 3500
rect 30716 3556 30772 3566
rect 30716 3462 30772 3500
rect 31276 3556 31332 3566
rect 31388 3556 31444 3726
rect 31276 3554 31444 3556
rect 31276 3502 31278 3554
rect 31330 3502 31444 3554
rect 31276 3500 31444 3502
rect 31276 3490 31332 3500
rect 31388 3444 31444 3500
rect 31948 3556 32004 4284
rect 31948 3462 32004 3500
rect 32284 4284 32396 4340
rect 31388 3378 31444 3388
rect 32060 3444 32116 3454
rect 32284 3444 32340 4284
rect 32396 4208 32452 4284
rect 32620 4228 32676 4844
rect 33068 4900 33124 4910
rect 33068 4340 33124 4844
rect 33964 4900 34020 4910
rect 33964 4806 34020 4844
rect 34412 4898 34468 4956
rect 34412 4846 34414 4898
rect 34466 4846 34468 4898
rect 33068 4274 33124 4284
rect 32620 4162 32676 4172
rect 33516 4228 33572 4238
rect 33516 4134 33572 4172
rect 33964 4228 34020 4238
rect 33964 4134 34020 4172
rect 34412 4228 34468 4846
rect 34860 4900 34916 4910
rect 34860 4562 34916 4844
rect 34860 4510 34862 4562
rect 34914 4510 34916 4562
rect 34860 4498 34916 4510
rect 35308 4900 35364 4910
rect 34860 4228 34916 4238
rect 34412 4226 34580 4228
rect 34412 4174 34414 4226
rect 34466 4174 34580 4226
rect 34412 4172 34580 4174
rect 34412 4162 34468 4172
rect 32116 3388 32340 3444
rect 32060 3312 32116 3388
rect 29184 3164 29448 3174
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29184 3098 29448 3108
rect 27244 1820 27412 1876
rect 27356 800 27412 1820
rect 32284 800 32340 3388
rect 32508 4114 32564 4126
rect 32508 4062 32510 4114
rect 32562 4062 32564 4114
rect 32508 3444 32564 4062
rect 33846 3948 34110 3958
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 33846 3882 34110 3892
rect 34412 3668 34468 3678
rect 34412 3574 34468 3612
rect 32508 3378 32564 3388
rect 33180 3444 33236 3454
rect 33292 3444 33348 3454
rect 33180 3442 33292 3444
rect 33180 3390 33182 3442
rect 33234 3390 33292 3442
rect 33180 3388 33292 3390
rect 33180 3378 33236 3388
rect 33292 3350 33348 3388
rect 33852 3444 33908 3454
rect 33964 3444 34020 3454
rect 33852 3442 33964 3444
rect 33852 3390 33854 3442
rect 33906 3390 33964 3442
rect 33852 3388 33964 3390
rect 33852 3378 33908 3388
rect 33964 3350 34020 3388
rect 34524 3444 34580 4172
rect 34860 3666 34916 4172
rect 34860 3614 34862 3666
rect 34914 3614 34916 3666
rect 34860 3602 34916 3614
rect 35308 3666 35364 4844
rect 38508 4732 38772 4742
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38508 4666 38772 4676
rect 35308 3614 35310 3666
rect 35362 3614 35364 3666
rect 35308 3602 35364 3614
rect 34524 3378 34580 3388
rect 35756 3444 35812 3454
rect 35756 3350 35812 3388
rect 37212 3444 37268 3454
rect 37212 800 37268 3388
rect 38508 3164 38772 3174
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38508 3098 38772 3108
rect 22764 700 23492 756
rect 27328 0 27440 800
rect 32256 0 32368 800
rect 37184 0 37296 800
<< via2 >>
rect 5874 36874 5930 36876
rect 5874 36822 5876 36874
rect 5876 36822 5928 36874
rect 5928 36822 5930 36874
rect 5874 36820 5930 36822
rect 5978 36874 6034 36876
rect 5978 36822 5980 36874
rect 5980 36822 6032 36874
rect 6032 36822 6034 36874
rect 5978 36820 6034 36822
rect 6082 36874 6138 36876
rect 6082 36822 6084 36874
rect 6084 36822 6136 36874
rect 6136 36822 6138 36874
rect 6082 36820 6138 36822
rect 15198 36874 15254 36876
rect 15198 36822 15200 36874
rect 15200 36822 15252 36874
rect 15252 36822 15254 36874
rect 15198 36820 15254 36822
rect 15302 36874 15358 36876
rect 15302 36822 15304 36874
rect 15304 36822 15356 36874
rect 15356 36822 15358 36874
rect 15302 36820 15358 36822
rect 15406 36874 15462 36876
rect 15406 36822 15408 36874
rect 15408 36822 15460 36874
rect 15460 36822 15462 36874
rect 15406 36820 15462 36822
rect 24522 36874 24578 36876
rect 24522 36822 24524 36874
rect 24524 36822 24576 36874
rect 24576 36822 24578 36874
rect 24522 36820 24578 36822
rect 24626 36874 24682 36876
rect 24626 36822 24628 36874
rect 24628 36822 24680 36874
rect 24680 36822 24682 36874
rect 24626 36820 24682 36822
rect 24730 36874 24786 36876
rect 24730 36822 24732 36874
rect 24732 36822 24784 36874
rect 24784 36822 24786 36874
rect 24730 36820 24786 36822
rect 33846 36874 33902 36876
rect 33846 36822 33848 36874
rect 33848 36822 33900 36874
rect 33900 36822 33902 36874
rect 33846 36820 33902 36822
rect 33950 36874 34006 36876
rect 33950 36822 33952 36874
rect 33952 36822 34004 36874
rect 34004 36822 34006 36874
rect 33950 36820 34006 36822
rect 34054 36874 34110 36876
rect 34054 36822 34056 36874
rect 34056 36822 34108 36874
rect 34108 36822 34110 36874
rect 34054 36820 34110 36822
rect 10536 36090 10592 36092
rect 10536 36038 10538 36090
rect 10538 36038 10590 36090
rect 10590 36038 10592 36090
rect 10536 36036 10592 36038
rect 10640 36090 10696 36092
rect 10640 36038 10642 36090
rect 10642 36038 10694 36090
rect 10694 36038 10696 36090
rect 10640 36036 10696 36038
rect 10744 36090 10800 36092
rect 10744 36038 10746 36090
rect 10746 36038 10798 36090
rect 10798 36038 10800 36090
rect 10744 36036 10800 36038
rect 19860 36090 19916 36092
rect 19860 36038 19862 36090
rect 19862 36038 19914 36090
rect 19914 36038 19916 36090
rect 19860 36036 19916 36038
rect 19964 36090 20020 36092
rect 19964 36038 19966 36090
rect 19966 36038 20018 36090
rect 20018 36038 20020 36090
rect 19964 36036 20020 36038
rect 20068 36090 20124 36092
rect 20068 36038 20070 36090
rect 20070 36038 20122 36090
rect 20122 36038 20124 36090
rect 20068 36036 20124 36038
rect 29184 36090 29240 36092
rect 29184 36038 29186 36090
rect 29186 36038 29238 36090
rect 29238 36038 29240 36090
rect 29184 36036 29240 36038
rect 29288 36090 29344 36092
rect 29288 36038 29290 36090
rect 29290 36038 29342 36090
rect 29342 36038 29344 36090
rect 29288 36036 29344 36038
rect 29392 36090 29448 36092
rect 29392 36038 29394 36090
rect 29394 36038 29446 36090
rect 29446 36038 29448 36090
rect 29392 36036 29448 36038
rect 38508 36090 38564 36092
rect 38508 36038 38510 36090
rect 38510 36038 38562 36090
rect 38562 36038 38564 36090
rect 38508 36036 38564 36038
rect 38612 36090 38668 36092
rect 38612 36038 38614 36090
rect 38614 36038 38666 36090
rect 38666 36038 38668 36090
rect 38612 36036 38668 36038
rect 38716 36090 38772 36092
rect 38716 36038 38718 36090
rect 38718 36038 38770 36090
rect 38770 36038 38772 36090
rect 38716 36036 38772 36038
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 10536 34522 10592 34524
rect 10536 34470 10538 34522
rect 10538 34470 10590 34522
rect 10590 34470 10592 34522
rect 10536 34468 10592 34470
rect 10640 34522 10696 34524
rect 10640 34470 10642 34522
rect 10642 34470 10694 34522
rect 10694 34470 10696 34522
rect 10640 34468 10696 34470
rect 10744 34522 10800 34524
rect 10744 34470 10746 34522
rect 10746 34470 10798 34522
rect 10798 34470 10800 34522
rect 10744 34468 10800 34470
rect 19860 34522 19916 34524
rect 19860 34470 19862 34522
rect 19862 34470 19914 34522
rect 19914 34470 19916 34522
rect 19860 34468 19916 34470
rect 19964 34522 20020 34524
rect 19964 34470 19966 34522
rect 19966 34470 20018 34522
rect 20018 34470 20020 34522
rect 19964 34468 20020 34470
rect 20068 34522 20124 34524
rect 20068 34470 20070 34522
rect 20070 34470 20122 34522
rect 20122 34470 20124 34522
rect 20068 34468 20124 34470
rect 29184 34522 29240 34524
rect 29184 34470 29186 34522
rect 29186 34470 29238 34522
rect 29238 34470 29240 34522
rect 29184 34468 29240 34470
rect 29288 34522 29344 34524
rect 29288 34470 29290 34522
rect 29290 34470 29342 34522
rect 29342 34470 29344 34522
rect 29288 34468 29344 34470
rect 29392 34522 29448 34524
rect 29392 34470 29394 34522
rect 29394 34470 29446 34522
rect 29446 34470 29448 34522
rect 29392 34468 29448 34470
rect 38508 34522 38564 34524
rect 38508 34470 38510 34522
rect 38510 34470 38562 34522
rect 38562 34470 38564 34522
rect 38508 34468 38564 34470
rect 38612 34522 38668 34524
rect 38612 34470 38614 34522
rect 38614 34470 38666 34522
rect 38666 34470 38668 34522
rect 38612 34468 38668 34470
rect 38716 34522 38772 34524
rect 38716 34470 38718 34522
rect 38718 34470 38770 34522
rect 38770 34470 38772 34522
rect 38716 34468 38772 34470
rect 5874 33738 5930 33740
rect 5874 33686 5876 33738
rect 5876 33686 5928 33738
rect 5928 33686 5930 33738
rect 5874 33684 5930 33686
rect 5978 33738 6034 33740
rect 5978 33686 5980 33738
rect 5980 33686 6032 33738
rect 6032 33686 6034 33738
rect 5978 33684 6034 33686
rect 6082 33738 6138 33740
rect 6082 33686 6084 33738
rect 6084 33686 6136 33738
rect 6136 33686 6138 33738
rect 6082 33684 6138 33686
rect 15198 33738 15254 33740
rect 15198 33686 15200 33738
rect 15200 33686 15252 33738
rect 15252 33686 15254 33738
rect 15198 33684 15254 33686
rect 15302 33738 15358 33740
rect 15302 33686 15304 33738
rect 15304 33686 15356 33738
rect 15356 33686 15358 33738
rect 15302 33684 15358 33686
rect 15406 33738 15462 33740
rect 15406 33686 15408 33738
rect 15408 33686 15460 33738
rect 15460 33686 15462 33738
rect 15406 33684 15462 33686
rect 24522 33738 24578 33740
rect 24522 33686 24524 33738
rect 24524 33686 24576 33738
rect 24576 33686 24578 33738
rect 24522 33684 24578 33686
rect 24626 33738 24682 33740
rect 24626 33686 24628 33738
rect 24628 33686 24680 33738
rect 24680 33686 24682 33738
rect 24626 33684 24682 33686
rect 24730 33738 24786 33740
rect 24730 33686 24732 33738
rect 24732 33686 24784 33738
rect 24784 33686 24786 33738
rect 24730 33684 24786 33686
rect 33846 33738 33902 33740
rect 33846 33686 33848 33738
rect 33848 33686 33900 33738
rect 33900 33686 33902 33738
rect 33846 33684 33902 33686
rect 33950 33738 34006 33740
rect 33950 33686 33952 33738
rect 33952 33686 34004 33738
rect 34004 33686 34006 33738
rect 33950 33684 34006 33686
rect 34054 33738 34110 33740
rect 34054 33686 34056 33738
rect 34056 33686 34108 33738
rect 34108 33686 34110 33738
rect 34054 33684 34110 33686
rect 10536 32954 10592 32956
rect 10536 32902 10538 32954
rect 10538 32902 10590 32954
rect 10590 32902 10592 32954
rect 10536 32900 10592 32902
rect 10640 32954 10696 32956
rect 10640 32902 10642 32954
rect 10642 32902 10694 32954
rect 10694 32902 10696 32954
rect 10640 32900 10696 32902
rect 10744 32954 10800 32956
rect 10744 32902 10746 32954
rect 10746 32902 10798 32954
rect 10798 32902 10800 32954
rect 10744 32900 10800 32902
rect 19860 32954 19916 32956
rect 19860 32902 19862 32954
rect 19862 32902 19914 32954
rect 19914 32902 19916 32954
rect 19860 32900 19916 32902
rect 19964 32954 20020 32956
rect 19964 32902 19966 32954
rect 19966 32902 20018 32954
rect 20018 32902 20020 32954
rect 19964 32900 20020 32902
rect 20068 32954 20124 32956
rect 20068 32902 20070 32954
rect 20070 32902 20122 32954
rect 20122 32902 20124 32954
rect 20068 32900 20124 32902
rect 29184 32954 29240 32956
rect 29184 32902 29186 32954
rect 29186 32902 29238 32954
rect 29238 32902 29240 32954
rect 29184 32900 29240 32902
rect 29288 32954 29344 32956
rect 29288 32902 29290 32954
rect 29290 32902 29342 32954
rect 29342 32902 29344 32954
rect 29288 32900 29344 32902
rect 29392 32954 29448 32956
rect 29392 32902 29394 32954
rect 29394 32902 29446 32954
rect 29446 32902 29448 32954
rect 29392 32900 29448 32902
rect 38508 32954 38564 32956
rect 38508 32902 38510 32954
rect 38510 32902 38562 32954
rect 38562 32902 38564 32954
rect 38508 32900 38564 32902
rect 38612 32954 38668 32956
rect 38612 32902 38614 32954
rect 38614 32902 38666 32954
rect 38666 32902 38668 32954
rect 38612 32900 38668 32902
rect 38716 32954 38772 32956
rect 38716 32902 38718 32954
rect 38718 32902 38770 32954
rect 38770 32902 38772 32954
rect 38716 32900 38772 32902
rect 5874 32170 5930 32172
rect 5874 32118 5876 32170
rect 5876 32118 5928 32170
rect 5928 32118 5930 32170
rect 5874 32116 5930 32118
rect 5978 32170 6034 32172
rect 5978 32118 5980 32170
rect 5980 32118 6032 32170
rect 6032 32118 6034 32170
rect 5978 32116 6034 32118
rect 6082 32170 6138 32172
rect 6082 32118 6084 32170
rect 6084 32118 6136 32170
rect 6136 32118 6138 32170
rect 6082 32116 6138 32118
rect 15198 32170 15254 32172
rect 15198 32118 15200 32170
rect 15200 32118 15252 32170
rect 15252 32118 15254 32170
rect 15198 32116 15254 32118
rect 15302 32170 15358 32172
rect 15302 32118 15304 32170
rect 15304 32118 15356 32170
rect 15356 32118 15358 32170
rect 15302 32116 15358 32118
rect 15406 32170 15462 32172
rect 15406 32118 15408 32170
rect 15408 32118 15460 32170
rect 15460 32118 15462 32170
rect 15406 32116 15462 32118
rect 24522 32170 24578 32172
rect 24522 32118 24524 32170
rect 24524 32118 24576 32170
rect 24576 32118 24578 32170
rect 24522 32116 24578 32118
rect 24626 32170 24682 32172
rect 24626 32118 24628 32170
rect 24628 32118 24680 32170
rect 24680 32118 24682 32170
rect 24626 32116 24682 32118
rect 24730 32170 24786 32172
rect 24730 32118 24732 32170
rect 24732 32118 24784 32170
rect 24784 32118 24786 32170
rect 24730 32116 24786 32118
rect 33846 32170 33902 32172
rect 33846 32118 33848 32170
rect 33848 32118 33900 32170
rect 33900 32118 33902 32170
rect 33846 32116 33902 32118
rect 33950 32170 34006 32172
rect 33950 32118 33952 32170
rect 33952 32118 34004 32170
rect 34004 32118 34006 32170
rect 33950 32116 34006 32118
rect 34054 32170 34110 32172
rect 34054 32118 34056 32170
rect 34056 32118 34108 32170
rect 34108 32118 34110 32170
rect 34054 32116 34110 32118
rect 10536 31386 10592 31388
rect 10536 31334 10538 31386
rect 10538 31334 10590 31386
rect 10590 31334 10592 31386
rect 10536 31332 10592 31334
rect 10640 31386 10696 31388
rect 10640 31334 10642 31386
rect 10642 31334 10694 31386
rect 10694 31334 10696 31386
rect 10640 31332 10696 31334
rect 10744 31386 10800 31388
rect 10744 31334 10746 31386
rect 10746 31334 10798 31386
rect 10798 31334 10800 31386
rect 10744 31332 10800 31334
rect 19860 31386 19916 31388
rect 19860 31334 19862 31386
rect 19862 31334 19914 31386
rect 19914 31334 19916 31386
rect 19860 31332 19916 31334
rect 19964 31386 20020 31388
rect 19964 31334 19966 31386
rect 19966 31334 20018 31386
rect 20018 31334 20020 31386
rect 19964 31332 20020 31334
rect 20068 31386 20124 31388
rect 20068 31334 20070 31386
rect 20070 31334 20122 31386
rect 20122 31334 20124 31386
rect 20068 31332 20124 31334
rect 29184 31386 29240 31388
rect 29184 31334 29186 31386
rect 29186 31334 29238 31386
rect 29238 31334 29240 31386
rect 29184 31332 29240 31334
rect 29288 31386 29344 31388
rect 29288 31334 29290 31386
rect 29290 31334 29342 31386
rect 29342 31334 29344 31386
rect 29288 31332 29344 31334
rect 29392 31386 29448 31388
rect 29392 31334 29394 31386
rect 29394 31334 29446 31386
rect 29446 31334 29448 31386
rect 29392 31332 29448 31334
rect 38508 31386 38564 31388
rect 38508 31334 38510 31386
rect 38510 31334 38562 31386
rect 38562 31334 38564 31386
rect 38508 31332 38564 31334
rect 38612 31386 38668 31388
rect 38612 31334 38614 31386
rect 38614 31334 38666 31386
rect 38666 31334 38668 31386
rect 38612 31332 38668 31334
rect 38716 31386 38772 31388
rect 38716 31334 38718 31386
rect 38718 31334 38770 31386
rect 38770 31334 38772 31386
rect 38716 31332 38772 31334
rect 5874 30602 5930 30604
rect 5874 30550 5876 30602
rect 5876 30550 5928 30602
rect 5928 30550 5930 30602
rect 5874 30548 5930 30550
rect 5978 30602 6034 30604
rect 5978 30550 5980 30602
rect 5980 30550 6032 30602
rect 6032 30550 6034 30602
rect 5978 30548 6034 30550
rect 6082 30602 6138 30604
rect 6082 30550 6084 30602
rect 6084 30550 6136 30602
rect 6136 30550 6138 30602
rect 6082 30548 6138 30550
rect 15198 30602 15254 30604
rect 15198 30550 15200 30602
rect 15200 30550 15252 30602
rect 15252 30550 15254 30602
rect 15198 30548 15254 30550
rect 15302 30602 15358 30604
rect 15302 30550 15304 30602
rect 15304 30550 15356 30602
rect 15356 30550 15358 30602
rect 15302 30548 15358 30550
rect 15406 30602 15462 30604
rect 15406 30550 15408 30602
rect 15408 30550 15460 30602
rect 15460 30550 15462 30602
rect 15406 30548 15462 30550
rect 24522 30602 24578 30604
rect 24522 30550 24524 30602
rect 24524 30550 24576 30602
rect 24576 30550 24578 30602
rect 24522 30548 24578 30550
rect 24626 30602 24682 30604
rect 24626 30550 24628 30602
rect 24628 30550 24680 30602
rect 24680 30550 24682 30602
rect 24626 30548 24682 30550
rect 24730 30602 24786 30604
rect 24730 30550 24732 30602
rect 24732 30550 24784 30602
rect 24784 30550 24786 30602
rect 24730 30548 24786 30550
rect 33846 30602 33902 30604
rect 33846 30550 33848 30602
rect 33848 30550 33900 30602
rect 33900 30550 33902 30602
rect 33846 30548 33902 30550
rect 33950 30602 34006 30604
rect 33950 30550 33952 30602
rect 33952 30550 34004 30602
rect 34004 30550 34006 30602
rect 33950 30548 34006 30550
rect 34054 30602 34110 30604
rect 34054 30550 34056 30602
rect 34056 30550 34108 30602
rect 34108 30550 34110 30602
rect 34054 30548 34110 30550
rect 10536 29818 10592 29820
rect 10536 29766 10538 29818
rect 10538 29766 10590 29818
rect 10590 29766 10592 29818
rect 10536 29764 10592 29766
rect 10640 29818 10696 29820
rect 10640 29766 10642 29818
rect 10642 29766 10694 29818
rect 10694 29766 10696 29818
rect 10640 29764 10696 29766
rect 10744 29818 10800 29820
rect 10744 29766 10746 29818
rect 10746 29766 10798 29818
rect 10798 29766 10800 29818
rect 10744 29764 10800 29766
rect 19860 29818 19916 29820
rect 19860 29766 19862 29818
rect 19862 29766 19914 29818
rect 19914 29766 19916 29818
rect 19860 29764 19916 29766
rect 19964 29818 20020 29820
rect 19964 29766 19966 29818
rect 19966 29766 20018 29818
rect 20018 29766 20020 29818
rect 19964 29764 20020 29766
rect 20068 29818 20124 29820
rect 20068 29766 20070 29818
rect 20070 29766 20122 29818
rect 20122 29766 20124 29818
rect 20068 29764 20124 29766
rect 29184 29818 29240 29820
rect 29184 29766 29186 29818
rect 29186 29766 29238 29818
rect 29238 29766 29240 29818
rect 29184 29764 29240 29766
rect 29288 29818 29344 29820
rect 29288 29766 29290 29818
rect 29290 29766 29342 29818
rect 29342 29766 29344 29818
rect 29288 29764 29344 29766
rect 29392 29818 29448 29820
rect 29392 29766 29394 29818
rect 29394 29766 29446 29818
rect 29446 29766 29448 29818
rect 29392 29764 29448 29766
rect 38508 29818 38564 29820
rect 38508 29766 38510 29818
rect 38510 29766 38562 29818
rect 38562 29766 38564 29818
rect 38508 29764 38564 29766
rect 38612 29818 38668 29820
rect 38612 29766 38614 29818
rect 38614 29766 38666 29818
rect 38666 29766 38668 29818
rect 38612 29764 38668 29766
rect 38716 29818 38772 29820
rect 38716 29766 38718 29818
rect 38718 29766 38770 29818
rect 38770 29766 38772 29818
rect 38716 29764 38772 29766
rect 5874 29034 5930 29036
rect 5874 28982 5876 29034
rect 5876 28982 5928 29034
rect 5928 28982 5930 29034
rect 5874 28980 5930 28982
rect 5978 29034 6034 29036
rect 5978 28982 5980 29034
rect 5980 28982 6032 29034
rect 6032 28982 6034 29034
rect 5978 28980 6034 28982
rect 6082 29034 6138 29036
rect 6082 28982 6084 29034
rect 6084 28982 6136 29034
rect 6136 28982 6138 29034
rect 6082 28980 6138 28982
rect 15198 29034 15254 29036
rect 15198 28982 15200 29034
rect 15200 28982 15252 29034
rect 15252 28982 15254 29034
rect 15198 28980 15254 28982
rect 15302 29034 15358 29036
rect 15302 28982 15304 29034
rect 15304 28982 15356 29034
rect 15356 28982 15358 29034
rect 15302 28980 15358 28982
rect 15406 29034 15462 29036
rect 15406 28982 15408 29034
rect 15408 28982 15460 29034
rect 15460 28982 15462 29034
rect 15406 28980 15462 28982
rect 24522 29034 24578 29036
rect 24522 28982 24524 29034
rect 24524 28982 24576 29034
rect 24576 28982 24578 29034
rect 24522 28980 24578 28982
rect 24626 29034 24682 29036
rect 24626 28982 24628 29034
rect 24628 28982 24680 29034
rect 24680 28982 24682 29034
rect 24626 28980 24682 28982
rect 24730 29034 24786 29036
rect 24730 28982 24732 29034
rect 24732 28982 24784 29034
rect 24784 28982 24786 29034
rect 24730 28980 24786 28982
rect 33846 29034 33902 29036
rect 33846 28982 33848 29034
rect 33848 28982 33900 29034
rect 33900 28982 33902 29034
rect 33846 28980 33902 28982
rect 33950 29034 34006 29036
rect 33950 28982 33952 29034
rect 33952 28982 34004 29034
rect 34004 28982 34006 29034
rect 33950 28980 34006 28982
rect 34054 29034 34110 29036
rect 34054 28982 34056 29034
rect 34056 28982 34108 29034
rect 34108 28982 34110 29034
rect 34054 28980 34110 28982
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 5874 27466 5930 27468
rect 5874 27414 5876 27466
rect 5876 27414 5928 27466
rect 5928 27414 5930 27466
rect 5874 27412 5930 27414
rect 5978 27466 6034 27468
rect 5978 27414 5980 27466
rect 5980 27414 6032 27466
rect 6032 27414 6034 27466
rect 5978 27412 6034 27414
rect 6082 27466 6138 27468
rect 6082 27414 6084 27466
rect 6084 27414 6136 27466
rect 6136 27414 6138 27466
rect 6082 27412 6138 27414
rect 15198 27466 15254 27468
rect 15198 27414 15200 27466
rect 15200 27414 15252 27466
rect 15252 27414 15254 27466
rect 15198 27412 15254 27414
rect 15302 27466 15358 27468
rect 15302 27414 15304 27466
rect 15304 27414 15356 27466
rect 15356 27414 15358 27466
rect 15302 27412 15358 27414
rect 15406 27466 15462 27468
rect 15406 27414 15408 27466
rect 15408 27414 15460 27466
rect 15460 27414 15462 27466
rect 15406 27412 15462 27414
rect 24522 27466 24578 27468
rect 24522 27414 24524 27466
rect 24524 27414 24576 27466
rect 24576 27414 24578 27466
rect 24522 27412 24578 27414
rect 24626 27466 24682 27468
rect 24626 27414 24628 27466
rect 24628 27414 24680 27466
rect 24680 27414 24682 27466
rect 24626 27412 24682 27414
rect 24730 27466 24786 27468
rect 24730 27414 24732 27466
rect 24732 27414 24784 27466
rect 24784 27414 24786 27466
rect 24730 27412 24786 27414
rect 33846 27466 33902 27468
rect 33846 27414 33848 27466
rect 33848 27414 33900 27466
rect 33900 27414 33902 27466
rect 33846 27412 33902 27414
rect 33950 27466 34006 27468
rect 33950 27414 33952 27466
rect 33952 27414 34004 27466
rect 34004 27414 34006 27466
rect 33950 27412 34006 27414
rect 34054 27466 34110 27468
rect 34054 27414 34056 27466
rect 34056 27414 34108 27466
rect 34108 27414 34110 27466
rect 34054 27412 34110 27414
rect 10536 26682 10592 26684
rect 10536 26630 10538 26682
rect 10538 26630 10590 26682
rect 10590 26630 10592 26682
rect 10536 26628 10592 26630
rect 10640 26682 10696 26684
rect 10640 26630 10642 26682
rect 10642 26630 10694 26682
rect 10694 26630 10696 26682
rect 10640 26628 10696 26630
rect 10744 26682 10800 26684
rect 10744 26630 10746 26682
rect 10746 26630 10798 26682
rect 10798 26630 10800 26682
rect 10744 26628 10800 26630
rect 19860 26682 19916 26684
rect 19860 26630 19862 26682
rect 19862 26630 19914 26682
rect 19914 26630 19916 26682
rect 19860 26628 19916 26630
rect 19964 26682 20020 26684
rect 19964 26630 19966 26682
rect 19966 26630 20018 26682
rect 20018 26630 20020 26682
rect 19964 26628 20020 26630
rect 20068 26682 20124 26684
rect 20068 26630 20070 26682
rect 20070 26630 20122 26682
rect 20122 26630 20124 26682
rect 20068 26628 20124 26630
rect 29184 26682 29240 26684
rect 29184 26630 29186 26682
rect 29186 26630 29238 26682
rect 29238 26630 29240 26682
rect 29184 26628 29240 26630
rect 29288 26682 29344 26684
rect 29288 26630 29290 26682
rect 29290 26630 29342 26682
rect 29342 26630 29344 26682
rect 29288 26628 29344 26630
rect 29392 26682 29448 26684
rect 29392 26630 29394 26682
rect 29394 26630 29446 26682
rect 29446 26630 29448 26682
rect 29392 26628 29448 26630
rect 38508 26682 38564 26684
rect 38508 26630 38510 26682
rect 38510 26630 38562 26682
rect 38562 26630 38564 26682
rect 38508 26628 38564 26630
rect 38612 26682 38668 26684
rect 38612 26630 38614 26682
rect 38614 26630 38666 26682
rect 38666 26630 38668 26682
rect 38612 26628 38668 26630
rect 38716 26682 38772 26684
rect 38716 26630 38718 26682
rect 38718 26630 38770 26682
rect 38770 26630 38772 26682
rect 38716 26628 38772 26630
rect 5874 25898 5930 25900
rect 5874 25846 5876 25898
rect 5876 25846 5928 25898
rect 5928 25846 5930 25898
rect 5874 25844 5930 25846
rect 5978 25898 6034 25900
rect 5978 25846 5980 25898
rect 5980 25846 6032 25898
rect 6032 25846 6034 25898
rect 5978 25844 6034 25846
rect 6082 25898 6138 25900
rect 6082 25846 6084 25898
rect 6084 25846 6136 25898
rect 6136 25846 6138 25898
rect 6082 25844 6138 25846
rect 15198 25898 15254 25900
rect 15198 25846 15200 25898
rect 15200 25846 15252 25898
rect 15252 25846 15254 25898
rect 15198 25844 15254 25846
rect 15302 25898 15358 25900
rect 15302 25846 15304 25898
rect 15304 25846 15356 25898
rect 15356 25846 15358 25898
rect 15302 25844 15358 25846
rect 15406 25898 15462 25900
rect 15406 25846 15408 25898
rect 15408 25846 15460 25898
rect 15460 25846 15462 25898
rect 15406 25844 15462 25846
rect 24522 25898 24578 25900
rect 24522 25846 24524 25898
rect 24524 25846 24576 25898
rect 24576 25846 24578 25898
rect 24522 25844 24578 25846
rect 24626 25898 24682 25900
rect 24626 25846 24628 25898
rect 24628 25846 24680 25898
rect 24680 25846 24682 25898
rect 24626 25844 24682 25846
rect 24730 25898 24786 25900
rect 24730 25846 24732 25898
rect 24732 25846 24784 25898
rect 24784 25846 24786 25898
rect 24730 25844 24786 25846
rect 33846 25898 33902 25900
rect 33846 25846 33848 25898
rect 33848 25846 33900 25898
rect 33900 25846 33902 25898
rect 33846 25844 33902 25846
rect 33950 25898 34006 25900
rect 33950 25846 33952 25898
rect 33952 25846 34004 25898
rect 34004 25846 34006 25898
rect 33950 25844 34006 25846
rect 34054 25898 34110 25900
rect 34054 25846 34056 25898
rect 34056 25846 34108 25898
rect 34108 25846 34110 25898
rect 34054 25844 34110 25846
rect 10536 25114 10592 25116
rect 10536 25062 10538 25114
rect 10538 25062 10590 25114
rect 10590 25062 10592 25114
rect 10536 25060 10592 25062
rect 10640 25114 10696 25116
rect 10640 25062 10642 25114
rect 10642 25062 10694 25114
rect 10694 25062 10696 25114
rect 10640 25060 10696 25062
rect 10744 25114 10800 25116
rect 10744 25062 10746 25114
rect 10746 25062 10798 25114
rect 10798 25062 10800 25114
rect 10744 25060 10800 25062
rect 19860 25114 19916 25116
rect 19860 25062 19862 25114
rect 19862 25062 19914 25114
rect 19914 25062 19916 25114
rect 19860 25060 19916 25062
rect 19964 25114 20020 25116
rect 19964 25062 19966 25114
rect 19966 25062 20018 25114
rect 20018 25062 20020 25114
rect 19964 25060 20020 25062
rect 20068 25114 20124 25116
rect 20068 25062 20070 25114
rect 20070 25062 20122 25114
rect 20122 25062 20124 25114
rect 20068 25060 20124 25062
rect 29184 25114 29240 25116
rect 29184 25062 29186 25114
rect 29186 25062 29238 25114
rect 29238 25062 29240 25114
rect 29184 25060 29240 25062
rect 29288 25114 29344 25116
rect 29288 25062 29290 25114
rect 29290 25062 29342 25114
rect 29342 25062 29344 25114
rect 29288 25060 29344 25062
rect 29392 25114 29448 25116
rect 29392 25062 29394 25114
rect 29394 25062 29446 25114
rect 29446 25062 29448 25114
rect 29392 25060 29448 25062
rect 38508 25114 38564 25116
rect 38508 25062 38510 25114
rect 38510 25062 38562 25114
rect 38562 25062 38564 25114
rect 38508 25060 38564 25062
rect 38612 25114 38668 25116
rect 38612 25062 38614 25114
rect 38614 25062 38666 25114
rect 38666 25062 38668 25114
rect 38612 25060 38668 25062
rect 38716 25114 38772 25116
rect 38716 25062 38718 25114
rect 38718 25062 38770 25114
rect 38770 25062 38772 25114
rect 38716 25060 38772 25062
rect 5874 24330 5930 24332
rect 5874 24278 5876 24330
rect 5876 24278 5928 24330
rect 5928 24278 5930 24330
rect 5874 24276 5930 24278
rect 5978 24330 6034 24332
rect 5978 24278 5980 24330
rect 5980 24278 6032 24330
rect 6032 24278 6034 24330
rect 5978 24276 6034 24278
rect 6082 24330 6138 24332
rect 6082 24278 6084 24330
rect 6084 24278 6136 24330
rect 6136 24278 6138 24330
rect 6082 24276 6138 24278
rect 15198 24330 15254 24332
rect 15198 24278 15200 24330
rect 15200 24278 15252 24330
rect 15252 24278 15254 24330
rect 15198 24276 15254 24278
rect 15302 24330 15358 24332
rect 15302 24278 15304 24330
rect 15304 24278 15356 24330
rect 15356 24278 15358 24330
rect 15302 24276 15358 24278
rect 15406 24330 15462 24332
rect 15406 24278 15408 24330
rect 15408 24278 15460 24330
rect 15460 24278 15462 24330
rect 15406 24276 15462 24278
rect 24522 24330 24578 24332
rect 24522 24278 24524 24330
rect 24524 24278 24576 24330
rect 24576 24278 24578 24330
rect 24522 24276 24578 24278
rect 24626 24330 24682 24332
rect 24626 24278 24628 24330
rect 24628 24278 24680 24330
rect 24680 24278 24682 24330
rect 24626 24276 24682 24278
rect 24730 24330 24786 24332
rect 24730 24278 24732 24330
rect 24732 24278 24784 24330
rect 24784 24278 24786 24330
rect 24730 24276 24786 24278
rect 33846 24330 33902 24332
rect 33846 24278 33848 24330
rect 33848 24278 33900 24330
rect 33900 24278 33902 24330
rect 33846 24276 33902 24278
rect 33950 24330 34006 24332
rect 33950 24278 33952 24330
rect 33952 24278 34004 24330
rect 34004 24278 34006 24330
rect 33950 24276 34006 24278
rect 34054 24330 34110 24332
rect 34054 24278 34056 24330
rect 34056 24278 34108 24330
rect 34108 24278 34110 24330
rect 34054 24276 34110 24278
rect 10536 23546 10592 23548
rect 10536 23494 10538 23546
rect 10538 23494 10590 23546
rect 10590 23494 10592 23546
rect 10536 23492 10592 23494
rect 10640 23546 10696 23548
rect 10640 23494 10642 23546
rect 10642 23494 10694 23546
rect 10694 23494 10696 23546
rect 10640 23492 10696 23494
rect 10744 23546 10800 23548
rect 10744 23494 10746 23546
rect 10746 23494 10798 23546
rect 10798 23494 10800 23546
rect 10744 23492 10800 23494
rect 19860 23546 19916 23548
rect 19860 23494 19862 23546
rect 19862 23494 19914 23546
rect 19914 23494 19916 23546
rect 19860 23492 19916 23494
rect 19964 23546 20020 23548
rect 19964 23494 19966 23546
rect 19966 23494 20018 23546
rect 20018 23494 20020 23546
rect 19964 23492 20020 23494
rect 20068 23546 20124 23548
rect 20068 23494 20070 23546
rect 20070 23494 20122 23546
rect 20122 23494 20124 23546
rect 20068 23492 20124 23494
rect 29184 23546 29240 23548
rect 29184 23494 29186 23546
rect 29186 23494 29238 23546
rect 29238 23494 29240 23546
rect 29184 23492 29240 23494
rect 29288 23546 29344 23548
rect 29288 23494 29290 23546
rect 29290 23494 29342 23546
rect 29342 23494 29344 23546
rect 29288 23492 29344 23494
rect 29392 23546 29448 23548
rect 29392 23494 29394 23546
rect 29394 23494 29446 23546
rect 29446 23494 29448 23546
rect 29392 23492 29448 23494
rect 38508 23546 38564 23548
rect 38508 23494 38510 23546
rect 38510 23494 38562 23546
rect 38562 23494 38564 23546
rect 38508 23492 38564 23494
rect 38612 23546 38668 23548
rect 38612 23494 38614 23546
rect 38614 23494 38666 23546
rect 38666 23494 38668 23546
rect 38612 23492 38668 23494
rect 38716 23546 38772 23548
rect 38716 23494 38718 23546
rect 38718 23494 38770 23546
rect 38770 23494 38772 23546
rect 38716 23492 38772 23494
rect 5874 22762 5930 22764
rect 5874 22710 5876 22762
rect 5876 22710 5928 22762
rect 5928 22710 5930 22762
rect 5874 22708 5930 22710
rect 5978 22762 6034 22764
rect 5978 22710 5980 22762
rect 5980 22710 6032 22762
rect 6032 22710 6034 22762
rect 5978 22708 6034 22710
rect 6082 22762 6138 22764
rect 6082 22710 6084 22762
rect 6084 22710 6136 22762
rect 6136 22710 6138 22762
rect 6082 22708 6138 22710
rect 15198 22762 15254 22764
rect 15198 22710 15200 22762
rect 15200 22710 15252 22762
rect 15252 22710 15254 22762
rect 15198 22708 15254 22710
rect 15302 22762 15358 22764
rect 15302 22710 15304 22762
rect 15304 22710 15356 22762
rect 15356 22710 15358 22762
rect 15302 22708 15358 22710
rect 15406 22762 15462 22764
rect 15406 22710 15408 22762
rect 15408 22710 15460 22762
rect 15460 22710 15462 22762
rect 15406 22708 15462 22710
rect 24522 22762 24578 22764
rect 24522 22710 24524 22762
rect 24524 22710 24576 22762
rect 24576 22710 24578 22762
rect 24522 22708 24578 22710
rect 24626 22762 24682 22764
rect 24626 22710 24628 22762
rect 24628 22710 24680 22762
rect 24680 22710 24682 22762
rect 24626 22708 24682 22710
rect 24730 22762 24786 22764
rect 24730 22710 24732 22762
rect 24732 22710 24784 22762
rect 24784 22710 24786 22762
rect 24730 22708 24786 22710
rect 33846 22762 33902 22764
rect 33846 22710 33848 22762
rect 33848 22710 33900 22762
rect 33900 22710 33902 22762
rect 33846 22708 33902 22710
rect 33950 22762 34006 22764
rect 33950 22710 33952 22762
rect 33952 22710 34004 22762
rect 34004 22710 34006 22762
rect 33950 22708 34006 22710
rect 34054 22762 34110 22764
rect 34054 22710 34056 22762
rect 34056 22710 34108 22762
rect 34108 22710 34110 22762
rect 34054 22708 34110 22710
rect 10536 21978 10592 21980
rect 10536 21926 10538 21978
rect 10538 21926 10590 21978
rect 10590 21926 10592 21978
rect 10536 21924 10592 21926
rect 10640 21978 10696 21980
rect 10640 21926 10642 21978
rect 10642 21926 10694 21978
rect 10694 21926 10696 21978
rect 10640 21924 10696 21926
rect 10744 21978 10800 21980
rect 10744 21926 10746 21978
rect 10746 21926 10798 21978
rect 10798 21926 10800 21978
rect 10744 21924 10800 21926
rect 19860 21978 19916 21980
rect 19860 21926 19862 21978
rect 19862 21926 19914 21978
rect 19914 21926 19916 21978
rect 19860 21924 19916 21926
rect 19964 21978 20020 21980
rect 19964 21926 19966 21978
rect 19966 21926 20018 21978
rect 20018 21926 20020 21978
rect 19964 21924 20020 21926
rect 20068 21978 20124 21980
rect 20068 21926 20070 21978
rect 20070 21926 20122 21978
rect 20122 21926 20124 21978
rect 20068 21924 20124 21926
rect 29184 21978 29240 21980
rect 29184 21926 29186 21978
rect 29186 21926 29238 21978
rect 29238 21926 29240 21978
rect 29184 21924 29240 21926
rect 29288 21978 29344 21980
rect 29288 21926 29290 21978
rect 29290 21926 29342 21978
rect 29342 21926 29344 21978
rect 29288 21924 29344 21926
rect 29392 21978 29448 21980
rect 29392 21926 29394 21978
rect 29394 21926 29446 21978
rect 29446 21926 29448 21978
rect 29392 21924 29448 21926
rect 38508 21978 38564 21980
rect 38508 21926 38510 21978
rect 38510 21926 38562 21978
rect 38562 21926 38564 21978
rect 38508 21924 38564 21926
rect 38612 21978 38668 21980
rect 38612 21926 38614 21978
rect 38614 21926 38666 21978
rect 38666 21926 38668 21978
rect 38612 21924 38668 21926
rect 38716 21978 38772 21980
rect 38716 21926 38718 21978
rect 38718 21926 38770 21978
rect 38770 21926 38772 21978
rect 38716 21924 38772 21926
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 10536 20410 10592 20412
rect 10536 20358 10538 20410
rect 10538 20358 10590 20410
rect 10590 20358 10592 20410
rect 10536 20356 10592 20358
rect 10640 20410 10696 20412
rect 10640 20358 10642 20410
rect 10642 20358 10694 20410
rect 10694 20358 10696 20410
rect 10640 20356 10696 20358
rect 10744 20410 10800 20412
rect 10744 20358 10746 20410
rect 10746 20358 10798 20410
rect 10798 20358 10800 20410
rect 10744 20356 10800 20358
rect 19860 20410 19916 20412
rect 19860 20358 19862 20410
rect 19862 20358 19914 20410
rect 19914 20358 19916 20410
rect 19860 20356 19916 20358
rect 19964 20410 20020 20412
rect 19964 20358 19966 20410
rect 19966 20358 20018 20410
rect 20018 20358 20020 20410
rect 19964 20356 20020 20358
rect 20068 20410 20124 20412
rect 20068 20358 20070 20410
rect 20070 20358 20122 20410
rect 20122 20358 20124 20410
rect 20068 20356 20124 20358
rect 29184 20410 29240 20412
rect 29184 20358 29186 20410
rect 29186 20358 29238 20410
rect 29238 20358 29240 20410
rect 29184 20356 29240 20358
rect 29288 20410 29344 20412
rect 29288 20358 29290 20410
rect 29290 20358 29342 20410
rect 29342 20358 29344 20410
rect 29288 20356 29344 20358
rect 29392 20410 29448 20412
rect 29392 20358 29394 20410
rect 29394 20358 29446 20410
rect 29446 20358 29448 20410
rect 29392 20356 29448 20358
rect 38508 20410 38564 20412
rect 38508 20358 38510 20410
rect 38510 20358 38562 20410
rect 38562 20358 38564 20410
rect 38508 20356 38564 20358
rect 38612 20410 38668 20412
rect 38612 20358 38614 20410
rect 38614 20358 38666 20410
rect 38666 20358 38668 20410
rect 38612 20356 38668 20358
rect 38716 20410 38772 20412
rect 38716 20358 38718 20410
rect 38718 20358 38770 20410
rect 38770 20358 38772 20410
rect 38716 20356 38772 20358
rect 5874 19626 5930 19628
rect 5874 19574 5876 19626
rect 5876 19574 5928 19626
rect 5928 19574 5930 19626
rect 5874 19572 5930 19574
rect 5978 19626 6034 19628
rect 5978 19574 5980 19626
rect 5980 19574 6032 19626
rect 6032 19574 6034 19626
rect 5978 19572 6034 19574
rect 6082 19626 6138 19628
rect 6082 19574 6084 19626
rect 6084 19574 6136 19626
rect 6136 19574 6138 19626
rect 6082 19572 6138 19574
rect 15198 19626 15254 19628
rect 15198 19574 15200 19626
rect 15200 19574 15252 19626
rect 15252 19574 15254 19626
rect 15198 19572 15254 19574
rect 15302 19626 15358 19628
rect 15302 19574 15304 19626
rect 15304 19574 15356 19626
rect 15356 19574 15358 19626
rect 15302 19572 15358 19574
rect 15406 19626 15462 19628
rect 15406 19574 15408 19626
rect 15408 19574 15460 19626
rect 15460 19574 15462 19626
rect 15406 19572 15462 19574
rect 24522 19626 24578 19628
rect 24522 19574 24524 19626
rect 24524 19574 24576 19626
rect 24576 19574 24578 19626
rect 24522 19572 24578 19574
rect 24626 19626 24682 19628
rect 24626 19574 24628 19626
rect 24628 19574 24680 19626
rect 24680 19574 24682 19626
rect 24626 19572 24682 19574
rect 24730 19626 24786 19628
rect 24730 19574 24732 19626
rect 24732 19574 24784 19626
rect 24784 19574 24786 19626
rect 24730 19572 24786 19574
rect 33846 19626 33902 19628
rect 33846 19574 33848 19626
rect 33848 19574 33900 19626
rect 33900 19574 33902 19626
rect 33846 19572 33902 19574
rect 33950 19626 34006 19628
rect 33950 19574 33952 19626
rect 33952 19574 34004 19626
rect 34004 19574 34006 19626
rect 33950 19572 34006 19574
rect 34054 19626 34110 19628
rect 34054 19574 34056 19626
rect 34056 19574 34108 19626
rect 34108 19574 34110 19626
rect 34054 19572 34110 19574
rect 10536 18842 10592 18844
rect 10536 18790 10538 18842
rect 10538 18790 10590 18842
rect 10590 18790 10592 18842
rect 10536 18788 10592 18790
rect 10640 18842 10696 18844
rect 10640 18790 10642 18842
rect 10642 18790 10694 18842
rect 10694 18790 10696 18842
rect 10640 18788 10696 18790
rect 10744 18842 10800 18844
rect 10744 18790 10746 18842
rect 10746 18790 10798 18842
rect 10798 18790 10800 18842
rect 10744 18788 10800 18790
rect 19860 18842 19916 18844
rect 19860 18790 19862 18842
rect 19862 18790 19914 18842
rect 19914 18790 19916 18842
rect 19860 18788 19916 18790
rect 19964 18842 20020 18844
rect 19964 18790 19966 18842
rect 19966 18790 20018 18842
rect 20018 18790 20020 18842
rect 19964 18788 20020 18790
rect 20068 18842 20124 18844
rect 20068 18790 20070 18842
rect 20070 18790 20122 18842
rect 20122 18790 20124 18842
rect 20068 18788 20124 18790
rect 29184 18842 29240 18844
rect 29184 18790 29186 18842
rect 29186 18790 29238 18842
rect 29238 18790 29240 18842
rect 29184 18788 29240 18790
rect 29288 18842 29344 18844
rect 29288 18790 29290 18842
rect 29290 18790 29342 18842
rect 29342 18790 29344 18842
rect 29288 18788 29344 18790
rect 29392 18842 29448 18844
rect 29392 18790 29394 18842
rect 29394 18790 29446 18842
rect 29446 18790 29448 18842
rect 29392 18788 29448 18790
rect 38508 18842 38564 18844
rect 38508 18790 38510 18842
rect 38510 18790 38562 18842
rect 38562 18790 38564 18842
rect 38508 18788 38564 18790
rect 38612 18842 38668 18844
rect 38612 18790 38614 18842
rect 38614 18790 38666 18842
rect 38666 18790 38668 18842
rect 38612 18788 38668 18790
rect 38716 18842 38772 18844
rect 38716 18790 38718 18842
rect 38718 18790 38770 18842
rect 38770 18790 38772 18842
rect 38716 18788 38772 18790
rect 5874 18058 5930 18060
rect 5874 18006 5876 18058
rect 5876 18006 5928 18058
rect 5928 18006 5930 18058
rect 5874 18004 5930 18006
rect 5978 18058 6034 18060
rect 5978 18006 5980 18058
rect 5980 18006 6032 18058
rect 6032 18006 6034 18058
rect 5978 18004 6034 18006
rect 6082 18058 6138 18060
rect 6082 18006 6084 18058
rect 6084 18006 6136 18058
rect 6136 18006 6138 18058
rect 6082 18004 6138 18006
rect 15198 18058 15254 18060
rect 15198 18006 15200 18058
rect 15200 18006 15252 18058
rect 15252 18006 15254 18058
rect 15198 18004 15254 18006
rect 15302 18058 15358 18060
rect 15302 18006 15304 18058
rect 15304 18006 15356 18058
rect 15356 18006 15358 18058
rect 15302 18004 15358 18006
rect 15406 18058 15462 18060
rect 15406 18006 15408 18058
rect 15408 18006 15460 18058
rect 15460 18006 15462 18058
rect 15406 18004 15462 18006
rect 24522 18058 24578 18060
rect 24522 18006 24524 18058
rect 24524 18006 24576 18058
rect 24576 18006 24578 18058
rect 24522 18004 24578 18006
rect 24626 18058 24682 18060
rect 24626 18006 24628 18058
rect 24628 18006 24680 18058
rect 24680 18006 24682 18058
rect 24626 18004 24682 18006
rect 24730 18058 24786 18060
rect 24730 18006 24732 18058
rect 24732 18006 24784 18058
rect 24784 18006 24786 18058
rect 24730 18004 24786 18006
rect 33846 18058 33902 18060
rect 33846 18006 33848 18058
rect 33848 18006 33900 18058
rect 33900 18006 33902 18058
rect 33846 18004 33902 18006
rect 33950 18058 34006 18060
rect 33950 18006 33952 18058
rect 33952 18006 34004 18058
rect 34004 18006 34006 18058
rect 33950 18004 34006 18006
rect 34054 18058 34110 18060
rect 34054 18006 34056 18058
rect 34056 18006 34108 18058
rect 34108 18006 34110 18058
rect 34054 18004 34110 18006
rect 10536 17274 10592 17276
rect 10536 17222 10538 17274
rect 10538 17222 10590 17274
rect 10590 17222 10592 17274
rect 10536 17220 10592 17222
rect 10640 17274 10696 17276
rect 10640 17222 10642 17274
rect 10642 17222 10694 17274
rect 10694 17222 10696 17274
rect 10640 17220 10696 17222
rect 10744 17274 10800 17276
rect 10744 17222 10746 17274
rect 10746 17222 10798 17274
rect 10798 17222 10800 17274
rect 10744 17220 10800 17222
rect 19860 17274 19916 17276
rect 19860 17222 19862 17274
rect 19862 17222 19914 17274
rect 19914 17222 19916 17274
rect 19860 17220 19916 17222
rect 19964 17274 20020 17276
rect 19964 17222 19966 17274
rect 19966 17222 20018 17274
rect 20018 17222 20020 17274
rect 19964 17220 20020 17222
rect 20068 17274 20124 17276
rect 20068 17222 20070 17274
rect 20070 17222 20122 17274
rect 20122 17222 20124 17274
rect 20068 17220 20124 17222
rect 29184 17274 29240 17276
rect 29184 17222 29186 17274
rect 29186 17222 29238 17274
rect 29238 17222 29240 17274
rect 29184 17220 29240 17222
rect 29288 17274 29344 17276
rect 29288 17222 29290 17274
rect 29290 17222 29342 17274
rect 29342 17222 29344 17274
rect 29288 17220 29344 17222
rect 29392 17274 29448 17276
rect 29392 17222 29394 17274
rect 29394 17222 29446 17274
rect 29446 17222 29448 17274
rect 29392 17220 29448 17222
rect 38508 17274 38564 17276
rect 38508 17222 38510 17274
rect 38510 17222 38562 17274
rect 38562 17222 38564 17274
rect 38508 17220 38564 17222
rect 38612 17274 38668 17276
rect 38612 17222 38614 17274
rect 38614 17222 38666 17274
rect 38666 17222 38668 17274
rect 38612 17220 38668 17222
rect 38716 17274 38772 17276
rect 38716 17222 38718 17274
rect 38718 17222 38770 17274
rect 38770 17222 38772 17274
rect 38716 17220 38772 17222
rect 5874 16490 5930 16492
rect 5874 16438 5876 16490
rect 5876 16438 5928 16490
rect 5928 16438 5930 16490
rect 5874 16436 5930 16438
rect 5978 16490 6034 16492
rect 5978 16438 5980 16490
rect 5980 16438 6032 16490
rect 6032 16438 6034 16490
rect 5978 16436 6034 16438
rect 6082 16490 6138 16492
rect 6082 16438 6084 16490
rect 6084 16438 6136 16490
rect 6136 16438 6138 16490
rect 6082 16436 6138 16438
rect 15198 16490 15254 16492
rect 15198 16438 15200 16490
rect 15200 16438 15252 16490
rect 15252 16438 15254 16490
rect 15198 16436 15254 16438
rect 15302 16490 15358 16492
rect 15302 16438 15304 16490
rect 15304 16438 15356 16490
rect 15356 16438 15358 16490
rect 15302 16436 15358 16438
rect 15406 16490 15462 16492
rect 15406 16438 15408 16490
rect 15408 16438 15460 16490
rect 15460 16438 15462 16490
rect 15406 16436 15462 16438
rect 24522 16490 24578 16492
rect 24522 16438 24524 16490
rect 24524 16438 24576 16490
rect 24576 16438 24578 16490
rect 24522 16436 24578 16438
rect 24626 16490 24682 16492
rect 24626 16438 24628 16490
rect 24628 16438 24680 16490
rect 24680 16438 24682 16490
rect 24626 16436 24682 16438
rect 24730 16490 24786 16492
rect 24730 16438 24732 16490
rect 24732 16438 24784 16490
rect 24784 16438 24786 16490
rect 24730 16436 24786 16438
rect 33846 16490 33902 16492
rect 33846 16438 33848 16490
rect 33848 16438 33900 16490
rect 33900 16438 33902 16490
rect 33846 16436 33902 16438
rect 33950 16490 34006 16492
rect 33950 16438 33952 16490
rect 33952 16438 34004 16490
rect 34004 16438 34006 16490
rect 33950 16436 34006 16438
rect 34054 16490 34110 16492
rect 34054 16438 34056 16490
rect 34056 16438 34108 16490
rect 34108 16438 34110 16490
rect 34054 16436 34110 16438
rect 10536 15706 10592 15708
rect 10536 15654 10538 15706
rect 10538 15654 10590 15706
rect 10590 15654 10592 15706
rect 10536 15652 10592 15654
rect 10640 15706 10696 15708
rect 10640 15654 10642 15706
rect 10642 15654 10694 15706
rect 10694 15654 10696 15706
rect 10640 15652 10696 15654
rect 10744 15706 10800 15708
rect 10744 15654 10746 15706
rect 10746 15654 10798 15706
rect 10798 15654 10800 15706
rect 10744 15652 10800 15654
rect 19860 15706 19916 15708
rect 19860 15654 19862 15706
rect 19862 15654 19914 15706
rect 19914 15654 19916 15706
rect 19860 15652 19916 15654
rect 19964 15706 20020 15708
rect 19964 15654 19966 15706
rect 19966 15654 20018 15706
rect 20018 15654 20020 15706
rect 19964 15652 20020 15654
rect 20068 15706 20124 15708
rect 20068 15654 20070 15706
rect 20070 15654 20122 15706
rect 20122 15654 20124 15706
rect 20068 15652 20124 15654
rect 29184 15706 29240 15708
rect 29184 15654 29186 15706
rect 29186 15654 29238 15706
rect 29238 15654 29240 15706
rect 29184 15652 29240 15654
rect 29288 15706 29344 15708
rect 29288 15654 29290 15706
rect 29290 15654 29342 15706
rect 29342 15654 29344 15706
rect 29288 15652 29344 15654
rect 29392 15706 29448 15708
rect 29392 15654 29394 15706
rect 29394 15654 29446 15706
rect 29446 15654 29448 15706
rect 29392 15652 29448 15654
rect 38508 15706 38564 15708
rect 38508 15654 38510 15706
rect 38510 15654 38562 15706
rect 38562 15654 38564 15706
rect 38508 15652 38564 15654
rect 38612 15706 38668 15708
rect 38612 15654 38614 15706
rect 38614 15654 38666 15706
rect 38666 15654 38668 15706
rect 38612 15652 38668 15654
rect 38716 15706 38772 15708
rect 38716 15654 38718 15706
rect 38718 15654 38770 15706
rect 38770 15654 38772 15706
rect 38716 15652 38772 15654
rect 5874 14922 5930 14924
rect 5874 14870 5876 14922
rect 5876 14870 5928 14922
rect 5928 14870 5930 14922
rect 5874 14868 5930 14870
rect 5978 14922 6034 14924
rect 5978 14870 5980 14922
rect 5980 14870 6032 14922
rect 6032 14870 6034 14922
rect 5978 14868 6034 14870
rect 6082 14922 6138 14924
rect 6082 14870 6084 14922
rect 6084 14870 6136 14922
rect 6136 14870 6138 14922
rect 6082 14868 6138 14870
rect 15198 14922 15254 14924
rect 15198 14870 15200 14922
rect 15200 14870 15252 14922
rect 15252 14870 15254 14922
rect 15198 14868 15254 14870
rect 15302 14922 15358 14924
rect 15302 14870 15304 14922
rect 15304 14870 15356 14922
rect 15356 14870 15358 14922
rect 15302 14868 15358 14870
rect 15406 14922 15462 14924
rect 15406 14870 15408 14922
rect 15408 14870 15460 14922
rect 15460 14870 15462 14922
rect 15406 14868 15462 14870
rect 24522 14922 24578 14924
rect 24522 14870 24524 14922
rect 24524 14870 24576 14922
rect 24576 14870 24578 14922
rect 24522 14868 24578 14870
rect 24626 14922 24682 14924
rect 24626 14870 24628 14922
rect 24628 14870 24680 14922
rect 24680 14870 24682 14922
rect 24626 14868 24682 14870
rect 24730 14922 24786 14924
rect 24730 14870 24732 14922
rect 24732 14870 24784 14922
rect 24784 14870 24786 14922
rect 24730 14868 24786 14870
rect 33846 14922 33902 14924
rect 33846 14870 33848 14922
rect 33848 14870 33900 14922
rect 33900 14870 33902 14922
rect 33846 14868 33902 14870
rect 33950 14922 34006 14924
rect 33950 14870 33952 14922
rect 33952 14870 34004 14922
rect 34004 14870 34006 14922
rect 33950 14868 34006 14870
rect 34054 14922 34110 14924
rect 34054 14870 34056 14922
rect 34056 14870 34108 14922
rect 34108 14870 34110 14922
rect 34054 14868 34110 14870
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 5874 13354 5930 13356
rect 5874 13302 5876 13354
rect 5876 13302 5928 13354
rect 5928 13302 5930 13354
rect 5874 13300 5930 13302
rect 5978 13354 6034 13356
rect 5978 13302 5980 13354
rect 5980 13302 6032 13354
rect 6032 13302 6034 13354
rect 5978 13300 6034 13302
rect 6082 13354 6138 13356
rect 6082 13302 6084 13354
rect 6084 13302 6136 13354
rect 6136 13302 6138 13354
rect 6082 13300 6138 13302
rect 15198 13354 15254 13356
rect 15198 13302 15200 13354
rect 15200 13302 15252 13354
rect 15252 13302 15254 13354
rect 15198 13300 15254 13302
rect 15302 13354 15358 13356
rect 15302 13302 15304 13354
rect 15304 13302 15356 13354
rect 15356 13302 15358 13354
rect 15302 13300 15358 13302
rect 15406 13354 15462 13356
rect 15406 13302 15408 13354
rect 15408 13302 15460 13354
rect 15460 13302 15462 13354
rect 15406 13300 15462 13302
rect 24522 13354 24578 13356
rect 24522 13302 24524 13354
rect 24524 13302 24576 13354
rect 24576 13302 24578 13354
rect 24522 13300 24578 13302
rect 24626 13354 24682 13356
rect 24626 13302 24628 13354
rect 24628 13302 24680 13354
rect 24680 13302 24682 13354
rect 24626 13300 24682 13302
rect 24730 13354 24786 13356
rect 24730 13302 24732 13354
rect 24732 13302 24784 13354
rect 24784 13302 24786 13354
rect 24730 13300 24786 13302
rect 33846 13354 33902 13356
rect 33846 13302 33848 13354
rect 33848 13302 33900 13354
rect 33900 13302 33902 13354
rect 33846 13300 33902 13302
rect 33950 13354 34006 13356
rect 33950 13302 33952 13354
rect 33952 13302 34004 13354
rect 34004 13302 34006 13354
rect 33950 13300 34006 13302
rect 34054 13354 34110 13356
rect 34054 13302 34056 13354
rect 34056 13302 34108 13354
rect 34108 13302 34110 13354
rect 34054 13300 34110 13302
rect 10536 12570 10592 12572
rect 10536 12518 10538 12570
rect 10538 12518 10590 12570
rect 10590 12518 10592 12570
rect 10536 12516 10592 12518
rect 10640 12570 10696 12572
rect 10640 12518 10642 12570
rect 10642 12518 10694 12570
rect 10694 12518 10696 12570
rect 10640 12516 10696 12518
rect 10744 12570 10800 12572
rect 10744 12518 10746 12570
rect 10746 12518 10798 12570
rect 10798 12518 10800 12570
rect 10744 12516 10800 12518
rect 19860 12570 19916 12572
rect 19860 12518 19862 12570
rect 19862 12518 19914 12570
rect 19914 12518 19916 12570
rect 19860 12516 19916 12518
rect 19964 12570 20020 12572
rect 19964 12518 19966 12570
rect 19966 12518 20018 12570
rect 20018 12518 20020 12570
rect 19964 12516 20020 12518
rect 20068 12570 20124 12572
rect 20068 12518 20070 12570
rect 20070 12518 20122 12570
rect 20122 12518 20124 12570
rect 20068 12516 20124 12518
rect 29184 12570 29240 12572
rect 29184 12518 29186 12570
rect 29186 12518 29238 12570
rect 29238 12518 29240 12570
rect 29184 12516 29240 12518
rect 29288 12570 29344 12572
rect 29288 12518 29290 12570
rect 29290 12518 29342 12570
rect 29342 12518 29344 12570
rect 29288 12516 29344 12518
rect 29392 12570 29448 12572
rect 29392 12518 29394 12570
rect 29394 12518 29446 12570
rect 29446 12518 29448 12570
rect 29392 12516 29448 12518
rect 38508 12570 38564 12572
rect 38508 12518 38510 12570
rect 38510 12518 38562 12570
rect 38562 12518 38564 12570
rect 38508 12516 38564 12518
rect 38612 12570 38668 12572
rect 38612 12518 38614 12570
rect 38614 12518 38666 12570
rect 38666 12518 38668 12570
rect 38612 12516 38668 12518
rect 38716 12570 38772 12572
rect 38716 12518 38718 12570
rect 38718 12518 38770 12570
rect 38770 12518 38772 12570
rect 38716 12516 38772 12518
rect 5874 11786 5930 11788
rect 5874 11734 5876 11786
rect 5876 11734 5928 11786
rect 5928 11734 5930 11786
rect 5874 11732 5930 11734
rect 5978 11786 6034 11788
rect 5978 11734 5980 11786
rect 5980 11734 6032 11786
rect 6032 11734 6034 11786
rect 5978 11732 6034 11734
rect 6082 11786 6138 11788
rect 6082 11734 6084 11786
rect 6084 11734 6136 11786
rect 6136 11734 6138 11786
rect 6082 11732 6138 11734
rect 15198 11786 15254 11788
rect 15198 11734 15200 11786
rect 15200 11734 15252 11786
rect 15252 11734 15254 11786
rect 15198 11732 15254 11734
rect 15302 11786 15358 11788
rect 15302 11734 15304 11786
rect 15304 11734 15356 11786
rect 15356 11734 15358 11786
rect 15302 11732 15358 11734
rect 15406 11786 15462 11788
rect 15406 11734 15408 11786
rect 15408 11734 15460 11786
rect 15460 11734 15462 11786
rect 15406 11732 15462 11734
rect 24522 11786 24578 11788
rect 24522 11734 24524 11786
rect 24524 11734 24576 11786
rect 24576 11734 24578 11786
rect 24522 11732 24578 11734
rect 24626 11786 24682 11788
rect 24626 11734 24628 11786
rect 24628 11734 24680 11786
rect 24680 11734 24682 11786
rect 24626 11732 24682 11734
rect 24730 11786 24786 11788
rect 24730 11734 24732 11786
rect 24732 11734 24784 11786
rect 24784 11734 24786 11786
rect 24730 11732 24786 11734
rect 33846 11786 33902 11788
rect 33846 11734 33848 11786
rect 33848 11734 33900 11786
rect 33900 11734 33902 11786
rect 33846 11732 33902 11734
rect 33950 11786 34006 11788
rect 33950 11734 33952 11786
rect 33952 11734 34004 11786
rect 34004 11734 34006 11786
rect 33950 11732 34006 11734
rect 34054 11786 34110 11788
rect 34054 11734 34056 11786
rect 34056 11734 34108 11786
rect 34108 11734 34110 11786
rect 34054 11732 34110 11734
rect 10536 11002 10592 11004
rect 10536 10950 10538 11002
rect 10538 10950 10590 11002
rect 10590 10950 10592 11002
rect 10536 10948 10592 10950
rect 10640 11002 10696 11004
rect 10640 10950 10642 11002
rect 10642 10950 10694 11002
rect 10694 10950 10696 11002
rect 10640 10948 10696 10950
rect 10744 11002 10800 11004
rect 10744 10950 10746 11002
rect 10746 10950 10798 11002
rect 10798 10950 10800 11002
rect 10744 10948 10800 10950
rect 19860 11002 19916 11004
rect 19860 10950 19862 11002
rect 19862 10950 19914 11002
rect 19914 10950 19916 11002
rect 19860 10948 19916 10950
rect 19964 11002 20020 11004
rect 19964 10950 19966 11002
rect 19966 10950 20018 11002
rect 20018 10950 20020 11002
rect 19964 10948 20020 10950
rect 20068 11002 20124 11004
rect 20068 10950 20070 11002
rect 20070 10950 20122 11002
rect 20122 10950 20124 11002
rect 20068 10948 20124 10950
rect 29184 11002 29240 11004
rect 29184 10950 29186 11002
rect 29186 10950 29238 11002
rect 29238 10950 29240 11002
rect 29184 10948 29240 10950
rect 29288 11002 29344 11004
rect 29288 10950 29290 11002
rect 29290 10950 29342 11002
rect 29342 10950 29344 11002
rect 29288 10948 29344 10950
rect 29392 11002 29448 11004
rect 29392 10950 29394 11002
rect 29394 10950 29446 11002
rect 29446 10950 29448 11002
rect 29392 10948 29448 10950
rect 38508 11002 38564 11004
rect 38508 10950 38510 11002
rect 38510 10950 38562 11002
rect 38562 10950 38564 11002
rect 38508 10948 38564 10950
rect 38612 11002 38668 11004
rect 38612 10950 38614 11002
rect 38614 10950 38666 11002
rect 38666 10950 38668 11002
rect 38612 10948 38668 10950
rect 38716 11002 38772 11004
rect 38716 10950 38718 11002
rect 38718 10950 38770 11002
rect 38770 10950 38772 11002
rect 38716 10948 38772 10950
rect 5874 10218 5930 10220
rect 5874 10166 5876 10218
rect 5876 10166 5928 10218
rect 5928 10166 5930 10218
rect 5874 10164 5930 10166
rect 5978 10218 6034 10220
rect 5978 10166 5980 10218
rect 5980 10166 6032 10218
rect 6032 10166 6034 10218
rect 5978 10164 6034 10166
rect 6082 10218 6138 10220
rect 6082 10166 6084 10218
rect 6084 10166 6136 10218
rect 6136 10166 6138 10218
rect 6082 10164 6138 10166
rect 15198 10218 15254 10220
rect 15198 10166 15200 10218
rect 15200 10166 15252 10218
rect 15252 10166 15254 10218
rect 15198 10164 15254 10166
rect 15302 10218 15358 10220
rect 15302 10166 15304 10218
rect 15304 10166 15356 10218
rect 15356 10166 15358 10218
rect 15302 10164 15358 10166
rect 15406 10218 15462 10220
rect 15406 10166 15408 10218
rect 15408 10166 15460 10218
rect 15460 10166 15462 10218
rect 15406 10164 15462 10166
rect 24522 10218 24578 10220
rect 24522 10166 24524 10218
rect 24524 10166 24576 10218
rect 24576 10166 24578 10218
rect 24522 10164 24578 10166
rect 24626 10218 24682 10220
rect 24626 10166 24628 10218
rect 24628 10166 24680 10218
rect 24680 10166 24682 10218
rect 24626 10164 24682 10166
rect 24730 10218 24786 10220
rect 24730 10166 24732 10218
rect 24732 10166 24784 10218
rect 24784 10166 24786 10218
rect 24730 10164 24786 10166
rect 33846 10218 33902 10220
rect 33846 10166 33848 10218
rect 33848 10166 33900 10218
rect 33900 10166 33902 10218
rect 33846 10164 33902 10166
rect 33950 10218 34006 10220
rect 33950 10166 33952 10218
rect 33952 10166 34004 10218
rect 34004 10166 34006 10218
rect 33950 10164 34006 10166
rect 34054 10218 34110 10220
rect 34054 10166 34056 10218
rect 34056 10166 34108 10218
rect 34108 10166 34110 10218
rect 34054 10164 34110 10166
rect 10536 9434 10592 9436
rect 10536 9382 10538 9434
rect 10538 9382 10590 9434
rect 10590 9382 10592 9434
rect 10536 9380 10592 9382
rect 10640 9434 10696 9436
rect 10640 9382 10642 9434
rect 10642 9382 10694 9434
rect 10694 9382 10696 9434
rect 10640 9380 10696 9382
rect 10744 9434 10800 9436
rect 10744 9382 10746 9434
rect 10746 9382 10798 9434
rect 10798 9382 10800 9434
rect 10744 9380 10800 9382
rect 19860 9434 19916 9436
rect 19860 9382 19862 9434
rect 19862 9382 19914 9434
rect 19914 9382 19916 9434
rect 19860 9380 19916 9382
rect 19964 9434 20020 9436
rect 19964 9382 19966 9434
rect 19966 9382 20018 9434
rect 20018 9382 20020 9434
rect 19964 9380 20020 9382
rect 20068 9434 20124 9436
rect 20068 9382 20070 9434
rect 20070 9382 20122 9434
rect 20122 9382 20124 9434
rect 20068 9380 20124 9382
rect 29184 9434 29240 9436
rect 29184 9382 29186 9434
rect 29186 9382 29238 9434
rect 29238 9382 29240 9434
rect 29184 9380 29240 9382
rect 29288 9434 29344 9436
rect 29288 9382 29290 9434
rect 29290 9382 29342 9434
rect 29342 9382 29344 9434
rect 29288 9380 29344 9382
rect 29392 9434 29448 9436
rect 29392 9382 29394 9434
rect 29394 9382 29446 9434
rect 29446 9382 29448 9434
rect 29392 9380 29448 9382
rect 38508 9434 38564 9436
rect 38508 9382 38510 9434
rect 38510 9382 38562 9434
rect 38562 9382 38564 9434
rect 38508 9380 38564 9382
rect 38612 9434 38668 9436
rect 38612 9382 38614 9434
rect 38614 9382 38666 9434
rect 38666 9382 38668 9434
rect 38612 9380 38668 9382
rect 38716 9434 38772 9436
rect 38716 9382 38718 9434
rect 38718 9382 38770 9434
rect 38770 9382 38772 9434
rect 38716 9380 38772 9382
rect 24220 8930 24276 8932
rect 24220 8878 24222 8930
rect 24222 8878 24274 8930
rect 24274 8878 24276 8930
rect 24220 8876 24276 8878
rect 5874 8650 5930 8652
rect 5874 8598 5876 8650
rect 5876 8598 5928 8650
rect 5928 8598 5930 8650
rect 5874 8596 5930 8598
rect 5978 8650 6034 8652
rect 5978 8598 5980 8650
rect 5980 8598 6032 8650
rect 6032 8598 6034 8650
rect 5978 8596 6034 8598
rect 6082 8650 6138 8652
rect 6082 8598 6084 8650
rect 6084 8598 6136 8650
rect 6136 8598 6138 8650
rect 6082 8596 6138 8598
rect 15198 8650 15254 8652
rect 15198 8598 15200 8650
rect 15200 8598 15252 8650
rect 15252 8598 15254 8650
rect 15198 8596 15254 8598
rect 15302 8650 15358 8652
rect 15302 8598 15304 8650
rect 15304 8598 15356 8650
rect 15356 8598 15358 8650
rect 15302 8596 15358 8598
rect 15406 8650 15462 8652
rect 15406 8598 15408 8650
rect 15408 8598 15460 8650
rect 15460 8598 15462 8650
rect 15406 8596 15462 8598
rect 23212 8034 23268 8036
rect 23212 7982 23214 8034
rect 23214 7982 23266 8034
rect 23266 7982 23268 8034
rect 23212 7980 23268 7982
rect 10536 7866 10592 7868
rect 10536 7814 10538 7866
rect 10538 7814 10590 7866
rect 10590 7814 10592 7866
rect 10536 7812 10592 7814
rect 10640 7866 10696 7868
rect 10640 7814 10642 7866
rect 10642 7814 10694 7866
rect 10694 7814 10696 7866
rect 10640 7812 10696 7814
rect 10744 7866 10800 7868
rect 10744 7814 10746 7866
rect 10746 7814 10798 7866
rect 10798 7814 10800 7866
rect 10744 7812 10800 7814
rect 19860 7866 19916 7868
rect 19860 7814 19862 7866
rect 19862 7814 19914 7866
rect 19914 7814 19916 7866
rect 19860 7812 19916 7814
rect 19964 7866 20020 7868
rect 19964 7814 19966 7866
rect 19966 7814 20018 7866
rect 20018 7814 20020 7866
rect 19964 7812 20020 7814
rect 20068 7866 20124 7868
rect 20068 7814 20070 7866
rect 20070 7814 20122 7866
rect 20122 7814 20124 7866
rect 20068 7812 20124 7814
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 19628 6748 19684 6804
rect 10536 6298 10592 6300
rect 10536 6246 10538 6298
rect 10538 6246 10590 6298
rect 10590 6246 10592 6298
rect 10536 6244 10592 6246
rect 10640 6298 10696 6300
rect 10640 6246 10642 6298
rect 10642 6246 10694 6298
rect 10694 6246 10696 6298
rect 10640 6244 10696 6246
rect 10744 6298 10800 6300
rect 10744 6246 10746 6298
rect 10746 6246 10798 6298
rect 10798 6246 10800 6298
rect 10744 6244 10800 6246
rect 5874 5514 5930 5516
rect 5874 5462 5876 5514
rect 5876 5462 5928 5514
rect 5928 5462 5930 5514
rect 5874 5460 5930 5462
rect 5978 5514 6034 5516
rect 5978 5462 5980 5514
rect 5980 5462 6032 5514
rect 6032 5462 6034 5514
rect 5978 5460 6034 5462
rect 6082 5514 6138 5516
rect 6082 5462 6084 5514
rect 6084 5462 6136 5514
rect 6136 5462 6138 5514
rect 6082 5460 6138 5462
rect 15198 5514 15254 5516
rect 15198 5462 15200 5514
rect 15200 5462 15252 5514
rect 15252 5462 15254 5514
rect 15198 5460 15254 5462
rect 15302 5514 15358 5516
rect 15302 5462 15304 5514
rect 15304 5462 15356 5514
rect 15356 5462 15358 5514
rect 15302 5460 15358 5462
rect 15406 5514 15462 5516
rect 15406 5462 15408 5514
rect 15408 5462 15460 5514
rect 15460 5462 15462 5514
rect 15406 5460 15462 5462
rect 21980 6748 22036 6804
rect 19860 6298 19916 6300
rect 19860 6246 19862 6298
rect 19862 6246 19914 6298
rect 19914 6246 19916 6298
rect 19860 6244 19916 6246
rect 19964 6298 20020 6300
rect 19964 6246 19966 6298
rect 19966 6246 20018 6298
rect 20018 6246 20020 6298
rect 19964 6244 20020 6246
rect 20068 6298 20124 6300
rect 20068 6246 20070 6298
rect 20070 6246 20122 6298
rect 20122 6246 20124 6298
rect 20068 6244 20124 6246
rect 21420 5852 21476 5908
rect 10536 4730 10592 4732
rect 10536 4678 10538 4730
rect 10538 4678 10590 4730
rect 10590 4678 10592 4730
rect 10536 4676 10592 4678
rect 10640 4730 10696 4732
rect 10640 4678 10642 4730
rect 10642 4678 10694 4730
rect 10694 4678 10696 4730
rect 10640 4676 10696 4678
rect 10744 4730 10800 4732
rect 10744 4678 10746 4730
rect 10746 4678 10798 4730
rect 10798 4678 10800 4730
rect 10744 4676 10800 4678
rect 18844 4562 18900 4564
rect 18844 4510 18846 4562
rect 18846 4510 18898 4562
rect 18898 4510 18900 4562
rect 18844 4508 18900 4510
rect 19180 4562 19236 4564
rect 19180 4510 19182 4562
rect 19182 4510 19234 4562
rect 19234 4510 19236 4562
rect 19180 4508 19236 4510
rect 5874 3946 5930 3948
rect 5874 3894 5876 3946
rect 5876 3894 5928 3946
rect 5928 3894 5930 3946
rect 5874 3892 5930 3894
rect 5978 3946 6034 3948
rect 5978 3894 5980 3946
rect 5980 3894 6032 3946
rect 6032 3894 6034 3946
rect 5978 3892 6034 3894
rect 6082 3946 6138 3948
rect 6082 3894 6084 3946
rect 6084 3894 6136 3946
rect 6136 3894 6138 3946
rect 6082 3892 6138 3894
rect 15198 3946 15254 3948
rect 15198 3894 15200 3946
rect 15200 3894 15252 3946
rect 15252 3894 15254 3946
rect 15198 3892 15254 3894
rect 15302 3946 15358 3948
rect 15302 3894 15304 3946
rect 15304 3894 15356 3946
rect 15356 3894 15358 3946
rect 15302 3892 15358 3894
rect 15406 3946 15462 3948
rect 15406 3894 15408 3946
rect 15408 3894 15460 3946
rect 15460 3894 15462 3946
rect 15406 3892 15462 3894
rect 16604 3778 16660 3780
rect 16604 3726 16606 3778
rect 16606 3726 16658 3778
rect 16658 3726 16660 3778
rect 16604 3724 16660 3726
rect 12572 3500 12628 3556
rect 2716 3388 2772 3444
rect 10536 3162 10592 3164
rect 10536 3110 10538 3162
rect 10538 3110 10590 3162
rect 10590 3110 10592 3162
rect 10536 3108 10592 3110
rect 10640 3162 10696 3164
rect 10640 3110 10642 3162
rect 10642 3110 10694 3162
rect 10694 3110 10696 3162
rect 10640 3108 10696 3110
rect 10744 3162 10800 3164
rect 10744 3110 10746 3162
rect 10746 3110 10798 3162
rect 10798 3110 10800 3162
rect 10744 3108 10800 3110
rect 17724 3554 17780 3556
rect 17724 3502 17726 3554
rect 17726 3502 17778 3554
rect 17778 3502 17780 3554
rect 17724 3500 17780 3502
rect 18172 3554 18228 3556
rect 18172 3502 18174 3554
rect 18174 3502 18226 3554
rect 18226 3502 18228 3554
rect 18172 3500 18228 3502
rect 18620 3554 18676 3556
rect 18620 3502 18622 3554
rect 18622 3502 18674 3554
rect 18674 3502 18676 3554
rect 18620 3500 18676 3502
rect 19860 4730 19916 4732
rect 19860 4678 19862 4730
rect 19862 4678 19914 4730
rect 19914 4678 19916 4730
rect 19860 4676 19916 4678
rect 19964 4730 20020 4732
rect 19964 4678 19966 4730
rect 19966 4678 20018 4730
rect 20018 4678 20020 4730
rect 19964 4676 20020 4678
rect 20068 4730 20124 4732
rect 20068 4678 20070 4730
rect 20070 4678 20122 4730
rect 20122 4678 20124 4730
rect 20068 4676 20124 4678
rect 20188 4508 20244 4564
rect 19292 4060 19348 4116
rect 20300 4114 20356 4116
rect 20300 4062 20302 4114
rect 20302 4062 20354 4114
rect 20354 4062 20356 4114
rect 20300 4060 20356 4062
rect 20188 3612 20244 3668
rect 20636 3666 20692 3668
rect 20636 3614 20638 3666
rect 20638 3614 20690 3666
rect 20690 3614 20692 3666
rect 20636 3612 20692 3614
rect 21980 5906 22036 5908
rect 21980 5854 21982 5906
rect 21982 5854 22034 5906
rect 22034 5854 22036 5906
rect 21980 5852 22036 5854
rect 24522 8650 24578 8652
rect 24522 8598 24524 8650
rect 24524 8598 24576 8650
rect 24576 8598 24578 8650
rect 24522 8596 24578 8598
rect 24626 8650 24682 8652
rect 24626 8598 24628 8650
rect 24628 8598 24680 8650
rect 24680 8598 24682 8650
rect 24626 8596 24682 8598
rect 24730 8650 24786 8652
rect 24730 8598 24732 8650
rect 24732 8598 24784 8650
rect 24784 8598 24786 8650
rect 24730 8596 24786 8598
rect 24220 7980 24276 8036
rect 24444 8034 24500 8036
rect 24444 7982 24446 8034
rect 24446 7982 24498 8034
rect 24498 7982 24500 8034
rect 24444 7980 24500 7982
rect 25676 8930 25732 8932
rect 25676 8878 25678 8930
rect 25678 8878 25730 8930
rect 25730 8878 25732 8930
rect 25676 8876 25732 8878
rect 26124 8930 26180 8932
rect 26124 8878 26126 8930
rect 26126 8878 26178 8930
rect 26178 8878 26180 8930
rect 26124 8876 26180 8878
rect 26572 8930 26628 8932
rect 26572 8878 26574 8930
rect 26574 8878 26626 8930
rect 26626 8878 26628 8930
rect 26572 8876 26628 8878
rect 26908 8930 26964 8932
rect 26908 8878 26910 8930
rect 26910 8878 26962 8930
rect 26962 8878 26964 8930
rect 26908 8876 26964 8878
rect 33846 8650 33902 8652
rect 33846 8598 33848 8650
rect 33848 8598 33900 8650
rect 33900 8598 33902 8650
rect 33846 8596 33902 8598
rect 33950 8650 34006 8652
rect 33950 8598 33952 8650
rect 33952 8598 34004 8650
rect 34004 8598 34006 8650
rect 33950 8596 34006 8598
rect 34054 8650 34110 8652
rect 34054 8598 34056 8650
rect 34056 8598 34108 8650
rect 34108 8598 34110 8650
rect 34054 8596 34110 8598
rect 22988 6466 23044 6468
rect 22988 6414 22990 6466
rect 22990 6414 23042 6466
rect 23042 6414 23044 6466
rect 22988 6412 23044 6414
rect 23660 6466 23716 6468
rect 23660 6414 23662 6466
rect 23662 6414 23714 6466
rect 23714 6414 23716 6466
rect 23660 6412 23716 6414
rect 22764 5682 22820 5684
rect 22764 5630 22766 5682
rect 22766 5630 22818 5682
rect 22818 5630 22820 5682
rect 22764 5628 22820 5630
rect 23212 5628 23268 5684
rect 21420 4060 21476 4116
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 25340 8034 25396 8036
rect 25340 7982 25342 8034
rect 25342 7982 25394 8034
rect 25394 7982 25396 8034
rect 25340 7980 25396 7982
rect 25564 7362 25620 7364
rect 25564 7310 25566 7362
rect 25566 7310 25618 7362
rect 25618 7310 25620 7362
rect 25564 7308 25620 7310
rect 26012 7362 26068 7364
rect 26012 7310 26014 7362
rect 26014 7310 26066 7362
rect 26066 7310 26068 7362
rect 26012 7308 26068 7310
rect 23436 5682 23492 5684
rect 23436 5630 23438 5682
rect 23438 5630 23490 5682
rect 23490 5630 23492 5682
rect 23436 5628 23492 5630
rect 21532 4450 21588 4452
rect 21532 4398 21534 4450
rect 21534 4398 21586 4450
rect 21586 4398 21588 4450
rect 21532 4396 21588 4398
rect 20972 3612 21028 3668
rect 19628 3500 19684 3556
rect 19852 3554 19908 3556
rect 19852 3502 19854 3554
rect 19854 3502 19906 3554
rect 19906 3502 19908 3554
rect 19852 3500 19908 3502
rect 20524 3554 20580 3556
rect 20524 3502 20526 3554
rect 20526 3502 20578 3554
rect 20578 3502 20580 3554
rect 20524 3500 20580 3502
rect 22204 4450 22260 4452
rect 22204 4398 22206 4450
rect 22206 4398 22258 4450
rect 22258 4398 22260 4450
rect 22204 4396 22260 4398
rect 21644 3666 21700 3668
rect 21644 3614 21646 3666
rect 21646 3614 21698 3666
rect 21698 3614 21700 3666
rect 21644 3612 21700 3614
rect 21532 3554 21588 3556
rect 21532 3502 21534 3554
rect 21534 3502 21586 3554
rect 21586 3502 21588 3554
rect 21532 3500 21588 3502
rect 16044 3442 16100 3444
rect 16044 3390 16046 3442
rect 16046 3390 16098 3442
rect 16098 3390 16100 3442
rect 16044 3388 16100 3390
rect 16492 3442 16548 3444
rect 16492 3390 16494 3442
rect 16494 3390 16546 3442
rect 16546 3390 16548 3442
rect 25004 6466 25060 6468
rect 25004 6414 25006 6466
rect 25006 6414 25058 6466
rect 25058 6414 25060 6466
rect 25004 6412 25060 6414
rect 24108 5682 24164 5684
rect 24108 5630 24110 5682
rect 24110 5630 24162 5682
rect 24162 5630 24164 5682
rect 24108 5628 24164 5630
rect 23996 4956 24052 5012
rect 24522 5514 24578 5516
rect 24522 5462 24524 5514
rect 24524 5462 24576 5514
rect 24576 5462 24578 5514
rect 24522 5460 24578 5462
rect 24626 5514 24682 5516
rect 24626 5462 24628 5514
rect 24628 5462 24680 5514
rect 24680 5462 24682 5514
rect 24626 5460 24682 5462
rect 24730 5514 24786 5516
rect 24730 5462 24732 5514
rect 24732 5462 24784 5514
rect 24784 5462 24786 5514
rect 24730 5460 24786 5462
rect 26236 6748 26292 6804
rect 26460 6748 26516 6804
rect 27356 8034 27412 8036
rect 27356 7982 27358 8034
rect 27358 7982 27410 8034
rect 27410 7982 27412 8034
rect 27356 7980 27412 7982
rect 26908 7362 26964 7364
rect 26908 7310 26910 7362
rect 26910 7310 26962 7362
rect 26962 7310 26964 7362
rect 26908 7308 26964 7310
rect 25676 6466 25732 6468
rect 25676 6414 25678 6466
rect 25678 6414 25730 6466
rect 25730 6414 25732 6466
rect 25676 6412 25732 6414
rect 25788 6130 25844 6132
rect 25788 6078 25790 6130
rect 25790 6078 25842 6130
rect 25842 6078 25844 6130
rect 25788 6076 25844 6078
rect 24332 5068 24388 5124
rect 22316 3666 22372 3668
rect 22316 3614 22318 3666
rect 22318 3614 22370 3666
rect 22370 3614 22372 3666
rect 22316 3612 22372 3614
rect 22988 3666 23044 3668
rect 22988 3614 22990 3666
rect 22990 3614 23042 3666
rect 23042 3614 23044 3666
rect 22988 3612 23044 3614
rect 23548 4338 23604 4340
rect 23548 4286 23550 4338
rect 23550 4286 23602 4338
rect 23602 4286 23604 4338
rect 23548 4284 23604 4286
rect 22204 3554 22260 3556
rect 22204 3502 22206 3554
rect 22206 3502 22258 3554
rect 22258 3502 22260 3554
rect 22204 3500 22260 3502
rect 22876 3554 22932 3556
rect 22876 3502 22878 3554
rect 22878 3502 22930 3554
rect 22930 3502 22932 3554
rect 22876 3500 22932 3502
rect 16492 3388 16548 3390
rect 19860 3162 19916 3164
rect 19860 3110 19862 3162
rect 19862 3110 19914 3162
rect 19914 3110 19916 3162
rect 19860 3108 19916 3110
rect 19964 3162 20020 3164
rect 19964 3110 19966 3162
rect 19966 3110 20018 3162
rect 20018 3110 20020 3162
rect 19964 3108 20020 3110
rect 20068 3162 20124 3164
rect 20068 3110 20070 3162
rect 20070 3110 20122 3162
rect 20122 3110 20124 3162
rect 20068 3108 20124 3110
rect 24220 4338 24276 4340
rect 24220 4286 24222 4338
rect 24222 4286 24274 4338
rect 24274 4286 24276 4338
rect 24220 4284 24276 4286
rect 25116 5122 25172 5124
rect 25116 5070 25118 5122
rect 25118 5070 25170 5122
rect 25170 5070 25172 5122
rect 25116 5068 25172 5070
rect 25676 5068 25732 5124
rect 24780 4956 24836 5012
rect 28252 8034 28308 8036
rect 28252 7982 28254 8034
rect 28254 7982 28306 8034
rect 28306 7982 28308 8034
rect 28252 7980 28308 7982
rect 28700 8034 28756 8036
rect 28700 7982 28702 8034
rect 28702 7982 28754 8034
rect 28754 7982 28756 8034
rect 28700 7980 28756 7982
rect 29184 7866 29240 7868
rect 29184 7814 29186 7866
rect 29186 7814 29238 7866
rect 29238 7814 29240 7866
rect 29184 7812 29240 7814
rect 29288 7866 29344 7868
rect 29288 7814 29290 7866
rect 29290 7814 29342 7866
rect 29342 7814 29344 7866
rect 29288 7812 29344 7814
rect 29392 7866 29448 7868
rect 29392 7814 29394 7866
rect 29394 7814 29446 7866
rect 29446 7814 29448 7866
rect 29392 7812 29448 7814
rect 38508 7866 38564 7868
rect 38508 7814 38510 7866
rect 38510 7814 38562 7866
rect 38562 7814 38564 7866
rect 38508 7812 38564 7814
rect 38612 7866 38668 7868
rect 38612 7814 38614 7866
rect 38614 7814 38666 7866
rect 38666 7814 38668 7866
rect 38612 7812 38668 7814
rect 38716 7866 38772 7868
rect 38716 7814 38718 7866
rect 38718 7814 38770 7866
rect 38770 7814 38772 7866
rect 38716 7812 38772 7814
rect 27468 6802 27524 6804
rect 27468 6750 27470 6802
rect 27470 6750 27522 6802
rect 27522 6750 27524 6802
rect 27468 6748 27524 6750
rect 26348 6076 26404 6132
rect 26460 6412 26516 6468
rect 27020 6466 27076 6468
rect 27020 6414 27022 6466
rect 27022 6414 27074 6466
rect 27074 6414 27076 6466
rect 27020 6412 27076 6414
rect 27132 4844 27188 4900
rect 25340 4284 25396 4340
rect 24522 3946 24578 3948
rect 24522 3894 24524 3946
rect 24524 3894 24576 3946
rect 24576 3894 24578 3946
rect 24522 3892 24578 3894
rect 24626 3946 24682 3948
rect 24626 3894 24628 3946
rect 24628 3894 24680 3946
rect 24680 3894 24682 3946
rect 24626 3892 24682 3894
rect 24730 3946 24786 3948
rect 24730 3894 24732 3946
rect 24732 3894 24784 3946
rect 24784 3894 24786 3946
rect 24730 3892 24786 3894
rect 23660 3666 23716 3668
rect 23660 3614 23662 3666
rect 23662 3614 23714 3666
rect 23714 3614 23716 3666
rect 23660 3612 23716 3614
rect 24332 3612 24388 3668
rect 23548 3554 23604 3556
rect 23548 3502 23550 3554
rect 23550 3502 23602 3554
rect 23602 3502 23604 3554
rect 23548 3500 23604 3502
rect 25676 4338 25732 4340
rect 25676 4286 25678 4338
rect 25678 4286 25730 4338
rect 25730 4286 25732 4338
rect 25676 4284 25732 4286
rect 27804 6130 27860 6132
rect 27804 6078 27806 6130
rect 27806 6078 27858 6130
rect 27858 6078 27860 6130
rect 27804 6076 27860 6078
rect 28812 6802 28868 6804
rect 28812 6750 28814 6802
rect 28814 6750 28866 6802
rect 28866 6750 28868 6802
rect 28812 6748 28868 6750
rect 28588 6524 28644 6580
rect 28364 6466 28420 6468
rect 28364 6414 28366 6466
rect 28366 6414 28418 6466
rect 28418 6414 28420 6466
rect 28364 6412 28420 6414
rect 28252 6076 28308 6132
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 30044 6748 30100 6804
rect 30940 6636 30996 6692
rect 29596 6578 29652 6580
rect 29596 6526 29598 6578
rect 29598 6526 29650 6578
rect 29650 6526 29652 6578
rect 29596 6524 29652 6526
rect 29036 6412 29092 6468
rect 29184 6298 29240 6300
rect 29184 6246 29186 6298
rect 29186 6246 29238 6298
rect 29238 6246 29240 6298
rect 29184 6244 29240 6246
rect 29288 6298 29344 6300
rect 29288 6246 29290 6298
rect 29290 6246 29342 6298
rect 29342 6246 29344 6298
rect 29288 6244 29344 6246
rect 29392 6298 29448 6300
rect 29392 6246 29394 6298
rect 29394 6246 29446 6298
rect 29446 6246 29448 6298
rect 29392 6244 29448 6246
rect 30156 6578 30212 6580
rect 30156 6526 30158 6578
rect 30158 6526 30210 6578
rect 30210 6526 30212 6578
rect 30156 6524 30212 6526
rect 29820 4956 29876 5012
rect 27244 4508 27300 4564
rect 27692 4844 27748 4900
rect 27132 4114 27188 4116
rect 27132 4062 27134 4114
rect 27134 4062 27186 4114
rect 27186 4062 27188 4114
rect 27132 4060 27188 4062
rect 27244 3724 27300 3780
rect 25340 3554 25396 3556
rect 25340 3502 25342 3554
rect 25342 3502 25394 3554
rect 25394 3502 25396 3554
rect 25340 3500 25396 3502
rect 26012 3554 26068 3556
rect 26012 3502 26014 3554
rect 26014 3502 26066 3554
rect 26066 3502 26068 3554
rect 26012 3500 26068 3502
rect 26684 3554 26740 3556
rect 26684 3502 26686 3554
rect 26686 3502 26738 3554
rect 26738 3502 26740 3554
rect 26684 3500 26740 3502
rect 29184 4730 29240 4732
rect 29184 4678 29186 4730
rect 29186 4678 29238 4730
rect 29238 4678 29240 4730
rect 29184 4676 29240 4678
rect 29288 4730 29344 4732
rect 29288 4678 29290 4730
rect 29290 4678 29342 4730
rect 29342 4678 29344 4730
rect 29288 4676 29344 4678
rect 29392 4730 29448 4732
rect 29392 4678 29394 4730
rect 29394 4678 29446 4730
rect 29446 4678 29448 4730
rect 29392 4676 29448 4678
rect 27804 4562 27860 4564
rect 27804 4510 27806 4562
rect 27806 4510 27858 4562
rect 27858 4510 27860 4562
rect 27804 4508 27860 4510
rect 28476 4562 28532 4564
rect 28476 4510 28478 4562
rect 28478 4510 28530 4562
rect 28530 4510 28532 4562
rect 28476 4508 28532 4510
rect 29148 4562 29204 4564
rect 29148 4510 29150 4562
rect 29150 4510 29202 4562
rect 29202 4510 29204 4562
rect 29148 4508 29204 4510
rect 29820 4562 29876 4564
rect 29820 4510 29822 4562
rect 29822 4510 29874 4562
rect 29874 4510 29876 4562
rect 29820 4508 29876 4510
rect 29260 4396 29316 4452
rect 27692 4060 27748 4116
rect 27692 3612 27748 3668
rect 28028 3666 28084 3668
rect 28028 3614 28030 3666
rect 28030 3614 28082 3666
rect 28082 3614 28084 3666
rect 28028 3612 28084 3614
rect 28364 3612 28420 3668
rect 29036 4338 29092 4340
rect 29036 4286 29038 4338
rect 29038 4286 29090 4338
rect 29090 4286 29092 4338
rect 29036 4284 29092 4286
rect 27468 3554 27524 3556
rect 27468 3502 27470 3554
rect 27470 3502 27522 3554
rect 27522 3502 27524 3554
rect 27468 3500 27524 3502
rect 28140 3554 28196 3556
rect 28140 3502 28142 3554
rect 28142 3502 28194 3554
rect 28194 3502 28196 3554
rect 28140 3500 28196 3502
rect 29708 4338 29764 4340
rect 29708 4286 29710 4338
rect 29710 4286 29762 4338
rect 29762 4286 29764 4338
rect 29708 4284 29764 4286
rect 30380 4956 30436 5012
rect 31052 5010 31108 5012
rect 31052 4958 31054 5010
rect 31054 4958 31106 5010
rect 31106 4958 31108 5010
rect 31052 4956 31108 4958
rect 38508 6298 38564 6300
rect 38508 6246 38510 6298
rect 38510 6246 38562 6298
rect 38562 6246 38564 6298
rect 38508 6244 38564 6246
rect 38612 6298 38668 6300
rect 38612 6246 38614 6298
rect 38614 6246 38666 6298
rect 38666 6246 38668 6298
rect 38612 6244 38668 6246
rect 38716 6298 38772 6300
rect 38716 6246 38718 6298
rect 38718 6246 38770 6298
rect 38770 6246 38772 6298
rect 38716 6244 38772 6246
rect 31836 5068 31892 5124
rect 31500 4956 31556 5012
rect 31164 4844 31220 4900
rect 31612 4844 31668 4900
rect 31724 5010 31780 5012
rect 31724 4958 31726 5010
rect 31726 4958 31778 5010
rect 31778 4958 31780 5010
rect 31724 4956 31780 4958
rect 29932 3778 29988 3780
rect 29932 3726 29934 3778
rect 29934 3726 29986 3778
rect 29986 3726 29988 3778
rect 29932 3724 29988 3726
rect 29036 3500 29092 3556
rect 29372 3612 29428 3668
rect 30604 3778 30660 3780
rect 30604 3726 30606 3778
rect 30606 3726 30658 3778
rect 30658 3726 30660 3778
rect 30604 3724 30660 3726
rect 31836 4844 31892 4900
rect 32172 4898 32228 4900
rect 32172 4846 32174 4898
rect 32174 4846 32226 4898
rect 32226 4846 32228 4898
rect 32172 4844 32228 4846
rect 33846 5514 33902 5516
rect 33846 5462 33848 5514
rect 33848 5462 33900 5514
rect 33900 5462 33902 5514
rect 33846 5460 33902 5462
rect 33950 5514 34006 5516
rect 33950 5462 33952 5514
rect 33952 5462 34004 5514
rect 34004 5462 34006 5514
rect 33950 5460 34006 5462
rect 34054 5514 34110 5516
rect 34054 5462 34056 5514
rect 34056 5462 34108 5514
rect 34108 5462 34110 5514
rect 34054 5460 34110 5462
rect 33516 5010 33572 5012
rect 33516 4958 33518 5010
rect 33518 4958 33570 5010
rect 33570 4958 33572 5010
rect 33516 4956 33572 4958
rect 34412 4956 34468 5012
rect 32620 4898 32676 4900
rect 32620 4846 32622 4898
rect 32622 4846 32674 4898
rect 32674 4846 32676 4898
rect 32620 4844 32676 4846
rect 30044 3554 30100 3556
rect 30044 3502 30046 3554
rect 30046 3502 30098 3554
rect 30098 3502 30100 3554
rect 30044 3500 30100 3502
rect 30716 3554 30772 3556
rect 30716 3502 30718 3554
rect 30718 3502 30770 3554
rect 30770 3502 30772 3554
rect 30716 3500 30772 3502
rect 31948 3554 32004 3556
rect 31948 3502 31950 3554
rect 31950 3502 32002 3554
rect 32002 3502 32004 3554
rect 31948 3500 32004 3502
rect 32396 4338 32452 4340
rect 32396 4286 32398 4338
rect 32398 4286 32450 4338
rect 32450 4286 32452 4338
rect 32396 4284 32452 4286
rect 31388 3388 31444 3444
rect 33068 4898 33124 4900
rect 33068 4846 33070 4898
rect 33070 4846 33122 4898
rect 33122 4846 33124 4898
rect 33068 4844 33124 4846
rect 33964 4898 34020 4900
rect 33964 4846 33966 4898
rect 33966 4846 34018 4898
rect 34018 4846 34020 4898
rect 33964 4844 34020 4846
rect 33068 4284 33124 4340
rect 32620 4172 32676 4228
rect 33516 4226 33572 4228
rect 33516 4174 33518 4226
rect 33518 4174 33570 4226
rect 33570 4174 33572 4226
rect 33516 4172 33572 4174
rect 33964 4226 34020 4228
rect 33964 4174 33966 4226
rect 33966 4174 34018 4226
rect 34018 4174 34020 4226
rect 33964 4172 34020 4174
rect 34860 4844 34916 4900
rect 35308 4844 35364 4900
rect 32060 3442 32116 3444
rect 32060 3390 32062 3442
rect 32062 3390 32114 3442
rect 32114 3390 32116 3442
rect 32060 3388 32116 3390
rect 29184 3162 29240 3164
rect 29184 3110 29186 3162
rect 29186 3110 29238 3162
rect 29238 3110 29240 3162
rect 29184 3108 29240 3110
rect 29288 3162 29344 3164
rect 29288 3110 29290 3162
rect 29290 3110 29342 3162
rect 29342 3110 29344 3162
rect 29288 3108 29344 3110
rect 29392 3162 29448 3164
rect 29392 3110 29394 3162
rect 29394 3110 29446 3162
rect 29446 3110 29448 3162
rect 29392 3108 29448 3110
rect 33846 3946 33902 3948
rect 33846 3894 33848 3946
rect 33848 3894 33900 3946
rect 33900 3894 33902 3946
rect 33846 3892 33902 3894
rect 33950 3946 34006 3948
rect 33950 3894 33952 3946
rect 33952 3894 34004 3946
rect 34004 3894 34006 3946
rect 33950 3892 34006 3894
rect 34054 3946 34110 3948
rect 34054 3894 34056 3946
rect 34056 3894 34108 3946
rect 34108 3894 34110 3946
rect 34054 3892 34110 3894
rect 34412 3666 34468 3668
rect 34412 3614 34414 3666
rect 34414 3614 34466 3666
rect 34466 3614 34468 3666
rect 34412 3612 34468 3614
rect 32508 3388 32564 3444
rect 33292 3442 33348 3444
rect 33292 3390 33294 3442
rect 33294 3390 33346 3442
rect 33346 3390 33348 3442
rect 33292 3388 33348 3390
rect 33964 3442 34020 3444
rect 33964 3390 33966 3442
rect 33966 3390 34018 3442
rect 34018 3390 34020 3442
rect 33964 3388 34020 3390
rect 34860 4172 34916 4228
rect 38508 4730 38564 4732
rect 38508 4678 38510 4730
rect 38510 4678 38562 4730
rect 38562 4678 38564 4730
rect 38508 4676 38564 4678
rect 38612 4730 38668 4732
rect 38612 4678 38614 4730
rect 38614 4678 38666 4730
rect 38666 4678 38668 4730
rect 38612 4676 38668 4678
rect 38716 4730 38772 4732
rect 38716 4678 38718 4730
rect 38718 4678 38770 4730
rect 38770 4678 38772 4730
rect 38716 4676 38772 4678
rect 34524 3388 34580 3444
rect 35756 3442 35812 3444
rect 35756 3390 35758 3442
rect 35758 3390 35810 3442
rect 35810 3390 35812 3442
rect 35756 3388 35812 3390
rect 37212 3388 37268 3444
rect 38508 3162 38564 3164
rect 38508 3110 38510 3162
rect 38510 3110 38562 3162
rect 38562 3110 38564 3162
rect 38508 3108 38564 3110
rect 38612 3162 38668 3164
rect 38612 3110 38614 3162
rect 38614 3110 38666 3162
rect 38666 3110 38668 3162
rect 38612 3108 38668 3110
rect 38716 3162 38772 3164
rect 38716 3110 38718 3162
rect 38718 3110 38770 3162
rect 38770 3110 38772 3162
rect 38716 3108 38772 3110
<< metal3 >>
rect 5864 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6148 36876
rect 15188 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15472 36876
rect 24512 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24796 36876
rect 33836 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34120 36876
rect 10526 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10810 36092
rect 19850 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20134 36092
rect 29174 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29458 36092
rect 38498 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38782 36092
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 10526 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10810 34524
rect 19850 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20134 34524
rect 29174 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29458 34524
rect 38498 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38782 34524
rect 5864 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6148 33740
rect 15188 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15472 33740
rect 24512 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24796 33740
rect 33836 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34120 33740
rect 10526 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10810 32956
rect 19850 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20134 32956
rect 29174 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29458 32956
rect 38498 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38782 32956
rect 5864 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6148 32172
rect 15188 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15472 32172
rect 24512 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24796 32172
rect 33836 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34120 32172
rect 10526 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10810 31388
rect 19850 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20134 31388
rect 29174 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29458 31388
rect 38498 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38782 31388
rect 5864 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6148 30604
rect 15188 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15472 30604
rect 24512 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24796 30604
rect 33836 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34120 30604
rect 10526 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10810 29820
rect 19850 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20134 29820
rect 29174 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29458 29820
rect 38498 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38782 29820
rect 5864 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6148 29036
rect 15188 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15472 29036
rect 24512 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24796 29036
rect 33836 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34120 29036
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 5864 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6148 27468
rect 15188 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15472 27468
rect 24512 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24796 27468
rect 33836 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34120 27468
rect 10526 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10810 26684
rect 19850 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20134 26684
rect 29174 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29458 26684
rect 38498 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38782 26684
rect 5864 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6148 25900
rect 15188 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15472 25900
rect 24512 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24796 25900
rect 33836 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34120 25900
rect 10526 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10810 25116
rect 19850 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20134 25116
rect 29174 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29458 25116
rect 38498 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38782 25116
rect 5864 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6148 24332
rect 15188 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15472 24332
rect 24512 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24796 24332
rect 33836 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34120 24332
rect 10526 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10810 23548
rect 19850 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20134 23548
rect 29174 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29458 23548
rect 38498 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38782 23548
rect 5864 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6148 22764
rect 15188 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15472 22764
rect 24512 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24796 22764
rect 33836 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34120 22764
rect 10526 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10810 21980
rect 19850 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20134 21980
rect 29174 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29458 21980
rect 38498 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38782 21980
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 10526 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10810 20412
rect 19850 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20134 20412
rect 29174 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29458 20412
rect 38498 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38782 20412
rect 5864 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6148 19628
rect 15188 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15472 19628
rect 24512 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24796 19628
rect 33836 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34120 19628
rect 10526 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10810 18844
rect 19850 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20134 18844
rect 29174 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29458 18844
rect 38498 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38782 18844
rect 5864 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6148 18060
rect 15188 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15472 18060
rect 24512 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24796 18060
rect 33836 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34120 18060
rect 10526 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10810 17276
rect 19850 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20134 17276
rect 29174 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29458 17276
rect 38498 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38782 17276
rect 5864 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6148 16492
rect 15188 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15472 16492
rect 24512 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24796 16492
rect 33836 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34120 16492
rect 10526 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10810 15708
rect 19850 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20134 15708
rect 29174 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29458 15708
rect 38498 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38782 15708
rect 5864 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6148 14924
rect 15188 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15472 14924
rect 24512 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24796 14924
rect 33836 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34120 14924
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 5864 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6148 13356
rect 15188 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15472 13356
rect 24512 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24796 13356
rect 33836 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34120 13356
rect 10526 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10810 12572
rect 19850 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20134 12572
rect 29174 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29458 12572
rect 38498 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38782 12572
rect 5864 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6148 11788
rect 15188 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15472 11788
rect 24512 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24796 11788
rect 33836 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34120 11788
rect 10526 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10810 11004
rect 19850 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20134 11004
rect 29174 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29458 11004
rect 38498 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38782 11004
rect 5864 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6148 10220
rect 15188 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15472 10220
rect 24512 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24796 10220
rect 33836 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34120 10220
rect 10526 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10810 9436
rect 19850 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20134 9436
rect 29174 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29458 9436
rect 38498 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38782 9436
rect 24210 8876 24220 8932
rect 24276 8876 25676 8932
rect 25732 8876 26124 8932
rect 26180 8876 26572 8932
rect 26628 8876 26908 8932
rect 26964 8876 26974 8932
rect 5864 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6148 8652
rect 15188 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15472 8652
rect 24512 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24796 8652
rect 33836 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34120 8652
rect 23202 7980 23212 8036
rect 23268 7980 24220 8036
rect 24276 7980 24286 8036
rect 24434 7980 24444 8036
rect 24500 7980 25340 8036
rect 25396 7980 25406 8036
rect 27346 7980 27356 8036
rect 27412 7980 28252 8036
rect 28308 7980 28700 8036
rect 28756 7980 28766 8036
rect 10526 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10810 7868
rect 19850 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20134 7868
rect 29174 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29458 7868
rect 38498 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38782 7868
rect 25554 7308 25564 7364
rect 25620 7308 26012 7364
rect 26068 7308 26908 7364
rect 26964 7308 26974 7364
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 19618 6748 19628 6804
rect 19684 6748 21980 6804
rect 22036 6748 22046 6804
rect 26226 6748 26236 6804
rect 26292 6748 26460 6804
rect 26516 6748 27468 6804
rect 27524 6748 28812 6804
rect 28868 6748 30044 6804
rect 30100 6748 30996 6804
rect 30940 6692 30996 6748
rect 30930 6636 30940 6692
rect 30996 6636 31006 6692
rect 28578 6524 28588 6580
rect 28644 6524 29596 6580
rect 29652 6524 30156 6580
rect 30212 6524 30222 6580
rect 22978 6412 22988 6468
rect 23044 6412 23660 6468
rect 23716 6412 23726 6468
rect 24994 6412 25004 6468
rect 25060 6412 25676 6468
rect 25732 6412 26460 6468
rect 26516 6412 27020 6468
rect 27076 6412 28364 6468
rect 28420 6412 29036 6468
rect 29092 6412 29102 6468
rect 10526 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10810 6300
rect 19850 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20134 6300
rect 29174 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29458 6300
rect 38498 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38782 6300
rect 25778 6076 25788 6132
rect 25844 6076 26348 6132
rect 26404 6076 27804 6132
rect 27860 6076 28252 6132
rect 28308 6076 28318 6132
rect 21410 5852 21420 5908
rect 21476 5852 21980 5908
rect 22036 5852 22046 5908
rect 21980 5684 22036 5852
rect 21980 5628 22764 5684
rect 22820 5628 23212 5684
rect 23268 5628 23436 5684
rect 23492 5628 24108 5684
rect 24164 5628 24174 5684
rect 5864 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6148 5516
rect 15188 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15472 5516
rect 24512 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24796 5516
rect 33836 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34120 5516
rect 24322 5068 24332 5124
rect 24388 5068 25116 5124
rect 25172 5068 25676 5124
rect 25732 5068 25742 5124
rect 31826 5068 31836 5124
rect 31892 5012 31948 5124
rect 23986 4956 23996 5012
rect 24052 4956 24780 5012
rect 24836 4956 24846 5012
rect 29810 4956 29820 5012
rect 29876 4956 30380 5012
rect 30436 4956 31052 5012
rect 31108 4956 31500 5012
rect 31556 4956 31724 5012
rect 31780 4956 31790 5012
rect 31892 4956 32228 5012
rect 33506 4956 33516 5012
rect 33572 4956 34412 5012
rect 34468 4956 34478 5012
rect 32172 4900 32228 4956
rect 27122 4844 27132 4900
rect 27188 4844 27692 4900
rect 27748 4844 27758 4900
rect 31154 4844 31164 4900
rect 31220 4844 31612 4900
rect 31668 4844 31836 4900
rect 31892 4844 31902 4900
rect 32162 4844 32172 4900
rect 32228 4844 32620 4900
rect 32676 4844 32686 4900
rect 33058 4844 33068 4900
rect 33124 4844 33964 4900
rect 34020 4844 34860 4900
rect 34916 4844 35308 4900
rect 35364 4844 35374 4900
rect 10526 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10810 4732
rect 19850 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20134 4732
rect 29174 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29458 4732
rect 38498 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38782 4732
rect 18834 4508 18844 4564
rect 18900 4508 19180 4564
rect 19236 4508 20188 4564
rect 20244 4508 20254 4564
rect 27234 4508 27244 4564
rect 27300 4508 27804 4564
rect 27860 4508 28476 4564
rect 28532 4508 28542 4564
rect 29138 4508 29148 4564
rect 29204 4508 29820 4564
rect 29876 4508 29886 4564
rect 28476 4452 28532 4508
rect 21522 4396 21532 4452
rect 21588 4396 22204 4452
rect 22260 4396 22270 4452
rect 28476 4396 29260 4452
rect 29316 4396 29326 4452
rect 23538 4284 23548 4340
rect 23604 4284 24220 4340
rect 24276 4284 25340 4340
rect 25396 4284 25676 4340
rect 25732 4284 25742 4340
rect 29026 4284 29036 4340
rect 29092 4284 29708 4340
rect 29764 4284 29774 4340
rect 32386 4284 32396 4340
rect 32452 4284 33068 4340
rect 33124 4284 33134 4340
rect 32610 4172 32620 4228
rect 32676 4172 33516 4228
rect 33572 4172 33964 4228
rect 34020 4172 34860 4228
rect 34916 4172 34926 4228
rect 19282 4060 19292 4116
rect 19348 4060 20300 4116
rect 20356 4060 21420 4116
rect 21476 4060 21486 4116
rect 27122 4060 27132 4116
rect 27188 4060 27692 4116
rect 27748 4060 27758 4116
rect 5864 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6148 3948
rect 15188 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15472 3948
rect 24512 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24796 3948
rect 33836 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34120 3948
rect 16594 3724 16604 3780
rect 16660 3724 27244 3780
rect 27300 3724 27310 3780
rect 29922 3724 29932 3780
rect 29988 3724 30604 3780
rect 30660 3724 30670 3780
rect 20178 3612 20188 3668
rect 20244 3612 20636 3668
rect 20692 3612 20972 3668
rect 21028 3612 21644 3668
rect 21700 3612 22316 3668
rect 22372 3612 22988 3668
rect 23044 3612 23660 3668
rect 23716 3612 24332 3668
rect 24388 3612 24398 3668
rect 27682 3612 27692 3668
rect 27748 3612 28028 3668
rect 28084 3612 28364 3668
rect 28420 3612 29372 3668
rect 29428 3612 34412 3668
rect 34468 3612 34478 3668
rect 12562 3500 12572 3556
rect 12628 3500 17724 3556
rect 17780 3500 18172 3556
rect 18228 3500 18620 3556
rect 18676 3500 19628 3556
rect 19684 3500 19852 3556
rect 19908 3500 20524 3556
rect 20580 3500 21532 3556
rect 21588 3500 21598 3556
rect 22194 3500 22204 3556
rect 22260 3500 22876 3556
rect 22932 3500 23548 3556
rect 23604 3500 23614 3556
rect 25330 3500 25340 3556
rect 25396 3500 26012 3556
rect 26068 3500 26684 3556
rect 26740 3500 26750 3556
rect 27458 3500 27468 3556
rect 27524 3500 28140 3556
rect 28196 3500 29036 3556
rect 29092 3500 30044 3556
rect 30100 3500 30716 3556
rect 30772 3500 30782 3556
rect 31938 3500 31948 3556
rect 32004 3500 32564 3556
rect 32508 3444 32564 3500
rect 2706 3388 2716 3444
rect 2772 3388 16044 3444
rect 16100 3388 16492 3444
rect 16548 3388 16558 3444
rect 31378 3388 31388 3444
rect 31444 3388 32060 3444
rect 32116 3388 32126 3444
rect 32498 3388 32508 3444
rect 32564 3388 33292 3444
rect 33348 3388 33964 3444
rect 34020 3388 34524 3444
rect 34580 3388 35756 3444
rect 35812 3388 37212 3444
rect 37268 3388 37278 3444
rect 10526 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10810 3164
rect 19850 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20134 3164
rect 29174 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29458 3164
rect 38498 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38782 3164
<< via3 >>
rect 5874 36820 5930 36876
rect 5978 36820 6034 36876
rect 6082 36820 6138 36876
rect 15198 36820 15254 36876
rect 15302 36820 15358 36876
rect 15406 36820 15462 36876
rect 24522 36820 24578 36876
rect 24626 36820 24682 36876
rect 24730 36820 24786 36876
rect 33846 36820 33902 36876
rect 33950 36820 34006 36876
rect 34054 36820 34110 36876
rect 10536 36036 10592 36092
rect 10640 36036 10696 36092
rect 10744 36036 10800 36092
rect 19860 36036 19916 36092
rect 19964 36036 20020 36092
rect 20068 36036 20124 36092
rect 29184 36036 29240 36092
rect 29288 36036 29344 36092
rect 29392 36036 29448 36092
rect 38508 36036 38564 36092
rect 38612 36036 38668 36092
rect 38716 36036 38772 36092
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 10536 34468 10592 34524
rect 10640 34468 10696 34524
rect 10744 34468 10800 34524
rect 19860 34468 19916 34524
rect 19964 34468 20020 34524
rect 20068 34468 20124 34524
rect 29184 34468 29240 34524
rect 29288 34468 29344 34524
rect 29392 34468 29448 34524
rect 38508 34468 38564 34524
rect 38612 34468 38668 34524
rect 38716 34468 38772 34524
rect 5874 33684 5930 33740
rect 5978 33684 6034 33740
rect 6082 33684 6138 33740
rect 15198 33684 15254 33740
rect 15302 33684 15358 33740
rect 15406 33684 15462 33740
rect 24522 33684 24578 33740
rect 24626 33684 24682 33740
rect 24730 33684 24786 33740
rect 33846 33684 33902 33740
rect 33950 33684 34006 33740
rect 34054 33684 34110 33740
rect 10536 32900 10592 32956
rect 10640 32900 10696 32956
rect 10744 32900 10800 32956
rect 19860 32900 19916 32956
rect 19964 32900 20020 32956
rect 20068 32900 20124 32956
rect 29184 32900 29240 32956
rect 29288 32900 29344 32956
rect 29392 32900 29448 32956
rect 38508 32900 38564 32956
rect 38612 32900 38668 32956
rect 38716 32900 38772 32956
rect 5874 32116 5930 32172
rect 5978 32116 6034 32172
rect 6082 32116 6138 32172
rect 15198 32116 15254 32172
rect 15302 32116 15358 32172
rect 15406 32116 15462 32172
rect 24522 32116 24578 32172
rect 24626 32116 24682 32172
rect 24730 32116 24786 32172
rect 33846 32116 33902 32172
rect 33950 32116 34006 32172
rect 34054 32116 34110 32172
rect 10536 31332 10592 31388
rect 10640 31332 10696 31388
rect 10744 31332 10800 31388
rect 19860 31332 19916 31388
rect 19964 31332 20020 31388
rect 20068 31332 20124 31388
rect 29184 31332 29240 31388
rect 29288 31332 29344 31388
rect 29392 31332 29448 31388
rect 38508 31332 38564 31388
rect 38612 31332 38668 31388
rect 38716 31332 38772 31388
rect 5874 30548 5930 30604
rect 5978 30548 6034 30604
rect 6082 30548 6138 30604
rect 15198 30548 15254 30604
rect 15302 30548 15358 30604
rect 15406 30548 15462 30604
rect 24522 30548 24578 30604
rect 24626 30548 24682 30604
rect 24730 30548 24786 30604
rect 33846 30548 33902 30604
rect 33950 30548 34006 30604
rect 34054 30548 34110 30604
rect 10536 29764 10592 29820
rect 10640 29764 10696 29820
rect 10744 29764 10800 29820
rect 19860 29764 19916 29820
rect 19964 29764 20020 29820
rect 20068 29764 20124 29820
rect 29184 29764 29240 29820
rect 29288 29764 29344 29820
rect 29392 29764 29448 29820
rect 38508 29764 38564 29820
rect 38612 29764 38668 29820
rect 38716 29764 38772 29820
rect 5874 28980 5930 29036
rect 5978 28980 6034 29036
rect 6082 28980 6138 29036
rect 15198 28980 15254 29036
rect 15302 28980 15358 29036
rect 15406 28980 15462 29036
rect 24522 28980 24578 29036
rect 24626 28980 24682 29036
rect 24730 28980 24786 29036
rect 33846 28980 33902 29036
rect 33950 28980 34006 29036
rect 34054 28980 34110 29036
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 5874 27412 5930 27468
rect 5978 27412 6034 27468
rect 6082 27412 6138 27468
rect 15198 27412 15254 27468
rect 15302 27412 15358 27468
rect 15406 27412 15462 27468
rect 24522 27412 24578 27468
rect 24626 27412 24682 27468
rect 24730 27412 24786 27468
rect 33846 27412 33902 27468
rect 33950 27412 34006 27468
rect 34054 27412 34110 27468
rect 10536 26628 10592 26684
rect 10640 26628 10696 26684
rect 10744 26628 10800 26684
rect 19860 26628 19916 26684
rect 19964 26628 20020 26684
rect 20068 26628 20124 26684
rect 29184 26628 29240 26684
rect 29288 26628 29344 26684
rect 29392 26628 29448 26684
rect 38508 26628 38564 26684
rect 38612 26628 38668 26684
rect 38716 26628 38772 26684
rect 5874 25844 5930 25900
rect 5978 25844 6034 25900
rect 6082 25844 6138 25900
rect 15198 25844 15254 25900
rect 15302 25844 15358 25900
rect 15406 25844 15462 25900
rect 24522 25844 24578 25900
rect 24626 25844 24682 25900
rect 24730 25844 24786 25900
rect 33846 25844 33902 25900
rect 33950 25844 34006 25900
rect 34054 25844 34110 25900
rect 10536 25060 10592 25116
rect 10640 25060 10696 25116
rect 10744 25060 10800 25116
rect 19860 25060 19916 25116
rect 19964 25060 20020 25116
rect 20068 25060 20124 25116
rect 29184 25060 29240 25116
rect 29288 25060 29344 25116
rect 29392 25060 29448 25116
rect 38508 25060 38564 25116
rect 38612 25060 38668 25116
rect 38716 25060 38772 25116
rect 5874 24276 5930 24332
rect 5978 24276 6034 24332
rect 6082 24276 6138 24332
rect 15198 24276 15254 24332
rect 15302 24276 15358 24332
rect 15406 24276 15462 24332
rect 24522 24276 24578 24332
rect 24626 24276 24682 24332
rect 24730 24276 24786 24332
rect 33846 24276 33902 24332
rect 33950 24276 34006 24332
rect 34054 24276 34110 24332
rect 10536 23492 10592 23548
rect 10640 23492 10696 23548
rect 10744 23492 10800 23548
rect 19860 23492 19916 23548
rect 19964 23492 20020 23548
rect 20068 23492 20124 23548
rect 29184 23492 29240 23548
rect 29288 23492 29344 23548
rect 29392 23492 29448 23548
rect 38508 23492 38564 23548
rect 38612 23492 38668 23548
rect 38716 23492 38772 23548
rect 5874 22708 5930 22764
rect 5978 22708 6034 22764
rect 6082 22708 6138 22764
rect 15198 22708 15254 22764
rect 15302 22708 15358 22764
rect 15406 22708 15462 22764
rect 24522 22708 24578 22764
rect 24626 22708 24682 22764
rect 24730 22708 24786 22764
rect 33846 22708 33902 22764
rect 33950 22708 34006 22764
rect 34054 22708 34110 22764
rect 10536 21924 10592 21980
rect 10640 21924 10696 21980
rect 10744 21924 10800 21980
rect 19860 21924 19916 21980
rect 19964 21924 20020 21980
rect 20068 21924 20124 21980
rect 29184 21924 29240 21980
rect 29288 21924 29344 21980
rect 29392 21924 29448 21980
rect 38508 21924 38564 21980
rect 38612 21924 38668 21980
rect 38716 21924 38772 21980
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20356 10592 20412
rect 10640 20356 10696 20412
rect 10744 20356 10800 20412
rect 19860 20356 19916 20412
rect 19964 20356 20020 20412
rect 20068 20356 20124 20412
rect 29184 20356 29240 20412
rect 29288 20356 29344 20412
rect 29392 20356 29448 20412
rect 38508 20356 38564 20412
rect 38612 20356 38668 20412
rect 38716 20356 38772 20412
rect 5874 19572 5930 19628
rect 5978 19572 6034 19628
rect 6082 19572 6138 19628
rect 15198 19572 15254 19628
rect 15302 19572 15358 19628
rect 15406 19572 15462 19628
rect 24522 19572 24578 19628
rect 24626 19572 24682 19628
rect 24730 19572 24786 19628
rect 33846 19572 33902 19628
rect 33950 19572 34006 19628
rect 34054 19572 34110 19628
rect 10536 18788 10592 18844
rect 10640 18788 10696 18844
rect 10744 18788 10800 18844
rect 19860 18788 19916 18844
rect 19964 18788 20020 18844
rect 20068 18788 20124 18844
rect 29184 18788 29240 18844
rect 29288 18788 29344 18844
rect 29392 18788 29448 18844
rect 38508 18788 38564 18844
rect 38612 18788 38668 18844
rect 38716 18788 38772 18844
rect 5874 18004 5930 18060
rect 5978 18004 6034 18060
rect 6082 18004 6138 18060
rect 15198 18004 15254 18060
rect 15302 18004 15358 18060
rect 15406 18004 15462 18060
rect 24522 18004 24578 18060
rect 24626 18004 24682 18060
rect 24730 18004 24786 18060
rect 33846 18004 33902 18060
rect 33950 18004 34006 18060
rect 34054 18004 34110 18060
rect 10536 17220 10592 17276
rect 10640 17220 10696 17276
rect 10744 17220 10800 17276
rect 19860 17220 19916 17276
rect 19964 17220 20020 17276
rect 20068 17220 20124 17276
rect 29184 17220 29240 17276
rect 29288 17220 29344 17276
rect 29392 17220 29448 17276
rect 38508 17220 38564 17276
rect 38612 17220 38668 17276
rect 38716 17220 38772 17276
rect 5874 16436 5930 16492
rect 5978 16436 6034 16492
rect 6082 16436 6138 16492
rect 15198 16436 15254 16492
rect 15302 16436 15358 16492
rect 15406 16436 15462 16492
rect 24522 16436 24578 16492
rect 24626 16436 24682 16492
rect 24730 16436 24786 16492
rect 33846 16436 33902 16492
rect 33950 16436 34006 16492
rect 34054 16436 34110 16492
rect 10536 15652 10592 15708
rect 10640 15652 10696 15708
rect 10744 15652 10800 15708
rect 19860 15652 19916 15708
rect 19964 15652 20020 15708
rect 20068 15652 20124 15708
rect 29184 15652 29240 15708
rect 29288 15652 29344 15708
rect 29392 15652 29448 15708
rect 38508 15652 38564 15708
rect 38612 15652 38668 15708
rect 38716 15652 38772 15708
rect 5874 14868 5930 14924
rect 5978 14868 6034 14924
rect 6082 14868 6138 14924
rect 15198 14868 15254 14924
rect 15302 14868 15358 14924
rect 15406 14868 15462 14924
rect 24522 14868 24578 14924
rect 24626 14868 24682 14924
rect 24730 14868 24786 14924
rect 33846 14868 33902 14924
rect 33950 14868 34006 14924
rect 34054 14868 34110 14924
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 5874 13300 5930 13356
rect 5978 13300 6034 13356
rect 6082 13300 6138 13356
rect 15198 13300 15254 13356
rect 15302 13300 15358 13356
rect 15406 13300 15462 13356
rect 24522 13300 24578 13356
rect 24626 13300 24682 13356
rect 24730 13300 24786 13356
rect 33846 13300 33902 13356
rect 33950 13300 34006 13356
rect 34054 13300 34110 13356
rect 10536 12516 10592 12572
rect 10640 12516 10696 12572
rect 10744 12516 10800 12572
rect 19860 12516 19916 12572
rect 19964 12516 20020 12572
rect 20068 12516 20124 12572
rect 29184 12516 29240 12572
rect 29288 12516 29344 12572
rect 29392 12516 29448 12572
rect 38508 12516 38564 12572
rect 38612 12516 38668 12572
rect 38716 12516 38772 12572
rect 5874 11732 5930 11788
rect 5978 11732 6034 11788
rect 6082 11732 6138 11788
rect 15198 11732 15254 11788
rect 15302 11732 15358 11788
rect 15406 11732 15462 11788
rect 24522 11732 24578 11788
rect 24626 11732 24682 11788
rect 24730 11732 24786 11788
rect 33846 11732 33902 11788
rect 33950 11732 34006 11788
rect 34054 11732 34110 11788
rect 10536 10948 10592 11004
rect 10640 10948 10696 11004
rect 10744 10948 10800 11004
rect 19860 10948 19916 11004
rect 19964 10948 20020 11004
rect 20068 10948 20124 11004
rect 29184 10948 29240 11004
rect 29288 10948 29344 11004
rect 29392 10948 29448 11004
rect 38508 10948 38564 11004
rect 38612 10948 38668 11004
rect 38716 10948 38772 11004
rect 5874 10164 5930 10220
rect 5978 10164 6034 10220
rect 6082 10164 6138 10220
rect 15198 10164 15254 10220
rect 15302 10164 15358 10220
rect 15406 10164 15462 10220
rect 24522 10164 24578 10220
rect 24626 10164 24682 10220
rect 24730 10164 24786 10220
rect 33846 10164 33902 10220
rect 33950 10164 34006 10220
rect 34054 10164 34110 10220
rect 10536 9380 10592 9436
rect 10640 9380 10696 9436
rect 10744 9380 10800 9436
rect 19860 9380 19916 9436
rect 19964 9380 20020 9436
rect 20068 9380 20124 9436
rect 29184 9380 29240 9436
rect 29288 9380 29344 9436
rect 29392 9380 29448 9436
rect 38508 9380 38564 9436
rect 38612 9380 38668 9436
rect 38716 9380 38772 9436
rect 5874 8596 5930 8652
rect 5978 8596 6034 8652
rect 6082 8596 6138 8652
rect 15198 8596 15254 8652
rect 15302 8596 15358 8652
rect 15406 8596 15462 8652
rect 24522 8596 24578 8652
rect 24626 8596 24682 8652
rect 24730 8596 24786 8652
rect 33846 8596 33902 8652
rect 33950 8596 34006 8652
rect 34054 8596 34110 8652
rect 10536 7812 10592 7868
rect 10640 7812 10696 7868
rect 10744 7812 10800 7868
rect 19860 7812 19916 7868
rect 19964 7812 20020 7868
rect 20068 7812 20124 7868
rect 29184 7812 29240 7868
rect 29288 7812 29344 7868
rect 29392 7812 29448 7868
rect 38508 7812 38564 7868
rect 38612 7812 38668 7868
rect 38716 7812 38772 7868
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6244 10592 6300
rect 10640 6244 10696 6300
rect 10744 6244 10800 6300
rect 19860 6244 19916 6300
rect 19964 6244 20020 6300
rect 20068 6244 20124 6300
rect 29184 6244 29240 6300
rect 29288 6244 29344 6300
rect 29392 6244 29448 6300
rect 38508 6244 38564 6300
rect 38612 6244 38668 6300
rect 38716 6244 38772 6300
rect 5874 5460 5930 5516
rect 5978 5460 6034 5516
rect 6082 5460 6138 5516
rect 15198 5460 15254 5516
rect 15302 5460 15358 5516
rect 15406 5460 15462 5516
rect 24522 5460 24578 5516
rect 24626 5460 24682 5516
rect 24730 5460 24786 5516
rect 33846 5460 33902 5516
rect 33950 5460 34006 5516
rect 34054 5460 34110 5516
rect 10536 4676 10592 4732
rect 10640 4676 10696 4732
rect 10744 4676 10800 4732
rect 19860 4676 19916 4732
rect 19964 4676 20020 4732
rect 20068 4676 20124 4732
rect 29184 4676 29240 4732
rect 29288 4676 29344 4732
rect 29392 4676 29448 4732
rect 38508 4676 38564 4732
rect 38612 4676 38668 4732
rect 38716 4676 38772 4732
rect 5874 3892 5930 3948
rect 5978 3892 6034 3948
rect 6082 3892 6138 3948
rect 15198 3892 15254 3948
rect 15302 3892 15358 3948
rect 15406 3892 15462 3948
rect 24522 3892 24578 3948
rect 24626 3892 24682 3948
rect 24730 3892 24786 3948
rect 33846 3892 33902 3948
rect 33950 3892 34006 3948
rect 34054 3892 34110 3948
rect 10536 3108 10592 3164
rect 10640 3108 10696 3164
rect 10744 3108 10800 3164
rect 19860 3108 19916 3164
rect 19964 3108 20020 3164
rect 20068 3108 20124 3164
rect 29184 3108 29240 3164
rect 29288 3108 29344 3164
rect 29392 3108 29448 3164
rect 38508 3108 38564 3164
rect 38612 3108 38668 3164
rect 38716 3108 38772 3164
<< metal4 >>
rect 5846 36876 6166 36908
rect 5846 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6166 36876
rect 5846 35308 6166 36820
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33740 6166 35252
rect 5846 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6166 33740
rect 5846 32172 6166 33684
rect 5846 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6166 32172
rect 5846 30604 6166 32116
rect 5846 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6166 30604
rect 5846 29036 6166 30548
rect 5846 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6166 29036
rect 5846 27468 6166 28980
rect 5846 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6166 27468
rect 5846 25900 6166 27412
rect 5846 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6166 25900
rect 5846 24332 6166 25844
rect 5846 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6166 24332
rect 5846 22764 6166 24276
rect 5846 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6166 22764
rect 5846 21196 6166 22708
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19628 6166 21140
rect 5846 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6166 19628
rect 5846 18060 6166 19572
rect 5846 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6166 18060
rect 5846 16492 6166 18004
rect 5846 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6166 16492
rect 5846 14924 6166 16436
rect 5846 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6166 14924
rect 5846 13356 6166 14868
rect 5846 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6166 13356
rect 5846 11788 6166 13300
rect 5846 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6166 11788
rect 5846 10220 6166 11732
rect 5846 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6166 10220
rect 5846 8652 6166 10164
rect 5846 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6166 8652
rect 5846 7084 6166 8596
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5516 6166 7028
rect 5846 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6166 5516
rect 5846 3948 6166 5460
rect 5846 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6166 3948
rect 5846 3076 6166 3892
rect 10508 36092 10828 36908
rect 10508 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10828 36092
rect 10508 34524 10828 36036
rect 10508 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10828 34524
rect 10508 32956 10828 34468
rect 10508 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10828 32956
rect 10508 31388 10828 32900
rect 10508 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10828 31388
rect 10508 29820 10828 31332
rect 10508 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10828 29820
rect 10508 28252 10828 29764
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26684 10828 28196
rect 10508 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10828 26684
rect 10508 25116 10828 26628
rect 10508 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10828 25116
rect 10508 23548 10828 25060
rect 10508 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10828 23548
rect 10508 21980 10828 23492
rect 10508 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10828 21980
rect 10508 20412 10828 21924
rect 10508 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10828 20412
rect 10508 18844 10828 20356
rect 10508 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10828 18844
rect 10508 17276 10828 18788
rect 10508 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10828 17276
rect 10508 15708 10828 17220
rect 10508 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10828 15708
rect 10508 14140 10828 15652
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 10508 12572 10828 14084
rect 10508 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10828 12572
rect 10508 11004 10828 12516
rect 10508 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10828 11004
rect 10508 9436 10828 10948
rect 10508 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10828 9436
rect 10508 7868 10828 9380
rect 10508 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10828 7868
rect 10508 6300 10828 7812
rect 10508 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10828 6300
rect 10508 4732 10828 6244
rect 10508 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10828 4732
rect 10508 3164 10828 4676
rect 10508 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10828 3164
rect 10508 3076 10828 3108
rect 15170 36876 15490 36908
rect 15170 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15490 36876
rect 15170 35308 15490 36820
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33740 15490 35252
rect 15170 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15490 33740
rect 15170 32172 15490 33684
rect 15170 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15490 32172
rect 15170 30604 15490 32116
rect 15170 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15490 30604
rect 15170 29036 15490 30548
rect 15170 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15490 29036
rect 15170 27468 15490 28980
rect 15170 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15490 27468
rect 15170 25900 15490 27412
rect 15170 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15490 25900
rect 15170 24332 15490 25844
rect 15170 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15490 24332
rect 15170 22764 15490 24276
rect 15170 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15490 22764
rect 15170 21196 15490 22708
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19628 15490 21140
rect 15170 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15490 19628
rect 15170 18060 15490 19572
rect 15170 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15490 18060
rect 15170 16492 15490 18004
rect 15170 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15490 16492
rect 15170 14924 15490 16436
rect 15170 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15490 14924
rect 15170 13356 15490 14868
rect 15170 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15490 13356
rect 15170 11788 15490 13300
rect 15170 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15490 11788
rect 15170 10220 15490 11732
rect 15170 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15490 10220
rect 15170 8652 15490 10164
rect 15170 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15490 8652
rect 15170 7084 15490 8596
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5516 15490 7028
rect 15170 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15490 5516
rect 15170 3948 15490 5460
rect 15170 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15490 3948
rect 15170 3076 15490 3892
rect 19832 36092 20152 36908
rect 19832 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20152 36092
rect 19832 34524 20152 36036
rect 19832 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20152 34524
rect 19832 32956 20152 34468
rect 19832 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20152 32956
rect 19832 31388 20152 32900
rect 19832 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20152 31388
rect 19832 29820 20152 31332
rect 19832 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20152 29820
rect 19832 28252 20152 29764
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26684 20152 28196
rect 19832 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20152 26684
rect 19832 25116 20152 26628
rect 19832 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20152 25116
rect 19832 23548 20152 25060
rect 19832 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20152 23548
rect 19832 21980 20152 23492
rect 19832 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20152 21980
rect 19832 20412 20152 21924
rect 19832 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20152 20412
rect 19832 18844 20152 20356
rect 19832 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20152 18844
rect 19832 17276 20152 18788
rect 19832 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20152 17276
rect 19832 15708 20152 17220
rect 19832 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20152 15708
rect 19832 14140 20152 15652
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12572 20152 14084
rect 19832 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20152 12572
rect 19832 11004 20152 12516
rect 19832 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20152 11004
rect 19832 9436 20152 10948
rect 19832 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20152 9436
rect 19832 7868 20152 9380
rect 19832 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20152 7868
rect 19832 6300 20152 7812
rect 19832 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20152 6300
rect 19832 4732 20152 6244
rect 19832 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20152 4732
rect 19832 3164 20152 4676
rect 19832 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20152 3164
rect 19832 3076 20152 3108
rect 24494 36876 24814 36908
rect 24494 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24814 36876
rect 24494 35308 24814 36820
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33740 24814 35252
rect 24494 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24814 33740
rect 24494 32172 24814 33684
rect 24494 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24814 32172
rect 24494 30604 24814 32116
rect 24494 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24814 30604
rect 24494 29036 24814 30548
rect 24494 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24814 29036
rect 24494 27468 24814 28980
rect 24494 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24814 27468
rect 24494 25900 24814 27412
rect 24494 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24814 25900
rect 24494 24332 24814 25844
rect 24494 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24814 24332
rect 24494 22764 24814 24276
rect 24494 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24814 22764
rect 24494 21196 24814 22708
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19628 24814 21140
rect 24494 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24814 19628
rect 24494 18060 24814 19572
rect 24494 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24814 18060
rect 24494 16492 24814 18004
rect 24494 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24814 16492
rect 24494 14924 24814 16436
rect 24494 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24814 14924
rect 24494 13356 24814 14868
rect 24494 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24814 13356
rect 24494 11788 24814 13300
rect 24494 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24814 11788
rect 24494 10220 24814 11732
rect 24494 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24814 10220
rect 24494 8652 24814 10164
rect 24494 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24814 8652
rect 24494 7084 24814 8596
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5516 24814 7028
rect 24494 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24814 5516
rect 24494 3948 24814 5460
rect 24494 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24814 3948
rect 24494 3076 24814 3892
rect 29156 36092 29476 36908
rect 29156 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29476 36092
rect 29156 34524 29476 36036
rect 29156 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29476 34524
rect 29156 32956 29476 34468
rect 29156 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29476 32956
rect 29156 31388 29476 32900
rect 29156 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29476 31388
rect 29156 29820 29476 31332
rect 29156 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29476 29820
rect 29156 28252 29476 29764
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26684 29476 28196
rect 29156 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29476 26684
rect 29156 25116 29476 26628
rect 29156 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29476 25116
rect 29156 23548 29476 25060
rect 29156 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29476 23548
rect 29156 21980 29476 23492
rect 29156 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29476 21980
rect 29156 20412 29476 21924
rect 29156 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29476 20412
rect 29156 18844 29476 20356
rect 29156 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29476 18844
rect 29156 17276 29476 18788
rect 29156 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29476 17276
rect 29156 15708 29476 17220
rect 29156 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29476 15708
rect 29156 14140 29476 15652
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12572 29476 14084
rect 29156 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29476 12572
rect 29156 11004 29476 12516
rect 29156 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29476 11004
rect 29156 9436 29476 10948
rect 29156 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29476 9436
rect 29156 7868 29476 9380
rect 29156 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29476 7868
rect 29156 6300 29476 7812
rect 29156 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29476 6300
rect 29156 4732 29476 6244
rect 29156 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29476 4732
rect 29156 3164 29476 4676
rect 29156 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29476 3164
rect 29156 3076 29476 3108
rect 33818 36876 34138 36908
rect 33818 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34138 36876
rect 33818 35308 34138 36820
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33740 34138 35252
rect 33818 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34138 33740
rect 33818 32172 34138 33684
rect 33818 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34138 32172
rect 33818 30604 34138 32116
rect 33818 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34138 30604
rect 33818 29036 34138 30548
rect 33818 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34138 29036
rect 33818 27468 34138 28980
rect 33818 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34138 27468
rect 33818 25900 34138 27412
rect 33818 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34138 25900
rect 33818 24332 34138 25844
rect 33818 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34138 24332
rect 33818 22764 34138 24276
rect 33818 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34138 22764
rect 33818 21196 34138 22708
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19628 34138 21140
rect 33818 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34138 19628
rect 33818 18060 34138 19572
rect 33818 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34138 18060
rect 33818 16492 34138 18004
rect 33818 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34138 16492
rect 33818 14924 34138 16436
rect 33818 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34138 14924
rect 33818 13356 34138 14868
rect 33818 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34138 13356
rect 33818 11788 34138 13300
rect 33818 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34138 11788
rect 33818 10220 34138 11732
rect 33818 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34138 10220
rect 33818 8652 34138 10164
rect 33818 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34138 8652
rect 33818 7084 34138 8596
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5516 34138 7028
rect 33818 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34138 5516
rect 33818 3948 34138 5460
rect 33818 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34138 3948
rect 33818 3076 34138 3892
rect 38480 36092 38800 36908
rect 38480 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38800 36092
rect 38480 34524 38800 36036
rect 38480 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38800 34524
rect 38480 32956 38800 34468
rect 38480 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38800 32956
rect 38480 31388 38800 32900
rect 38480 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38800 31388
rect 38480 29820 38800 31332
rect 38480 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38800 29820
rect 38480 28252 38800 29764
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26684 38800 28196
rect 38480 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38800 26684
rect 38480 25116 38800 26628
rect 38480 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38800 25116
rect 38480 23548 38800 25060
rect 38480 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38800 23548
rect 38480 21980 38800 23492
rect 38480 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38800 21980
rect 38480 20412 38800 21924
rect 38480 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38800 20412
rect 38480 18844 38800 20356
rect 38480 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38800 18844
rect 38480 17276 38800 18788
rect 38480 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38800 17276
rect 38480 15708 38800 17220
rect 38480 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38800 15708
rect 38480 14140 38800 15652
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 38480 12572 38800 14084
rect 38480 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38800 12572
rect 38480 11004 38800 12516
rect 38480 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38800 11004
rect 38480 9436 38800 10948
rect 38480 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38800 9436
rect 38480 7868 38800 9380
rect 38480 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38800 7868
rect 38480 6300 38800 7812
rect 38480 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38800 6300
rect 38480 4732 38800 6244
rect 38480 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38800 4732
rect 38480 3164 38800 4676
rect 38480 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38800 3164
rect 38480 3076 38800 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0__I pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[0\].fbn_I
timestamp 1667941163
transform -1 0 24752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[0\].fbp_I
timestamp 1667941163
transform -1 0 26656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[1\].fbn_I
timestamp 1667941163
transform 1 0 23856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[1\].fbp_I
timestamp 1667941163
transform 1 0 24528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[2\].fbn_I
timestamp 1667941163
transform 1 0 24752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[2\].fbp_I
timestamp 1667941163
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[3\].fbn_I
timestamp 1667941163
transform -1 0 18928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_FB\[3\].fbp_I
timestamp 1667941163
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[0\].thrun_I
timestamp 1667941163
transform 1 0 19600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[0\].thrup_I
timestamp 1667941163
transform 1 0 23184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[1\].thrun_I
timestamp 1667941163
transform 1 0 18144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[1\].thrup_I
timestamp 1667941163
transform 1 0 21840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[2\].thrun_I
timestamp 1667941163
transform 1 0 17696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[2\].thrup_I
timestamp 1667941163
transform 1 0 22288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[3\].thrun_I
timestamp 1667941163
transform 1 0 19936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[3\].thrup_I
timestamp 1667941163
transform -1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[4\].thrun_I
timestamp 1667941163
transform 1 0 20496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[4\].thrup_I
timestamp 1667941163
transform -1 0 26208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[5\].thrun_I
timestamp 1667941163
transform 1 0 20384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[5\].thrup_I
timestamp 1667941163
transform -1 0 24304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[6\].thrun_I
timestamp 1667941163
transform 1 0 20832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[6\].thrup_I
timestamp 1667941163
transform 1 0 22736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[7\].thrun_I
timestamp 1667941163
transform -1 0 22512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[7\].thrup_I
timestamp 1667941163
transform -1 0 26656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[8\].thrun_I
timestamp 1667941163
transform 1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[8\].thrup_I
timestamp 1667941163
transform 1 0 26880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[9\].thrun_I
timestamp 1667941163
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_T\[9\].thrup_I
timestamp 1667941163
transform -1 0 19712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[0\].crossn_I
timestamp 1667941163
transform 1 0 21392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[0\].crossp_I
timestamp 1667941163
transform 1 0 23184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[1\].crossn_I
timestamp 1667941163
transform 1 0 31808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[1\].crossp_I
timestamp 1667941163
transform 1 0 23856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[2\].crossn_I
timestamp 1667941163
transform -1 0 24528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[2\].crossp_I
timestamp 1667941163
transform 1 0 19152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[3\].crossn_I
timestamp 1667941163
transform 1 0 32144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[3\].crossp_I
timestamp 1667941163
transform 1 0 19040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[4\].crossn_I
timestamp 1667941163
transform -1 0 25424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans0p.gen_X\[4\].crossp_I
timestamp 1667941163
transform 1 0 24752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[0\].fbn_I
timestamp 1667941163
transform 1 0 29120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[0\].fbp_I
timestamp 1667941163
transform -1 0 29792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[1\].fbn_I
timestamp 1667941163
transform 1 0 34384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[1\].fbp_I
timestamp 1667941163
transform 1 0 33040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[2\].fbn_I
timestamp 1667941163
transform 1 0 33488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[2\].fbp_I
timestamp 1667941163
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[3\].fbn_I
timestamp 1667941163
transform 1 0 30576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_FB\[3\].fbp_I
timestamp 1667941163
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[0\].thrun_I
timestamp 1667941163
transform 1 0 33936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[0\].thrup_I
timestamp 1667941163
transform 1 0 25984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[1\].thrun_I
timestamp 1667941163
transform 1 0 31360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[1\].thrup_I
timestamp 1667941163
transform 1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[2\].thrun_I
timestamp 1667941163
transform 1 0 32592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[2\].thrup_I
timestamp 1667941163
transform 1 0 27328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[3\].thrun_I
timestamp 1667941163
transform -1 0 28000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[3\].thrup_I
timestamp 1667941163
transform 1 0 28672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[4\].thrun_I
timestamp 1667941163
transform 1 0 34832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[4\].thrup_I
timestamp 1667941163
transform 1 0 34384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[5\].thrun_I
timestamp 1667941163
transform 1 0 30016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[5\].thrup_I
timestamp 1667941163
transform 1 0 27328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[6\].thrun_I
timestamp 1667941163
transform 1 0 26432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[6\].thrup_I
timestamp 1667941163
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[7\].thrun_I
timestamp 1667941163
transform 1 0 27776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[7\].thrup_I
timestamp 1667941163
transform 1 0 28224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[8\].thrun_I
timestamp 1667941163
transform 1 0 30912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[8\].thrup_I
timestamp 1667941163
transform 1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[9\].thrun_I
timestamp 1667941163
transform 1 0 27440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_T\[9\].thrup_I
timestamp 1667941163
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[0\].crossn_I
timestamp 1667941163
transform 1 0 31920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[0\].crossp_I
timestamp 1667941163
transform 1 0 33488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[1\].crossn_I
timestamp 1667941163
transform 1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[1\].crossp_I
timestamp 1667941163
transform 1 0 31472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[2\].crossn_I
timestamp 1667941163
transform 1 0 33936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[2\].crossp_I
timestamp 1667941163
transform 1 0 35728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[3\].crossn_I
timestamp 1667941163
transform 1 0 34832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[3\].crossp_I
timestamp 1667941163
transform 1 0 30128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[4\].crossn_I
timestamp 1667941163
transform 1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_trans1p.gen_X\[4\].crossp_I
timestamp 1667941163
transform 1 0 34384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37
timestamp 1667941163
transform 1 0 5488 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72
timestamp 1667941163
transform 1 0 9408 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 13328 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 15120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 15568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129
timestamp 1667941163
transform 1 0 15792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132
timestamp 1667941163
transform 1 0 16128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 16800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142
timestamp 1667941163
transform 1 0 17248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148
timestamp 1667941163
transform 1 0 17920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_152
timestamp 1667941163
transform 1 0 18368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_156
timestamp 1667941163
transform 1 0 18816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_162
timestamp 1667941163
transform 1 0 19488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168
timestamp 1667941163
transform 1 0 20160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_177
timestamp 1667941163
transform 1 0 21168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_183
timestamp 1667941163
transform 1 0 21840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_189
timestamp 1667941163
transform 1 0 22512 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195
timestamp 1667941163
transform 1 0 23184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_201
timestamp 1667941163
transform 1 0 23856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_207
timestamp 1667941163
transform 1 0 24528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1667941163
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1667941163
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_217
timestamp 1667941163
transform 1 0 25648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_223
timestamp 1667941163
transform 1 0 26320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_229
timestamp 1667941163
transform 1 0 26992 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_235
timestamp 1667941163
transform 1 0 27664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_241
timestamp 1667941163
transform 1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1667941163
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_252
timestamp 1667941163
transform 1 0 29568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_258
timestamp 1667941163
transform 1 0 30240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_264
timestamp 1667941163
transform 1 0 30912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_270
timestamp 1667941163
transform 1 0 31584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_276
timestamp 1667941163
transform 1 0 32256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1667941163
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_287
timestamp 1667941163
transform 1 0 33488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_293
timestamp 1667941163
transform 1 0 34160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_297
timestamp 1667941163
transform 1 0 34608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_301
timestamp 1667941163
transform 1 0 35056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_305
timestamp 1667941163
transform 1 0 35504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_309
timestamp 1667941163
transform 1 0 35952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1667941163
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_317 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 36848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_325
timestamp 1667941163
transform 1 0 37744 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329
timestamp 1667941163
transform 1 0 38192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1667941163
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_144
timestamp 1667941163
transform 1 0 17472 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_152
timestamp 1667941163
transform 1 0 18368 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_154
timestamp 1667941163
transform 1 0 18592 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_157
timestamp 1667941163
transform 1 0 18928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_161
timestamp 1667941163
transform 1 0 19376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_165
timestamp 1667941163
transform 1 0 19824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_171
timestamp 1667941163
transform 1 0 20496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_177
timestamp 1667941163
transform 1 0 21168 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_183
timestamp 1667941163
transform 1 0 21840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_189
timestamp 1667941163
transform 1 0 22512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_195
timestamp 1667941163
transform 1 0 23184 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_201
timestamp 1667941163
transform 1 0 23856 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_207
timestamp 1667941163
transform 1 0 24528 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_211
timestamp 1667941163
transform 1 0 24976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1667941163
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_220
timestamp 1667941163
transform 1 0 25984 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_226
timestamp 1667941163
transform 1 0 26656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_232
timestamp 1667941163
transform 1 0 27328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_238
timestamp 1667941163
transform 1 0 28000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_244
timestamp 1667941163
transform 1 0 28672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_250
timestamp 1667941163
transform 1 0 29344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_256
timestamp 1667941163
transform 1 0 30016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_262
timestamp 1667941163
transform 1 0 30688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_268
timestamp 1667941163
transform 1 0 31360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_274
timestamp 1667941163
transform 1 0 32032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_280
timestamp 1667941163
transform 1 0 32704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1667941163
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_289
timestamp 1667941163
transform 1 0 33712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_293
timestamp 1667941163
transform 1 0 34160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_297
timestamp 1667941163
transform 1 0 34608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_301
timestamp 1667941163
transform 1 0 35056 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_317
timestamp 1667941163
transform 1 0 36848 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_325
timestamp 1667941163
transform 1 0 37744 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_329
timestamp 1667941163
transform 1 0 38192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1667941163
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1667941163
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1667941163
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_108
timestamp 1667941163
transform 1 0 13440 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_140
timestamp 1667941163
transform 1 0 17024 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_156
timestamp 1667941163
transform 1 0 18816 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_160
timestamp 1667941163
transform 1 0 19264 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_164
timestamp 1667941163
transform 1 0 19712 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_168
timestamp 1667941163
transform 1 0 20160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_172
timestamp 1667941163
transform 1 0 20608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_179
timestamp 1667941163
transform 1 0 21392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_185
timestamp 1667941163
transform 1 0 22064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_191
timestamp 1667941163
transform 1 0 22736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 23408 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_203
timestamp 1667941163
transform 1 0 24080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_209
timestamp 1667941163
transform 1 0 24752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_215
timestamp 1667941163
transform 1 0 25424 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_221
timestamp 1667941163
transform 1 0 26096 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_227
timestamp 1667941163
transform 1 0 26768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_233
timestamp 1667941163
transform 1 0 27440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_239
timestamp 1667941163
transform 1 0 28112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_245
timestamp 1667941163
transform 1 0 28784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1667941163
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1667941163
transform 1 0 29344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_255
timestamp 1667941163
transform 1 0 29904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_261
timestamp 1667941163
transform 1 0 30576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_267
timestamp 1667941163
transform 1 0 31248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_273
timestamp 1667941163
transform 1 0 31920 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_277
timestamp 1667941163
transform 1 0 32368 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_281
timestamp 1667941163
transform 1 0 32816 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_285
timestamp 1667941163
transform 1 0 33264 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_289
timestamp 1667941163
transform 1 0 33712 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_293
timestamp 1667941163
transform 1 0 34160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_297
timestamp 1667941163
transform 1 0 34608 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_313
timestamp 1667941163
transform 1 0 36400 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_317
timestamp 1667941163
transform 1 0 36848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_321
timestamp 1667941163
transform 1 0 37296 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_329
timestamp 1667941163
transform 1 0 38192 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1667941163
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_144
timestamp 1667941163
transform 1 0 17472 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_160
timestamp 1667941163
transform 1 0 19264 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_168
timestamp 1667941163
transform 1 0 20160 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_170
timestamp 1667941163
transform 1 0 20384 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_173
timestamp 1667941163
transform 1 0 20720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_177
timestamp 1667941163
transform 1 0 21168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_181
timestamp 1667941163
transform 1 0 21616 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_187
timestamp 1667941163
transform 1 0 22288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_193
timestamp 1667941163
transform 1 0 22960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_199
timestamp 1667941163
transform 1 0 23632 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_205
timestamp 1667941163
transform 1 0 24304 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_211
timestamp 1667941163
transform 1 0 24976 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1667941163
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_220
timestamp 1667941163
transform 1 0 25984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_226
timestamp 1667941163
transform 1 0 26656 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_232
timestamp 1667941163
transform 1 0 27328 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_238
timestamp 1667941163
transform 1 0 28000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_244
timestamp 1667941163
transform 1 0 28672 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_250
timestamp 1667941163
transform 1 0 29344 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_256
timestamp 1667941163
transform 1 0 30016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_262
timestamp 1667941163
transform 1 0 30688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_266
timestamp 1667941163
transform 1 0 31136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_270
timestamp 1667941163
transform 1 0 31584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_274
timestamp 1667941163
transform 1 0 32032 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 32480 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1667941163
transform 1 0 32928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1667941163
transform 1 0 33376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_289
timestamp 1667941163
transform 1 0 33712 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_321
timestamp 1667941163
transform 1 0 37296 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_329
timestamp 1667941163
transform 1 0 38192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1667941163
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1667941163
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1667941163
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1667941163
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1667941163
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_179
timestamp 1667941163
transform 1 0 21392 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_185
timestamp 1667941163
transform 1 0 22064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_189
timestamp 1667941163
transform 1 0 22512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_195
timestamp 1667941163
transform 1 0 23184 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_201
timestamp 1667941163
transform 1 0 23856 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_207
timestamp 1667941163
transform 1 0 24528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_213
timestamp 1667941163
transform 1 0 25200 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_219
timestamp 1667941163
transform 1 0 25872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_225
timestamp 1667941163
transform 1 0 26544 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_231
timestamp 1667941163
transform 1 0 27216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_235
timestamp 1667941163
transform 1 0 27664 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_243
timestamp 1667941163
transform 1 0 28560 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1667941163
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1667941163
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_255
timestamp 1667941163
transform 1 0 29904 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_259
timestamp 1667941163
transform 1 0 30352 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_263
timestamp 1667941163
transform 1 0 30800 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_267
timestamp 1667941163
transform 1 0 31248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_271
timestamp 1667941163
transform 1 0 31696 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_275
timestamp 1667941163
transform 1 0 32144 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_307
timestamp 1667941163
transform 1 0 35728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_315
timestamp 1667941163
transform 1 0 36624 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_321
timestamp 1667941163
transform 1 0 37296 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_329
timestamp 1667941163
transform 1 0 38192 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1667941163
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1667941163
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_144
timestamp 1667941163
transform 1 0 17472 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_176
timestamp 1667941163
transform 1 0 21056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_184
timestamp 1667941163
transform 1 0 21952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_186
timestamp 1667941163
transform 1 0 22176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_189
timestamp 1667941163
transform 1 0 22512 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_193
timestamp 1667941163
transform 1 0 22960 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_197
timestamp 1667941163
transform 1 0 23408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_203
timestamp 1667941163
transform 1 0 24080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_209
timestamp 1667941163
transform 1 0 24752 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1667941163
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_218
timestamp 1667941163
transform 1 0 25760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 26208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_226
timestamp 1667941163
transform 1 0 26656 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_230
timestamp 1667941163
transform 1 0 27104 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_234
timestamp 1667941163
transform 1 0 27552 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_238
timestamp 1667941163
transform 1 0 28000 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_246
timestamp 1667941163
transform 1 0 28896 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_250
timestamp 1667941163
transform 1 0 29344 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_254
timestamp 1667941163
transform 1 0 29792 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_258
timestamp 1667941163
transform 1 0 30240 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_274
timestamp 1667941163
transform 1 0 32032 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1667941163
transform 1 0 32928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_286
timestamp 1667941163
transform 1 0 33376 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_318
timestamp 1667941163
transform 1 0 36960 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_326
timestamp 1667941163
transform 1 0 37856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_330
timestamp 1667941163
transform 1 0 38304 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1667941163
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1667941163
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1667941163
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1667941163
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1667941163
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_179
timestamp 1667941163
transform 1 0 21392 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_197
timestamp 1667941163
transform 1 0 23408 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_203
timestamp 1667941163
transform 1 0 24080 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_207
timestamp 1667941163
transform 1 0 24528 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_211
timestamp 1667941163
transform 1 0 24976 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_215
timestamp 1667941163
transform 1 0 25424 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_219
timestamp 1667941163
transform 1 0 25872 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_222
timestamp 1667941163
transform 1 0 26208 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_226
timestamp 1667941163
transform 1 0 26656 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_230
timestamp 1667941163
transform 1 0 27104 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_234
timestamp 1667941163
transform 1 0 27552 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_238
timestamp 1667941163
transform 1 0 28000 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1667941163
transform 1 0 28448 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_246
timestamp 1667941163
transform 1 0 28896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1667941163
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1667941163
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1667941163
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_321
timestamp 1667941163
transform 1 0 37296 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_329
timestamp 1667941163
transform 1 0 38192 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1667941163
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1667941163
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_144
timestamp 1667941163
transform 1 0 17472 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_176
timestamp 1667941163
transform 1 0 21056 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_192
timestamp 1667941163
transform 1 0 22848 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_200
timestamp 1667941163
transform 1 0 23744 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_202
timestamp 1667941163
transform 1 0 23968 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_205
timestamp 1667941163
transform 1 0 24304 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_209
timestamp 1667941163
transform 1 0 24752 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_215
timestamp 1667941163
transform 1 0 25424 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_218
timestamp 1667941163
transform 1 0 25760 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 26208 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_226
timestamp 1667941163
transform 1 0 26656 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_230
timestamp 1667941163
transform 1 0 27104 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_262
timestamp 1667941163
transform 1 0 30688 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_278
timestamp 1667941163
transform 1 0 32480 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_282
timestamp 1667941163
transform 1 0 32928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_286
timestamp 1667941163
transform 1 0 33376 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_318
timestamp 1667941163
transform 1 0 36960 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_326
timestamp 1667941163
transform 1 0 37856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_330
timestamp 1667941163
transform 1 0 38304 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1667941163
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1667941163
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1667941163
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1667941163
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1667941163
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1667941163
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1667941163
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1667941163
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1667941163
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1667941163
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_321
timestamp 1667941163
transform 1 0 37296 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_329
timestamp 1667941163
transform 1 0 38192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1667941163
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1667941163
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1667941163
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1667941163
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1667941163
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1667941163
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1667941163
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1667941163
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_286
timestamp 1667941163
transform 1 0 33376 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_318
timestamp 1667941163
transform 1 0 36960 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_326
timestamp 1667941163
transform 1 0 37856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_330
timestamp 1667941163
transform 1 0 38304 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1667941163
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1667941163
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1667941163
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1667941163
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1667941163
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1667941163
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1667941163
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1667941163
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1667941163
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_321
timestamp 1667941163
transform 1 0 37296 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_329
timestamp 1667941163
transform 1 0 38192 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1667941163
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1667941163
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1667941163
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1667941163
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1667941163
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1667941163
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1667941163
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1667941163
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_286
timestamp 1667941163
transform 1 0 33376 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_318
timestamp 1667941163
transform 1 0 36960 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_326
timestamp 1667941163
transform 1 0 37856 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_330
timestamp 1667941163
transform 1 0 38304 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1667941163
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1667941163
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1667941163
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1667941163
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1667941163
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1667941163
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1667941163
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1667941163
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1667941163
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1667941163
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1667941163
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_321
timestamp 1667941163
transform 1 0 37296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_329
timestamp 1667941163
transform 1 0 38192 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1667941163
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1667941163
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1667941163
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1667941163
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1667941163
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1667941163
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1667941163
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_286
timestamp 1667941163
transform 1 0 33376 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_318
timestamp 1667941163
transform 1 0 36960 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_326
timestamp 1667941163
transform 1 0 37856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_330
timestamp 1667941163
transform 1 0 38304 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1667941163
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1667941163
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1667941163
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1667941163
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1667941163
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1667941163
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1667941163
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1667941163
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1667941163
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1667941163
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1667941163
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1667941163
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_321
timestamp 1667941163
transform 1 0 37296 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_329
timestamp 1667941163
transform 1 0 38192 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1667941163
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1667941163
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1667941163
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1667941163
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1667941163
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1667941163
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1667941163
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1667941163
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_286
timestamp 1667941163
transform 1 0 33376 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_318
timestamp 1667941163
transform 1 0 36960 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_326
timestamp 1667941163
transform 1 0 37856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_330
timestamp 1667941163
transform 1 0 38304 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1667941163
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1667941163
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1667941163
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1667941163
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1667941163
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1667941163
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1667941163
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1667941163
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1667941163
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1667941163
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1667941163
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1667941163
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1667941163
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_321
timestamp 1667941163
transform 1 0 37296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_329
timestamp 1667941163
transform 1 0 38192 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1667941163
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1667941163
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1667941163
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1667941163
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1667941163
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1667941163
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1667941163
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1667941163
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1667941163
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1667941163
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1667941163
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1667941163
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_286
timestamp 1667941163
transform 1 0 33376 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_318
timestamp 1667941163
transform 1 0 36960 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_326
timestamp 1667941163
transform 1 0 37856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_330
timestamp 1667941163
transform 1 0 38304 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1667941163
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1667941163
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1667941163
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1667941163
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1667941163
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1667941163
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1667941163
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1667941163
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1667941163
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1667941163
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1667941163
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1667941163
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1667941163
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1667941163
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_321
timestamp 1667941163
transform 1 0 37296 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_329
timestamp 1667941163
transform 1 0 38192 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1667941163
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1667941163
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1667941163
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1667941163
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1667941163
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1667941163
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1667941163
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1667941163
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1667941163
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1667941163
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1667941163
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1667941163
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_286
timestamp 1667941163
transform 1 0 33376 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_318
timestamp 1667941163
transform 1 0 36960 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_326
timestamp 1667941163
transform 1 0 37856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_330
timestamp 1667941163
transform 1 0 38304 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1667941163
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1667941163
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1667941163
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1667941163
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1667941163
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_108
timestamp 1667941163
transform 1 0 13440 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_140
timestamp 1667941163
transform 1 0 17024 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_156
timestamp 1667941163
transform 1 0 18816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_164
timestamp 1667941163
transform 1 0 19712 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_169
timestamp 1667941163
transform 1 0 20272 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_175
timestamp 1667941163
transform 1 0 20944 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1667941163
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1667941163
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1667941163
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1667941163
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1667941163
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1667941163
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_321
timestamp 1667941163
transform 1 0 37296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_329
timestamp 1667941163
transform 1 0 38192 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1667941163
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1667941163
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1667941163
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1667941163
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1667941163
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1667941163
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_144
timestamp 1667941163
transform 1 0 17472 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_152
timestamp 1667941163
transform 1 0 18368 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_158
timestamp 1667941163
transform 1 0 19040 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_164
timestamp 1667941163
transform 1 0 19712 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_170
timestamp 1667941163
transform 1 0 20384 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_176
timestamp 1667941163
transform 1 0 21056 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1667941163
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1667941163
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1667941163
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1667941163
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1667941163
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_286
timestamp 1667941163
transform 1 0 33376 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_318
timestamp 1667941163
transform 1 0 36960 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_326
timestamp 1667941163
transform 1 0 37856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_330
timestamp 1667941163
transform 1 0 38304 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1667941163
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1667941163
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1667941163
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1667941163
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1667941163
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_108
timestamp 1667941163
transform 1 0 13440 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_140
timestamp 1667941163
transform 1 0 17024 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_156
timestamp 1667941163
transform 1 0 18816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_160
timestamp 1667941163
transform 1 0 19264 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_162
timestamp 1667941163
transform 1 0 19488 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_167
timestamp 1667941163
transform 1 0 20048 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_173
timestamp 1667941163
transform 1 0 20720 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1667941163
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1667941163
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1667941163
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1667941163
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1667941163
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_321
timestamp 1667941163
transform 1 0 37296 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_329
timestamp 1667941163
transform 1 0 38192 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1667941163
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1667941163
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1667941163
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1667941163
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1667941163
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1667941163
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1667941163
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1667941163
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1667941163
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1667941163
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1667941163
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1667941163
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_286
timestamp 1667941163
transform 1 0 33376 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_318
timestamp 1667941163
transform 1 0 36960 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_326
timestamp 1667941163
transform 1 0 37856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_330
timestamp 1667941163
transform 1 0 38304 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1667941163
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1667941163
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1667941163
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1667941163
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1667941163
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1667941163
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1667941163
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1667941163
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1667941163
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1667941163
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1667941163
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1667941163
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1667941163
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_321
timestamp 1667941163
transform 1 0 37296 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_329
timestamp 1667941163
transform 1 0 38192 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1667941163
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1667941163
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1667941163
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1667941163
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1667941163
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1667941163
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1667941163
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1667941163
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1667941163
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1667941163
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1667941163
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1667941163
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_286
timestamp 1667941163
transform 1 0 33376 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_318
timestamp 1667941163
transform 1 0 36960 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_326
timestamp 1667941163
transform 1 0 37856 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_330
timestamp 1667941163
transform 1 0 38304 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1667941163
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1667941163
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1667941163
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1667941163
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1667941163
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1667941163
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1667941163
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1667941163
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1667941163
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1667941163
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1667941163
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1667941163
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1667941163
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1667941163
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_321
timestamp 1667941163
transform 1 0 37296 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_329
timestamp 1667941163
transform 1 0 38192 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1667941163
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1667941163
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1667941163
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1667941163
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1667941163
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1667941163
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1667941163
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1667941163
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1667941163
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1667941163
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1667941163
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1667941163
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_286
timestamp 1667941163
transform 1 0 33376 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_318
timestamp 1667941163
transform 1 0 36960 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_326
timestamp 1667941163
transform 1 0 37856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_330
timestamp 1667941163
transform 1 0 38304 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1667941163
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1667941163
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1667941163
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1667941163
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1667941163
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1667941163
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1667941163
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1667941163
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1667941163
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1667941163
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1667941163
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1667941163
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1667941163
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1667941163
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_321
timestamp 1667941163
transform 1 0 37296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_329
timestamp 1667941163
transform 1 0 38192 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1667941163
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1667941163
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1667941163
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1667941163
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1667941163
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1667941163
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1667941163
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1667941163
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1667941163
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1667941163
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1667941163
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1667941163
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_286
timestamp 1667941163
transform 1 0 33376 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_318
timestamp 1667941163
transform 1 0 36960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_326
timestamp 1667941163
transform 1 0 37856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_330
timestamp 1667941163
transform 1 0 38304 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1667941163
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1667941163
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1667941163
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1667941163
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1667941163
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1667941163
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1667941163
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1667941163
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1667941163
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1667941163
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1667941163
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1667941163
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1667941163
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1667941163
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_321
timestamp 1667941163
transform 1 0 37296 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_329
timestamp 1667941163
transform 1 0 38192 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1667941163
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1667941163
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1667941163
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1667941163
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1667941163
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1667941163
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1667941163
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1667941163
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1667941163
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1667941163
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1667941163
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1667941163
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_286
timestamp 1667941163
transform 1 0 33376 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_318
timestamp 1667941163
transform 1 0 36960 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_326
timestamp 1667941163
transform 1 0 37856 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_330
timestamp 1667941163
transform 1 0 38304 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1667941163
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1667941163
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1667941163
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1667941163
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1667941163
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1667941163
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1667941163
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1667941163
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1667941163
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1667941163
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1667941163
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1667941163
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1667941163
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1667941163
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_321
timestamp 1667941163
transform 1 0 37296 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_329
timestamp 1667941163
transform 1 0 38192 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1667941163
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1667941163
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1667941163
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1667941163
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1667941163
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1667941163
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1667941163
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1667941163
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1667941163
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1667941163
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1667941163
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1667941163
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_286
timestamp 1667941163
transform 1 0 33376 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_318
timestamp 1667941163
transform 1 0 36960 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_326
timestamp 1667941163
transform 1 0 37856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_330
timestamp 1667941163
transform 1 0 38304 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1667941163
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1667941163
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1667941163
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1667941163
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1667941163
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1667941163
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1667941163
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1667941163
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1667941163
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1667941163
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1667941163
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1667941163
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1667941163
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1667941163
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_321
timestamp 1667941163
transform 1 0 37296 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_329
timestamp 1667941163
transform 1 0 38192 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1667941163
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1667941163
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1667941163
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1667941163
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1667941163
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1667941163
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1667941163
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1667941163
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1667941163
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1667941163
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1667941163
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1667941163
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_286
timestamp 1667941163
transform 1 0 33376 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_318
timestamp 1667941163
transform 1 0 36960 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_326
timestamp 1667941163
transform 1 0 37856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_330
timestamp 1667941163
transform 1 0 38304 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1667941163
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1667941163
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1667941163
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1667941163
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1667941163
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1667941163
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1667941163
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1667941163
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1667941163
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1667941163
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1667941163
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1667941163
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1667941163
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1667941163
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_321
timestamp 1667941163
transform 1 0 37296 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_329
timestamp 1667941163
transform 1 0 38192 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1667941163
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1667941163
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1667941163
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1667941163
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1667941163
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1667941163
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1667941163
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1667941163
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1667941163
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1667941163
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1667941163
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1667941163
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_286
timestamp 1667941163
transform 1 0 33376 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_318
timestamp 1667941163
transform 1 0 36960 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_326
timestamp 1667941163
transform 1 0 37856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_330
timestamp 1667941163
transform 1 0 38304 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1667941163
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1667941163
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1667941163
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1667941163
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1667941163
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1667941163
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1667941163
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1667941163
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1667941163
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1667941163
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1667941163
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1667941163
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1667941163
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1667941163
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_321
timestamp 1667941163
transform 1 0 37296 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_329
timestamp 1667941163
transform 1 0 38192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1667941163
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1667941163
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1667941163
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1667941163
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1667941163
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1667941163
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1667941163
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1667941163
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1667941163
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1667941163
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1667941163
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1667941163
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_286
timestamp 1667941163
transform 1 0 33376 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_318
timestamp 1667941163
transform 1 0 36960 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_326
timestamp 1667941163
transform 1 0 37856 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_330
timestamp 1667941163
transform 1 0 38304 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1667941163
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1667941163
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1667941163
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1667941163
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1667941163
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1667941163
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1667941163
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1667941163
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1667941163
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1667941163
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1667941163
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1667941163
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1667941163
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1667941163
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_321
timestamp 1667941163
transform 1 0 37296 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_329
timestamp 1667941163
transform 1 0 38192 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1667941163
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1667941163
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1667941163
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1667941163
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1667941163
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1667941163
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1667941163
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1667941163
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1667941163
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1667941163
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1667941163
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1667941163
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_286
timestamp 1667941163
transform 1 0 33376 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_318
timestamp 1667941163
transform 1 0 36960 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_326
timestamp 1667941163
transform 1 0 37856 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_330
timestamp 1667941163
transform 1 0 38304 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1667941163
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1667941163
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_37
timestamp 1667941163
transform 1 0 5488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_69
timestamp 1667941163
transform 1 0 9072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_72
timestamp 1667941163
transform 1 0 9408 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1667941163
transform 1 0 12992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_107
timestamp 1667941163
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 16912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_142
timestamp 1667941163
transform 1 0 17248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1667941163
transform 1 0 20832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1667941163
transform 1 0 21168 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1667941163
transform 1 0 24752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_212
timestamp 1667941163
transform 1 0 25088 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1667941163
transform 1 0 28672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_247
timestamp 1667941163
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_279
timestamp 1667941163
transform 1 0 32592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_282
timestamp 1667941163
transform 1 0 32928 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1667941163
transform 1 0 36512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_317
timestamp 1667941163
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_325
timestamp 1667941163
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_329
timestamp 1667941163
transform 1 0 38192 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1667941163
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1667941163
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1667941163
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1667941163
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1667941163
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1667941163
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1667941163
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1667941163
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1667941163
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1667941163
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1667941163
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1667941163
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1667941163
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1667941163
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1667941163
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1667941163
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1667941163
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1667941163
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1667941163
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1667941163
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1667941163
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1667941163
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1667941163
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1667941163
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1667941163
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1667941163
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1667941163
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1667941163
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1667941163
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1667941163
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1667941163
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1667941163
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1667941163
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1667941163
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1667941163
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1667941163
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1667941163
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1667941163
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1667941163
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1667941163
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1667941163
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1667941163
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1667941163
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1667941163
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1667941163
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1667941163
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1667941163
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1667941163
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1667941163
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1667941163
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1667941163
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1667941163
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1667941163
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1667941163
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1667941163
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1667941163
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1667941163
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1667941163
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1667941163
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1667941163
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1667941163
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1667941163
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1667941163
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1667941163
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1667941163
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1667941163
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1667941163
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1667941163
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1667941163
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1667941163
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1667941163
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1667941163
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1667941163
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1667941163
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1667941163
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1667941163
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1667941163
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1667941163
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1667941163
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1667941163
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1667941163
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1667941163
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1667941163
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1667941163
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1667941163
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1667941163
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1667941163
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1667941163
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1667941163
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1667941163
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1667941163
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1667941163
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1667941163
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1667941163
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1667941163
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1667941163
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1667941163
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1667941163
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1667941163
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1667941163
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1667941163
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1667941163
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1667941163
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1667941163
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1667941163
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1667941163
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1667941163
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1667941163
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1667941163
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1667941163
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1667941163
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1667941163
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1667941163
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1667941163
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1667941163
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1667941163
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1667941163
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1667941163
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1667941163
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1667941163
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1667941163
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1667941163
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1667941163
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1667941163
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1667941163
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1667941163
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 17024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 16352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 19040 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _2_
timestamp 1667941163
transform -1 0 20272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _3_
timestamp 1667941163
transform -1 0 19712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _4_
timestamp 1667941163
transform -1 0 20048 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _5_
timestamp 1667941163
transform -1 0 20384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _6_
timestamp 1667941163
transform -1 0 21056 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _7_
timestamp 1667941163
transform -1 0 20720 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _8_
timestamp 1667941163
transform -1 0 20944 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[0\].fbn
timestamp 1667941163
transform -1 0 24528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 25648 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 23632 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 24080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 22288 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[2\].fbp
timestamp 1667941163
transform -1 0 27664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 22736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 26208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 22064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 23408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 20384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 23184 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 19712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 22512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 20720 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 25536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 22736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 25200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 21392 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 24304 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 21616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 25872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 21392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 26544 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 21840 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 22736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[1\].crossn
timestamp 1667941163
transform -1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 23408 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 24528 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 20048 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 26880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 19040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 24976 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans0p.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 23856 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[0\].fbn
timestamp 1667941163
transform -1 0 28896 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 28896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 33712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 29456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 33040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 29456 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 30240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[0\].thrun
timestamp 1667941163
transform -1 0 30240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 26208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 26320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 28896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 26992 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 27664 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 28224 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[4\].thrun
timestamp 1667941163
transform -1 0 30912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[4\].thrup
timestamp 1667941163
transform -1 0 29568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 29568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 26880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 26096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 25424 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 27552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 27552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 28224 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 26768 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 25536 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 24752 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 30800 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 30912 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 29568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 30240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 31472 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 31808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 28112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 30128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_trans1p.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 31584 0 -1 4704
box -86 -86 534 870
<< labels >>
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 27328 0 27440 800 0 FreeSans 448 90 0 0 clko
port 1 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 latch
port 2 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 on
port 3 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 op
port 4 nsew signal tristate
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 rst
port 5 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 sdi
port 6 nsew signal input
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 sig
port 7 nsew signal input
flabel metal4 s 5846 3076 6166 36908 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 15170 3076 15490 36908 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 24494 3076 24814 36908 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 33818 3076 34138 36908 0 FreeSans 1280 90 0 0 vdd
port 8 nsew power bidirectional
flabel metal4 s 10508 3076 10828 36908 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
flabel metal4 s 19832 3076 20152 36908 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
flabel metal4 s 29156 3076 29476 36908 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
flabel metal4 s 38480 3076 38800 36908 0 FreeSans 1280 90 0 0 vss
port 9 nsew ground bidirectional
rlabel metal1 19992 36848 19992 36848 0 vdd
rlabel via1 20072 36064 20072 36064 0 vss
rlabel metal2 2744 2086 2744 2086 0 clk
rlabel metal2 27384 1302 27384 1302 0 clko
rlabel metal3 26096 6104 26096 6104 0 on
rlabel metal3 25368 6440 25368 6440 0 op
rlabel metal2 21000 5712 21000 5712 0 sdi
rlabel metal2 23520 4312 23520 4312 0 sig
rlabel metal2 29400 3584 29400 3584 0 u_trans0p.outn
rlabel metal2 21448 4928 21448 4928 0 u_trans0p.outp
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
