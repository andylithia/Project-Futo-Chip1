* NGSPICE file created from caparray_s1_flat.ext - technology: gf180mcuC

.subckt caparray_s1_flat cap_series_gygyn cap_series_gygyp cap_series_gyn cap_series_gyp
+ cap_shunt_gyn cap_shunt_gyp cap_shunt_n cap_shunt_p tune_series_gy[0] tune_series_gy[1]
+ tune_series_gy[2] tune_series_gy[3] tune_series_gy[4] tune_series_gy[5] tune_series_gygy[0]
+ tune_series_gygy[1] tune_series_gygy[2] tune_series_gygy[3] tune_series_gygy[4]
+ tune_series_gygy[5] tune_shunt[0] tune_shunt[1] tune_shunt[2] tune_shunt[3] tune_shunt[4]
+ tune_shunt[5] tune_shunt[6] tune_shunt[7] tune_shunt_gy[0] tune_shunt_gy[1] tune_shunt_gy[2]
+ tune_shunt_gy[3] tune_shunt_gy[4] tune_shunt_gy[5] tune_shunt_gy[6] vss vdd

X0 a_32604_48983# a_32516_49080# vss vss nmos_6p0 w=0.82u l=1u
X1 a_3828_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2 a_2500_50652# cap_shunt_n a_2708_50306# vdd pmos_6p0 w=1.2u l=0.5u
X3 a_24452_36540# cap_shunt_p a_24660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X4 a_9428_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5 a_16500_42812# cap_shunt_n a_16708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X6 a_19524_10260# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7 vss tune_shunt[5] a_9876_53080# vss nmos_6p0 w=0.51u l=0.6u
X8 vss cap_shunt_n a_19936_27992# vss nmos_6p0 w=0.82u l=0.6u
X9 a_6760_7124# cap_series_gyp a_6784_7608# vss nmos_6p0 w=0.82u l=0.6u
X10 a_7748_33058# cap_shunt_n a_7540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X11 vdd a_33500_25896# a_33412_25940# vdd pmos_6p0 w=1.22u l=1u
X12 a_6292_15810# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13 a_31904_45944# cap_shunt_gyp a_31904_45540# vdd pmos_6p0 w=1.215u l=0.5u
X14 a_25572_27508# cap_shunt_p a_25780_27992# vdd pmos_6p0 w=1.2u l=0.5u
X15 vdd a_28124_5079# a_28036_5176# vdd pmos_6p0 w=1.22u l=1u
X16 a_31624_8316# cap_series_gygyn a_31436_8316# vdd pmos_6p0 w=1.2u l=0.5u
X17 vdd a_28572_31735# a_28484_31832# vdd pmos_6p0 w=1.22u l=1u
X18 a_33732_27992# cap_shunt_p a_34664_27992# vss nmos_6p0 w=0.82u l=0.6u
X19 a_24452_33404# cap_shunt_p a_24660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X20 a_34308_19292# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X21 a_35692_14964# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X22 a_35292_52119# a_35204_52216# vss vss nmos_6p0 w=0.82u l=1u
X23 a_3620_43188# cap_shunt_p a_3828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X24 vss cap_shunt_n a_19936_24856# vss nmos_6p0 w=0.82u l=0.6u
X25 vdd a_9644_7080# a_9556_7124# vdd pmos_6p0 w=1.22u l=1u
X26 vdd a_33500_22760# a_33412_22804# vdd pmos_6p0 w=1.22u l=1u
X27 a_19544_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X28 a_22064_23288# cap_shunt_p a_20740_23288# vss nmos_6p0 w=0.82u l=0.6u
X29 a_8968_6340# cap_series_gyp a_7768_6748# vss nmos_6p0 w=0.82u l=0.6u
X30 a_34308_16156# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X31 a_21316_3988# cap_series_gyn a_21524_4472# vdd pmos_6p0 w=1.2u l=0.5u
X32 a_35692_11828# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X33 a_24660_11106# cap_series_gyp a_24452_11452# vdd pmos_6p0 w=1.2u l=0.5u
X34 vdd a_8860_11351# a_8772_11448# vdd pmos_6p0 w=1.22u l=1u
X35 vdd a_36636_40008# a_36548_40052# vdd pmos_6p0 w=1.22u l=1u
X36 vdd a_20620_45847# a_20532_45944# vdd pmos_6p0 w=1.22u l=1u
X37 vss tune_series_gy[3] a_29720_9884# vss nmos_6p0 w=0.51u l=0.6u
X38 a_19276_23895# a_19188_23992# vss vss nmos_6p0 w=0.82u l=1u
X39 a_10548_27992# cap_shunt_n a_12264_27992# vss nmos_6p0 w=0.82u l=0.6u
X40 vdd a_37868_23895# a_37780_23992# vdd pmos_6p0 w=1.22u l=1u
X41 a_7580_8316# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X42 a_7952_14180# cap_shunt_p a_6628_14242# vss nmos_6p0 w=0.82u l=0.6u
X43 a_13460_26424# cap_shunt_n a_13252_25940# vdd pmos_6p0 w=1.2u l=0.5u
X44 a_7748_42466# cap_shunt_n a_7540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X45 vdd tune_shunt[7] a_9668_19668# vdd pmos_6p0 w=1.2u l=0.5u
X46 vss tune_shunt[4] a_17828_48376# vss nmos_6p0 w=0.51u l=0.6u
X47 a_32612_37762# cap_shunt_p a_32404_38108# vdd pmos_6p0 w=1.2u l=0.5u
X48 a_25572_36916# cap_shunt_p a_25780_37400# vdd pmos_6p0 w=1.2u l=0.5u
X49 a_3036_29032# a_2948_29076# vss vss nmos_6p0 w=0.82u l=1u
X50 a_3620_19668# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X51 a_38092_35304# a_38004_35348# vss vss nmos_6p0 w=0.82u l=1u
X52 vss cap_shunt_p a_23856_23588# vss nmos_6p0 w=0.82u l=0.6u
X53 vss cap_shunt_p a_11200_17016# vss nmos_6p0 w=0.82u l=0.6u
X54 vdd a_20620_42711# a_20532_42808# vdd pmos_6p0 w=1.22u l=1u
X55 a_9204_51874# cap_shunt_n a_10920_51812# vss nmos_6p0 w=0.82u l=0.6u
X56 a_10548_24856# cap_shunt_n a_12264_24856# vss nmos_6p0 w=0.82u l=0.6u
X57 a_7952_11044# cap_shunt_n a_5844_11106# vss nmos_6p0 w=0.82u l=0.6u
X58 vdd a_37868_20759# a_37780_20856# vdd pmos_6p0 w=1.22u l=1u
X59 a_13460_23288# cap_shunt_n a_13252_22804# vdd pmos_6p0 w=1.2u l=0.5u
X60 a_11800_8692# cap_series_gyp a_11612_8692# vdd pmos_6p0 w=1.2u l=0.5u
X61 a_4704_49944# cap_shunt_p a_3380_49944# vss nmos_6p0 w=0.82u l=0.6u
X62 a_3036_25896# a_2948_25940# vss vss nmos_6p0 w=0.82u l=1u
X63 a_25780_15448# cap_series_gyp a_25572_14964# vdd pmos_6p0 w=1.2u l=0.5u
X64 a_13796_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X65 vdd tune_shunt[6] a_11460_44756# vdd pmos_6p0 w=1.2u l=0.5u
X66 a_24452_14588# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X67 a_35740_53687# a_35652_53784# vss vss nmos_6p0 w=0.82u l=1u
X68 vdd tune_shunt[6] a_10452_45948# vdd pmos_6p0 w=1.2u l=0.5u
X69 a_10660_6402# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X70 a_2724_8692# cap_shunt_n a_2932_9176# vdd pmos_6p0 w=1.2u l=0.5u
X71 vdd a_35628_33303# a_35540_33400# vdd pmos_6p0 w=1.22u l=1u
X72 a_3828_27992# cap_shunt_n a_3620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X73 a_24452_8316# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X74 a_4828_52119# a_4740_52216# vss vss nmos_6p0 w=0.82u l=1u
X75 a_25780_12312# cap_series_gyp a_25572_11828# vdd pmos_6p0 w=1.2u l=0.5u
X76 a_7540_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X77 vdd a_5612_44279# a_5524_44376# vdd pmos_6p0 w=1.22u l=1u
X78 a_22436_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X79 a_17596_50984# a_17508_51028# vss vss nmos_6p0 w=0.82u l=1u
X80 a_35740_50551# a_35652_50648# vss vss nmos_6p0 w=0.82u l=1u
X81 a_17828_48376# cap_shunt_p a_18760_48376# vss nmos_6p0 w=0.82u l=0.6u
X82 a_6740_23288# cap_shunt_p a_8456_23288# vss nmos_6p0 w=0.82u l=0.6u
X83 a_21748_45602# cap_shunt_p a_21540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X84 a_2500_44380# cap_shunt_p a_2708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X85 a_16500_36540# cap_shunt_n a_16708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X86 a_10452_6748# cap_series_gyn a_10660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X87 a_6740_20152# cap_shunt_p a_6532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X88 a_7748_26786# cap_shunt_n a_7540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X89 a_28692_9176# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X90 vdd a_28572_25463# a_28484_25560# vdd pmos_6p0 w=1.22u l=1u
X91 a_3828_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X92 a_17620_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X93 vdd a_26444_53687# a_26356_53784# vdd pmos_6p0 w=1.22u l=1u
X94 a_21516_53687# a_21428_53784# vss vss nmos_6p0 w=0.82u l=1u
X95 a_2500_41244# cap_shunt_p a_2708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X96 a_16500_33404# cap_shunt_n a_16708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X97 a_24452_27132# cap_shunt_p a_24660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X98 a_18612_9538# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X99 a_29700_29922# cap_shunt_p a_31416_29860# vss nmos_6p0 w=0.82u l=0.6u
X100 a_5844_9538# cap_shunt_p a_5636_9884# vdd pmos_6p0 w=1.2u l=0.5u
X101 vdd a_1692_23895# a_1604_23992# vdd pmos_6p0 w=1.22u l=1u
X102 vss cap_shunt_p a_19936_18584# vss nmos_6p0 w=0.82u l=0.6u
X103 a_6292_18584# cap_shunt_p a_8008_18584# vss nmos_6p0 w=0.82u l=0.6u
X104 vdd a_33500_16488# a_33412_16532# vdd pmos_6p0 w=1.22u l=1u
X105 a_29700_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X106 a_31260_38440# a_31172_38484# vss vss nmos_6p0 w=0.82u l=1u
X107 a_10452_30268# cap_shunt_n a_10660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X108 a_28484_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X109 vdd a_28572_22327# a_28484_22424# vdd pmos_6p0 w=1.22u l=1u
X110 a_10316_53687# a_10228_53784# vss vss nmos_6p0 w=0.82u l=1u
X111 vdd a_26444_50551# a_26356_50648# vdd pmos_6p0 w=1.22u l=1u
X112 a_21516_50551# a_21428_50648# vss vss nmos_6p0 w=0.82u l=1u
X113 a_29700_26786# cap_shunt_p a_31416_26724# vss nmos_6p0 w=0.82u l=0.6u
X114 vdd tune_shunt[5] a_13588_49084# vdd pmos_6p0 w=1.2u l=0.5u
X115 a_17620_33780# cap_shunt_n a_17828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X116 vss cap_shunt_p a_19936_15448# vss nmos_6p0 w=0.82u l=0.6u
X117 vdd a_1692_20759# a_1604_20856# vdd pmos_6p0 w=1.22u l=1u
X118 a_12788_49944# cap_shunt_n a_12580_49460# vdd pmos_6p0 w=1.2u l=0.5u
X119 vdd a_20620_39575# a_20532_39672# vdd pmos_6p0 w=1.22u l=1u
X120 a_28484_22804# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X121 a_20532_41620# cap_shunt_p a_20740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X122 a_7748_36194# cap_shunt_n a_7540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X123 a_17620_30644# cap_shunt_n a_17828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X124 a_25780_7608# cap_series_gyn a_25572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X125 a_14692_10744# cap_series_gyn a_14484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X126 a_38092_29032# a_38004_29076# vss vss nmos_6p0 w=0.82u l=1u
X127 vdd a_11884_54120# a_11796_54164# vdd pmos_6p0 w=1.22u l=1u
X128 vdd a_20620_36439# a_20532_36536# vdd pmos_6p0 w=1.22u l=1u
X129 a_34348_8316# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X130 a_15700_7970# cap_series_gyn a_15492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X131 vdd a_37084_54120# a_36996_54164# vdd pmos_6p0 w=1.22u l=1u
X132 a_16500_42812# cap_shunt_n a_16708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X133 vdd a_37868_14487# a_37780_14584# vdd pmos_6p0 w=1.22u l=1u
X134 a_21316_3612# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X135 a_7748_33058# cap_shunt_n a_7540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X136 a_20532_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X137 a_25572_27508# cap_shunt_p a_25780_27992# vdd pmos_6p0 w=1.2u l=0.5u
X138 vdd a_13452_55688# a_13364_55732# vdd pmos_6p0 w=1.22u l=1u
X139 vdd a_37868_11351# a_37780_11448# vdd pmos_6p0 w=1.22u l=1u
X140 a_36160_44757# tune_shunt_gy[3] vdd vdd pmos_6p0 w=1.215u l=0.5u
X141 vss cap_shunt_n a_22848_35832# vss nmos_6p0 w=0.82u l=0.6u
X142 a_24660_44034# cap_shunt_p a_24452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X143 vdd tune_series_gy[1] a_10340_3612# vdd pmos_6p0 w=1.2u l=0.5u
X144 a_16708_20514# cap_shunt_p a_16500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X145 vdd tune_shunt[6] a_10452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X146 a_6572_7124# cap_series_gyp a_6760_7124# vdd pmos_6p0 w=1.2u l=0.5u
X147 a_20740_18584# cap_shunt_p a_20532_18100# vdd pmos_6p0 w=1.2u l=0.5u
X148 a_13564_11351# a_13476_11448# vss vss nmos_6p0 w=0.82u l=1u
X149 a_7540_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X150 vdd a_10428_55688# a_10340_55732# vdd pmos_6p0 w=1.22u l=1u
X151 a_14728_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X152 a_4424_12612# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X153 a_24660_40898# cap_shunt_n a_24452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X154 a_15512_20452# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X155 a_28796_41576# a_28708_41620# vss vss nmos_6p0 w=0.82u l=1u
X156 vss tune_shunt[7] a_6740_20152# vss nmos_6p0 w=0.51u l=0.6u
X157 a_21748_39330# cap_shunt_p a_21540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X158 a_6740_38968# cap_shunt_n a_7672_38968# vss nmos_6p0 w=0.82u l=0.6u
X159 vss cap_series_gyn a_16800_6040# vss nmos_6p0 w=0.82u l=0.6u
X160 a_36524_33303# a_36436_33400# vss vss nmos_6p0 w=0.82u l=1u
X161 a_28684_52119# a_28596_52216# vss vss nmos_6p0 w=0.82u l=1u
X162 vdd a_9644_54120# a_9556_54164# vdd pmos_6p0 w=1.22u l=1u
X163 vss tune_shunt[4] a_32612_31490# vss nmos_6p0 w=0.51u l=0.6u
X164 a_5836_5512# a_5748_5556# vss vss nmos_6p0 w=0.82u l=1u
X165 vdd tune_shunt[3] a_2724_11828# vdd pmos_6p0 w=1.2u l=0.5u
X166 a_24660_4834# cap_series_gyp a_24452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X167 a_7748_45602# cap_shunt_p a_8680_45540# vss nmos_6p0 w=0.82u l=0.6u
X168 a_32612_37762# cap_shunt_p a_32404_38108# vdd pmos_6p0 w=1.2u l=0.5u
X169 a_16500_27132# cap_shunt_n a_16708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X170 a_12108_12919# a_12020_13016# vss vss nmos_6p0 w=0.82u l=1u
X171 vdd a_28572_16055# a_28484_16152# vdd pmos_6p0 w=1.22u l=1u
X172 a_7748_42466# cap_shunt_n a_8680_42404# vss nmos_6p0 w=0.82u l=0.6u
X173 vdd a_1692_14487# a_1604_14584# vdd pmos_6p0 w=1.22u l=1u
X174 vdd tune_shunt[6] a_11460_44756# vdd pmos_6p0 w=1.2u l=0.5u
X175 a_17828_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X176 vss cap_series_gygyp a_36624_22020# vss nmos_6p0 w=0.82u l=0.6u
X177 a_7768_5180# cap_series_gyn a_7580_5180# vdd pmos_6p0 w=1.2u l=0.5u
X178 a_29916_8215# a_29828_8312# vss vss nmos_6p0 w=0.82u l=1u
X179 a_29700_17378# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X180 a_28484_16532# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X181 vdd a_28572_12919# a_28484_13016# vdd pmos_6p0 w=1.22u l=1u
X182 a_29700_17378# cap_series_gyp a_31416_17316# vss nmos_6p0 w=0.82u l=0.6u
X183 a_3380_49944# cap_shunt_p a_3172_49460# vdd pmos_6p0 w=1.2u l=0.5u
X184 a_17620_24372# cap_shunt_n a_17828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X185 a_25592_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X186 vdd a_1692_11351# a_1604_11448# vdd pmos_6p0 w=1.22u l=1u
X187 vss tune_series_gy[5] a_19732_12312# vss nmos_6p0 w=0.51u l=0.6u
X188 a_17828_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X189 a_25780_6040# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X190 a_19544_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X191 a_14484_3988# cap_series_gyp a_14692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X192 a_21748_45602# cap_shunt_p a_21540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X193 a_16500_36540# cap_shunt_n a_16708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X194 vss cap_series_gyp a_23856_9476# vss nmos_6p0 w=0.82u l=0.6u
X195 vss cap_shunt_n a_11984_39268# vss nmos_6p0 w=0.82u l=0.6u
X196 a_13796_37762# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X197 a_7748_26786# cap_shunt_n a_7540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X198 vdd a_10092_40008# a_10004_40052# vdd pmos_6p0 w=1.22u l=1u
X199 a_20532_32212# cap_shunt_n a_20740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X200 a_16136_11044# cap_series_gyp a_15720_11452# vss nmos_6p0 w=0.82u l=0.6u
X201 vdd a_2588_19624# a_2500_19668# vdd pmos_6p0 w=1.22u l=1u
X202 vdd a_31036_41576# a_30948_41620# vdd pmos_6p0 w=1.22u l=1u
X203 vss cap_shunt_n a_30016_38968# vss nmos_6p0 w=0.82u l=0.6u
X204 a_17620_21236# cap_shunt_p a_17828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X205 vdd a_20620_27031# a_20532_27128# vdd pmos_6p0 w=1.22u l=1u
X206 vdd tune_shunt[7] a_7540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X207 vdd a_24652_46280# a_24564_46324# vdd pmos_6p0 w=1.22u l=1u
X208 a_13796_37762# cap_shunt_n a_15512_37700# vss nmos_6p0 w=0.82u l=0.6u
X209 vdd a_18044_13352# a_17956_13396# vdd pmos_6p0 w=1.22u l=1u
X210 vdd a_21628_49416# a_21540_49460# vdd pmos_6p0 w=1.22u l=1u
X211 a_34144_48676# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X212 a_23856_37700# cap_shunt_n a_21748_37762# vss nmos_6p0 w=0.82u l=0.6u
X213 a_16500_33404# cap_shunt_n a_16708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X214 vss cap_shunt_n a_22848_29560# vss nmos_6p0 w=0.82u l=0.6u
X215 a_21540_23996# cap_shunt_p a_21748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X216 a_23072_4772# cap_series_gyp a_21748_4834# vss nmos_6p0 w=0.82u l=0.6u
X217 a_6292_51874# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X218 vss tune_shunt[6] a_3828_43672# vss nmos_6p0 w=0.51u l=0.6u
X219 a_13796_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X220 a_10660_6402# cap_series_gyn a_10452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X221 a_2724_8692# cap_shunt_n a_2932_9176# vdd pmos_6p0 w=1.2u l=0.5u
X222 vss tune_shunt[7] a_12788_17016# vss nmos_6p0 w=0.51u l=0.6u
X223 a_20532_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X224 vss tune_shunt[7] a_20740_32696# vss nmos_6p0 w=0.51u l=0.6u
X225 vss tune_shunt[2] a_1924_6040# vss nmos_6p0 w=0.51u l=0.6u
X226 vdd a_23756_18056# a_23668_18100# vdd pmos_6p0 w=1.22u l=1u
X227 vss cap_shunt_n a_22848_26424# vss nmos_6p0 w=0.82u l=0.6u
X228 vdd a_31708_10216# a_31620_10260# vdd pmos_6p0 w=1.22u l=1u
X229 a_3620_47892# cap_shunt_p a_3828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X230 a_15512_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X231 a_7404_55688# a_7316_55732# vss vss nmos_6p0 w=0.82u l=1u
X232 vss tune_shunt[6] a_3828_40536# vss nmos_6p0 w=0.51u l=0.6u
X233 vdd a_32156_33736# a_32068_33780# vdd pmos_6p0 w=1.22u l=1u
X234 vss cap_shunt_p a_25984_43972# vss nmos_6p0 w=0.82u l=0.6u
X235 a_29744_15748# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X236 vdd tune_shunt[6] a_6532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X237 vdd a_19836_53687# a_19748_53784# vdd pmos_6p0 w=1.22u l=1u
X238 a_14908_53687# a_14820_53784# vss vss nmos_6p0 w=0.82u l=1u
X239 vdd a_33948_38440# a_33860_38484# vdd pmos_6p0 w=1.22u l=1u
X240 vdd tune_shunt[7] a_9668_21236# vdd pmos_6p0 w=1.2u l=0.5u
X241 vdd tune_shunt[6] a_28484_33780# vdd pmos_6p0 w=1.2u l=0.5u
X242 a_2500_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X243 a_6084_51028# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X244 a_20532_41620# cap_shunt_p a_20740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X245 a_15700_4834# cap_series_gyn a_16632_4772# vss nmos_6p0 w=0.82u l=0.6u
X246 a_3620_44756# cap_shunt_p a_3828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X247 a_14692_10744# cap_series_gyn a_14484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X248 a_24652_38440# a_24564_38484# vss vss nmos_6p0 w=0.82u l=1u
X249 vdd a_32156_30600# a_32068_30644# vdd pmos_6p0 w=1.22u l=1u
X250 vss cap_shunt_n a_14784_27992# vss nmos_6p0 w=0.82u l=0.6u
X251 vss cap_shunt_n a_25984_40836# vss nmos_6p0 w=0.82u l=0.6u
X252 a_32612_29922# cap_shunt_p a_32404_30268# vdd pmos_6p0 w=1.2u l=0.5u
X253 a_2500_49084# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X254 vdd tune_shunt[5] a_25572_40052# vdd pmos_6p0 w=1.2u l=0.5u
X255 a_10660_44034# cap_shunt_n a_10452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X256 a_8456_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X257 a_3828_43672# cap_shunt_p a_4760_43672# vss nmos_6p0 w=0.82u l=0.6u
X258 vdd tune_shunt[5] a_28484_30644# vdd pmos_6p0 w=1.2u l=0.5u
X259 vdd a_2140_17623# a_2052_17720# vdd pmos_6p0 w=1.22u l=1u
X260 vdd tune_shunt[4] a_13588_50652# vdd pmos_6p0 w=1.2u l=0.5u
X261 vdd a_36076_38007# a_35988_38104# vdd pmos_6p0 w=1.22u l=1u
X262 a_12788_17016# cap_shunt_p a_13720_17016# vss nmos_6p0 w=0.82u l=0.6u
X263 a_7748_36194# cap_shunt_n a_8680_36132# vss nmos_6p0 w=0.82u l=0.6u
X264 a_32612_36194# cap_shunt_n a_32404_36540# vdd pmos_6p0 w=1.2u l=0.5u
X265 vss cap_shunt_n a_14784_24856# vss nmos_6p0 w=0.82u l=0.6u
X266 a_7540_44380# cap_shunt_p a_7748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X267 a_11668_40536# cap_shunt_n a_11460_40052# vdd pmos_6p0 w=1.2u l=0.5u
X268 vdd tune_shunt[6] a_24452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X269 vdd a_34844_3944# a_34756_3988# vdd pmos_6p0 w=1.22u l=1u
X270 a_10660_40898# cap_shunt_n a_10452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X271 vdd a_14908_5079# a_14820_5176# vdd pmos_6p0 w=1.22u l=1u
X272 a_5636_3612# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X273 a_24660_44034# cap_shunt_p a_24452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X274 a_3828_40536# cap_shunt_n a_4760_40536# vss nmos_6p0 w=0.82u l=0.6u
X275 vdd tune_shunt[7] a_9332_9884# vdd pmos_6p0 w=1.2u l=0.5u
X276 a_3620_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X277 a_23632_4472# cap_series_gyn a_21524_4472# vss nmos_6p0 w=0.82u l=0.6u
X278 a_20740_18584# cap_shunt_p a_20532_18100# vdd pmos_6p0 w=1.2u l=0.5u
X279 a_32612_33058# cap_shunt_n a_32404_33404# vdd pmos_6p0 w=1.2u l=0.5u
X280 a_7540_41244# cap_shunt_n a_7748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X281 vdd tune_shunt[7] a_24452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X282 a_10548_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X283 a_30812_6647# a_30724_6744# vss vss nmos_6p0 w=0.82u l=1u
X284 vss cap_shunt_n a_5936_13880# vss nmos_6p0 w=0.82u l=0.6u
X285 vdd tune_series_gy[5] a_20532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X286 a_30812_20759# a_30724_20856# vss vss nmos_6p0 w=0.82u l=1u
X287 vdd a_32716_23895# a_32628_23992# vdd pmos_6p0 w=1.22u l=1u
X288 a_24660_40898# cap_shunt_n a_24452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X289 a_17828_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X290 a_31260_44279# a_31172_44376# vss vss nmos_6p0 w=0.82u l=1u
X291 a_17828_21720# cap_shunt_p a_19544_21720# vss nmos_6p0 w=0.82u l=0.6u
X292 vdd a_29916_55255# a_29828_55352# vdd pmos_6p0 w=1.22u l=1u
X293 a_21748_39330# cap_shunt_p a_21540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X294 vdd tune_shunt[2] a_1716_7124# vdd pmos_6p0 w=1.2u l=0.5u
X295 a_6760_7124# cap_series_gyp a_6572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X296 vss tune_series_gy[2] a_11780_4472# vss nmos_6p0 w=0.51u l=0.6u
X297 vdd tune_series_gy[0] a_28484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X298 a_27888_21720# cap_shunt_p a_25780_21720# vss nmos_6p0 w=0.82u l=0.6u
X299 a_33732_34264# cap_shunt_n a_33524_33780# vdd pmos_6p0 w=1.2u l=0.5u
X300 a_13796_18946# cap_shunt_p a_14728_18884# vss nmos_6p0 w=0.82u l=0.6u
X301 a_21672_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X302 a_11872_3204# cap_series_gyn a_10548_3266# vss nmos_6p0 w=0.82u l=0.6u
X303 vss tune_series_gy[5] a_21748_12674# vss nmos_6p0 w=0.51u l=0.6u
X304 a_9428_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X305 a_17828_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X306 a_35880_5556# cap_series_gygyn a_36688_6040# vss nmos_6p0 w=0.82u l=0.6u
X307 a_31260_41143# a_31172_41240# vss vss nmos_6p0 w=0.82u l=1u
X308 a_24452_9884# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X309 vdd a_29916_52119# a_29828_52216# vdd pmos_6p0 w=1.22u l=1u
X310 a_34844_50984# a_34756_51028# vss vss nmos_6p0 w=0.82u l=1u
X311 a_16500_27132# cap_shunt_n a_16708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X312 vss cap_series_gygyn a_34952_9476# vss nmos_6p0 w=0.82u l=0.6u
X313 a_29700_31490# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X314 a_33732_31128# cap_shunt_n a_33524_30644# vdd pmos_6p0 w=1.2u l=0.5u
X315 a_13796_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X316 a_6784_6040# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X317 a_13796_15810# cap_shunt_p a_14728_15748# vss nmos_6p0 w=0.82u l=0.6u
X318 a_21316_3988# cap_series_gyn a_21524_4472# vdd pmos_6p0 w=1.2u l=0.5u
X319 vss cap_shunt_p a_33936_29860# vss nmos_6p0 w=0.82u l=0.6u
X320 a_24452_6748# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X321 a_33732_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X322 a_21748_20514# cap_shunt_p a_23464_20452# vss nmos_6p0 w=0.82u l=0.6u
X323 a_13796_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X324 a_24540_3511# a_24452_3608# vss vss nmos_6p0 w=0.82u l=1u
X325 a_13788_10216# a_13700_10260# vss vss nmos_6p0 w=0.82u l=1u
X326 a_21540_14588# cap_series_gyn a_21748_14242# vdd pmos_6p0 w=1.2u l=0.5u
X327 vdd a_29468_47415# a_29380_47512# vdd pmos_6p0 w=1.22u l=1u
X328 vss tune_shunt[6] a_3828_34264# vss nmos_6p0 w=0.51u l=0.6u
X329 vdd tune_shunt[5] a_6084_18100# vdd pmos_6p0 w=1.2u l=0.5u
X330 a_31424_20152# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X331 vss cap_shunt_p a_33936_26724# vss nmos_6p0 w=0.82u l=0.6u
X332 a_12444_50984# a_12356_51028# vss vss nmos_6p0 w=0.82u l=1u
X333 vss tune_shunt[7] a_20740_23288# vss nmos_6p0 w=0.51u l=0.6u
X334 a_24360_13880# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X335 vss cap_shunt_n a_14112_49944# vss nmos_6p0 w=0.82u l=0.6u
X336 vss cap_shunt_p a_22848_17016# vss nmos_6p0 w=0.82u l=0.6u
X337 a_3620_38484# cap_shunt_n a_3828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X338 vss cap_shunt_p a_25984_34564# vss nmos_6p0 w=0.82u l=0.6u
X339 vss tune_shunt[7] a_3828_31128# vss nmos_6p0 w=0.51u l=0.6u
X340 vdd a_32156_24328# a_32068_24372# vdd pmos_6p0 w=1.22u l=1u
X341 vdd a_30028_52552# a_29940_52596# vdd pmos_6p0 w=1.22u l=1u
X342 vdd tune_shunt[7] a_6532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X343 a_34328_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X344 a_34308_13020# cap_series_gygyp a_34516_12674# vdd pmos_6p0 w=1.2u l=0.5u
X345 a_4380_54120# a_4292_54164# vss vss nmos_6p0 w=0.82u l=1u
X346 vdd tune_shunt[7] a_28484_24372# vdd pmos_6p0 w=1.2u l=0.5u
X347 a_24360_10744# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X348 vdd tune_shunt[6] a_13588_44380# vdd pmos_6p0 w=1.2u l=0.5u
X349 a_20532_32212# cap_shunt_n a_20740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X350 a_22456_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X351 a_3620_35348# cap_shunt_n a_3828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X352 vss cap_shunt_p a_25984_31428# vss nmos_6p0 w=0.82u l=0.6u
X353 a_22436_8692# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X354 vss cap_shunt_p a_8064_20152# vss nmos_6p0 w=0.82u l=0.6u
X355 a_34328_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X356 a_29492_36540# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X357 vss cap_shunt_n a_18816_22020# vss nmos_6p0 w=0.82u l=0.6u
X358 vdd tune_shunt[6] a_13588_41244# vdd pmos_6p0 w=1.2u l=0.5u
X359 a_20740_37400# cap_shunt_n a_21672_37400# vss nmos_6p0 w=0.82u l=0.6u
X360 a_3828_34264# cap_shunt_n a_4760_34264# vss nmos_6p0 w=0.82u l=0.6u
X361 a_6740_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X362 a_25572_25940# cap_shunt_p a_25780_26424# vdd pmos_6p0 w=1.2u l=0.5u
X363 a_32612_26786# cap_shunt_p a_32404_27132# vdd pmos_6p0 w=1.2u l=0.5u
X364 a_24452_8316# cap_series_gyp a_24660_7970# vdd pmos_6p0 w=1.2u l=0.5u
X365 vdd tune_shunt[7] a_24452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X366 a_3828_13880# cap_shunt_n a_3620_13396# vdd pmos_6p0 w=1.2u l=0.5u
X367 a_29492_33404# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X368 vss tune_series_gy[5] a_21748_15810# vss nmos_6p0 w=0.51u l=0.6u
X369 a_3828_31128# cap_shunt_n a_4760_31128# vss nmos_6p0 w=0.82u l=0.6u
X370 a_6740_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X371 a_25572_22804# cap_shunt_p a_25780_23288# vdd pmos_6p0 w=1.2u l=0.5u
X372 a_31436_22428# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X373 vdd a_29916_48983# a_29828_49080# vdd pmos_6p0 w=1.22u l=1u
X374 a_27228_38007# a_27140_38104# vss vss nmos_6p0 w=0.82u l=1u
X375 vss tune_shunt[6] a_25780_32696# vss nmos_6p0 w=0.51u l=0.6u
X376 a_35448_23588# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X377 vdd tune_shunt[7] a_24452_22428# vdd pmos_6p0 w=1.2u l=0.5u
X378 a_11780_4472# cap_series_gyp a_11572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X379 a_6084_51028# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X380 a_20532_41620# cap_shunt_p a_20740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X381 vdd tune_shunt[6] a_28484_33780# vdd pmos_6p0 w=1.2u l=0.5u
X382 a_12788_12312# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X383 vdd a_28124_41143# a_28036_41240# vdd pmos_6p0 w=1.22u l=1u
X384 vdd a_36748_33736# a_36660_33780# vdd pmos_6p0 w=1.22u l=1u
X385 a_9464_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X386 a_15804_13352# a_15716_13396# vss vss nmos_6p0 w=0.82u l=1u
X387 vss tune_series_gygy[5] a_35880_24372# vss nmos_6p0 w=0.51u l=0.6u
X388 a_17828_48376# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X389 a_4760_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X390 a_27888_12312# cap_series_gyp a_25780_12312# vss nmos_6p0 w=0.82u l=0.6u
X391 vdd a_31820_47848# a_31732_47892# vdd pmos_6p0 w=1.22u l=1u
X392 a_10660_44034# cap_shunt_n a_10452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X393 vdd tune_shunt[6] a_3620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X394 vdd a_26892_53687# a_26804_53784# vdd pmos_6p0 w=1.22u l=1u
X395 vdd tune_shunt[5] a_28484_30644# vdd pmos_6p0 w=1.2u l=0.5u
X396 vss cap_series_gyn a_19936_11044# vss nmos_6p0 w=0.82u l=0.6u
X397 a_21964_53687# a_21876_53784# vss vss nmos_6p0 w=0.82u l=1u
X398 vdd a_36748_30600# a_36660_30644# vdd pmos_6p0 w=1.22u l=1u
X399 a_17620_36916# cap_shunt_n a_17828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X400 a_9464_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X401 vdd tune_shunt[5] a_6084_52220# vdd pmos_6p0 w=1.2u l=0.5u
X402 a_7540_44380# cap_shunt_p a_7748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X403 a_21748_14242# cap_series_gyn a_23464_14180# vss nmos_6p0 w=0.82u l=0.6u
X404 a_4760_42104# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X405 a_34844_41576# a_34756_41620# vss vss nmos_6p0 w=0.82u l=1u
X406 a_11668_40536# cap_shunt_n a_11460_40052# vdd pmos_6p0 w=1.2u l=0.5u
X407 a_10660_40898# cap_shunt_n a_10452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X408 a_35736_6340# cap_series_gygyp a_34536_6748# vss nmos_6p0 w=0.82u l=0.6u
X409 vdd a_26892_50551# a_26804_50648# vdd pmos_6p0 w=1.22u l=1u
X410 a_33732_27992# cap_shunt_p a_33524_27508# vdd pmos_6p0 w=1.2u l=0.5u
X411 a_9220_20860# cap_shunt_p a_9428_20514# vdd pmos_6p0 w=1.2u l=0.5u
X412 a_10764_53687# a_10676_53784# vss vss nmos_6p0 w=0.82u l=1u
X413 a_21964_50551# a_21876_50648# vss vss nmos_6p0 w=0.82u l=1u
X414 a_18044_55255# a_17956_55352# vss vss nmos_6p0 w=0.82u l=1u
X415 a_10360_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X416 a_7540_41244# cap_shunt_n a_7748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X417 a_21748_11106# cap_series_gyn a_23464_11044# vss nmos_6p0 w=0.82u l=0.6u
X418 a_2140_19624# a_2052_19668# vss vss nmos_6p0 w=0.82u l=1u
X419 vdd tune_shunt[5] a_20532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X420 a_9540_11106# cap_shunt_p a_9332_11452# vdd pmos_6p0 w=1.2u l=0.5u
X421 a_34396_36872# a_34308_36916# vss vss nmos_6p0 w=0.82u l=1u
X422 vss cap_shunt_n a_25984_28292# vss nmos_6p0 w=0.82u l=0.6u
X423 a_34328_28292# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X424 vss tune_shunt[5] a_3828_48376# vss nmos_6p0 w=0.51u l=0.6u
X425 a_17828_42104# cap_shunt_n a_17620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X426 a_31708_52119# a_31620_52216# vss vss nmos_6p0 w=0.82u l=1u
X427 a_27228_6647# a_27140_6744# vss vss nmos_6p0 w=0.82u l=1u
X428 a_36688_13880# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X429 a_13588_17724# cap_shunt_p a_13796_17378# vdd pmos_6p0 w=1.2u l=0.5u
X430 vss cap_shunt_n a_22064_32696# vss nmos_6p0 w=0.82u l=0.6u
X431 a_3620_29076# cap_shunt_n a_3828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X432 a_34144_49080# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X433 a_14580_45240# cap_shunt_p a_16296_45240# vss nmos_6p0 w=0.82u l=0.6u
X434 a_25780_42104# cap_shunt_n a_27496_42104# vss nmos_6p0 w=0.82u l=0.6u
X435 vss cap_shunt_p a_25984_25156# vss nmos_6p0 w=0.82u l=0.6u
X436 vss tune_series_gy[2] a_10660_6402# vss nmos_6p0 w=0.51u l=0.6u
X437 a_29468_19191# a_29380_19288# vss vss nmos_6p0 w=0.82u l=1u
X438 a_11460_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X439 a_34328_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X440 a_31260_8648# a_31172_8692# vss vss nmos_6p0 w=0.82u l=1u
X441 a_6740_48376# cap_shunt_p a_6532_47892# vdd pmos_6p0 w=1.2u l=0.5u
X442 a_21748_39330# cap_shunt_p a_22680_39268# vss nmos_6p0 w=0.82u l=0.6u
X443 a_26712_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X444 vdd tune_shunt[7] a_17620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X445 a_13588_23996# cap_shunt_n a_13796_23650# vdd pmos_6p0 w=1.2u l=0.5u
X446 a_34516_23650# cap_series_gygyp a_36232_23588# vss nmos_6p0 w=0.82u l=0.6u
X447 a_36688_10744# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X448 a_31436_19292# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X449 a_9316_50306# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X450 a_34412_45540# cap_shunt_gyn a_34144_45540# vss nmos_6p0 w=0.82u l=0.6u
X451 vdd a_33612_5079# a_33524_5176# vdd pmos_6p0 w=1.22u l=1u
X452 a_14580_42104# cap_shunt_n a_16296_42104# vss nmos_6p0 w=0.82u l=0.6u
X453 vdd tune_series_gy[4] a_24452_19292# vdd pmos_6p0 w=1.2u l=0.5u
X454 vss cap_shunt_n a_11200_51512# vss nmos_6p0 w=0.82u l=0.6u
X455 a_13796_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X456 vss tune_shunt[6] a_25780_35832# vss nmos_6p0 w=0.51u l=0.6u
X457 vss tune_shunt[7] a_13460_34264# vss nmos_6p0 w=0.51u l=0.6u
X458 a_29492_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X459 vss cap_shunt_p a_11536_17316# vss nmos_6p0 w=0.82u l=0.6u
X460 vss cap_shunt_p a_14896_20152# vss nmos_6p0 w=0.82u l=0.6u
X461 a_6740_45240# cap_shunt_p a_6532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X462 vss tune_shunt[7] a_3380_17016# vss nmos_6p0 w=0.51u l=0.6u
X463 a_15512_43672# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X464 vdd tune_shunt[5] a_6084_18100# vdd pmos_6p0 w=1.2u l=0.5u
X465 a_6292_18584# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X466 vdd a_33948_55255# a_33860_55352# vdd pmos_6p0 w=1.22u l=1u
X467 a_18424_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X468 a_34412_42404# cap_shunt_gyn a_34144_42404# vss nmos_6p0 w=0.82u l=0.6u
X469 a_26712_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X470 a_25572_16532# cap_series_gyp a_25780_17016# vdd pmos_6p0 w=1.2u l=0.5u
X471 vdd a_10876_55688# a_10788_55732# vdd pmos_6p0 w=1.22u l=1u
X472 a_2500_13020# cap_shunt_n a_2708_12674# vdd pmos_6p0 w=1.2u l=0.5u
X473 vdd tune_series_gy[5] a_24452_16156# vdd pmos_6p0 w=1.2u l=0.5u
X474 vss tune_shunt[7] a_13460_31128# vss nmos_6p0 w=0.51u l=0.6u
X475 a_23308_35304# a_23220_35348# vss vss nmos_6p0 w=0.82u l=1u
X476 a_15512_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X477 vss tune_series_gygy[5] a_35880_18100# vss nmos_6p0 w=0.51u l=0.6u
X478 vdd a_33948_52119# a_33860_52216# vdd pmos_6p0 w=1.22u l=1u
X479 a_18424_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X480 a_6740_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X481 a_14372_46324# cap_shunt_p a_14580_46808# vdd pmos_6p0 w=1.2u l=0.5u
X482 a_34308_13020# cap_series_gygyp a_34516_12674# vdd pmos_6p0 w=1.2u l=0.5u
X483 vss tune_shunt[7] a_25780_23288# vss nmos_6p0 w=0.51u l=0.6u
X484 vss tune_shunt[4] a_13796_50306# vss nmos_6p0 w=0.51u l=0.6u
X485 a_33920_44757# cap_shunt_gyn a_33920_45302# vdd pmos_6p0 w=1.215u l=0.5u
X486 vdd tune_shunt[7] a_28484_24372# vdd pmos_6p0 w=1.2u l=0.5u
X487 a_2708_18946# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X488 vdd a_26444_52552# a_26356_52596# vdd pmos_6p0 w=1.22u l=1u
X489 a_20532_32212# cap_shunt_n a_20740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X490 a_5544_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X491 a_9540_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X492 vss cap_shunt_n a_35840_32696# vss nmos_6p0 w=0.82u l=0.6u
X493 a_19152_35832# cap_shunt_n a_17828_35832# vss nmos_6p0 w=0.82u l=0.6u
X494 vss tune_series_gygy[4] a_35880_14964# vss nmos_6p0 w=0.51u l=0.6u
X495 a_12556_12919# a_12468_13016# vss vss nmos_6p0 w=0.82u l=1u
X496 vdd tune_shunt[7] a_3620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X497 a_31024_29860# cap_shunt_p a_29700_29922# vss nmos_6p0 w=0.82u l=0.6u
X498 vdd tune_series_gy[1] a_7580_5180# vdd pmos_6p0 w=1.2u l=0.5u
X499 a_5544_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X500 a_9540_11106# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X501 a_12788_18584# cap_shunt_p a_12580_18100# vdd pmos_6p0 w=1.2u l=0.5u
X502 a_17620_27508# cap_shunt_n a_17828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X503 a_21748_45602# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X504 vdd tune_shunt[6] a_20532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X505 a_29700_23650# cap_shunt_p a_29492_23996# vdd pmos_6p0 w=1.2u l=0.5u
X506 a_35292_55688# a_35204_55732# vss vss nmos_6p0 w=0.82u l=1u
X507 a_31024_26724# cap_shunt_p a_29700_26786# vss nmos_6p0 w=0.82u l=0.6u
X508 a_21840_9176# cap_series_gyp a_19732_9176# vss nmos_6p0 w=0.82u l=0.6u
X509 a_31436_22428# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X510 a_9876_17016# cap_shunt_p a_11592_17016# vss nmos_6p0 w=0.82u l=0.6u
X511 a_9220_17724# cap_shunt_p a_9428_17378# vdd pmos_6p0 w=1.2u l=0.5u
X512 a_18612_4834# cap_series_gyp a_20328_4772# vss nmos_6p0 w=0.82u l=0.6u
X513 vss cap_shunt_p a_31808_39268# vss nmos_6p0 w=0.82u l=0.6u
X514 a_25780_34264# cap_shunt_p a_25572_33780# vdd pmos_6p0 w=1.2u l=0.5u
X515 a_3172_51028# cap_shunt_n a_3380_51512# vdd pmos_6p0 w=1.2u l=0.5u
X516 a_9316_47170# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X517 vdd tune_shunt[6] a_20532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X518 a_24660_7970# cap_series_gyp a_24452_8316# vdd pmos_6p0 w=1.2u l=0.5u
X519 a_16708_33058# cap_shunt_n a_18424_32996# vss nmos_6p0 w=0.82u l=0.6u
X520 a_8412_8648# a_8324_8692# vss vss nmos_6p0 w=0.82u l=1u
X521 vdd tune_series_gy[5] a_21540_13020# vdd pmos_6p0 w=1.2u l=0.5u
X522 a_10540_8648# a_10452_8692# vss vss nmos_6p0 w=0.82u l=1u
X523 a_10548_37400# cap_shunt_n a_10340_36916# vdd pmos_6p0 w=1.2u l=0.5u
X524 a_26768_32996# cap_shunt_p a_24660_33058# vss nmos_6p0 w=0.82u l=0.6u
X525 a_32268_55688# a_32180_55732# vss vss nmos_6p0 w=0.82u l=1u
X526 vdd tune_shunt_gy[4] a_31060_44757# vdd pmos_6p0 w=1.215u l=0.5u
X527 vdd a_34396_7080# a_34308_7124# vdd pmos_6p0 w=1.22u l=1u
X528 a_31708_42711# a_31620_42808# vss vss nmos_6p0 w=0.82u l=1u
X529 a_17828_32696# cap_shunt_n a_17620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X530 a_32464_46325# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X531 vdd a_31484_41576# a_31396_41620# vdd pmos_6p0 w=1.22u l=1u
X532 vss tune_shunt[7] a_13460_37400# vss nmos_6p0 w=0.51u l=0.6u
X533 a_25780_31128# cap_shunt_p a_25572_30644# vdd pmos_6p0 w=1.2u l=0.5u
X534 vdd tune_shunt[6] a_9668_47892# vdd pmos_6p0 w=1.2u l=0.5u
X535 a_35600_47893# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X536 vss cap_shunt_n a_4032_37700# vss nmos_6p0 w=0.82u l=0.6u
X537 vss cap_shunt_p a_22064_23288# vss nmos_6p0 w=0.82u l=0.6u
X538 vdd a_18492_13352# a_18404_13396# vdd pmos_6p0 w=1.22u l=1u
X539 a_3620_47892# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X540 vdd tune_shunt[5] a_6084_52220# vdd pmos_6p0 w=1.2u l=0.5u
X541 a_21748_34626# cap_shunt_p a_21540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X542 vss tune_series_gy[4] a_22644_7608# vss nmos_6p0 w=0.51u l=0.6u
X543 a_33164_5079# a_33076_5176# vss vss nmos_6p0 w=0.82u l=1u
X544 vss tune_shunt[7] a_25780_29560# vss nmos_6p0 w=0.51u l=0.6u
X545 a_6740_38968# cap_shunt_n a_6532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X546 a_13588_14588# cap_shunt_p a_13796_14242# vdd pmos_6p0 w=1.2u l=0.5u
X547 a_26712_34264# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X548 vdd tune_shunt[7] a_17620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X549 a_33732_27992# cap_shunt_p a_33524_27508# vdd pmos_6p0 w=1.2u l=0.5u
X550 vss cap_shunt_p a_7952_14180# vss nmos_6p0 w=0.82u l=0.6u
X551 a_3620_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X552 vdd tune_shunt[2] a_1716_5556# vdd pmos_6p0 w=1.2u l=0.5u
X553 a_7852_55688# a_7764_55732# vss vss nmos_6p0 w=0.82u l=1u
X554 vss tune_shunt[6] a_13796_47170# vss nmos_6p0 w=0.51u l=0.6u
X555 a_21748_31490# cap_shunt_n a_21540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X556 vss tune_shunt[7] a_25780_26424# vss nmos_6p0 w=0.51u l=0.6u
X557 a_11612_7124# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X558 a_1924_3266# cap_shunt_n a_1716_3612# vdd pmos_6p0 w=1.2u l=0.5u
X559 a_13460_21720# cap_shunt_n a_14392_21720# vss nmos_6p0 w=0.82u l=0.6u
X560 vdd a_32156_41143# a_32068_41240# vdd pmos_6p0 w=1.22u l=1u
X561 a_6740_35832# cap_shunt_n a_6532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X562 a_12216_9176# cap_series_gyp a_11800_8692# vss nmos_6p0 w=0.82u l=0.6u
X563 a_23308_29032# a_23220_29076# vss vss nmos_6p0 w=0.82u l=1u
X564 vdd a_14124_54120# a_14036_54164# vdd pmos_6p0 w=1.22u l=1u
X565 a_18424_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X566 a_26712_31128# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X567 vdd tune_shunt[7] a_2500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X568 a_11780_6040# cap_series_gyn a_13496_6040# vss nmos_6p0 w=0.82u l=0.6u
X569 a_32604_5512# a_32516_5556# vss vss nmos_6p0 w=0.82u l=1u
X570 vss cap_shunt_n a_7952_11044# vss nmos_6p0 w=0.82u l=0.6u
X571 a_22188_47848# a_22100_47892# vss vss nmos_6p0 w=0.82u l=1u
X572 vdd tune_shunt[4] a_32404_36540# vdd pmos_6p0 w=1.2u l=0.5u
X573 vdd a_2140_25896# a_2052_25940# vdd pmos_6p0 w=1.22u l=1u
X574 a_25780_13880# cap_series_gyn a_26712_13880# vss nmos_6p0 w=0.82u l=0.6u
X575 vss tune_shunt[6] a_13796_44034# vss nmos_6p0 w=0.51u l=0.6u
X576 a_4828_55688# a_4740_55732# vss vss nmos_6p0 w=0.82u l=1u
X577 a_16500_47516# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X578 a_13588_17724# cap_shunt_p a_13796_17378# vdd pmos_6p0 w=1.2u l=0.5u
X579 vdd a_27340_47415# a_27252_47512# vdd pmos_6p0 w=1.22u l=1u
X580 a_23308_25896# a_23220_25940# vss vss nmos_6p0 w=0.82u l=1u
X581 vdd a_14908_11351# a_14820_11448# vdd pmos_6p0 w=1.22u l=1u
X582 a_19152_29560# cap_shunt_n a_17828_29560# vss nmos_6p0 w=0.82u l=0.6u
X583 vdd tune_shunt[7] a_9332_9884# vdd pmos_6p0 w=1.2u l=0.5u
X584 vdd tune_shunt[4] a_32404_33404# vdd pmos_6p0 w=1.2u l=0.5u
X585 vdd a_2140_22760# a_2052_22804# vdd pmos_6p0 w=1.22u l=1u
X586 a_25780_10744# cap_series_gyn a_26712_10744# vss nmos_6p0 w=0.82u l=0.6u
X587 a_6740_48376# cap_shunt_p a_6532_47892# vdd pmos_6p0 w=1.2u l=0.5u
X588 a_35692_13396# cap_series_gygyn a_35880_13396# vdd pmos_6p0 w=1.2u l=0.5u
X589 a_31436_19292# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X590 a_3828_20152# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X591 a_21540_38108# cap_shunt_n a_21748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X592 a_35692_19668# cap_series_gygyp a_35880_19668# vdd pmos_6p0 w=1.2u l=0.5u
X593 a_12376_43972# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X594 a_17620_25940# cap_shunt_n a_17828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X595 vss tune_series_gy[3] a_25780_6040# vss nmos_6p0 w=0.51u l=0.6u
X596 a_7168_3204# cap_shunt_n a_5844_3266# vss nmos_6p0 w=0.82u l=0.6u
X597 vdd a_1692_13352# a_1604_13396# vdd pmos_6p0 w=1.22u l=1u
X598 a_6292_17378# cap_shunt_p a_7224_17316# vss nmos_6p0 w=0.82u l=0.6u
X599 a_31624_20860# cap_series_gygyn a_31648_20452# vss nmos_6p0 w=0.82u l=0.6u
X600 a_17620_47892# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X601 a_3828_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X602 a_21748_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X603 a_19152_26424# cap_shunt_n a_17828_26424# vss nmos_6p0 w=0.82u l=0.6u
X604 a_16252_18056# a_16164_18100# vss vss nmos_6p0 w=0.82u l=1u
X605 a_6740_45240# cap_shunt_p a_6532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X606 a_13776_46808# cap_shunt_n a_11668_46808# vss nmos_6p0 w=0.82u l=0.6u
X607 a_21316_3612# cap_series_gyp a_21524_3266# vdd pmos_6p0 w=1.2u l=0.5u
X608 a_5544_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X609 a_3380_18584# cap_shunt_p a_3172_18100# vdd pmos_6p0 w=1.2u l=0.5u
X610 a_10548_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X611 a_1924_7608# cap_shunt_n a_1716_7124# vdd pmos_6p0 w=1.2u l=0.5u
X612 a_12376_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X613 a_17620_22804# cap_shunt_n a_17828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X614 vdd tune_series_gy[2] a_6572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X615 a_19524_11828# cap_series_gyn a_19732_12312# vdd pmos_6p0 w=1.2u l=0.5u
X616 a_2500_13020# cap_shunt_n a_2708_12674# vdd pmos_6p0 w=1.2u l=0.5u
X617 a_32632_14588# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X618 a_17620_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X619 a_3828_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X620 a_18156_50551# a_18068_50648# vss vss nmos_6p0 w=0.82u l=1u
X621 vdd a_37196_35304# a_37108_35348# vdd pmos_6p0 w=1.22u l=1u
X622 a_29700_14242# cap_series_gyp a_29492_14588# vdd pmos_6p0 w=1.2u l=0.5u
X623 vdd tune_shunt[7] a_20532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X624 a_16252_14920# a_16164_14964# vss vss nmos_6p0 w=0.82u l=1u
X625 vss cap_shunt_p a_19936_43672# vss nmos_6p0 w=0.82u l=0.6u
X626 a_13460_32696# cap_shunt_n a_13252_32212# vdd pmos_6p0 w=1.2u l=0.5u
X627 vdd a_33500_41576# a_33412_41620# vdd pmos_6p0 w=1.22u l=1u
X628 a_31024_17316# cap_series_gyp a_29700_17378# vss nmos_6p0 w=0.82u l=0.6u
X629 a_6532_52596# cap_shunt_n a_6740_53080# vdd pmos_6p0 w=1.2u l=0.5u
X630 a_14372_46324# cap_shunt_p a_14580_46808# vdd pmos_6p0 w=1.2u l=0.5u
X631 a_32632_11452# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X632 a_15176_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X633 vdd tune_shunt[1] a_25236_3612# vdd pmos_6p0 w=1.2u l=0.5u
X634 a_20720_9476# cap_series_gyp a_18612_9538# vss nmos_6p0 w=0.82u l=0.6u
X635 a_25780_24856# cap_shunt_p a_25572_24372# vdd pmos_6p0 w=1.2u l=0.5u
X636 vdd tune_shunt[4] a_29492_39676# vdd pmos_6p0 w=1.2u l=0.5u
X637 vdd a_16812_12919# a_16724_13016# vdd pmos_6p0 w=1.22u l=1u
X638 vss cap_shunt_n a_19936_40536# vss nmos_6p0 w=0.82u l=0.6u
X639 a_16708_23650# cap_shunt_n a_18424_23588# vss nmos_6p0 w=0.82u l=0.6u
X640 a_10548_27992# cap_shunt_n a_10340_27508# vdd pmos_6p0 w=1.2u l=0.5u
X641 a_26768_23588# cap_shunt_p a_24660_23650# vss nmos_6p0 w=0.82u l=0.6u
X642 a_13796_34626# cap_shunt_n a_13588_34972# vdd pmos_6p0 w=1.2u l=0.5u
X643 a_4380_53687# a_4292_53784# vss vss nmos_6p0 w=0.82u l=1u
X644 a_10548_3266# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X645 vss cap_shunt_p a_5152_48376# vss nmos_6p0 w=0.82u l=0.6u
X646 a_15176_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X647 a_24452_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X648 a_14260_3612# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X649 a_25780_21720# cap_shunt_p a_25572_21236# vdd pmos_6p0 w=1.2u l=0.5u
X650 a_22644_9176# cap_series_gyp a_24360_9176# vss nmos_6p0 w=0.82u l=0.6u
X651 a_3620_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X652 a_37420_30167# a_37332_30264# vss vss nmos_6p0 w=0.82u l=1u
X653 vdd tune_series_gy[4] a_25572_19668# vdd pmos_6p0 w=1.2u l=0.5u
X654 a_21748_25218# cap_shunt_n a_21540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X655 a_13796_31490# cap_shunt_n a_13588_31836# vdd pmos_6p0 w=1.2u l=0.5u
X656 vdd a_18268_55688# a_18180_55732# vdd pmos_6p0 w=1.22u l=1u
X657 a_3828_43672# cap_shunt_p a_3620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X658 a_6740_29560# cap_shunt_n a_6532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X659 a_29700_23650# cap_shunt_p a_29492_23996# vdd pmos_6p0 w=1.2u l=0.5u
X660 a_31624_8316# tune_series_gygy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X661 vdd a_19836_52552# a_19748_52596# vdd pmos_6p0 w=1.22u l=1u
X662 vss tune_shunt_gy[4] a_31248_44757# vss nmos_6p0 w=0.51u l=0.6u
X663 a_28484_10260# cap_series_gyp a_28692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X664 a_9220_17724# cap_shunt_p a_9428_17378# vdd pmos_6p0 w=1.2u l=0.5u
X665 a_12892_50984# a_12804_51028# vss vss nmos_6p0 w=0.82u l=1u
X666 a_3036_44712# a_2948_44756# vss vss nmos_6p0 w=0.82u l=1u
X667 a_3620_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X668 a_37420_27031# a_37332_27128# vss vss nmos_6p0 w=0.82u l=1u
X669 vss tune_shunt[3] a_5844_9176# vss nmos_6p0 w=0.51u l=0.6u
X670 vss cap_shunt_p a_15904_47108# vss nmos_6p0 w=0.82u l=0.6u
X671 a_21748_22082# cap_shunt_p a_21540_22428# vdd pmos_6p0 w=1.2u l=0.5u
X672 vss cap_series_gygyn a_32824_6340# vss nmos_6p0 w=0.82u l=0.6u
X673 a_25780_34264# cap_shunt_p a_25572_33780# vdd pmos_6p0 w=1.2u l=0.5u
X674 a_3172_51028# cap_shunt_n a_3380_51512# vdd pmos_6p0 w=1.2u l=0.5u
X675 vss tune_series_gy[5] a_25780_17016# vss nmos_6p0 w=0.51u l=0.6u
X676 vdd a_30476_52552# a_30388_52596# vdd pmos_6p0 w=1.22u l=1u
X677 a_21748_12674# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X678 a_8400_50244# cap_shunt_p a_6292_50306# vss nmos_6p0 w=0.82u l=0.6u
X679 a_10548_37400# cap_shunt_n a_10340_36916# vdd pmos_6p0 w=1.2u l=0.5u
X680 a_25780_9176# cap_series_gyp a_25572_8692# vdd pmos_6p0 w=1.2u l=0.5u
X681 a_22436_8692# cap_series_gyp a_22644_9176# vdd pmos_6p0 w=1.2u l=0.5u
X682 a_3036_41576# a_2948_41620# vss vss nmos_6p0 w=0.82u l=1u
X683 vdd tune_shunt[7] a_32404_27132# vdd pmos_6p0 w=1.2u l=0.5u
X684 vdd a_2140_16488# a_2052_16532# vdd pmos_6p0 w=1.22u l=1u
X685 a_3828_46808# cap_shunt_p a_3620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X686 a_15700_9538# cap_series_gyn a_15492_9884# vdd pmos_6p0 w=1.2u l=0.5u
X687 a_25780_31128# cap_shunt_p a_25572_30644# vdd pmos_6p0 w=1.2u l=0.5u
X688 a_10660_6402# cap_series_gyn a_12376_6340# vss nmos_6p0 w=0.82u l=0.6u
X689 a_16500_38108# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X690 a_24452_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X691 a_23308_16488# a_23220_16532# vss vss nmos_6p0 w=0.82u l=1u
X692 a_6404_22082# cap_shunt_p a_7336_22020# vss nmos_6p0 w=0.82u l=0.6u
X693 a_25780_6040# cap_series_gyp a_25572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X694 vss tune_shunt[7] a_16708_18946# vss nmos_6p0 w=0.51u l=0.6u
X695 a_6740_38968# cap_shunt_n a_6532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X696 a_15700_6402# cap_series_gyp a_15492_6748# vdd pmos_6p0 w=1.2u l=0.5u
X697 a_12376_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X698 a_17620_16532# cap_shunt_p a_17828_17016# vdd pmos_6p0 w=1.2u l=0.5u
X699 a_3828_34264# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X700 a_10988_43144# a_10900_43188# vss vss nmos_6p0 w=0.82u l=1u
X701 a_17620_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X702 a_19152_17016# cap_shunt_p a_17828_17016# vss nmos_6p0 w=0.82u l=0.6u
X703 vdd a_37196_29032# a_37108_29076# vdd pmos_6p0 w=1.22u l=1u
X704 a_27676_38007# a_27588_38104# vss vss nmos_6p0 w=0.82u l=1u
X705 a_6740_35832# cap_shunt_n a_6532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X706 a_17828_43672# cap_shunt_p a_17620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X707 vdd tune_shunt[7] a_2500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X708 vdd a_28572_5079# a_28484_5176# vdd pmos_6p0 w=1.22u l=1u
X709 vdd tune_shunt_gy[5] a_32740_45944# vdd pmos_6p0 w=1.215u l=0.5u
X710 a_12376_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X711 vdd a_28572_41143# a_28484_41240# vdd pmos_6p0 w=1.22u l=1u
X712 a_3828_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X713 a_9668_52596# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X714 a_10988_40008# a_10900_40052# vss vss nmos_6p0 w=0.82u l=1u
X715 a_17620_35348# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X716 a_35692_24372# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X717 a_36188_40008# a_36100_40052# vss vss nmos_6p0 w=0.82u l=1u
X718 vdd a_35292_14920# a_35204_14964# vdd pmos_6p0 w=1.22u l=1u
X719 a_29492_39676# cap_shunt_p a_29700_39330# vdd pmos_6p0 w=1.2u l=0.5u
X720 vss cap_shunt_n a_19936_34264# vss nmos_6p0 w=0.82u l=0.6u
X721 a_6532_43188# cap_shunt_p a_6740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X722 vdd tune_shunt[6] a_7540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X723 vdd a_21180_54120# a_21092_54164# vdd pmos_6p0 w=1.22u l=1u
X724 a_33732_34264# cap_shunt_n a_34664_34264# vss nmos_6p0 w=0.82u l=0.6u
X725 a_8064_27992# cap_shunt_n a_6740_27992# vss nmos_6p0 w=0.82u l=0.6u
X726 a_25780_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X727 a_27340_52552# a_27252_52596# vss vss nmos_6p0 w=0.82u l=1u
X728 a_35692_21236# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X729 a_37868_55255# a_37780_55352# vss vss nmos_6p0 w=0.82u l=1u
X730 vdd a_2588_47848# a_2500_47892# vdd pmos_6p0 w=1.22u l=1u
X731 vdd a_35292_11784# a_35204_11828# vdd pmos_6p0 w=1.22u l=1u
X732 vss cap_shunt_n a_5040_12312# vss nmos_6p0 w=0.82u l=0.6u
X733 vss cap_shunt_n a_19936_31128# vss nmos_6p0 w=0.82u l=0.6u
X734 a_1924_4472# cap_shunt_p a_2856_4472# vss nmos_6p0 w=0.82u l=0.6u
X735 vdd tune_shunt[7] a_13252_25940# vdd pmos_6p0 w=1.2u l=0.5u
X736 a_13796_25218# cap_shunt_n a_13588_25564# vdd pmos_6p0 w=1.2u l=0.5u
X737 vss tune_series_gy[3] a_10680_8316# vss nmos_6p0 w=0.51u l=0.6u
X738 a_21748_18946# cap_shunt_p a_21540_19292# vdd pmos_6p0 w=1.2u l=0.5u
X739 vdd a_18044_8648# a_17956_8692# vdd pmos_6p0 w=1.22u l=1u
X740 a_30428_21236# cap_series_gygyn a_30616_21236# vdd pmos_6p0 w=1.2u l=0.5u
X741 vdd a_21180_50984# a_21092_51028# vdd pmos_6p0 w=1.22u l=1u
X742 a_33732_31128# cap_shunt_n a_34664_31128# vss nmos_6p0 w=0.82u l=0.6u
X743 vdd tune_shunt[7] a_3620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X744 a_18492_55255# a_18404_55352# vss vss nmos_6p0 w=0.82u l=1u
X745 a_8064_24856# cap_shunt_p a_6740_24856# vss nmos_6p0 w=0.82u l=0.6u
X746 a_3380_18584# cap_shunt_p a_3172_18100# vdd pmos_6p0 w=1.2u l=0.5u
X747 a_24316_52552# a_24228_52596# vss vss nmos_6p0 w=0.82u l=1u
X748 a_32156_47415# a_32068_47512# vss vss nmos_6p0 w=0.82u l=1u
X749 vdd a_2588_44712# a_2500_44756# vdd pmos_6p0 w=1.22u l=1u
X750 a_33024_44376# cap_shunt_gyn a_33024_43972# vdd pmos_6p0 w=1.215u l=0.5u
X751 a_3620_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X752 vdd tune_shunt[7] a_13252_22804# vdd pmos_6p0 w=1.2u l=0.5u
X753 a_13796_22082# cap_shunt_n a_13588_22428# vdd pmos_6p0 w=1.2u l=0.5u
X754 vss tune_series_gy[3] a_14692_4472# vss nmos_6p0 w=0.51u l=0.6u
X755 a_21748_15810# cap_series_gyn a_21540_16156# vdd pmos_6p0 w=1.2u l=0.5u
X756 vdd a_18044_5512# a_17956_5556# vdd pmos_6p0 w=1.22u l=1u
X757 a_20664_12312# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X758 a_29700_14242# cap_series_gyp a_29492_14588# vdd pmos_6p0 w=1.2u l=0.5u
X759 a_10548_34264# cap_shunt_n a_12264_34264# vss nmos_6p0 w=0.82u l=0.6u
X760 vdd a_37868_30167# a_37780_30264# vdd pmos_6p0 w=1.22u l=1u
X761 vdd tune_shunt[7] a_3620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X762 a_7568_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X763 a_13460_32696# cap_shunt_n a_13252_32212# vdd pmos_6p0 w=1.2u l=0.5u
X764 a_9644_8648# a_9556_8692# vss vss nmos_6p0 w=0.82u l=1u
X765 a_13720_49944# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X766 a_33500_24328# a_33412_24372# vss vss nmos_6p0 w=0.82u l=1u
X767 a_6532_52596# cap_shunt_n a_6740_53080# vdd pmos_6p0 w=1.2u l=0.5u
X768 a_37420_17623# a_37332_17720# vss vss nmos_6p0 w=0.82u l=1u
X769 a_10452_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X770 a_19524_7124# cap_series_gyp a_19732_7608# vdd pmos_6p0 w=1.2u l=0.5u
X771 a_33832_14180# cap_series_gyp a_32632_14588# vss nmos_6p0 w=0.82u l=0.6u
X772 a_20620_33303# a_20532_33400# vss vss nmos_6p0 w=0.82u l=1u
X773 a_25780_24856# cap_shunt_p a_25572_24372# vdd pmos_6p0 w=1.2u l=0.5u
X774 a_28484_3988# cap_series_gyp a_28692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X775 a_10548_31128# cap_shunt_n a_12264_31128# vss nmos_6p0 w=0.82u l=0.6u
X776 a_12108_9783# a_12020_9880# vss vss nmos_6p0 w=0.82u l=1u
X777 vss tune_shunt[7] a_10548_27992# vss nmos_6p0 w=0.51u l=0.6u
X778 a_29700_4834# cap_shunt_p a_29492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X779 a_16800_9176# cap_series_gyn a_14692_9176# vss nmos_6p0 w=0.82u l=0.6u
X780 a_8008_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X781 vdd a_20172_47415# a_20084_47512# vdd pmos_6p0 w=1.22u l=1u
X782 a_13796_34626# cap_shunt_n a_13588_34972# vdd pmos_6p0 w=1.2u l=0.5u
X783 a_10548_27992# cap_shunt_n a_10340_27508# vdd pmos_6p0 w=1.2u l=0.5u
X784 a_11480_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X785 a_33832_11044# cap_series_gyp a_32632_11452# vss nmos_6p0 w=0.82u l=0.6u
X786 a_2500_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X787 a_21540_28700# cap_shunt_n a_21748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X788 a_1924_7608# cap_shunt_n a_1716_7124# vdd pmos_6p0 w=1.2u l=0.5u
X789 a_25780_21720# cap_shunt_p a_25572_21236# vdd pmos_6p0 w=1.2u l=0.5u
X790 a_12376_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X791 vss tune_shunt[7] a_10548_24856# vss nmos_6p0 w=0.51u l=0.6u
X792 a_8008_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X793 a_30408_27992# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X794 a_13796_31490# cap_shunt_n a_13588_31836# vdd pmos_6p0 w=1.2u l=0.5u
X795 a_9540_12674# cap_shunt_p a_11256_12612# vss nmos_6p0 w=0.82u l=0.6u
X796 vdd a_33612_17623# a_33524_17720# vdd pmos_6p0 w=1.22u l=1u
X797 a_6740_29560# cap_shunt_n a_6532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X798 a_30616_21236# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X799 a_1692_55255# a_1604_55352# vss vss nmos_6p0 w=0.82u l=1u
X800 vss tune_shunt[7] a_13796_23650# vss nmos_6p0 w=0.51u l=0.6u
X801 a_35880_5556# cap_series_gygyn a_35904_6040# vss nmos_6p0 w=0.82u l=0.6u
X802 vdd tune_series_gy[4] a_14484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X803 a_28484_10260# cap_series_gyp a_28692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X804 a_12376_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X805 a_5152_21720# cap_shunt_p a_3828_21720# vss nmos_6p0 w=0.82u l=0.6u
X806 a_12580_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X807 a_17620_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X808 a_30408_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X809 a_36100_39672# cap_shunt_gyn a_36288_39672# vdd pmos_6p0 w=1.215u l=0.5u
X810 a_23756_35304# a_23668_35348# vss vss nmos_6p0 w=0.82u l=1u
X811 a_29700_36194# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X812 a_6292_49944# cap_shunt_p a_7224_49944# vss nmos_6p0 w=0.82u l=0.6u
X813 vdd tune_series_gy[3] a_14484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X814 vss tune_shunt[7] a_13796_20514# vss nmos_6p0 w=0.51u l=0.6u
X815 vdd tune_series_gygy[5] a_34308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X816 vdd a_26892_52552# a_26804_52596# vdd pmos_6p0 w=1.22u l=1u
X817 a_32612_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X818 a_15624_6040# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X819 a_18612_12674# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X820 a_29700_36194# cap_shunt_n a_31416_36132# vss nmos_6p0 w=0.82u l=0.6u
X821 a_4816_29860# cap_shunt_n a_2708_29922# vss nmos_6p0 w=0.82u l=0.6u
X822 vss cap_shunt_p a_7616_48676# vss nmos_6p0 w=0.82u l=0.6u
X823 vdd a_1692_30167# a_1604_30264# vdd pmos_6p0 w=1.22u l=1u
X824 a_1924_7970# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X825 a_16708_48738# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X826 vdd a_20620_48983# a_20532_49080# vdd pmos_6p0 w=1.22u l=1u
X827 a_29700_33058# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X828 a_13796_18946# cap_shunt_p a_13588_19292# vdd pmos_6p0 w=1.2u l=0.5u
X829 a_28484_32212# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X830 a_25780_12312# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X831 a_35880_36916# cap_series_gygyp a_35692_36916# vdd pmos_6p0 w=1.2u l=0.5u
X832 a_32432_6340# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X833 vdd a_23868_52552# a_23780_52596# vdd pmos_6p0 w=1.22u l=1u
X834 a_13796_44034# cap_shunt_n a_14728_43972# vss nmos_6p0 w=0.82u l=0.6u
X835 a_29408_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X836 vdd a_2588_38440# a_2500_38484# vdd pmos_6p0 w=1.22u l=1u
X837 a_4816_26724# cap_shunt_p a_2708_26786# vss nmos_6p0 w=0.82u l=0.6u
X838 vdd a_16700_19624# a_16612_19668# vdd pmos_6p0 w=1.22u l=1u
X839 a_17620_40052# cap_shunt_n a_17828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X840 a_9856_39268# cap_shunt_n a_7748_39330# vss nmos_6p0 w=0.82u l=0.6u
X841 a_1924_4834# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X842 a_34720_34564# cap_shunt_n a_32612_34626# vss nmos_6p0 w=0.82u l=0.6u
X843 a_37868_9783# a_37780_9880# vss vss nmos_6p0 w=0.82u l=1u
X844 a_13796_15810# cap_shunt_p a_13588_16156# vdd pmos_6p0 w=1.2u l=0.5u
X845 a_10660_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X846 a_33948_7080# a_33860_7124# vss vss nmos_6p0 w=0.82u l=1u
X847 a_8064_15448# cap_shunt_p a_6740_15448# vss nmos_6p0 w=0.82u l=0.6u
X848 a_13796_40898# cap_shunt_n a_14728_40836# vss nmos_6p0 w=0.82u l=0.6u
X849 vss tune_series_gy[5] a_21748_9538# vss nmos_6p0 w=0.51u l=0.6u
X850 a_33500_18056# a_33412_18100# vss vss nmos_6p0 w=0.82u l=1u
X851 vdd a_2588_35304# a_2500_35348# vdd pmos_6p0 w=1.22u l=1u
X852 a_35692_14964# cap_series_gygyn a_35880_14964# vdd pmos_6p0 w=1.2u l=0.5u
X853 a_25780_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X854 a_20532_46324# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X855 a_34720_31428# cap_shunt_n a_32612_31490# vss nmos_6p0 w=0.82u l=0.6u
X856 a_9332_13020# cap_shunt_p a_9540_12674# vdd pmos_6p0 w=1.2u l=0.5u
X857 vdd tune_shunt[7] a_16500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X858 a_24204_53687# a_24116_53784# vss vss nmos_6p0 w=0.82u l=1u
X859 a_6292_48738# cap_shunt_p a_6084_49084# vdd pmos_6p0 w=1.2u l=0.5u
X860 a_19732_13880# cap_series_gyn a_19524_13396# vdd pmos_6p0 w=1.2u l=0.5u
X861 a_13588_47516# cap_shunt_p a_13796_47170# vdd pmos_6p0 w=1.2u l=0.5u
X862 vss cap_shunt_n a_22848_45240# vss nmos_6p0 w=0.82u l=0.6u
X863 a_13796_50306# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X864 a_31624_8316# cap_series_gygyn a_31648_7908# vss nmos_6p0 w=0.82u l=0.6u
X865 a_33500_14920# a_33412_14964# vss vss nmos_6p0 w=0.82u l=1u
X866 vdd tune_shunt[7] a_33524_27508# vdd pmos_6p0 w=1.2u l=0.5u
X867 a_35692_11828# cap_series_gygyp a_35880_11828# vdd pmos_6p0 w=1.2u l=0.5u
X868 a_6628_12674# cap_shunt_p a_6420_13020# vdd pmos_6p0 w=1.2u l=0.5u
X869 a_6532_43188# cap_shunt_p a_6740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X870 a_2500_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X871 a_20620_23895# a_20532_23992# vss vss nmos_6p0 w=0.82u l=1u
X872 a_24204_50551# a_24116_50648# vss vss nmos_6p0 w=0.82u l=1u
X873 vss cap_shunt_gyp a_34748_48376# vss nmos_6p0 w=0.82u l=0.6u
X874 vss cap_shunt_p a_22848_42104# vss nmos_6p0 w=0.82u l=0.6u
X875 a_4424_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X876 a_15700_9538# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X877 vdd a_20172_38007# a_20084_38104# vdd pmos_6p0 w=1.22u l=1u
X878 a_35840_23588# cap_series_gygyp a_34516_23650# vss nmos_6p0 w=0.82u l=0.6u
X879 a_6740_48376# cap_shunt_p a_7672_48376# vss nmos_6p0 w=0.82u l=0.6u
X880 a_14372_41620# cap_shunt_n a_14580_42104# vdd pmos_6p0 w=1.2u l=0.5u
X881 a_13796_25218# cap_shunt_n a_13588_25564# vdd pmos_6p0 w=1.2u l=0.5u
X882 a_11480_23288# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X883 a_28692_7608# cap_series_gyp a_28484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X884 vdd a_33948_54120# a_33860_54164# vdd pmos_6p0 w=1.22u l=1u
X885 a_2500_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X886 a_18612_7970# cap_series_gyp a_18404_8316# vdd pmos_6p0 w=1.2u l=0.5u
X887 vdd tune_series_gy[4] a_21540_5180# vdd pmos_6p0 w=1.2u l=0.5u
X888 a_1692_48983# a_1604_49080# vss vss nmos_6p0 w=0.82u l=1u
X889 a_30408_18584# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X890 a_20172_19191# a_20084_19288# vss vss nmos_6p0 w=0.82u l=1u
X891 a_23756_29032# a_23668_29076# vss vss nmos_6p0 w=0.82u l=1u
X892 vss tune_shunt[7] a_7748_26786# vss nmos_6p0 w=0.51u l=0.6u
X893 vdd a_14572_54120# a_14484_54164# vdd pmos_6p0 w=1.22u l=1u
X894 a_13796_22082# cap_shunt_n a_13588_22428# vdd pmos_6p0 w=1.2u l=0.5u
X895 a_13252_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X896 vss tune_shunt[5] a_3380_51512# vss nmos_6p0 w=0.51u l=0.6u
X897 vdd a_33948_50984# a_33860_51028# vdd pmos_6p0 w=1.22u l=1u
X898 a_37280_43189# tune_shunt_gy[3] vdd vdd pmos_6p0 w=1.215u l=0.5u
X899 a_35628_14487# a_35540_14584# vss vss nmos_6p0 w=0.82u l=1u
X900 a_3172_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X901 a_9108_47516# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X902 vdd a_2140_33303# a_2052_33400# vdd pmos_6p0 w=1.22u l=1u
X903 vss tune_shunt[7] a_13796_14242# vss nmos_6p0 w=0.51u l=0.6u
X904 a_3620_33780# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X905 a_35692_3988# cap_series_gygyp a_35880_3988# vdd pmos_6p0 w=1.2u l=0.5u
X906 a_6532_52596# cap_shunt_n a_6740_53080# vdd pmos_6p0 w=1.2u l=0.5u
X907 a_30408_15448# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X908 a_20172_16055# a_20084_16152# vss vss nmos_6p0 w=0.82u l=1u
X909 a_31372_52552# a_31284_52596# vss vss nmos_6p0 w=0.82u l=1u
X910 a_23756_25896# a_23668_25940# vss vss nmos_6p0 w=0.82u l=1u
X911 a_11984_21720# cap_shunt_p a_9876_21720# vss nmos_6p0 w=0.82u l=0.6u
X912 vdd a_16140_55688# a_16052_55732# vdd pmos_6p0 w=1.22u l=1u
X913 a_21628_54120# a_21540_54164# vss vss nmos_6p0 w=0.82u l=1u
X914 vdd tune_shunt[7] a_20532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X915 a_13252_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X916 a_34952_6340# cap_series_gygyp a_34536_6748# vss nmos_6p0 w=0.82u l=0.6u
X917 a_35628_11351# a_35540_11448# vss vss nmos_6p0 w=0.82u l=1u
X918 a_25548_47415# a_25460_47512# vss vss nmos_6p0 w=0.82u l=1u
X919 a_15492_5180# cap_series_gyn a_15700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X920 a_3620_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X921 a_18388_3266# cap_series_gyn a_18180_3612# vdd pmos_6p0 w=1.2u l=0.5u
X922 a_36076_34871# a_35988_34968# vss vss nmos_6p0 w=0.82u l=1u
X923 a_21316_3612# cap_series_gyp a_21524_3266# vdd pmos_6p0 w=1.2u l=0.5u
X924 a_19524_11828# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X925 a_10340_38484# cap_shunt_n a_10548_38968# vdd pmos_6p0 w=1.2u l=0.5u
X926 a_21540_28700# cap_shunt_n a_21748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X927 vss tune_shunt[7] a_21748_31490# vss nmos_6p0 w=0.51u l=0.6u
X928 vdd tune_shunt[7] a_20532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X929 a_34720_28292# cap_shunt_p a_32612_28354# vss nmos_6p0 w=0.82u l=0.6u
X930 a_19544_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X931 vss cap_shunt_p a_18032_20452# vss nmos_6p0 w=0.82u l=0.6u
X932 a_32444_11452# cap_series_gyp a_32632_11452# vdd pmos_6p0 w=1.2u l=0.5u
X933 a_37080_13880# cap_series_gygyn a_35880_13396# vss nmos_6p0 w=0.82u l=0.6u
X934 a_36076_31735# a_35988_31832# vss vss nmos_6p0 w=0.82u l=1u
X935 vdd a_33500_3944# a_33412_3988# vdd pmos_6p0 w=1.22u l=1u
X936 a_26376_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X937 a_10340_35348# cap_shunt_n a_10548_35832# vdd pmos_6p0 w=1.2u l=0.5u
X938 vdd tune_series_gy[4] a_29492_17724# vdd pmos_6p0 w=1.2u l=0.5u
X939 a_13796_47170# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X940 a_13796_34626# cap_shunt_n a_14728_34564# vss nmos_6p0 w=0.82u l=0.6u
X941 vdd a_2588_29032# a_2500_29076# vdd pmos_6p0 w=1.22u l=1u
X942 a_19524_7124# cap_series_gyp a_19732_7608# vdd pmos_6p0 w=1.2u l=0.5u
X943 a_28484_10260# cap_series_gyp a_28692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X944 a_4816_17316# cap_shunt_p a_2708_17378# vss nmos_6p0 w=0.82u l=0.6u
X945 a_34720_25156# cap_shunt_p a_32612_25218# vss nmos_6p0 w=0.82u l=0.6u
X946 vdd a_27900_45847# a_27812_45944# vdd pmos_6p0 w=1.22u l=1u
X947 a_8968_7908# cap_series_gyn a_7768_8316# vss nmos_6p0 w=0.82u l=0.6u
X948 a_37080_10744# cap_series_gygyp a_35880_10260# vss nmos_6p0 w=0.82u l=0.6u
X949 a_11096_7908# cap_series_gyp a_10680_8316# vss nmos_6p0 w=0.82u l=0.6u
X950 a_3932_52552# a_3844_52596# vss vss nmos_6p0 w=0.82u l=1u
X951 a_13796_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X952 a_13796_31490# cap_shunt_n a_14728_31428# vss nmos_6p0 w=0.82u l=0.6u
X953 a_1716_3988# cap_shunt_p a_1924_4472# vdd pmos_6p0 w=1.2u l=0.5u
X954 a_23532_55688# a_23444_55732# vss vss nmos_6p0 w=0.82u l=1u
X955 a_9876_51512# cap_shunt_n a_11592_51512# vss nmos_6p0 w=0.82u l=0.6u
X956 a_18032_32996# cap_shunt_n a_16708_33058# vss nmos_6p0 w=0.82u l=0.6u
X957 a_24452_23996# cap_shunt_p a_24660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X958 vss tune_shunt[7] a_6740_13880# vss nmos_6p0 w=0.51u l=0.6u
X959 vdd tune_shunt[7] a_7540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X960 vss tune_shunt[2] a_1924_6040# vss nmos_6p0 w=0.51u l=0.6u
X961 a_9540_14242# cap_shunt_p a_9332_14588# vdd pmos_6p0 w=1.2u l=0.5u
X962 a_13588_38108# cap_shunt_n a_13796_37762# vdd pmos_6p0 w=1.2u l=0.5u
X963 a_21540_30268# cap_shunt_n a_21748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X964 a_3640_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X965 a_13796_18946# cap_shunt_p a_13588_19292# vdd pmos_6p0 w=1.2u l=0.5u
X966 a_35880_13396# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X967 a_17148_52119# a_17060_52216# vss vss nmos_6p0 w=0.82u l=1u
X968 a_35880_36916# cap_series_gygyp a_35692_36916# vdd pmos_6p0 w=1.2u l=0.5u
X969 a_20508_55688# a_20420_55732# vss vss nmos_6p0 w=0.82u l=1u
X970 a_2500_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X971 a_13588_42812# cap_shunt_n a_13796_42466# vdd pmos_6p0 w=1.2u l=0.5u
X972 a_31036_43144# a_30948_43188# vss vss nmos_6p0 w=0.82u l=1u
X973 vdd tune_shunt[6] a_10452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X974 vdd a_32156_40008# a_32068_40052# vdd pmos_6p0 w=1.22u l=1u
X975 vss tune_shunt[7] a_24660_29922# vss nmos_6p0 w=0.51u l=0.6u
X976 a_37420_49416# a_37332_49460# vss vss nmos_6p0 w=0.82u l=1u
X977 a_29468_44279# a_29380_44376# vss vss nmos_6p0 w=0.82u l=1u
X978 a_6532_14964# cap_shunt_p a_6740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X979 a_13796_15810# cap_shunt_p a_13588_16156# vdd pmos_6p0 w=1.2u l=0.5u
X980 vdd a_27340_49416# a_27252_49460# vdd pmos_6p0 w=1.22u l=1u
X981 vdd a_32268_5079# a_32180_5176# vdd pmos_6p0 w=1.22u l=1u
X982 vss cap_shunt_p a_27888_4472# vss nmos_6p0 w=0.82u l=0.6u
X983 a_35880_10260# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X984 a_2708_47170# cap_shunt_p a_4424_47108# vss nmos_6p0 w=0.82u l=0.6u
X985 vdd tune_shunt[4] a_28484_40052# vdd pmos_6p0 w=1.2u l=0.5u
X986 a_25780_10744# cap_series_gyn a_25572_10260# vdd pmos_6p0 w=1.2u l=0.5u
X987 a_35740_55255# a_35652_55352# vss vss nmos_6p0 w=0.82u l=1u
X988 a_1692_39575# a_1604_39672# vss vss nmos_6p0 w=0.82u l=1u
X989 a_35040_45302# cap_shunt_gyp a_35040_44757# vdd pmos_6p0 w=1.215u l=0.5u
X990 vss cap_shunt_n a_14784_34264# vss nmos_6p0 w=0.82u l=0.6u
X991 a_37420_46280# a_37332_46324# vss vss nmos_6p0 w=0.82u l=1u
X992 vdd tune_shunt[3] a_24452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X993 a_29468_41143# a_29380_41240# vss vss nmos_6p0 w=0.82u l=1u
X994 a_6532_11828# cap_shunt_p a_6740_12312# vdd pmos_6p0 w=1.2u l=0.5u
X995 vss cap_shunt_p a_4704_17016# vss nmos_6p0 w=0.82u l=0.6u
X996 vdd tune_shunt[7] a_16500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X997 vdd a_27340_46280# a_27252_46324# vdd pmos_6p0 w=1.22u l=1u
X998 a_19732_13880# cap_series_gyn a_19524_13396# vdd pmos_6p0 w=1.2u l=0.5u
X999 vdd a_24316_49416# a_24228_49460# vdd pmos_6p0 w=1.22u l=1u
X1000 a_13252_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1001 a_24660_37762# cap_shunt_p a_26376_37700# vss nmos_6p0 w=0.82u l=0.6u
X1002 a_3620_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1003 vdd a_19388_55255# a_19300_55352# vdd pmos_6p0 w=1.22u l=1u
X1004 a_2500_45948# cap_shunt_p a_2708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X1005 a_6740_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1006 a_6532_43188# cap_shunt_p a_6740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X1007 a_25572_41620# cap_shunt_n a_25780_42104# vdd pmos_6p0 w=1.2u l=0.5u
X1008 a_36076_28599# a_35988_28696# vss vss nmos_6p0 w=0.82u l=1u
X1009 vss cap_shunt_n a_14784_31128# vss nmos_6p0 w=0.82u l=0.6u
X1010 a_17024_6340# cap_series_gyp a_15700_6402# vss nmos_6p0 w=0.82u l=0.6u
X1011 a_11984_12312# cap_shunt_p a_9876_12312# vss nmos_6p0 w=0.82u l=0.6u
X1012 vdd tune_shunt[5] a_24452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X1013 a_23756_16488# a_23668_16532# vss vss nmos_6p0 w=0.82u l=1u
X1014 vss tune_shunt[6] a_9876_48376# vss nmos_6p0 w=0.51u l=0.6u
X1015 vdd tune_shunt[5] a_20532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X1016 a_13252_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1017 a_32156_32168# a_32068_32212# vss vss nmos_6p0 w=0.82u l=1u
X1018 a_10548_26424# cap_shunt_n a_10340_25940# vdd pmos_6p0 w=1.2u l=0.5u
X1019 vss cap_shunt_p a_18032_14180# vss nmos_6p0 w=0.82u l=0.6u
X1020 a_31260_53687# a_31172_53784# vss vss nmos_6p0 w=0.82u l=1u
X1021 a_3620_21236# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1022 a_21516_55255# a_21428_55352# vss vss nmos_6p0 w=0.82u l=1u
X1023 vdd a_19388_52119# a_19300_52216# vdd pmos_6p0 w=1.22u l=1u
X1024 vss cap_shunt_gyp a_37548_43672# vss nmos_6p0 w=0.82u l=0.6u
X1025 a_14372_41620# cap_shunt_n a_14580_42104# vdd pmos_6p0 w=1.2u l=0.5u
X1026 a_6740_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1027 a_36076_25463# a_35988_25560# vss vss nmos_6p0 w=0.82u l=1u
X1028 a_26376_14180# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1029 a_14484_7124# cap_series_gyp a_14692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X1030 vdd a_36636_38440# a_36548_38484# vdd pmos_6p0 w=1.22u l=1u
X1031 a_10340_29076# cap_shunt_n a_10548_29560# vdd pmos_6p0 w=1.2u l=0.5u
X1032 a_13796_28354# cap_shunt_n a_14728_28292# vss nmos_6p0 w=0.82u l=0.6u
X1033 a_17416_4772# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1034 a_12580_19668# cap_shunt_p a_12788_20152# vdd pmos_6p0 w=1.2u l=0.5u
X1035 vss tune_series_gygy[5] a_34516_23650# vss nmos_6p0 w=0.51u l=0.6u
X1036 vss tune_shunt[7] a_21748_22082# vss nmos_6p0 w=0.51u l=0.6u
X1037 vss cap_shunt_p a_5936_20152# vss nmos_6p0 w=0.82u l=0.6u
X1038 vdd tune_shunt[7] a_20532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X1039 a_6292_51874# cap_shunt_p a_7224_51812# vss nmos_6p0 w=0.82u l=0.6u
X1040 a_10548_23288# cap_shunt_n a_10340_22804# vdd pmos_6p0 w=1.2u l=0.5u
X1041 a_31260_50551# a_31172_50648# vss vss nmos_6p0 w=0.82u l=1u
X1042 a_9464_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1043 a_26376_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X1044 a_19724_22327# a_19636_22424# vss vss nmos_6p0 w=0.82u l=1u
X1045 a_13252_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1046 a_13796_25218# cap_shunt_n a_14728_25156# vss nmos_6p0 w=0.82u l=0.6u
X1047 a_3172_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1048 vss tune_series_gygy[5] a_34516_20514# vss nmos_6p0 w=0.51u l=0.6u
X1049 a_7672_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1050 a_28348_45847# a_28260_45944# vss vss nmos_6p0 w=0.82u l=1u
X1051 a_9464_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1052 a_30364_22327# a_30276_22424# vss vss nmos_6p0 w=0.82u l=1u
X1053 a_9428_18946# cap_shunt_p a_9220_19292# vdd pmos_6p0 w=1.2u l=0.5u
X1054 vss tune_shunt[7] a_17828_21720# vss nmos_6p0 w=0.51u l=0.6u
X1055 a_13252_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1056 vdd a_5388_3944# a_5300_3988# vdd pmos_6p0 w=1.22u l=1u
X1057 vss tune_shunt[0] a_28692_6040# vss nmos_6p0 w=0.51u l=0.6u
X1058 a_34348_9884# cap_series_gygyn a_34536_9884# vdd pmos_6p0 w=1.2u l=0.5u
X1059 a_18032_23588# cap_shunt_n a_16708_23650# vss nmos_6p0 w=0.82u l=0.6u
X1060 a_7960_6040# cap_series_gyp a_6760_5556# vss nmos_6p0 w=0.82u l=0.6u
X1061 vdd tune_shunt_gy[2] a_37444_41240# vdd pmos_6p0 w=1.215u l=0.5u
X1062 vss cap_shunt_n a_33936_36132# vss nmos_6p0 w=0.82u l=0.6u
X1063 vss cap_shunt_n a_12768_32996# vss nmos_6p0 w=0.82u l=0.6u
X1064 a_5844_3266# cap_shunt_n a_5636_3612# vdd pmos_6p0 w=1.2u l=0.5u
X1065 a_24452_14588# cap_series_gyn a_24660_14242# vdd pmos_6p0 w=1.2u l=0.5u
X1066 vdd a_2588_55255# a_2500_55352# vdd pmos_6p0 w=1.22u l=1u
X1067 a_33732_34264# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1068 a_13588_36540# cap_shunt_n a_13796_36194# vdd pmos_6p0 w=1.2u l=0.5u
X1069 vss tune_shunt[7] a_6740_27992# vss nmos_6p0 w=0.51u l=0.6u
X1070 vss cap_series_gyp a_21056_9176# vss nmos_6p0 w=0.82u l=0.6u
X1071 vdd tune_shunt[7] a_10452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X1072 a_12580_49460# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1073 a_34348_6748# cap_series_gygyp a_34536_6748# vdd pmos_6p0 w=1.2u l=0.5u
X1074 a_11780_6040# cap_series_gyn a_12712_6040# vss nmos_6p0 w=0.82u l=0.6u
X1075 a_22436_13396# cap_series_gyn a_22644_13880# vdd pmos_6p0 w=1.2u l=0.5u
X1076 vdd a_31372_55688# a_31284_55732# vdd pmos_6p0 w=1.22u l=1u
X1077 a_24764_52552# a_24676_52596# vss vss nmos_6p0 w=0.82u l=1u
X1078 vdd tune_shunt[7] a_32404_28700# vdd pmos_6p0 w=1.2u l=0.5u
X1079 a_32444_11452# cap_series_gyp a_32632_11452# vdd pmos_6p0 w=1.2u l=0.5u
X1080 vdd a_2588_52119# a_2500_52216# vdd pmos_6p0 w=1.22u l=1u
X1081 a_35692_10260# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1082 a_35308_43672# cap_shunt_gyp a_35040_43734# vss nmos_6p0 w=0.82u l=0.6u
X1083 a_33732_31128# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1084 a_35692_3988# cap_series_gygyp a_35880_3988# vdd pmos_6p0 w=1.2u l=0.5u
X1085 a_17596_49416# a_17508_49460# vss vss nmos_6p0 w=0.82u l=1u
X1086 a_13588_33404# cap_shunt_n a_13796_33058# vdd pmos_6p0 w=1.2u l=0.5u
X1087 vss tune_shunt[7] a_6740_24856# vss nmos_6p0 w=0.51u l=0.6u
X1088 a_24660_12674# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1089 vdd tune_shunt[7] a_10452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X1090 a_9668_16532# cap_shunt_p a_9876_17016# vdd pmos_6p0 w=1.2u l=0.5u
X1091 a_9668_16532# cap_shunt_p a_9876_17016# vdd pmos_6p0 w=1.2u l=0.5u
X1092 a_24660_9538# cap_series_gyn a_24452_9884# vdd pmos_6p0 w=1.2u l=0.5u
X1093 a_2500_39676# cap_shunt_n a_2708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X1094 vss cap_series_gyp a_26768_4772# vss nmos_6p0 w=0.82u l=0.6u
X1095 vdd a_17596_10216# a_17508_10260# vdd pmos_6p0 w=1.22u l=1u
X1096 vss tune_shunt[6] a_10660_40898# vss nmos_6p0 w=0.51u l=0.6u
X1097 a_24452_23996# cap_shunt_p a_24660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X1098 vss cap_series_gyp a_16800_7608# vss nmos_6p0 w=0.82u l=0.6u
X1099 a_33524_33780# cap_shunt_n a_33732_34264# vdd pmos_6p0 w=1.2u l=0.5u
X1100 a_20740_35832# cap_shunt_n a_22456_35832# vss nmos_6p0 w=0.82u l=0.6u
X1101 a_25236_3612# cap_shunt_p a_25444_3266# vdd pmos_6p0 w=1.2u l=0.5u
X1102 a_5836_7080# a_5748_7124# vss vss nmos_6p0 w=0.82u l=1u
X1103 vdd a_13564_8215# a_13476_8312# vdd pmos_6p0 w=1.22u l=1u
X1104 a_24660_6402# cap_series_gyn a_24452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X1105 vss cap_series_gyp a_7960_6040# vss nmos_6p0 w=0.82u l=0.6u
X1106 a_23072_12612# cap_series_gyn a_21748_12674# vss nmos_6p0 w=0.82u l=0.6u
X1107 a_6740_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1108 a_25572_32212# cap_shunt_p a_25780_32696# vdd pmos_6p0 w=1.2u l=0.5u
X1109 a_21516_48983# a_21428_49080# vss vss nmos_6p0 w=0.82u l=1u
X1110 vdd a_21292_47848# a_21204_47892# vdd pmos_6p0 w=1.22u l=1u
X1111 a_33524_30644# cap_shunt_n a_33732_31128# vdd pmos_6p0 w=1.2u l=0.5u
X1112 a_25592_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1113 a_15132_50984# a_15044_51028# vss vss nmos_6p0 w=0.82u l=1u
X1114 a_2708_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1115 vdd tune_series_gy[3] a_28484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X1116 a_15120_20452# cap_shunt_n a_13796_20514# vss nmos_6p0 w=0.82u l=0.6u
X1117 vdd a_3932_55688# a_3844_55732# vdd pmos_6p0 w=1.22u l=1u
X1118 a_13588_42812# cap_shunt_n a_13796_42466# vdd pmos_6p0 w=1.2u l=0.5u
X1119 a_14468_3266# cap_series_gyn a_14260_3612# vdd pmos_6p0 w=1.2u l=0.5u
X1120 a_32156_22760# a_32068_22804# vss vss nmos_6p0 w=0.82u l=1u
X1121 a_30616_21236# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1122 a_6740_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1123 a_25592_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1124 a_17828_18584# cap_shunt_p a_17620_18100# vdd pmos_6p0 w=1.2u l=0.5u
X1125 a_9876_53080# cap_shunt_n a_9668_52596# vdd pmos_6p0 w=1.2u l=0.5u
X1126 vdd tune_shunt[6] a_3620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X1127 a_25780_10744# cap_series_gyn a_25572_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1128 a_5544_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1129 vdd tune_shunt[4] a_28484_40052# vdd pmos_6p0 w=1.2u l=0.5u
X1130 a_2708_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1131 a_7768_6748# cap_series_gyp a_7580_6748# vdd pmos_6p0 w=1.2u l=0.5u
X1132 a_6852_53442# cap_shunt_n a_6644_53788# vdd pmos_6p0 w=1.2u l=0.5u
X1133 a_14504_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1134 a_17620_46324# cap_shunt_n a_17828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X1135 a_9464_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1136 a_12444_17623# a_12356_17720# vss vss nmos_6p0 w=0.82u l=1u
X1137 a_15804_19624# a_15716_19668# vss vss nmos_6p0 w=0.82u l=1u
X1138 a_13796_20514# cap_shunt_n a_13588_20860# vdd pmos_6p0 w=1.2u l=0.5u
X1139 vdd a_10092_44712# a_10004_44756# vdd pmos_6p0 w=1.22u l=1u
X1140 a_29196_3612# cap_series_gyn a_29384_3612# vdd pmos_6p0 w=1.2u l=0.5u
X1141 vdd a_31820_54120# a_31732_54164# vdd pmos_6p0 w=1.22u l=1u
X1142 a_20532_36916# cap_shunt_n a_20740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X1143 a_13252_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1144 a_34188_45240# cap_shunt_gyn a_33920_45302# vss nmos_6p0 w=0.82u l=0.6u
X1145 a_25780_7608# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X1146 a_22644_9176# cap_series_gyp a_23576_9176# vss nmos_6p0 w=0.82u l=0.6u
X1147 a_7672_12312# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1148 a_5544_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1149 vdd tune_series_gy[5] a_18404_13020# vdd pmos_6p0 w=1.2u l=0.5u
X1150 a_29720_16156# cap_series_gyn a_29532_16156# vdd pmos_6p0 w=1.2u l=0.5u
X1151 a_5612_12919# a_5524_13016# vss vss nmos_6p0 w=0.82u l=1u
X1152 a_31436_8316# cap_series_gygyn a_31624_8316# vdd pmos_6p0 w=1.2u l=0.5u
X1153 a_24660_40898# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1154 a_33948_3511# a_33860_3608# vss vss nmos_6p0 w=0.82u l=1u
X1155 vdd a_32268_16055# a_32180_16152# vdd pmos_6p0 w=1.22u l=1u
X1156 a_35692_18100# cap_series_gygyn a_35880_18100# vdd pmos_6p0 w=1.2u l=0.5u
X1157 vdd a_31820_50984# a_31732_51028# vdd pmos_6p0 w=1.22u l=1u
X1158 a_13252_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1159 vdd a_31372_49416# a_31284_49460# vdd pmos_6p0 w=1.22u l=1u
X1160 a_4648_12312# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1161 vss cap_shunt_n a_12768_23588# vss nmos_6p0 w=0.82u l=0.6u
X1162 vdd a_31708_14920# a_31620_14964# vdd pmos_6p0 w=1.22u l=1u
X1163 a_24660_39330# cap_shunt_p a_24452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X1164 a_28692_32696# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1165 a_2708_23650# cap_shunt_p a_2500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X1166 a_9332_13020# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1167 a_25572_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1168 a_15512_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1169 a_13588_27132# cap_shunt_n a_13796_26786# vdd pmos_6p0 w=1.2u l=0.5u
X1170 a_27676_6647# a_27588_6744# vss vss nmos_6p0 w=0.82u l=1u
X1171 vdd a_32268_12919# a_32180_13016# vdd pmos_6p0 w=1.22u l=1u
X1172 a_36748_32168# a_36660_32212# vss vss nmos_6p0 w=0.82u l=1u
X1173 vdd tune_shunt[7] a_10452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X1174 a_15356_11784# a_15268_11828# vss vss nmos_6p0 w=0.82u l=1u
X1175 vdd a_31372_46280# a_31284_46324# vdd pmos_6p0 w=1.22u l=1u
X1176 vss tune_shunt[2] a_1924_7608# vss nmos_6p0 w=0.51u l=0.6u
X1177 a_10340_33780# cap_shunt_n a_10548_34264# vdd pmos_6p0 w=1.2u l=0.5u
X1178 vdd tune_series_gy[5] a_19524_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1179 vdd a_31708_11784# a_31620_11828# vdd pmos_6p0 w=1.22u l=1u
X1180 a_15512_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1181 vdd tune_shunt[5] a_17620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X1182 a_10660_6402# cap_series_gyn a_11592_6340# vss nmos_6p0 w=0.82u l=0.6u
X1183 vss tune_shunt[7] a_6740_15448# vss nmos_6p0 w=0.51u l=0.6u
X1184 a_36688_20152# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X1185 a_24652_53687# a_24564_53784# vss vss nmos_6p0 w=0.82u l=1u
X1186 vdd a_30812_47415# a_30724_47512# vdd pmos_6p0 w=1.22u l=1u
X1187 vdd tune_series_gy[4] a_21428_5556# vdd pmos_6p0 w=1.2u l=0.5u
X1188 a_14908_55255# a_14820_55352# vss vss nmos_6p0 w=0.82u l=1u
X1189 a_20740_29560# cap_shunt_n a_22456_29560# vss nmos_6p0 w=0.82u l=0.6u
X1190 a_37652_42104# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X1191 a_10340_30644# cap_shunt_n a_10548_31128# vdd pmos_6p0 w=1.2u l=0.5u
X1192 vss tune_shunt[7] a_32612_26786# vss nmos_6p0 w=0.51u l=0.6u
X1193 a_28692_7608# cap_series_gyp a_28484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X1194 a_19524_8692# cap_series_gyp a_19732_9176# vdd pmos_6p0 w=1.2u l=0.5u
X1195 a_13588_30268# cap_shunt_n a_13796_29922# vdd pmos_6p0 w=1.2u l=0.5u
X1196 a_11668_45240# cap_shunt_n a_11460_44756# vdd pmos_6p0 w=1.2u l=0.5u
X1197 a_32716_39575# a_32628_39672# vss vss nmos_6p0 w=0.82u l=1u
X1198 a_18612_7970# cap_series_gyp a_18404_8316# vdd pmos_6p0 w=1.2u l=0.5u
X1199 a_37420_52119# a_37332_52216# vss vss nmos_6p0 w=0.82u l=1u
X1200 a_24652_50551# a_24564_50648# vss vss nmos_6p0 w=0.82u l=1u
X1201 a_24452_14588# cap_series_gyn a_24660_14242# vdd pmos_6p0 w=1.2u l=0.5u
X1202 a_10660_45602# cap_shunt_n a_10452_45948# vdd pmos_6p0 w=1.2u l=0.5u
X1203 a_20740_26424# cap_shunt_n a_22456_26424# vss nmos_6p0 w=0.82u l=0.6u
X1204 a_15120_14180# cap_shunt_p a_13796_14242# vss nmos_6p0 w=0.82u l=0.6u
X1205 vss tune_shunt[6] a_14580_45240# vss nmos_6p0 w=0.51u l=0.6u
X1206 vss tune_shunt[4] a_25780_42104# vss nmos_6p0 w=0.51u l=0.6u
X1207 a_13588_36540# cap_shunt_n a_13796_36194# vdd pmos_6p0 w=1.2u l=0.5u
X1208 a_23308_44712# a_23220_44756# vss vss nmos_6p0 w=0.82u l=1u
X1209 vdd a_10540_43144# a_10452_43188# vdd pmos_6p0 w=1.22u l=1u
X1210 vss tune_shunt[7] a_16708_23650# vss nmos_6p0 w=0.51u l=0.6u
X1211 a_7540_45948# cap_shunt_p a_7748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X1212 a_21672_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1213 a_22436_13396# cap_series_gyn a_22644_13880# vdd pmos_6p0 w=1.2u l=0.5u
X1214 a_6292_49944# cap_shunt_p a_6084_49460# vdd pmos_6p0 w=1.2u l=0.5u
X1215 vdd a_2140_41576# a_2052_41620# vdd pmos_6p0 w=1.22u l=1u
X1216 a_29700_28354# cap_shunt_p a_29492_28700# vdd pmos_6p0 w=1.2u l=0.5u
X1217 a_32444_11452# cap_series_gyp a_32632_11452# vdd pmos_6p0 w=1.2u l=0.5u
X1218 vdd a_15356_53687# a_15268_53784# vdd pmos_6p0 w=1.22u l=1u
X1219 a_27104_37400# cap_shunt_p a_25780_37400# vss nmos_6p0 w=0.82u l=0.6u
X1220 vss cap_series_gygyn a_36624_17316# vss nmos_6p0 w=0.82u l=0.6u
X1221 a_17828_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1222 a_2708_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1223 vss tune_shunt[6] a_14580_42104# vss nmos_6p0 w=0.51u l=0.6u
X1224 a_13588_33404# cap_shunt_n a_13796_33058# vdd pmos_6p0 w=1.2u l=0.5u
X1225 a_23308_41576# a_23220_41620# vss vss nmos_6p0 w=0.82u l=1u
X1226 vss tune_shunt[7] a_16708_20514# vss nmos_6p0 w=0.51u l=0.6u
X1227 a_19152_45240# cap_shunt_p a_17828_45240# vss nmos_6p0 w=0.82u l=0.6u
X1228 a_21672_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1229 a_30812_8215# a_30724_8312# vss vss nmos_6p0 w=0.82u l=1u
X1230 a_25592_17316# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X1231 a_17620_19668# cap_shunt_p a_17828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X1232 a_2708_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1233 vdd tune_shunt[3] a_2724_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1234 a_5544_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1235 a_17620_41620# cap_shunt_n a_17828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X1236 a_24452_23996# cap_shunt_p a_24660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X1237 vss tune_series_gy[2] a_7768_8316# vss nmos_6p0 w=0.51u l=0.6u
X1238 a_9668_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1239 a_25996_47415# a_25908_47512# vss vss nmos_6p0 w=0.82u l=1u
X1240 a_19152_42104# cap_shunt_n a_17828_42104# vss nmos_6p0 w=0.82u l=0.6u
X1241 a_6060_30167# a_5972_30264# vss vss nmos_6p0 w=0.82u l=1u
X1242 vss tune_shunt_gy[5] a_37632_47512# vss nmos_6p0 w=0.51u l=0.6u
X1243 a_20532_27508# cap_shunt_n a_20740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X1244 a_28692_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1245 a_5636_9884# cap_shunt_p a_5844_9538# vdd pmos_6p0 w=1.2u l=0.5u
X1246 a_31024_36132# cap_shunt_n a_29700_36194# vss nmos_6p0 w=0.82u l=0.6u
X1247 a_35880_7124# cap_series_gygyp a_36688_7608# vss nmos_6p0 w=0.82u l=0.6u
X1248 vss tune_series_gy[4] a_18612_4472# vss nmos_6p0 w=0.51u l=0.6u
X1249 a_6292_17016# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1250 a_5544_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1251 a_35880_36916# cap_series_gygyp a_36688_37400# vss nmos_6p0 w=0.82u l=0.6u
X1252 vss tune_series_gy[1] a_7768_5180# vss nmos_6p0 w=0.51u l=0.6u
X1253 vdd a_36636_55255# a_36548_55352# vdd pmos_6p0 w=1.22u l=1u
X1254 a_35880_13396# cap_series_gygyn a_35692_13396# vdd pmos_6p0 w=1.2u l=0.5u
X1255 a_6060_27031# a_5972_27128# vss vss nmos_6p0 w=0.82u l=1u
X1256 a_6784_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X1257 a_7560_12612# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1258 a_35040_43189# cap_shunt_gyp a_35040_43734# vdd pmos_6p0 w=1.215u l=0.5u
X1259 vss tune_shunt[6] a_3828_38968# vss nmos_6p0 w=0.51u l=0.6u
X1260 a_9644_36872# a_9556_36916# vss vss nmos_6p0 w=0.82u l=1u
X1261 a_29700_29922# cap_shunt_p a_29492_30268# vdd pmos_6p0 w=1.2u l=0.5u
X1262 a_8860_8648# a_8772_8692# vss vss nmos_6p0 w=0.82u l=1u
X1263 vdd tune_shunt[7] a_9332_16156# vdd pmos_6p0 w=1.2u l=0.5u
X1264 vss cap_shunt_p a_19152_21720# vss nmos_6p0 w=0.82u l=0.6u
X1265 vdd tune_shunt[7] a_9668_19668# vdd pmos_6p0 w=1.2u l=0.5u
X1266 a_29492_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1267 vss tune_series_gy[5] a_21748_7970# vss nmos_6p0 w=0.51u l=0.6u
X1268 vdd a_36636_52119# a_36548_52216# vdd pmos_6p0 w=1.22u l=1u
X1269 a_2708_14242# cap_shunt_n a_2500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X1270 a_25780_40536# cap_shunt_n a_25572_40052# vdd pmos_6p0 w=1.2u l=0.5u
X1271 a_28692_23288# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1272 vdd a_29132_52552# a_29044_52596# vdd pmos_6p0 w=1.22u l=1u
X1273 vdd tune_shunt[6] a_25572_38484# vdd pmos_6p0 w=1.2u l=0.5u
X1274 vdd tune_shunt[6] a_6532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X1275 vss cap_shunt_n a_8064_27992# vss nmos_6p0 w=0.82u l=0.6u
X1276 vss tune_series_gy[4] a_15700_9538# vss nmos_6p0 w=0.51u l=0.6u
X1277 a_34308_17724# cap_series_gygyn a_34516_17378# vdd pmos_6p0 w=1.2u l=0.5u
X1278 a_18816_47108# cap_shunt_n a_16708_47170# vss nmos_6p0 w=0.82u l=0.6u
X1279 a_13796_50306# cap_shunt_p a_13588_50652# vdd pmos_6p0 w=1.2u l=0.5u
X1280 a_21748_44034# cap_shunt_n a_21540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X1281 vss tune_series_gy[4] a_21748_4834# vss nmos_6p0 w=0.51u l=0.6u
X1282 a_13796_20514# cap_shunt_n a_13588_20860# vdd pmos_6p0 w=1.2u l=0.5u
X1283 vss cap_shunt_n a_18816_29860# vss nmos_6p0 w=0.82u l=0.6u
X1284 a_20532_36916# cap_shunt_n a_20740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X1285 a_10340_24372# cap_shunt_n a_10548_24856# vdd pmos_6p0 w=1.2u l=0.5u
X1286 a_23980_55688# a_23892_55732# vss vss nmos_6p0 w=0.82u l=1u
X1287 a_14580_40536# cap_shunt_n a_14372_40052# vdd pmos_6p0 w=1.2u l=0.5u
X1288 a_30800_27992# cap_shunt_p a_28692_27992# vss nmos_6p0 w=0.82u l=0.6u
X1289 vss cap_shunt_p a_8064_24856# vss nmos_6p0 w=0.82u l=0.6u
X1290 vdd tune_shunt[6] a_25572_35348# vdd pmos_6p0 w=1.2u l=0.5u
X1291 a_21748_40898# cap_shunt_p a_21540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X1292 a_10660_39330# cap_shunt_n a_10452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X1293 a_27496_32696# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1294 vss cap_shunt_n a_18816_26724# vss nmos_6p0 w=0.82u l=0.6u
X1295 a_6532_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1296 vdd tune_shunt[6] a_13588_45948# vdd pmos_6p0 w=1.2u l=0.5u
X1297 a_3828_38968# cap_shunt_n a_4760_38968# vss nmos_6p0 w=0.82u l=0.6u
X1298 a_17596_52119# a_17508_52216# vss vss nmos_6p0 w=0.82u l=1u
X1299 a_7540_39676# cap_shunt_n a_7748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X1300 a_21748_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1301 a_30800_24856# cap_shunt_p a_28692_24856# vss nmos_6p0 w=0.82u l=0.6u
X1302 a_20740_15448# cap_series_gyn a_20532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X1303 vdd tune_shunt[5] a_9668_51028# vdd pmos_6p0 w=1.2u l=0.5u
X1304 a_34396_8648# a_34308_8692# vss vss nmos_6p0 w=0.82u l=1u
X1305 a_30812_19191# a_30724_19288# vss vss nmos_6p0 w=0.82u l=1u
X1306 a_31484_43144# a_31396_43188# vss vss nmos_6p0 w=0.82u l=1u
X1307 a_24660_39330# cap_shunt_p a_24452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X1308 a_20740_17016# cap_shunt_p a_22456_17016# vss nmos_6p0 w=0.82u l=0.6u
X1309 a_13588_27132# cap_shunt_n a_13796_26786# vdd pmos_6p0 w=1.2u l=0.5u
X1310 a_1924_3266# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X1311 a_21524_4472# cap_series_gyn a_21316_3988# vdd pmos_6p0 w=1.2u l=0.5u
X1312 a_6532_11828# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1313 vdd tune_series_gy[5] a_19524_13396# vdd pmos_6p0 w=1.2u l=0.5u
X1314 vss tune_shunt[7] a_16708_14242# vss nmos_6p0 w=0.51u l=0.6u
X1315 a_21672_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1316 vss tune_shunt[7] a_16708_37762# vss nmos_6p0 w=0.51u l=0.6u
X1317 a_13588_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1318 a_10340_33780# cap_shunt_n a_10548_34264# vdd pmos_6p0 w=1.2u l=0.5u
X1319 vdd a_2140_32168# a_2052_32212# vdd pmos_6p0 w=1.22u l=1u
X1320 a_6292_18946# cap_shunt_p a_8008_18884# vss nmos_6p0 w=0.82u l=0.6u
X1321 a_25780_20152# cap_series_gyp a_26712_20152# vss nmos_6p0 w=0.82u l=0.6u
X1322 a_23464_39268# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1323 vss cap_series_gyn a_16016_9176# vss nmos_6p0 w=0.82u l=0.6u
X1324 a_34844_49416# a_34756_49460# vss vss nmos_6p0 w=0.82u l=1u
X1325 vdd a_24764_49416# a_24676_49460# vdd pmos_6p0 w=1.22u l=1u
X1326 a_24452_5180# cap_series_gyp a_24660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X1327 a_21672_15448# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1328 vss tune_shunt[7] a_16708_34626# vss nmos_6p0 w=0.51u l=0.6u
X1329 a_10340_30644# cap_shunt_n a_10548_31128# vdd pmos_6p0 w=1.2u l=0.5u
X1330 a_28692_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1331 a_6740_13880# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1332 a_6292_15810# cap_shunt_p a_8008_15748# vss nmos_6p0 w=0.82u l=0.6u
X1333 vdd a_28124_42711# a_28036_42808# vdd pmos_6p0 w=1.22u l=1u
X1334 vdd a_27228_17623# a_27140_17720# vdd pmos_6p0 w=1.22u l=1u
X1335 a_10660_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1336 a_2140_27464# a_2052_27508# vss vss nmos_6p0 w=0.82u l=1u
X1337 a_21748_18946# cap_shunt_p a_23464_18884# vss nmos_6p0 w=0.82u l=0.6u
X1338 a_4760_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1339 a_11668_45240# cap_shunt_n a_11460_44756# vdd pmos_6p0 w=1.2u l=0.5u
X1340 a_17620_32212# cap_shunt_n a_17828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X1341 a_29700_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1342 vdd a_34844_10216# a_34756_10260# vdd pmos_6p0 w=1.22u l=1u
X1343 a_24452_14588# cap_series_gyn a_24660_14242# vdd pmos_6p0 w=1.2u l=0.5u
X1344 a_10660_45602# cap_shunt_n a_10452_45948# vdd pmos_6p0 w=1.2u l=0.5u
X1345 a_9876_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1346 a_21964_55255# a_21876_55352# vss vss nmos_6p0 w=0.82u l=1u
X1347 a_28692_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1348 vdd tune_series_gygy[5] a_34308_23996# vdd pmos_6p0 w=1.2u l=0.5u
X1349 a_9668_49460# cap_shunt_p a_9876_49944# vdd pmos_6p0 w=1.2u l=0.5u
X1350 a_7540_45948# cap_shunt_p a_7748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X1351 a_2140_24328# a_2052_24372# vss vss nmos_6p0 w=0.82u l=1u
X1352 a_22644_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1353 a_21748_15810# cap_series_gyn a_23464_15748# vss nmos_6p0 w=0.82u l=0.6u
X1354 a_29700_28354# cap_shunt_p a_29492_28700# vdd pmos_6p0 w=1.2u l=0.5u
X1355 a_22436_13396# cap_series_gyn a_22644_13880# vdd pmos_6p0 w=1.2u l=0.5u
X1356 a_17640_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1357 a_35736_7908# cap_series_gygyp a_34536_8316# vss nmos_6p0 w=0.82u l=0.6u
X1358 a_12768_37700# cap_shunt_n a_10660_37762# vss nmos_6p0 w=0.82u l=0.6u
X1359 a_14896_48376# cap_shunt_p a_12788_48376# vss nmos_6p0 w=0.82u l=0.6u
X1360 vdd a_16700_47848# a_16612_47892# vdd pmos_6p0 w=1.22u l=1u
X1361 a_10452_23996# cap_shunt_n a_10660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X1362 a_13796_44034# cap_shunt_n a_13588_44380# vdd pmos_6p0 w=1.2u l=0.5u
X1363 a_22644_10744# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1364 a_10548_3266# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X1365 vdd a_12444_10216# a_12356_10260# vdd pmos_6p0 w=1.22u l=1u
X1366 a_8064_43672# cap_shunt_p a_6740_43672# vss nmos_6p0 w=0.82u l=0.6u
X1367 a_15176_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1368 a_7748_23650# cap_shunt_p a_7540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X1369 vdd tune_shunt[7] a_12580_18100# vdd pmos_6p0 w=1.2u l=0.5u
X1370 a_28796_45847# a_28708_45944# vss vss nmos_6p0 w=0.82u l=1u
X1371 a_35904_26424# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X1372 vdd tune_shunt[7] a_25572_29076# vdd pmos_6p0 w=1.2u l=0.5u
X1373 vdd tune_shunt[7] a_6532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X1374 a_13796_40898# cap_shunt_n a_13588_41244# vdd pmos_6p0 w=1.2u l=0.5u
X1375 a_31624_8316# tune_series_gygy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X1376 vdd a_19948_50551# a_19860_50648# vdd pmos_6p0 w=1.22u l=1u
X1377 a_20532_27508# cap_shunt_n a_20740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X1378 a_27228_8215# a_27140_8312# vss vss nmos_6p0 w=0.82u l=1u
X1379 vdd tune_shunt[6] a_3620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X1380 a_8064_40536# cap_shunt_n a_6740_40536# vss nmos_6p0 w=0.82u l=0.6u
X1381 vdd tune_shunt[7] a_13588_39676# vdd pmos_6p0 w=1.2u l=0.5u
X1382 a_6508_38007# a_6420_38104# vss vss nmos_6p0 w=0.82u l=1u
X1383 a_15176_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1384 a_6740_13880# cap_shunt_p a_6532_13396# vdd pmos_6p0 w=1.2u l=0.5u
X1385 a_9332_16156# cap_shunt_p a_9540_15810# vdd pmos_6p0 w=1.2u l=0.5u
X1386 a_30800_18584# cap_series_gyp a_28692_18584# vss nmos_6p0 w=0.82u l=0.6u
X1387 a_14580_46808# cap_shunt_p a_16296_46808# vss nmos_6p0 w=0.82u l=0.6u
X1388 vdd a_15804_16488# a_15716_16532# vdd pmos_6p0 w=1.22u l=1u
X1389 a_37420_36439# a_37332_36536# vss vss nmos_6p0 w=0.82u l=1u
X1390 vss cap_shunt_p a_4032_6040# vss nmos_6p0 w=0.82u l=0.6u
X1391 vss cap_shunt_p a_8064_15448# vss nmos_6p0 w=0.82u l=0.6u
X1392 vss tune_shunt[7] a_13460_38968# vss nmos_6p0 w=0.51u l=0.6u
X1393 vss cap_shunt_p a_9856_43972# vss nmos_6p0 w=0.82u l=0.6u
X1394 a_27496_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1395 a_29700_29922# cap_shunt_p a_29492_30268# vdd pmos_6p0 w=1.2u l=0.5u
X1396 vss cap_shunt_p a_18816_17316# vss nmos_6p0 w=0.82u l=0.6u
X1397 a_33500_40008# a_33412_40052# vss vss nmos_6p0 w=0.82u l=1u
X1398 a_21748_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1399 a_30800_15448# cap_series_gyn a_28692_15448# vss nmos_6p0 w=0.82u l=0.6u
X1400 a_2500_17724# cap_shunt_p a_2708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X1401 a_6084_51028# cap_shunt_p a_6292_51512# vdd pmos_6p0 w=1.2u l=0.5u
X1402 a_34480_48438# cap_shunt_gyp a_34480_47893# vdd pmos_6p0 w=1.215u l=0.5u
X1403 vdd tune_series_gy[5] a_24452_13020# vdd pmos_6p0 w=1.2u l=0.5u
X1404 vdd a_28124_39575# a_28036_39672# vdd pmos_6p0 w=1.22u l=1u
X1405 vss cap_shunt_n a_9856_40836# vss nmos_6p0 w=0.82u l=0.6u
X1406 a_25780_40536# cap_shunt_n a_25572_40052# vdd pmos_6p0 w=1.2u l=0.5u
X1407 a_4032_47108# cap_shunt_p a_2708_47170# vss nmos_6p0 w=0.82u l=0.6u
X1408 a_25236_3612# cap_shunt_p a_25444_3266# vdd pmos_6p0 w=1.2u l=0.5u
X1409 a_34536_9884# cap_series_gygyn a_35344_9476# vss nmos_6p0 w=0.82u l=0.6u
X1410 a_37980_50984# a_37892_51028# vss vss nmos_6p0 w=0.82u l=1u
X1411 a_36288_39672# cap_shunt_gyn a_36308_39268# vss nmos_6p0 w=0.82u l=0.6u
X1412 a_32604_11784# a_32516_11828# vss vss nmos_6p0 w=0.82u l=1u
X1413 a_34308_17724# cap_series_gygyn a_34516_17378# vdd pmos_6p0 w=1.2u l=0.5u
X1414 vss cap_shunt_n a_12656_37400# vss nmos_6p0 w=0.82u l=0.6u
X1415 a_13588_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1416 a_13796_50306# cap_shunt_p a_13588_50652# vdd pmos_6p0 w=1.2u l=0.5u
X1417 vss tune_shunt[7] a_16708_28354# vss nmos_6p0 w=0.51u l=0.6u
X1418 vdd a_19388_54120# a_19300_54164# vdd pmos_6p0 w=1.22u l=1u
X1419 a_20532_36916# cap_shunt_n a_20740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X1420 vdd a_28124_36439# a_28036_36536# vdd pmos_6p0 w=1.22u l=1u
X1421 a_10340_24372# cap_shunt_n a_10548_24856# vdd pmos_6p0 w=1.2u l=0.5u
X1422 a_14580_40536# cap_shunt_n a_14372_40052# vdd pmos_6p0 w=1.2u l=0.5u
X1423 a_24660_34626# cap_shunt_p a_24452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X1424 a_31932_3511# a_31844_3608# vss vss nmos_6p0 w=0.82u l=1u
X1425 vss cap_series_gygyp a_37080_23288# vss nmos_6p0 w=0.82u l=0.6u
X1426 a_20172_44279# a_20084_44376# vss vss nmos_6p0 w=0.82u l=1u
X1427 a_14468_3266# cap_series_gyn a_14260_3612# vdd pmos_6p0 w=1.2u l=0.5u
X1428 a_10660_39330# cap_shunt_n a_10452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X1429 a_3620_14964# cap_shunt_p a_3828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X1430 a_36188_52552# a_36100_52596# vss vss nmos_6p0 w=0.82u l=1u
X1431 vss cap_shunt_n a_4704_51512# vss nmos_6p0 w=0.82u l=0.6u
X1432 vss tune_shunt[7] a_16708_25218# vss nmos_6p0 w=0.51u l=0.6u
X1433 vdd a_19388_50984# a_19300_51028# vdd pmos_6p0 w=1.22u l=1u
X1434 a_21964_48983# a_21876_49080# vss vss nmos_6p0 w=0.82u l=1u
X1435 a_24660_31490# cap_shunt_p a_24452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X1436 a_7540_39676# cap_shunt_n a_7748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X1437 a_11872_35832# cap_shunt_n a_10548_35832# vss nmos_6p0 w=0.82u l=0.6u
X1438 a_10360_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1439 a_2140_18056# a_2052_18100# vss vss nmos_6p0 w=0.82u l=1u
X1440 a_15580_50984# a_15492_51028# vss vss nmos_6p0 w=0.82u l=1u
X1441 a_20172_41143# a_20084_41240# vss vss nmos_6p0 w=0.82u l=1u
X1442 a_30408_40536# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1443 a_9876_12312# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1444 a_17640_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1445 a_29700_17378# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1446 a_25572_43188# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1447 vdd tune_series_gy[2] a_7580_6748# vdd pmos_6p0 w=1.2u l=0.5u
X1448 vdd a_35292_24328# a_35204_24372# vdd pmos_6p0 w=1.22u l=1u
X1449 a_28692_17016# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1450 vss cap_shunt_p a_11984_21720# vss nmos_6p0 w=0.82u l=0.6u
X1451 a_35488_41621# cap_shunt_gyn a_35488_42166# vdd pmos_6p0 w=1.215u l=0.5u
X1452 vdd a_10092_55255# a_10004_55352# vdd pmos_6p0 w=1.22u l=1u
X1453 a_2140_14920# a_2052_14964# vss vss nmos_6p0 w=0.82u l=1u
X1454 a_28484_3988# tune_series_gy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1455 vdd tune_shunt[4] a_21540_17724# vdd pmos_6p0 w=1.2u l=0.5u
X1456 vdd a_32604_53687# a_32516_53784# vdd pmos_6p0 w=1.22u l=1u
X1457 a_14372_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1458 a_12892_17623# a_12804_17720# vss vss nmos_6p0 w=0.82u l=1u
X1459 a_4816_45540# cap_shunt_p a_2708_45602# vss nmos_6p0 w=0.82u l=0.6u
X1460 vdd a_32156_3944# a_32068_3988# vdd pmos_6p0 w=1.22u l=1u
X1461 vdd a_35292_21192# a_35204_21236# vdd pmos_6p0 w=1.22u l=1u
X1462 a_17828_37400# cap_shunt_n a_17620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X1463 vss tune_series_gy[3] a_10680_8316# vss nmos_6p0 w=0.51u l=0.6u
X1464 vdd a_18492_8648# a_18404_8692# vdd pmos_6p0 w=1.22u l=1u
X1465 vdd tune_shunt[5] a_3172_18100# vdd pmos_6p0 w=1.2u l=0.5u
X1466 a_9316_48738# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1467 a_8064_34264# cap_shunt_n a_6740_34264# vss nmos_6p0 w=0.82u l=0.6u
X1468 vdd a_32604_50551# a_32516_50648# vdd pmos_6p0 w=1.22u l=1u
X1469 vdd a_2588_54120# a_2500_54164# vdd pmos_6p0 w=1.22u l=1u
X1470 vss cap_shunt_p a_11200_49944# vss nmos_6p0 w=0.82u l=0.6u
X1471 a_4816_42404# cap_shunt_p a_2708_42466# vss nmos_6p0 w=0.82u l=0.6u
X1472 a_21448_13880# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1473 a_35904_17016# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X1474 a_32612_37762# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X1475 vss cap_shunt_p a_14896_18584# vss nmos_6p0 w=0.82u l=0.6u
X1476 vdd tune_shunt[7] a_13252_32212# vdd pmos_6p0 w=1.2u l=0.5u
X1477 a_21524_4472# cap_series_gyn a_21316_3988# vdd pmos_6p0 w=1.2u l=0.5u
X1478 a_28348_55688# a_28260_55732# vss vss nmos_6p0 w=0.82u l=1u
X1479 a_23856_9476# cap_series_gyp a_21748_9538# vss nmos_6p0 w=0.82u l=0.6u
X1480 a_10660_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1481 a_26712_38968# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1482 vdd tune_shunt[7] a_3620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X1483 a_8064_31128# cap_shunt_n a_6740_31128# vss nmos_6p0 w=0.82u l=0.6u
X1484 vdd a_2588_50984# a_2500_51028# vdd pmos_6p0 w=1.22u l=1u
X1485 a_21448_10744# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1486 a_5636_11452# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1487 vss tune_shunt_gy[6] a_30688_45944# vss nmos_6p0 w=0.51u l=0.6u
X1488 a_32612_34626# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1489 vss cap_shunt_p a_14896_15448# vss nmos_6p0 w=0.82u l=0.6u
X1490 vdd a_5724_52552# a_5636_52596# vdd pmos_6p0 w=1.22u l=1u
X1491 vss cap_shunt_n a_9856_34564# vss nmos_6p0 w=0.82u l=0.6u
X1492 a_29384_3612# cap_series_gyn a_30192_3204# vss nmos_6p0 w=0.82u l=0.6u
X1493 vdd a_12332_22327# a_12244_22424# vdd pmos_6p0 w=1.22u l=1u
X1494 a_12556_9783# a_12468_9880# vss vss nmos_6p0 w=0.82u l=1u
X1495 a_18940_13352# a_18852_13396# vss vss nmos_6p0 w=0.82u l=1u
X1496 a_37980_44712# a_37892_44756# vss vss nmos_6p0 w=0.82u l=1u
X1497 vss tune_shunt[5] a_13796_48738# vss nmos_6p0 w=0.51u l=0.6u
X1498 a_13796_44034# cap_shunt_n a_13588_44380# vdd pmos_6p0 w=1.2u l=0.5u
X1499 a_3828_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1500 vss tune_series_gygy[3] a_34536_8316# vss nmos_6p0 w=0.51u l=0.6u
X1501 vdd a_32156_42711# a_32068_42808# vdd pmos_6p0 w=1.22u l=1u
X1502 vss cap_shunt_n a_9856_31428# vss nmos_6p0 w=0.82u l=0.6u
X1503 a_15700_9538# cap_series_gyn a_17416_9476# vss nmos_6p0 w=0.82u l=0.6u
X1504 a_32604_7080# a_32516_7124# vss vss nmos_6p0 w=0.82u l=1u
X1505 a_21748_4834# cap_series_gyp a_23464_4772# vss nmos_6p0 w=0.82u l=0.6u
X1506 a_18940_10216# a_18852_10260# vss vss nmos_6p0 w=0.82u l=1u
X1507 vss tune_shunt[7] a_10548_34264# vss nmos_6p0 w=0.51u l=0.6u
X1508 a_21540_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1509 a_13796_40898# cap_shunt_n a_13588_41244# vdd pmos_6p0 w=1.2u l=0.5u
X1510 a_9072_32996# cap_shunt_n a_7748_33058# vss nmos_6p0 w=0.82u l=0.6u
X1511 a_20532_27508# cap_shunt_n a_20740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X1512 a_3828_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1513 a_11424_22020# cap_shunt_p a_9316_22082# vss nmos_6p0 w=0.82u l=0.6u
X1514 vdd a_28124_27031# a_28036_27128# vdd pmos_6p0 w=1.22u l=1u
X1515 a_24660_25218# cap_shunt_p a_24452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X1516 a_20048_6040# cap_series_gyn a_18724_6040# vss nmos_6p0 w=0.82u l=0.6u
X1517 a_11872_29560# cap_shunt_n a_10548_29560# vss nmos_6p0 w=0.82u l=0.6u
X1518 a_30016_32696# cap_shunt_p a_28692_32696# vss nmos_6p0 w=0.82u l=0.6u
X1519 vss tune_shunt[7] a_10548_31128# vss nmos_6p0 w=0.51u l=0.6u
X1520 a_20172_34871# a_20084_34968# vss vss nmos_6p0 w=0.82u l=1u
X1521 a_30408_34264# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1522 a_21540_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1523 a_23756_44712# a_23668_44756# vss vss nmos_6p0 w=0.82u l=1u
X1524 vss tune_shunt[6] a_7748_42466# vss nmos_6p0 w=0.51u l=0.6u
X1525 a_24660_22082# cap_shunt_p a_24452_22428# vdd pmos_6p0 w=1.2u l=0.5u
X1526 vss tune_series_gy[3] a_25780_7608# vss nmos_6p0 w=0.51u l=0.6u
X1527 a_2500_17724# cap_shunt_p a_2708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X1528 a_34844_52119# a_34756_52216# vss vss nmos_6p0 w=0.82u l=1u
X1529 a_6084_51028# cap_shunt_p a_6292_51512# vdd pmos_6p0 w=1.2u l=0.5u
X1530 a_11872_26424# cap_shunt_n a_10548_26424# vss nmos_6p0 w=0.82u l=0.6u
X1531 a_32612_36194# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1532 a_20172_31735# a_20084_31832# vss vss nmos_6p0 w=0.82u l=1u
X1533 a_30408_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1534 a_12580_47892# cap_shunt_p a_12788_48376# vdd pmos_6p0 w=1.2u l=0.5u
X1535 a_23756_41576# a_23668_41620# vss vss nmos_6p0 w=0.82u l=1u
X1536 a_13460_37400# cap_shunt_n a_13252_36916# vdd pmos_6p0 w=1.2u l=0.5u
X1537 vss tune_shunt_gy[0] a_37632_33781# vss nmos_6p0 w=0.51u l=0.6u
X1538 a_28692_13880# cap_series_gyp a_30408_13880# vss nmos_6p0 w=0.82u l=0.6u
X1539 a_4940_5512# a_4852_5556# vss vss nmos_6p0 w=0.82u l=1u
X1540 vdd tune_series_gygy[0] a_35692_3988# vdd pmos_6p0 w=1.2u l=0.5u
X1541 a_11572_3988# cap_series_gyp a_11780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X1542 vss cap_shunt_p a_11984_12312# vss nmos_6p0 w=0.82u l=0.6u
X1543 a_8996_52220# cap_shunt_n a_9204_51874# vdd pmos_6p0 w=1.2u l=0.5u
X1544 a_1716_3612# cap_shunt_n a_1924_3266# vdd pmos_6p0 w=1.2u l=0.5u
X1545 a_25984_39268# cap_shunt_p a_24660_39330# vss nmos_6p0 w=0.82u l=0.6u
X1546 a_32612_33058# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1547 a_11200_13880# cap_shunt_p a_9876_13880# vss nmos_6p0 w=0.82u l=0.6u
X1548 vdd tune_shunt[5] a_29492_36540# vdd pmos_6p0 w=1.2u l=0.5u
X1549 a_24660_34626# cap_shunt_p a_24452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X1550 vdd tune_series_gy[5] a_21540_8316# vdd pmos_6p0 w=1.2u l=0.5u
X1551 a_33024_47512# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X1552 a_4816_36132# cap_shunt_n a_2708_36194# vss nmos_6p0 w=0.82u l=0.6u
X1553 a_28692_10744# cap_series_gyp a_30408_10744# vss nmos_6p0 w=0.82u l=0.6u
X1554 a_17828_27992# cap_shunt_n a_17620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X1555 a_6760_5556# cap_series_gyp a_6572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X1556 a_24660_15810# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1557 a_37644_35304# a_37556_35348# vss vss nmos_6p0 w=0.82u l=1u
X1558 a_10660_36194# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1559 a_11200_10744# cap_shunt_p a_9876_10744# vss nmos_6p0 w=0.82u l=0.6u
X1560 a_13796_50306# cap_shunt_p a_14728_50244# vss nmos_6p0 w=0.82u l=0.6u
X1561 vdd tune_shunt[5] a_29492_33404# vdd pmos_6p0 w=1.2u l=0.5u
X1562 a_24660_31490# cap_shunt_p a_24452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X1563 a_36688_6040# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X1564 a_31416_32996# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1565 a_35692_24372# cap_series_gygyp a_35880_24372# vdd pmos_6p0 w=1.2u l=0.5u
X1566 vdd a_35180_36439# a_35092_36536# vdd pmos_6p0 w=1.22u l=1u
X1567 a_32612_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1568 a_16708_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1569 a_4380_55255# a_4292_55352# vss vss nmos_6p0 w=0.82u l=1u
X1570 vss cap_shunt_n a_9856_28292# vss nmos_6p0 w=0.82u l=0.6u
X1571 vss cap_shunt_gyp a_36988_49944# vss nmos_6p0 w=0.82u l=0.6u
X1572 a_10660_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1573 vss cap_series_gyp a_19936_9476# vss nmos_6p0 w=0.82u l=0.6u
X1574 a_28484_14964# cap_series_gyn a_28692_15448# vdd pmos_6p0 w=1.2u l=0.5u
X1575 a_10548_3266# cap_series_gyn a_12264_3204# vss nmos_6p0 w=0.82u l=0.6u
X1576 a_16500_17724# cap_shunt_p a_16708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X1577 a_8232_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1578 a_35692_21236# cap_series_gygyp a_35880_21236# vdd pmos_6p0 w=1.2u l=0.5u
X1579 a_32612_25218# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1580 a_18404_8316# cap_series_gyp a_18612_7970# vdd pmos_6p0 w=1.2u l=0.5u
X1581 a_16708_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1582 vss cap_shunt_n a_4816_12612# vss nmos_6p0 w=0.82u l=0.6u
X1583 vdd a_36188_55688# a_36100_55732# vdd pmos_6p0 w=1.22u l=1u
X1584 vdd a_29580_52552# a_29492_52596# vdd pmos_6p0 w=1.22u l=1u
X1585 vss cap_shunt_n a_9856_25156# vss nmos_6p0 w=0.82u l=0.6u
X1586 a_11460_43188# cap_shunt_n a_11668_43672# vdd pmos_6p0 w=1.2u l=0.5u
X1587 a_9876_10744# cap_shunt_p a_9668_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1588 vss cap_shunt_gyp a_36988_46808# vss nmos_6p0 w=0.82u l=0.6u
X1589 a_28484_11828# cap_series_gyn a_28692_12312# vdd pmos_6p0 w=1.2u l=0.5u
X1590 a_3036_46280# a_2948_46324# vss vss nmos_6p0 w=0.82u l=1u
X1591 a_11612_7124# cap_series_gyp a_11800_7124# vdd pmos_6p0 w=1.2u l=0.5u
X1592 vss cap_series_gyp a_7176_6040# vss nmos_6p0 w=0.82u l=0.6u
X1593 vss cap_series_gygyn a_32824_7908# vss nmos_6p0 w=0.82u l=0.6u
X1594 a_36160_43734# tune_shunt_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X1595 a_6532_33780# cap_shunt_n a_6740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X1596 a_7616_17016# cap_shunt_p a_6292_17016# vss nmos_6p0 w=0.82u l=0.6u
X1597 a_3380_18584# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1598 a_31624_19292# cap_series_gygyn a_31648_18884# vss nmos_6p0 w=0.82u l=0.6u
X1599 a_24660_18946# cap_series_gyn a_24452_19292# vdd pmos_6p0 w=1.2u l=0.5u
X1600 a_10340_3612# cap_series_gyn a_10548_3266# vdd pmos_6p0 w=1.2u l=0.5u
X1601 a_20172_28599# a_20084_28696# vss vss nmos_6p0 w=0.82u l=1u
X1602 a_21540_25564# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1603 vss tune_shunt[7] a_2708_23650# vss nmos_6p0 w=0.51u l=0.6u
X1604 vss tune_shunt[6] a_7748_36194# vss nmos_6p0 w=0.51u l=0.6u
X1605 a_9072_23588# cap_shunt_p a_7748_23650# vss nmos_6p0 w=0.82u l=0.6u
X1606 a_6532_30644# cap_shunt_n a_6740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X1607 vdd a_24204_5512# a_24116_5556# vdd pmos_6p0 w=1.22u l=1u
X1608 a_3828_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1609 a_11460_46324# cap_shunt_n a_11668_46808# vdd pmos_6p0 w=1.2u l=0.5u
X1610 a_18180_3612# cap_series_gyn a_18388_3266# vdd pmos_6p0 w=1.2u l=0.5u
X1611 a_18612_12674# cap_series_gyn a_19544_12612# vss nmos_6p0 w=0.82u l=0.6u
X1612 a_24660_15810# cap_series_gyn a_24452_16156# vdd pmos_6p0 w=1.2u l=0.5u
X1613 a_3828_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1614 a_30016_23288# cap_shunt_p a_28692_23288# vss nmos_6p0 w=0.82u l=0.6u
X1615 a_20172_25463# a_20084_25560# vss vss nmos_6p0 w=0.82u l=1u
X1616 a_21540_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1617 a_10472_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1618 vss tune_shunt[5] a_2708_20514# vss nmos_6p0 w=0.51u l=0.6u
X1619 vss cap_shunt_p a_11424_47108# vss nmos_6p0 w=0.82u l=0.6u
X1620 vss tune_shunt[7] a_7748_33058# vss nmos_6p0 w=0.51u l=0.6u
X1621 a_10660_29922# cap_shunt_n a_11592_29860# vss nmos_6p0 w=0.82u l=0.6u
X1622 vdd a_8748_55688# a_8660_55732# vdd pmos_6p0 w=1.22u l=1u
X1623 a_3620_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1624 a_35880_21236# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1625 a_1924_4834# cap_shunt_p a_1716_5180# vdd pmos_6p0 w=1.2u l=0.5u
X1626 a_10472_11044# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1627 vss cap_series_gyn a_23072_12612# vss nmos_6p0 w=0.82u l=0.6u
X1628 a_13460_27992# cap_shunt_n a_13252_27508# vdd pmos_6p0 w=1.2u l=0.5u
X1629 a_9876_18584# cap_shunt_p a_9668_18100# vdd pmos_6p0 w=1.2u l=0.5u
X1630 vss cap_shunt_n a_19936_38968# vss nmos_6p0 w=0.82u l=0.6u
X1631 vdd tune_shunt[6] a_20532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X1632 vdd a_33500_36872# a_33412_36916# vdd pmos_6p0 w=1.22u l=1u
X1633 a_10660_26786# cap_shunt_n a_11592_26724# vss nmos_6p0 w=0.82u l=0.6u
X1634 a_5040_12312# cap_shunt_n a_2932_12312# vss nmos_6p0 w=0.82u l=0.6u
X1635 vdd a_28572_42711# a_28484_42808# vdd pmos_6p0 w=1.22u l=1u
X1636 a_2140_20759# a_2052_20856# vss vss nmos_6p0 w=0.82u l=1u
X1637 vdd a_16028_25896# a_15940_25940# vdd pmos_6p0 w=1.22u l=1u
X1638 a_18612_4472# cap_series_gyp a_19544_4472# vss nmos_6p0 w=0.82u l=0.6u
X1639 a_15720_11452# cap_series_gyp a_16528_11044# vss nmos_6p0 w=0.82u l=0.6u
X1640 vdd a_27676_17623# a_27588_17720# vdd pmos_6p0 w=1.22u l=1u
X1641 a_25780_20152# cap_series_gyp a_25572_19668# vdd pmos_6p0 w=1.2u l=0.5u
X1642 a_37644_29032# a_37556_29076# vss vss nmos_6p0 w=0.82u l=1u
X1643 vdd tune_shunt[7] a_29492_27132# vdd pmos_6p0 w=1.2u l=0.5u
X1644 a_24660_25218# cap_shunt_p a_24452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X1645 vdd a_36636_54120# a_36548_54164# vdd pmos_6p0 w=1.22u l=1u
X1646 a_27340_54120# a_27252_54164# vss vss nmos_6p0 w=0.82u l=1u
X1647 vdd a_35292_41143# a_35204_41240# vdd pmos_6p0 w=1.22u l=1u
X1648 vdd a_16028_22760# a_15940_22804# vdd pmos_6p0 w=1.22u l=1u
X1649 a_37080_20152# cap_series_gygyp a_35880_19668# vss nmos_6p0 w=0.82u l=0.6u
X1650 a_22644_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1651 vss tune_shunt[5] a_12788_49944# vss nmos_6p0 w=0.51u l=0.6u
X1652 a_24660_22082# cap_shunt_p a_24452_22428# vdd pmos_6p0 w=1.2u l=0.5u
X1653 a_6292_51512# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1654 vdd a_36636_50984# a_36548_51028# vdd pmos_6p0 w=1.22u l=1u
X1655 vdd a_35180_27031# a_35092_27128# vdd pmos_6p0 w=1.22u l=1u
X1656 a_31416_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1657 a_21748_12674# cap_series_gyn a_21540_13020# vdd pmos_6p0 w=1.2u l=0.5u
X1658 a_16708_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1659 vdd a_16700_55255# a_16612_55352# vdd pmos_6p0 w=1.22u l=1u
X1660 a_10548_38968# cap_shunt_n a_12264_38968# vss nmos_6p0 w=0.82u l=0.6u
X1661 vdd a_37868_34871# a_37780_34968# vdd pmos_6p0 w=1.22u l=1u
X1662 a_18404_5180# cap_series_gyp a_18612_4834# vdd pmos_6p0 w=1.2u l=0.5u
X1663 a_13460_37400# cap_shunt_n a_13252_36916# vdd pmos_6p0 w=1.2u l=0.5u
X1664 a_22644_10744# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1665 a_22848_21720# cap_shunt_p a_20740_21720# vss nmos_6p0 w=0.82u l=0.6u
X1666 a_24316_54120# a_24228_54164# vss vss nmos_6p0 w=0.82u l=1u
X1667 a_8400_48676# cap_shunt_p a_6292_48738# vss nmos_6p0 w=0.82u l=0.6u
X1668 a_9108_47516# cap_shunt_p a_9316_47170# vdd pmos_6p0 w=1.2u l=0.5u
X1669 vdd a_12892_10216# a_12804_10260# vdd pmos_6p0 w=1.22u l=1u
X1670 a_29700_14242# cap_series_gyp a_30632_14180# vss nmos_6p0 w=0.82u l=0.6u
X1671 vdd a_27004_55688# a_26916_55732# vdd pmos_6p0 w=1.22u l=1u
X1672 a_7540_34972# cap_shunt_n a_7748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X1673 a_28236_47415# a_28148_47512# vss vss nmos_6p0 w=0.82u l=1u
X1674 vdd a_10988_46280# a_10900_46324# vdd pmos_6p0 w=1.22u l=1u
X1675 a_24452_30268# cap_shunt_n a_24660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X1676 vss tune_shunt[7] a_6740_20152# vss nmos_6p0 w=0.51u l=0.6u
X1677 vdd a_16700_52119# a_16612_52216# vdd pmos_6p0 w=1.22u l=1u
X1678 a_15512_43972# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1679 a_24660_9538# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1680 vss tune_shunt[6] a_6740_43672# vss nmos_6p0 w=0.51u l=0.6u
X1681 a_5844_9176# cap_shunt_p a_5636_8692# vdd pmos_6p0 w=1.2u l=0.5u
X1682 vss cap_shunt_n a_8848_37400# vss nmos_6p0 w=0.82u l=0.6u
X1683 a_24660_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1684 a_29700_11106# cap_series_gyp a_30632_11044# vss nmos_6p0 w=0.82u l=0.6u
X1685 vdd a_14236_50984# a_14148_51028# vdd pmos_6p0 w=1.22u l=1u
X1686 vss tune_shunt[6] a_24660_39330# vss nmos_6p0 w=0.51u l=0.6u
X1687 a_7540_31836# cap_shunt_n a_7748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X1688 vss tune_shunt[4] a_32612_31490# vss nmos_6p0 w=0.51u l=0.6u
X1689 a_21540_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1690 a_29468_53687# a_29380_53784# vss vss nmos_6p0 w=0.82u l=1u
X1691 a_6956_38007# a_6868_38104# vss vss nmos_6p0 w=0.82u l=1u
X1692 a_6532_24372# cap_shunt_p a_6740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X1693 a_18760_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1694 a_35880_19668# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1695 a_23968_13880# cap_series_gyn a_22644_13880# vss nmos_6p0 w=0.82u l=0.6u
X1696 a_12788_49944# cap_shunt_n a_13720_49944# vss nmos_6p0 w=0.82u l=0.6u
X1697 a_15512_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1698 vss cap_shunt_p a_5488_18584# vss nmos_6p0 w=0.82u l=0.6u
X1699 vss tune_shunt[6] a_6740_40536# vss nmos_6p0 w=0.51u l=0.6u
X1700 vss tune_series_gy[4] a_24660_7970# vss nmos_6p0 w=0.51u l=0.6u
X1701 vss tune_shunt[4] a_2708_14242# vss nmos_6p0 w=0.51u l=0.6u
X1702 a_21540_16156# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1703 a_37420_55688# a_37332_55732# vss vss nmos_6p0 w=0.82u l=1u
X1704 a_29468_50551# a_29380_50648# vss vss nmos_6p0 w=0.82u l=1u
X1705 a_2708_28354# cap_shunt_n a_2500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X1706 a_1716_5556# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1707 a_10680_8316# cap_series_gyp a_10492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X1708 a_6532_21236# cap_shunt_p a_6740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X1709 a_9316_22082# cap_shunt_p a_9108_22428# vdd pmos_6p0 w=1.2u l=0.5u
X1710 a_14692_10744# cap_series_gyn a_15624_10744# vss nmos_6p0 w=0.82u l=0.6u
X1711 vss cap_shunt_n a_15568_32696# vss nmos_6p0 w=0.82u l=0.6u
X1712 a_23968_10744# cap_series_gyp a_22644_10744# vss nmos_6p0 w=0.82u l=0.6u
X1713 a_28484_14964# cap_series_gyn a_28692_15448# vdd pmos_6p0 w=1.2u l=0.5u
X1714 a_31624_20860# cap_series_gygyn a_31436_20860# vdd pmos_6p0 w=1.2u l=0.5u
X1715 a_6740_53080# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1716 vdd a_28572_39575# a_28484_39672# vdd pmos_6p0 w=1.22u l=1u
X1717 a_16500_47516# cap_shunt_n a_16708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X1718 vss tune_series_gy[3] a_24660_4834# vss nmos_6p0 w=0.51u l=0.6u
X1719 a_36188_38440# a_36100_38484# vss vss nmos_6p0 w=0.82u l=1u
X1720 vss tune_shunt[3] a_2708_11106# vss nmos_6p0 w=0.51u l=0.6u
X1721 a_11460_43188# cap_shunt_n a_11668_43672# vdd pmos_6p0 w=1.2u l=0.5u
X1722 a_7748_37762# cap_shunt_n a_7540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X1723 a_9876_10744# cap_shunt_p a_9668_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1724 a_35880_7124# cap_series_gygyp a_35904_7608# vss nmos_6p0 w=0.82u l=0.6u
X1725 a_28484_11828# cap_series_gyn a_28692_12312# vdd pmos_6p0 w=1.2u l=0.5u
X1726 a_24452_38108# cap_shunt_p a_24660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X1727 vdd a_28572_36439# a_28484_36536# vdd pmos_6p0 w=1.22u l=1u
X1728 a_18612_7970# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1729 a_2140_14487# a_2052_14584# vss vss nmos_6p0 w=0.82u l=1u
X1730 a_35880_11828# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1731 a_35692_19668# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1732 vdd a_1692_34871# a_1604_34968# vdd pmos_6p0 w=1.22u l=1u
X1733 vdd a_8860_19191# a_8772_19288# vdd pmos_6p0 w=1.22u l=1u
X1734 a_17620_47892# cap_shunt_p a_17828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X1735 a_24660_18946# cap_series_gyn a_24452_19292# vdd pmos_6p0 w=1.2u l=0.5u
X1736 vss cap_series_gyp a_30800_4472# vss nmos_6p0 w=0.82u l=0.6u
X1737 a_3828_26424# cap_shunt_p a_3620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X1738 vdd tune_shunt[7] a_6532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X1739 a_19544_9476# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X1740 vss cap_shunt_p a_27104_37400# vss nmos_6p0 w=0.82u l=0.6u
X1741 a_28484_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1742 a_10548_32696# cap_shunt_n a_10340_32212# vdd pmos_6p0 w=1.2u l=0.5u
X1743 a_13564_5079# a_13476_5176# vss vss nmos_6p0 w=0.82u l=1u
X1744 vdd a_31260_13352# a_31172_13396# vdd pmos_6p0 w=1.22u l=1u
X1745 a_30428_19668# cap_series_gygyn a_30616_19668# vdd pmos_6p0 w=1.2u l=0.5u
X1746 a_15624_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X1747 a_18612_4834# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1748 a_2140_11351# a_2052_11448# vss vss nmos_6p0 w=0.82u l=1u
X1749 a_27340_47848# a_27252_47892# vss vss nmos_6p0 w=0.82u l=1u
X1750 vdd a_29916_6647# a_29828_6744# vdd pmos_6p0 w=1.22u l=1u
X1751 a_8412_9783# a_8324_9880# vss vss nmos_6p0 w=0.82u l=1u
X1752 a_17620_44756# cap_shunt_p a_17828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X1753 a_25592_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1754 a_24660_15810# cap_series_gyn a_24452_16156# vdd pmos_6p0 w=1.2u l=0.5u
X1755 a_2708_50306# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1756 vss tune_shunt[7] a_7748_23650# vss nmos_6p0 w=0.51u l=0.6u
X1757 a_3828_23288# cap_shunt_p a_3620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X1758 vdd tune_shunt[7] a_6532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X1759 vdd a_37868_28599# a_37780_28696# vdd pmos_6p0 w=1.22u l=1u
X1760 a_32432_7908# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X1761 vdd tune_series_gy[4] a_29532_13020# vdd pmos_6p0 w=1.2u l=0.5u
X1762 vss cap_series_gygyn a_31816_20152# vss nmos_6p0 w=0.82u l=0.6u
X1763 vss tune_shunt[7] a_20740_32696# vss nmos_6p0 w=0.51u l=0.6u
X1764 a_10452_28700# cap_shunt_n a_10660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X1765 vdd tune_shunt[6] a_9668_47892# vdd pmos_6p0 w=1.2u l=0.5u
X1766 vdd a_31708_33736# a_31620_33780# vdd pmos_6p0 w=1.22u l=1u
X1767 a_4424_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1768 a_13460_27992# cap_shunt_n a_13252_27508# vdd pmos_6p0 w=1.2u l=0.5u
X1769 a_12788_12312# cap_shunt_p a_14504_12312# vss nmos_6p0 w=0.82u l=0.6u
X1770 a_16708_34626# cap_shunt_n a_16500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X1771 a_6508_6647# a_6420_6744# vss vss nmos_6p0 w=0.82u l=1u
X1772 a_12788_48376# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1773 vss cap_shunt_n a_34720_34564# vss nmos_6p0 w=0.82u l=0.6u
X1774 a_7768_6748# cap_series_gyp a_8576_6340# vss nmos_6p0 w=0.82u l=0.6u
X1775 a_7540_25564# cap_shunt_n a_7748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X1776 a_25780_20152# cap_series_gyp a_25572_19668# vdd pmos_6p0 w=1.2u l=0.5u
X1777 a_24204_55255# a_24116_55352# vss vss nmos_6p0 w=0.82u l=1u
X1778 vdd a_31708_30600# a_31620_30644# vdd pmos_6p0 w=1.22u l=1u
X1779 vss cap_shunt_p a_22848_46808# vss nmos_6p0 w=0.82u l=0.6u
X1780 a_4424_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1781 a_15512_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1782 a_16708_31490# cap_shunt_n a_16500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X1783 vss tune_shunt[7] a_6740_34264# vss nmos_6p0 w=0.51u l=0.6u
X1784 a_24660_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1785 a_3036_52119# a_2948_52216# vss vss nmos_6p0 w=0.82u l=1u
X1786 vss cap_shunt_n a_34720_31428# vss nmos_6p0 w=0.82u l=0.6u
X1787 a_33732_27992# cap_shunt_p a_35448_27992# vss nmos_6p0 w=0.82u l=0.6u
X1788 vdd a_31708_8648# a_31620_8692# vdd pmos_6p0 w=1.22u l=1u
X1789 vdd a_35628_38007# a_35540_38104# vdd pmos_6p0 w=1.22u l=1u
X1790 a_18760_23288# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1791 vdd tune_series_gy[5] a_21540_9884# vdd pmos_6p0 w=1.2u l=0.5u
X1792 a_15512_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1793 a_2500_49084# cap_shunt_p a_2708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X1794 vss tune_shunt[7] a_6740_31128# vss nmos_6p0 w=0.51u l=0.6u
X1795 a_12788_13880# cap_shunt_p a_12580_13396# vdd pmos_6p0 w=1.2u l=0.5u
X1796 vdd a_12780_22327# a_12692_22424# vdd pmos_6p0 w=1.22u l=1u
X1797 vdd a_31708_5512# a_31620_5556# vdd pmos_6p0 w=1.22u l=1u
X1798 a_20740_45240# cap_shunt_n a_22456_45240# vss nmos_6p0 w=0.82u l=0.6u
X1799 a_6420_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1800 vdd tune_series_gy[4] a_21540_6748# vdd pmos_6p0 w=1.2u l=0.5u
X1801 vss tune_shunt[7] a_13796_18946# vss nmos_6p0 w=0.51u l=0.6u
X1802 a_34516_20514# cap_series_gygyp a_34308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X1803 vss cap_series_gygyp a_35840_23588# vss nmos_6p0 w=0.82u l=0.6u
X1804 vss cap_shunt_n a_15568_23288# vss nmos_6p0 w=0.82u l=0.6u
X1805 a_9108_47516# cap_shunt_p a_9316_47170# vdd pmos_6p0 w=1.2u l=0.5u
X1806 a_23072_22020# cap_shunt_p a_21748_22082# vss nmos_6p0 w=0.82u l=0.6u
X1807 a_29244_21192# a_29156_21236# vss vss nmos_6p0 w=0.82u l=1u
X1808 a_16500_38108# cap_shunt_n a_16708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X1809 a_24452_30268# cap_shunt_n a_24660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X1810 a_30812_44279# a_30724_44376# vss vss nmos_6p0 w=0.82u l=1u
X1811 vdd a_1692_28599# a_1604_28696# vdd pmos_6p0 w=1.22u l=1u
X1812 a_7560_3204# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1813 a_25572_8692# cap_series_gyp a_25780_9176# vdd pmos_6p0 w=1.2u l=0.5u
X1814 a_20740_42104# cap_shunt_p a_22456_42104# vss nmos_6p0 w=0.82u l=0.6u
X1815 vdd tune_series_gygy[3] a_34348_9884# vdd pmos_6p0 w=1.2u l=0.5u
X1816 a_2708_47170# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1817 a_15492_9884# cap_series_gyn a_15700_9538# vdd pmos_6p0 w=1.2u l=0.5u
X1818 a_13496_6040# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1819 vdd tune_shunt[4] a_33524_32212# vdd pmos_6p0 w=1.2u l=0.5u
X1820 vdd a_28572_27031# a_28484_27128# vdd pmos_6p0 w=1.22u l=1u
X1821 a_31372_54120# a_31284_54164# vss vss nmos_6p0 w=0.82u l=1u
X1822 a_21672_43672# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1823 a_32404_34972# cap_shunt_n a_32612_34626# vdd pmos_6p0 w=1.2u l=0.5u
X1824 a_30812_41143# a_30724_41240# vss vss nmos_6p0 w=0.82u l=1u
X1825 a_17620_38484# cap_shunt_n a_17828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X1826 a_25592_36132# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1827 a_25572_5556# cap_series_gyp a_25780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X1828 a_34952_7908# cap_series_gygyp a_34536_8316# vss nmos_6p0 w=0.82u l=0.6u
X1829 vdd tune_series_gygy[2] a_34348_6748# vdd pmos_6p0 w=1.2u l=0.5u
X1830 a_2708_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1831 a_15492_6748# cap_series_gyp a_15700_6402# vdd pmos_6p0 w=1.2u l=0.5u
X1832 a_28484_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1833 a_8456_13880# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1834 vdd a_20732_55255# a_20644_55352# vdd pmos_6p0 w=1.22u l=1u
X1835 a_21672_40536# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1836 a_2708_28354# cap_shunt_n a_2500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X1837 vdd a_10092_54120# a_10004_54164# vdd pmos_6p0 w=1.22u l=1u
X1838 a_32404_31836# cap_shunt_n a_32612_31490# vdd pmos_6p0 w=1.2u l=0.5u
X1839 a_32824_22020# cap_series_gygyn a_31624_22428# vss nmos_6p0 w=0.82u l=0.6u
X1840 a_25572_18100# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1841 a_20532_46324# cap_shunt_p a_20740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X1842 a_17620_35348# cap_shunt_n a_17828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X1843 a_28484_14964# cap_series_gyn a_28692_15448# vdd pmos_6p0 w=1.2u l=0.5u
X1844 a_33732_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1845 vdd a_36076_14487# a_35988_14584# vdd pmos_6p0 w=1.22u l=1u
X1846 a_16500_47516# cap_shunt_n a_16708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X1847 a_21748_44034# cap_shunt_n a_23464_43972# vss nmos_6p0 w=0.82u l=0.6u
X1848 a_13588_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1849 a_5612_22327# a_5524_22424# vss vss nmos_6p0 w=0.82u l=1u
X1850 a_21540_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1851 vdd a_37868_19191# a_37780_19288# vdd pmos_6p0 w=1.22u l=1u
X1852 vdd a_20732_52119# a_20644_52216# vdd pmos_6p0 w=1.22u l=1u
X1853 a_6060_45847# a_5972_45944# vss vss nmos_6p0 w=0.82u l=1u
X1854 a_36384_45540# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1855 a_21748_7970# cap_series_gyp a_21540_8316# vdd pmos_6p0 w=1.2u l=0.5u
X1856 a_13796_48738# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1857 a_7748_37762# cap_shunt_n a_7540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X1858 a_9876_10744# cap_shunt_p a_9668_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1859 vss cap_shunt_p a_34720_28292# vss nmos_6p0 w=0.82u l=0.6u
X1860 vss tune_shunt[7] a_20740_23288# vss nmos_6p0 w=0.51u l=0.6u
X1861 vdd a_36076_11351# a_35988_11448# vdd pmos_6p0 w=1.22u l=1u
X1862 a_28484_11828# cap_series_gyn a_28692_12312# vdd pmos_6p0 w=1.2u l=0.5u
X1863 a_24660_12674# cap_series_gyn a_25592_12612# vss nmos_6p0 w=0.82u l=0.6u
X1864 a_21748_40898# cap_shunt_p a_23464_40836# vss nmos_6p0 w=0.82u l=0.6u
X1865 vdd a_31708_24328# a_31620_24372# vdd pmos_6p0 w=1.22u l=1u
X1866 vss cap_series_gyp a_24752_9176# vss nmos_6p0 w=0.82u l=0.6u
X1867 a_9540_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1868 a_24204_48983# a_24116_49080# vss vss nmos_6p0 w=0.82u l=1u
X1869 a_13460_26424# cap_shunt_n a_13252_25940# vdd pmos_6p0 w=1.2u l=0.5u
X1870 a_6060_42711# a_5972_42808# vss vss nmos_6p0 w=0.82u l=1u
X1871 a_36384_42404# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X1872 a_5936_37400# cap_shunt_n a_3828_37400# vss nmos_6p0 w=0.82u l=0.6u
X1873 vss cap_shunt_p a_30800_32696# vss nmos_6p0 w=0.82u l=0.6u
X1874 a_15512_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1875 a_16708_25218# cap_shunt_n a_16500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X1876 a_3932_54120# a_3844_54164# vss vss nmos_6p0 w=0.82u l=1u
X1877 vdd a_30588_43144# a_30500_43188# vdd pmos_6p0 w=1.22u l=1u
X1878 vss cap_shunt_p a_34720_25156# vss nmos_6p0 w=0.82u l=0.6u
X1879 vss tune_shunt[2] a_1924_7608# vss nmos_6p0 w=0.51u l=0.6u
X1880 a_19612_55688# a_19524_55732# vss vss nmos_6p0 w=0.82u l=1u
X1881 a_16500_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1882 a_13460_23288# cap_shunt_n a_13252_22804# vdd pmos_6p0 w=1.2u l=0.5u
X1883 a_2708_29922# cap_shunt_n a_2500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X1884 a_15512_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1885 a_16708_22082# cap_shunt_n a_16500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X1886 a_4424_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1887 a_21524_3266# cap_series_gyp a_21316_3612# vdd pmos_6p0 w=1.2u l=0.5u
X1888 vss cap_shunt_p a_8064_43672# vss nmos_6p0 w=0.82u l=0.6u
X1889 a_10988_5512# a_10900_5556# vss vss nmos_6p0 w=0.82u l=1u
X1890 vss tune_shunt[5] a_3380_49944# vss nmos_6p0 w=0.51u l=0.6u
X1891 a_6532_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1892 a_9332_9884# cap_shunt_p a_9540_9538# vdd pmos_6p0 w=1.2u l=0.5u
X1893 a_25780_15448# cap_series_gyp a_25572_14964# vdd pmos_6p0 w=1.2u l=0.5u
X1894 vss cap_shunt_p a_18816_45540# vss nmos_6p0 w=0.82u l=0.6u
X1895 vss tune_shunt[4] a_32612_36194# vss nmos_6p0 w=0.51u l=0.6u
X1896 a_16708_28354# cap_shunt_n a_16500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X1897 vdd tune_series_gy[4] a_29532_13020# vdd pmos_6p0 w=1.2u l=0.5u
X1898 a_2708_37762# cap_shunt_n a_3640_37700# vss nmos_6p0 w=0.82u l=0.6u
X1899 a_10452_28700# cap_shunt_n a_10660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X1900 vss cap_shunt_n a_14784_38968# vss nmos_6p0 w=0.82u l=0.6u
X1901 a_20740_34264# cap_shunt_n a_20532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X1902 a_16016_6040# cap_series_gyn a_14692_6040# vss nmos_6p0 w=0.82u l=0.6u
X1903 a_10340_3612# cap_series_gyn a_10548_3266# vdd pmos_6p0 w=1.2u l=0.5u
X1904 vss cap_shunt_n a_8064_40536# vss nmos_6p0 w=0.82u l=0.6u
X1905 a_6532_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1906 a_21524_4472# cap_series_gyn a_23240_4472# vss nmos_6p0 w=0.82u l=0.6u
X1907 a_25780_12312# cap_series_gyp a_25572_11828# vdd pmos_6p0 w=1.2u l=0.5u
X1908 vss cap_shunt_n a_18816_42404# vss nmos_6p0 w=0.82u l=0.6u
X1909 vss tune_shunt[4] a_32612_33058# vss nmos_6p0 w=0.51u l=0.6u
X1910 vdd tune_series_gygy[1] a_31436_8316# vdd pmos_6p0 w=1.2u l=0.5u
X1911 a_2500_42812# cap_shunt_p a_2708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X1912 a_30800_40536# cap_shunt_p a_28692_40536# vss nmos_6p0 w=0.82u l=0.6u
X1913 a_20740_31128# cap_shunt_n a_20532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X1914 a_5844_10744# cap_shunt_p a_5636_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1915 vss tune_series_gy[4] a_28692_12312# vss nmos_6p0 w=0.51u l=0.6u
X1916 a_6628_14242# cap_shunt_p a_7560_14180# vss nmos_6p0 w=0.82u l=0.6u
X1917 a_31372_47848# a_31284_47892# vss vss nmos_6p0 w=0.82u l=1u
X1918 vss cap_shunt_n a_5936_27992# vss nmos_6p0 w=0.82u l=0.6u
X1919 a_29720_9884# cap_series_gyn a_29532_9884# vdd pmos_6p0 w=1.2u l=0.5u
X1920 vdd a_1692_19191# a_1604_19288# vdd pmos_6p0 w=1.22u l=1u
X1921 a_17828_48376# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X1922 vss cap_shunt_p a_18032_18884# vss nmos_6p0 w=0.82u l=0.6u
X1923 a_17828_35832# cap_shunt_n a_19544_35832# vss nmos_6p0 w=0.82u l=0.6u
X1924 vdd a_29468_20759# a_29380_20856# vdd pmos_6p0 w=1.22u l=1u
X1925 a_27888_35832# cap_shunt_p a_25780_35832# vss nmos_6p0 w=0.82u l=0.6u
X1926 vdd a_16924_33736# a_16836_33780# vdd pmos_6p0 w=1.22u l=1u
X1927 a_26376_18884# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1928 a_19724_30167# a_19636_30264# vss vss nmos_6p0 w=0.82u l=1u
X1929 a_17024_7908# cap_series_gyn a_15700_7970# vss nmos_6p0 w=0.82u l=0.6u
X1930 a_5844_11106# cap_shunt_n a_7560_11044# vss nmos_6p0 w=0.82u l=0.6u
X1931 a_18044_11784# a_17956_11828# vss vss nmos_6p0 w=0.82u l=1u
X1932 a_21672_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1933 a_32404_25564# cap_shunt_p a_32612_25218# vdd pmos_6p0 w=1.2u l=0.5u
X1934 vss cap_shunt_p a_5936_24856# vss nmos_6p0 w=0.82u l=0.6u
X1935 vss tune_shunt[7] a_21748_26786# vss nmos_6p0 w=0.51u l=0.6u
X1936 a_12376_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1937 a_12580_16532# cap_shunt_p a_12788_17016# vdd pmos_6p0 w=1.2u l=0.5u
X1938 a_17620_29076# cap_shunt_n a_17828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X1939 a_29532_16156# cap_series_gyn a_29720_16156# vdd pmos_6p0 w=1.2u l=0.5u
X1940 vss cap_shunt_p a_18032_15748# vss nmos_6p0 w=0.82u l=0.6u
X1941 a_31260_55255# a_31172_55352# vss vss nmos_6p0 w=0.82u l=1u
X1942 vdd a_16924_30600# a_16836_30644# vdd pmos_6p0 w=1.22u l=1u
X1943 a_26376_15748# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X1944 a_27340_53687# a_27252_53784# vss vss nmos_6p0 w=0.82u l=1u
X1945 a_19724_27031# a_19636_27128# vss vss nmos_6p0 w=0.82u l=1u
X1946 a_21672_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1947 a_13460_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1948 a_21840_13880# cap_series_gyn a_19732_13880# vss nmos_6p0 w=0.82u l=0.6u
X1949 a_34516_20514# cap_series_gygyp a_34308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X1950 a_9876_49944# cap_shunt_p a_11592_49944# vss nmos_6p0 w=0.82u l=0.6u
X1951 a_1924_4834# cap_shunt_p a_2856_4772# vss nmos_6p0 w=0.82u l=0.6u
X1952 vdd a_27228_33303# a_27140_33400# vdd pmos_6p0 w=1.22u l=1u
X1953 a_10660_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X1954 a_2140_43144# a_2052_43188# vss vss nmos_6p0 w=0.82u l=1u
X1955 a_35404_39575# a_35316_39672# vss vss nmos_6p0 w=0.82u l=1u
X1956 a_16500_38108# cap_shunt_n a_16708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X1957 a_21748_34626# cap_shunt_p a_23464_34564# vss nmos_6p0 w=0.82u l=0.6u
X1958 a_24452_30268# cap_shunt_n a_24660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X1959 a_21540_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1960 a_27340_50551# a_27252_50648# vss vss nmos_6p0 w=0.82u l=1u
X1961 a_33948_36872# a_33860_36916# vss vss nmos_6p0 w=0.82u l=1u
X1962 a_23072_9476# cap_series_gyp a_21748_9538# vss nmos_6p0 w=0.82u l=0.6u
X1963 a_6060_36439# a_5972_36536# vss vss nmos_6p0 w=0.82u l=1u
X1964 a_13460_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X1965 a_16708_18946# cap_shunt_p a_16500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X1966 vss tune_shunt[5] a_3828_48376# vss nmos_6p0 w=0.51u l=0.6u
X1967 vdd a_16476_25896# a_16388_25940# vdd pmos_6p0 w=1.22u l=1u
X1968 a_21840_10744# cap_series_gyn a_19732_10744# vss nmos_6p0 w=0.82u l=0.6u
X1969 a_10340_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1970 a_29720_13020# cap_series_gyn a_29744_12612# vss nmos_6p0 w=0.82u l=0.6u
X1971 vdd tune_shunt_gy[3] a_37444_45944# vdd pmos_6p0 w=1.215u l=0.5u
X1972 a_2140_40008# a_2052_40052# vss vss nmos_6p0 w=0.82u l=1u
X1973 a_32404_34972# cap_shunt_n a_32612_34626# vdd pmos_6p0 w=1.2u l=0.5u
X1974 a_21748_31490# cap_shunt_n a_23464_31428# vss nmos_6p0 w=0.82u l=0.6u
X1975 vss cap_shunt_p a_30800_23288# vss nmos_6p0 w=0.82u l=0.6u
X1976 vdd a_18044_53687# a_17956_53784# vdd pmos_6p0 w=1.22u l=1u
X1977 vdd tune_shunt[5] a_21540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X1978 a_28692_37400# cap_shunt_p a_29624_37400# vss nmos_6p0 w=0.82u l=0.6u
X1979 a_16708_15810# cap_shunt_p a_16500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X1980 vdd a_32156_38440# a_32068_38484# vdd pmos_6p0 w=1.22u l=1u
X1981 vdd a_16476_22760# a_16388_22804# vdd pmos_6p0 w=1.22u l=1u
X1982 vss tune_series_gy[3] a_28692_7608# vss nmos_6p0 w=0.51u l=0.6u
X1983 vdd tune_shunt[6] a_6532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X1984 a_22680_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X1985 a_10340_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1986 a_7960_7608# cap_series_gyp a_6760_7124# vss nmos_6p0 w=0.82u l=0.6u
X1987 a_28692_10744# cap_series_gyp a_28484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X1988 vdd tune_shunt_gy[2] a_37444_42808# vdd pmos_6p0 w=1.215u l=0.5u
X1989 a_35692_14964# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X1990 vdd tune_shunt[5] a_28484_38484# vdd pmos_6p0 w=1.2u l=0.5u
X1991 a_32404_31836# cap_shunt_n a_32612_31490# vdd pmos_6p0 w=1.2u l=0.5u
X1992 a_20532_46324# cap_shunt_p a_20740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X1993 a_15700_9538# cap_series_gyn a_16632_9476# vss nmos_6p0 w=0.82u l=0.6u
X1994 a_16708_20514# cap_shunt_p a_16500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X1995 a_2856_4472# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X1996 vdd a_37420_8215# a_37332_8312# vdd pmos_6p0 w=1.22u l=1u
X1997 vdd a_32156_35304# a_32068_35348# vdd pmos_6p0 w=1.22u l=1u
X1998 vss cap_shunt_n a_8064_34264# vss nmos_6p0 w=0.82u l=0.6u
X1999 a_24764_54120# a_24676_54164# vss vss nmos_6p0 w=0.82u l=1u
X2000 a_32464_45302# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2001 a_31248_44757# cap_shunt_gyn a_31060_44757# vdd pmos_6p0 w=1.215u l=0.5u
X2002 vss tune_series_gy[3] a_21524_4472# vss nmos_6p0 w=0.51u l=0.6u
X2003 a_35692_11828# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2004 vdd a_27452_55688# a_27364_55732# vdd pmos_6p0 w=1.22u l=1u
X2005 a_28684_47415# a_28596_47512# vss vss nmos_6p0 w=0.82u l=1u
X2006 vss cap_shunt_n a_18816_36132# vss nmos_6p0 w=0.82u l=0.6u
X2007 vdd tune_shunt[6] a_28484_35348# vdd pmos_6p0 w=1.2u l=0.5u
X2008 a_6532_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2009 a_29384_3612# cap_series_gyn a_29196_3612# vdd pmos_6p0 w=1.2u l=0.5u
X2010 a_3828_48376# cap_shunt_p a_4760_48376# vss nmos_6p0 w=0.82u l=0.6u
X2011 a_2500_36540# cap_shunt_n a_2708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X2012 a_20740_24856# cap_shunt_n a_20532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X2013 vdd tune_shunt[6] a_24452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X2014 a_30800_34264# cap_shunt_p a_28692_34264# vss nmos_6p0 w=0.82u l=0.6u
X2015 a_15568_37400# cap_shunt_n a_13460_37400# vss nmos_6p0 w=0.82u l=0.6u
X2016 vss cap_shunt_n a_8064_31128# vss nmos_6p0 w=0.82u l=0.6u
X2017 vdd a_14684_50984# a_14596_51028# vdd pmos_6p0 w=1.22u l=1u
X2018 a_13460_26424# cap_shunt_n a_13252_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2019 a_35880_21236# cap_series_gygyp a_35904_21720# vss nmos_6p0 w=0.82u l=0.6u
X2020 a_7748_42466# cap_shunt_n a_7540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X2021 vss tune_shunt[7] a_21748_29922# vss nmos_6p0 w=0.51u l=0.6u
X2022 a_17828_29560# cap_shunt_n a_19544_29560# vss nmos_6p0 w=0.82u l=0.6u
X2023 a_10680_8316# cap_series_gyp a_10492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X2024 a_6532_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2025 vdd a_24428_55688# a_24340_55732# vdd pmos_6p0 w=1.22u l=1u
X2026 a_6740_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2027 a_25572_36916# cap_shunt_p a_25780_37400# vdd pmos_6p0 w=1.2u l=0.5u
X2028 vdd a_17596_11784# a_17508_11828# vdd pmos_6p0 w=1.22u l=1u
X2029 a_34396_13352# a_34308_13396# vss vss nmos_6p0 w=0.82u l=1u
X2030 vss tune_shunt[5] a_6292_17378# vss nmos_6p0 w=0.51u l=0.6u
X2031 a_3620_19668# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2032 a_32612_37762# cap_shunt_p a_32404_38108# vdd pmos_6p0 w=1.2u l=0.5u
X2033 a_2500_33404# cap_shunt_p a_2708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X2034 a_27888_29560# cap_shunt_p a_25780_29560# vss nmos_6p0 w=0.82u l=0.6u
X2035 a_30800_31128# cap_shunt_n a_28692_31128# vss nmos_6p0 w=0.82u l=0.6u
X2036 a_20740_21720# cap_shunt_p a_20532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X2037 vss tune_shunt[5] a_16708_47170# vss nmos_6p0 w=0.51u l=0.6u
X2038 a_20284_52552# a_20196_52596# vss vss nmos_6p0 w=0.82u l=1u
X2039 a_7616_51512# cap_shunt_p a_6292_51512# vss nmos_6p0 w=0.82u l=0.6u
X2040 vdd tune_shunt[7] a_20532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X2041 vss cap_shunt_n a_31024_37700# vss nmos_6p0 w=0.82u l=0.6u
X2042 a_13460_23288# cap_shunt_n a_13252_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2043 a_17828_26424# cap_shunt_n a_19544_26424# vss nmos_6p0 w=0.82u l=0.6u
X2044 vss cap_series_gyp a_7960_7608# vss nmos_6p0 w=0.82u l=0.6u
X2045 a_31260_48983# a_31172_49080# vss vss nmos_6p0 w=0.82u l=1u
X2046 a_13252_33780# cap_shunt_n a_13460_34264# vdd pmos_6p0 w=1.2u l=0.5u
X2047 a_34396_10216# a_34308_10260# vss vss nmos_6p0 w=0.82u l=1u
X2048 vss tune_series_gy[5] a_22644_13880# vss nmos_6p0 w=0.51u l=0.6u
X2049 a_8008_50244# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2050 a_27888_26424# cap_shunt_p a_25780_26424# vss nmos_6p0 w=0.82u l=0.6u
X2051 vdd a_16924_24328# a_16836_24372# vdd pmos_6p0 w=1.22u l=1u
X2052 a_3172_16532# cap_shunt_p a_3380_17016# vdd pmos_6p0 w=1.2u l=0.5u
X2053 a_28692_26424# cap_shunt_p a_28484_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2054 vss tune_shunt[6] a_16708_44034# vss nmos_6p0 w=0.51u l=0.6u
X2055 a_3620_33780# cap_shunt_n a_3828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X2056 a_13588_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2057 a_25780_15448# cap_series_gyp a_25572_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2058 vss cap_shunt_p a_5936_15448# vss nmos_6p0 w=0.82u l=0.6u
X2059 vss tune_shunt[4] a_21748_17378# vss nmos_6p0 w=0.51u l=0.6u
X2060 a_11032_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2061 a_35880_7124# cap_series_gygyp a_35692_7124# vdd pmos_6p0 w=1.2u l=0.5u
X2062 vss tune_series_gygy[5] a_34516_18946# vss nmos_6p0 w=0.51u l=0.6u
X2063 vdd a_25548_47848# a_25460_47892# vdd pmos_6p0 w=1.22u l=1u
X2064 vss cap_shunt_n a_9072_32996# vss nmos_6p0 w=0.82u l=0.6u
X2065 a_10452_28700# cap_shunt_n a_10660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X2066 vss tune_shunt[7] a_10660_31490# vss nmos_6p0 w=0.51u l=0.6u
X2067 vss tune_shunt[7] a_9876_13880# vss nmos_6p0 w=0.51u l=0.6u
X2068 a_10660_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2069 a_13252_30644# cap_shunt_n a_13460_31128# vdd pmos_6p0 w=1.2u l=0.5u
X2070 a_21748_28354# cap_shunt_n a_23464_28292# vss nmos_6p0 w=0.82u l=0.6u
X2071 vss tune_series_gy[5] a_22644_10744# vss nmos_6p0 w=0.51u l=0.6u
X2072 a_34844_55688# a_34756_55732# vss vss nmos_6p0 w=0.82u l=1u
X2073 a_29700_36194# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2074 a_19724_17623# a_19636_17720# vss vss nmos_6p0 w=0.82u l=1u
X2075 vdd a_16924_21192# a_16836_21236# vdd pmos_6p0 w=1.22u l=1u
X2076 a_28692_23288# cap_shunt_p a_28484_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2077 a_33732_35832# cap_shunt_n a_33524_35348# vdd pmos_6p0 w=1.2u l=0.5u
X2078 a_3620_30644# cap_shunt_n a_3828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X2079 a_25780_12312# cap_series_gyp a_25572_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2080 vss cap_shunt_n a_15120_20452# vss nmos_6p0 w=0.82u l=0.6u
X2081 a_35904_6040# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X2082 a_6740_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2083 vdd a_25548_44712# a_25460_44756# vdd pmos_6p0 w=1.22u l=1u
X2084 vdd tune_shunt_gy[1] a_37444_39672# vdd pmos_6p0 w=1.215u l=0.5u
X2085 a_28124_33303# a_28036_33400# vss vss nmos_6p0 w=0.82u l=1u
X2086 a_30028_50984# a_29940_51028# vss vss nmos_6p0 w=0.82u l=1u
X2087 a_2500_42812# cap_shunt_p a_2708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X2088 a_29800_3204# cap_series_gyn a_29384_3612# vss nmos_6p0 w=0.82u l=0.6u
X2089 vss tune_shunt[7] a_9876_10744# vss nmos_6p0 w=0.51u l=0.6u
X2090 vss cap_shunt_n a_13776_45240# vss nmos_6p0 w=0.82u l=0.6u
X2091 a_2140_33736# a_2052_33780# vss vss nmos_6p0 w=0.82u l=1u
X2092 a_21748_25218# cap_shunt_n a_23464_25156# vss nmos_6p0 w=0.82u l=0.6u
X2093 a_6420_13020# cap_shunt_p a_6628_12674# vdd pmos_6p0 w=1.2u l=0.5u
X2094 a_29700_33058# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2095 a_21524_3266# cap_series_gyp a_21316_3612# vdd pmos_6p0 w=1.2u l=0.5u
X2096 vdd tune_shunt[6] a_21540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X2097 vdd a_35292_40008# a_35204_40052# vdd pmos_6p0 w=1.22u l=1u
X2098 a_9332_9884# cap_shunt_p a_9540_9538# vdd pmos_6p0 w=1.2u l=0.5u
X2099 vss cap_shunt_n a_13776_42104# vss nmos_6p0 w=0.82u l=0.6u
X2100 a_2140_30600# a_2052_30644# vss vss nmos_6p0 w=0.82u l=1u
X2101 a_32404_25564# cap_shunt_p a_32612_25218# vdd pmos_6p0 w=1.2u l=0.5u
X2102 a_12580_16532# cap_shunt_p a_12788_17016# vdd pmos_6p0 w=1.2u l=0.5u
X2103 a_2708_20514# cap_shunt_p a_2500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X2104 a_8064_53080# cap_shunt_n a_6740_53080# vss nmos_6p0 w=0.82u l=0.6u
X2105 a_21540_23996# cap_shunt_p a_21748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X2106 vdd tune_shunt[7] a_21540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X2107 vdd a_32156_29032# a_32068_29076# vdd pmos_6p0 w=1.22u l=1u
X2108 vss cap_shunt_p a_25984_39268# vss nmos_6p0 w=0.82u l=0.6u
X2109 a_10452_30268# cap_shunt_n a_10660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X2110 a_22680_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2111 a_12992_43672# cap_shunt_n a_11668_43672# vss nmos_6p0 w=0.82u l=0.6u
X2112 a_9196_55255# a_9108_55352# vss vss nmos_6p0 w=0.82u l=1u
X2113 vdd tune_shunt[7] a_28484_29076# vdd pmos_6p0 w=1.2u l=0.5u
X2114 a_36688_24856# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X2115 a_27676_8215# a_27588_8312# vss vss nmos_6p0 w=0.82u l=1u
X2116 vdd tune_shunt[5] a_13588_49084# vdd pmos_6p0 w=1.2u l=0.5u
X2117 a_7748_29922# cap_shunt_n a_7540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X2118 a_33500_52552# a_33412_52596# vss vss nmos_6p0 w=0.82u l=1u
X2119 vdd a_31708_41143# a_31620_41240# vdd pmos_6p0 w=1.22u l=1u
X2120 a_12992_40536# cap_shunt_n a_11668_40536# vss nmos_6p0 w=0.82u l=0.6u
X2121 a_13796_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2122 vdd tune_series_gy[5] a_19524_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2123 vdd a_16252_49416# a_16164_49460# vdd pmos_6p0 w=1.22u l=1u
X2124 a_7748_36194# cap_shunt_n a_7540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X2125 a_14692_10744# cap_series_gyn a_14484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X2126 a_24652_55255# a_24564_55352# vss vss nmos_6p0 w=0.82u l=1u
X2127 a_2500_27132# cap_shunt_p a_2708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X2128 a_16500_42812# cap_shunt_n a_16708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X2129 a_11800_7124# cap_series_gyp a_12608_7608# vss nmos_6p0 w=0.82u l=0.6u
X2130 a_34516_20514# cap_series_gygyp a_35448_20452# vss nmos_6p0 w=0.82u l=0.6u
X2131 a_28692_13880# cap_series_gyp a_28484_13396# vdd pmos_6p0 w=1.2u l=0.5u
X2132 a_15120_18884# cap_shunt_p a_13796_18946# vss nmos_6p0 w=0.82u l=0.6u
X2133 a_3484_52119# a_3396_52216# vss vss nmos_6p0 w=0.82u l=1u
X2134 a_29492_38108# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2135 a_35880_11828# cap_series_gygyp a_35904_12312# vss nmos_6p0 w=0.82u l=0.6u
X2136 a_7748_33058# cap_shunt_n a_7540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X2137 a_25572_27508# cap_shunt_p a_25780_27992# vdd pmos_6p0 w=1.2u l=0.5u
X2138 a_28692_10744# cap_series_gyp a_28484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X2139 vdd tune_shunt[6] a_14372_40052# vdd pmos_6p0 w=1.2u l=0.5u
X2140 a_7748_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2141 vss tune_series_gy[5] a_18612_7970# vss nmos_6p0 w=0.51u l=0.6u
X2142 a_3828_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2143 vdd tune_shunt[5] a_28484_38484# vdd pmos_6p0 w=1.2u l=0.5u
X2144 a_15120_15748# cap_shunt_p a_13796_15810# vss nmos_6p0 w=0.82u l=0.6u
X2145 vss tune_shunt[6] a_14580_46808# vss nmos_6p0 w=0.51u l=0.6u
X2146 a_20532_46324# cap_shunt_p a_20740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X2147 a_12788_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2148 a_23308_46280# a_23220_46324# vss vss nmos_6p0 w=0.82u l=1u
X2149 a_24660_44034# cap_shunt_p a_24452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X2150 vdd a_37420_31735# a_37332_31832# vdd pmos_6p0 w=1.22u l=1u
X2151 vdd a_15356_18056# a_15268_18100# vdd pmos_6p0 w=1.22u l=1u
X2152 a_16708_20514# cap_shunt_p a_16500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X2153 vss tune_series_gygy[0] a_31624_6748# vss nmos_6p0 w=0.51u l=0.6u
X2154 a_17828_17016# cap_shunt_p a_19544_17016# vss nmos_6p0 w=0.82u l=0.6u
X2155 a_15804_18056# a_15716_18100# vss vss nmos_6p0 w=0.82u l=1u
X2156 a_20740_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2157 a_13252_24372# cap_shunt_n a_13460_24856# vdd pmos_6p0 w=1.2u l=0.5u
X2158 a_27888_17016# cap_series_gyp a_25780_17016# vss nmos_6p0 w=0.82u l=0.6u
X2159 a_28692_17016# cap_series_gyn a_28484_16532# vdd pmos_6p0 w=1.2u l=0.5u
X2160 a_33732_29560# cap_shunt_p a_33524_29076# vdd pmos_6p0 w=1.2u l=0.5u
X2161 a_3620_24372# cap_shunt_p a_3828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X2162 vss tune_series_gy[4] a_18612_4834# vss nmos_6p0 w=0.51u l=0.6u
X2163 vss cap_shunt_p a_15120_14180# vss nmos_6p0 w=0.82u l=0.6u
X2164 a_3828_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2165 vdd tune_shunt[6] a_28484_35348# vdd pmos_6p0 w=1.2u l=0.5u
X2166 a_29692_21192# a_29604_21236# vss vss nmos_6p0 w=0.82u l=1u
X2167 a_17708_50551# a_17620_50648# vss vss nmos_6p0 w=0.82u l=1u
X2168 a_5544_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2169 a_24660_40898# cap_shunt_n a_24452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X2170 a_2500_36540# cap_shunt_n a_2708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X2171 vdd a_36748_35304# a_36660_35348# vdd pmos_6p0 w=1.22u l=1u
X2172 vss cap_shunt_p a_9072_23588# vss nmos_6p0 w=0.82u l=0.6u
X2173 a_30028_44712# a_29940_44756# vss vss nmos_6p0 w=0.82u l=1u
X2174 vss cap_shunt_n a_15904_32996# vss nmos_6p0 w=0.82u l=0.6u
X2175 a_15804_14920# a_15716_14964# vss vss nmos_6p0 w=0.82u l=1u
X2176 a_19152_46808# cap_shunt_n a_17828_46808# vss nmos_6p0 w=0.82u l=0.6u
X2177 vdd a_6060_8215# a_5972_8312# vdd pmos_6p0 w=1.22u l=1u
X2178 a_13252_21236# cap_shunt_n a_13460_21720# vdd pmos_6p0 w=1.2u l=0.5u
X2179 a_19732_9176# cap_series_gyp a_21448_9176# vss nmos_6p0 w=0.82u l=0.6u
X2180 a_33024_47108# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2181 a_3620_21236# cap_shunt_p a_3828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X2182 vdd tune_shunt[3] a_2724_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2183 a_28124_23895# a_28036_23992# vss vss nmos_6p0 w=0.82u l=1u
X2184 a_2500_33404# cap_shunt_p a_2708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X2185 a_28484_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2186 a_25572_13396# cap_series_gyn a_25780_13880# vdd pmos_6p0 w=1.2u l=0.5u
X2187 a_19732_9176# cap_series_gyp a_19524_8692# vdd pmos_6p0 w=1.2u l=0.5u
X2188 a_3932_53687# a_3844_53784# vss vss nmos_6p0 w=0.82u l=1u
X2189 vdd tune_shunt[7] a_21540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X2190 a_16500_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2191 a_9540_15810# cap_shunt_p a_9332_16156# vdd pmos_6p0 w=1.2u l=0.5u
X2192 a_13252_33780# cap_shunt_n a_13460_34264# vdd pmos_6p0 w=1.2u l=0.5u
X2193 a_3172_16532# cap_shunt_p a_3380_17016# vdd pmos_6p0 w=1.2u l=0.5u
X2194 a_17828_46808# cap_shunt_n a_17620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X2195 a_2708_11106# cap_shunt_n a_2500_11452# vdd pmos_6p0 w=1.2u l=0.5u
X2196 a_36688_18584# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X2197 a_21540_14588# cap_series_gyn a_21748_14242# vdd pmos_6p0 w=1.2u l=0.5u
X2198 a_13252_30644# cap_shunt_n a_13460_31128# vdd pmos_6p0 w=1.2u l=0.5u
X2199 a_8848_32696# cap_shunt_n a_6740_32696# vss nmos_6p0 w=0.82u l=0.6u
X2200 a_6852_53442# cap_shunt_n a_7784_53380# vss nmos_6p0 w=0.82u l=0.6u
X2201 a_9668_49460# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2202 a_14580_45240# cap_shunt_p a_14372_44756# vdd pmos_6p0 w=1.2u l=0.5u
X2203 a_36688_15448# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X2204 a_24652_48983# a_24564_49080# vss vss nmos_6p0 w=0.82u l=1u
X2205 a_28484_33780# cap_shunt_p a_28692_34264# vdd pmos_6p0 w=1.2u l=0.5u
X2206 a_1716_5556# cap_shunt_p a_1924_6040# vdd pmos_6p0 w=1.2u l=0.5u
X2207 a_10092_3944# a_10004_3988# vss vss nmos_6p0 w=0.82u l=1u
X2208 a_21748_45602# cap_shunt_p a_21540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X2209 a_16500_36540# cap_shunt_n a_16708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X2210 a_13460_35832# cap_shunt_n a_14392_35832# vss nmos_6p0 w=0.82u l=0.6u
X2211 a_21748_12674# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2212 vdd a_32156_55255# a_32068_55352# vdd pmos_6p0 w=1.22u l=1u
X2213 a_7748_26786# cap_shunt_n a_7540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X2214 a_35292_22760# a_35204_22804# vss vss nmos_6p0 w=0.82u l=1u
X2215 a_33164_12919# a_33076_13016# vss vss nmos_6p0 w=0.82u l=1u
X2216 a_26444_50984# a_26356_51028# vss vss nmos_6p0 w=0.82u l=1u
X2217 a_34412_47108# cap_shunt_gyp a_34144_47108# vss nmos_6p0 w=0.82u l=0.6u
X2218 a_32612_28354# cap_shunt_p a_32404_28700# vdd pmos_6p0 w=1.2u l=0.5u
X2219 a_28484_30644# cap_shunt_n a_28692_31128# vdd pmos_6p0 w=1.2u l=0.5u
X2220 a_1692_21192# a_1604_21236# vss vss nmos_6p0 w=0.82u l=1u
X2221 a_25780_27992# cap_shunt_p a_26712_27992# vss nmos_6p0 w=0.82u l=0.6u
X2222 vdd tune_shunt[7] a_7540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X2223 vss tune_shunt[5] a_6292_15810# vss nmos_6p0 w=0.51u l=0.6u
X2224 a_16500_33404# cap_shunt_n a_16708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X2225 a_35056_27992# cap_shunt_p a_33732_27992# vss nmos_6p0 w=0.82u l=0.6u
X2226 vss cap_shunt_gyn a_34412_45540# vss nmos_6p0 w=0.82u l=0.6u
X2227 a_35180_33303# a_35092_33400# vss vss nmos_6p0 w=0.82u l=1u
X2228 vdd a_32156_52119# a_32068_52216# vdd pmos_6p0 w=1.22u l=1u
X2229 vss tune_shunt[7] a_16708_18946# vss nmos_6p0 w=0.51u l=0.6u
X2230 vdd a_37420_25463# a_37332_25560# vdd pmos_6p0 w=1.22u l=1u
X2231 a_18424_47108# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2232 a_10680_8316# cap_series_gyp a_11488_7908# vss nmos_6p0 w=0.82u l=0.6u
X2233 a_21540_44380# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2234 vdd a_2140_36872# a_2052_36916# vdd pmos_6p0 w=1.22u l=1u
X2235 a_25780_24856# cap_shunt_p a_26712_24856# vss nmos_6p0 w=0.82u l=0.6u
X2236 a_22644_7608# cap_series_gyp a_22436_7124# vdd pmos_6p0 w=1.2u l=0.5u
X2237 vdd tune_shunt[7] a_28484_29076# vdd pmos_6p0 w=1.2u l=0.5u
X2238 vdd tune_shunt[3] a_5636_10260# vdd pmos_6p0 w=1.2u l=0.5u
X2239 a_9316_50306# cap_shunt_p a_9108_50652# vdd pmos_6p0 w=1.2u l=0.5u
X2240 vss cap_shunt_gyn a_34412_42404# vss nmos_6p0 w=0.82u l=0.6u
X2241 a_20740_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2242 a_3828_34264# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2243 vdd a_36748_29032# a_36660_29076# vdd pmos_6p0 w=1.22u l=1u
X2244 a_3828_21720# cap_shunt_p a_5544_21720# vss nmos_6p0 w=0.82u l=0.6u
X2245 vdd a_37420_22327# a_37332_22424# vdd pmos_6p0 w=1.22u l=1u
X2246 a_24452_9884# cap_series_gyn a_24660_9538# vdd pmos_6p0 w=1.2u l=0.5u
X2247 vdd a_5276_54120# a_5188_54164# vdd pmos_6p0 w=1.22u l=1u
X2248 a_20740_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2249 a_27888_4472# cap_shunt_p a_25780_4472# vss nmos_6p0 w=0.82u l=0.6u
X2250 vss cap_series_gyn a_23968_13880# vss nmos_6p0 w=0.82u l=0.6u
X2251 a_21540_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2252 a_12656_27992# cap_shunt_n a_10548_27992# vss nmos_6p0 w=0.82u l=0.6u
X2253 a_3828_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2254 a_9220_19292# cap_shunt_p a_9428_18946# vdd pmos_6p0 w=1.2u l=0.5u
X2255 a_17620_36916# cap_shunt_n a_17828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X2256 a_2500_27132# cap_shunt_p a_2708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X2257 vss cap_shunt_n a_15904_23588# vss nmos_6p0 w=0.82u l=0.6u
X2258 vdd a_34844_14920# a_34756_14964# vdd pmos_6p0 w=1.22u l=1u
X2259 a_32612_29922# cap_shunt_p a_32404_30268# vdd pmos_6p0 w=1.2u l=0.5u
X2260 a_24452_6748# cap_series_gyn a_24660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X2261 vss cap_series_gyp a_23968_10744# vss nmos_6p0 w=0.82u l=0.6u
X2262 a_37280_51574# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2263 a_12656_24856# cap_shunt_n a_10548_24856# vss nmos_6p0 w=0.82u l=0.6u
X2264 a_18492_11784# a_18404_11828# vss vss nmos_6p0 w=0.82u l=1u
X2265 vdd a_33500_55688# a_33412_55732# vdd pmos_6p0 w=1.22u l=1u
X2266 vdd a_20732_54120# a_20644_54164# vdd pmos_6p0 w=1.22u l=1u
X2267 a_10660_45602# cap_shunt_n a_11592_45540# vss nmos_6p0 w=0.82u l=0.6u
X2268 a_18612_9538# cap_series_gyp a_20328_9476# vss nmos_6p0 w=0.82u l=0.6u
X2269 a_19936_20152# cap_shunt_p a_17828_20152# vss nmos_6p0 w=0.82u l=0.6u
X2270 vdd a_34844_11784# a_34756_11828# vdd pmos_6p0 w=1.22u l=1u
X2271 a_32612_37762# cap_shunt_p a_33544_37700# vss nmos_6p0 w=0.82u l=0.6u
X2272 a_5636_9884# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2273 a_25780_38968# cap_shunt_p a_25572_38484# vdd pmos_6p0 w=1.2u l=0.5u
X2274 a_17828_15448# cap_shunt_p a_17620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2275 a_24660_44034# cap_shunt_p a_24452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X2276 a_16500_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2277 vdd a_20732_50984# a_20644_51028# vdd pmos_6p0 w=1.22u l=1u
X2278 a_10660_42466# cap_shunt_n a_11592_42404# vss nmos_6p0 w=0.82u l=0.6u
X2279 a_7768_6748# cap_series_gyp a_7792_6340# vss nmos_6p0 w=0.82u l=0.6u
X2280 a_13252_24372# cap_shunt_n a_13460_24856# vdd pmos_6p0 w=1.2u l=0.5u
X2281 a_31708_47415# a_31620_47512# vss vss nmos_6p0 w=0.82u l=1u
X2282 a_15176_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2283 vdd a_20284_49416# a_20196_49460# vdd pmos_6p0 w=1.22u l=1u
X2284 vdd a_27676_33303# a_27588_33400# vdd pmos_6p0 w=1.22u l=1u
X2285 a_25780_35832# cap_shunt_p a_25572_35348# vdd pmos_6p0 w=1.2u l=0.5u
X2286 vdd tune_shunt[7] a_9220_20860# vdd pmos_6p0 w=1.2u l=0.5u
X2287 a_32404_34972# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2288 a_11200_20152# cap_shunt_p a_9876_20152# vss nmos_6p0 w=0.82u l=0.6u
X2289 a_24660_40898# cap_shunt_n a_24452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X2290 a_21748_39330# cap_shunt_p a_21540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X2291 a_33164_9783# a_33076_9880# vss vss nmos_6p0 w=0.82u l=1u
X2292 a_12332_47415# a_12244_47512# vss vss nmos_6p0 w=0.82u l=1u
X2293 a_13796_45602# cap_shunt_p a_13588_45948# vdd pmos_6p0 w=1.2u l=0.5u
X2294 a_13460_29560# cap_shunt_n a_14392_29560# vss nmos_6p0 w=0.82u l=0.6u
X2295 a_8848_23288# cap_shunt_p a_6740_23288# vss nmos_6p0 w=0.82u l=0.6u
X2296 a_16708_20514# cap_shunt_p a_17640_20452# vss nmos_6p0 w=0.82u l=0.6u
X2297 a_13252_21236# cap_shunt_n a_13460_21720# vdd pmos_6p0 w=1.2u l=0.5u
X2298 vdd a_37868_53687# a_37780_53784# vdd pmos_6p0 w=1.22u l=1u
X2299 vdd a_32156_48983# a_32068_49080# vdd pmos_6p0 w=1.22u l=1u
X2300 a_6292_17378# cap_shunt_p a_6084_17724# vdd pmos_6p0 w=1.2u l=0.5u
X2301 a_6060_55688# a_5972_55732# vss vss nmos_6p0 w=0.82u l=1u
X2302 a_26444_44712# a_26356_44756# vss vss nmos_6p0 w=0.82u l=1u
X2303 a_32404_31836# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2304 a_28484_24372# cap_shunt_p a_28692_24856# vdd pmos_6p0 w=1.2u l=0.5u
X2305 vss tune_shunt_gy[1] a_36288_39672# vss nmos_6p0 w=0.51u l=0.6u
X2306 a_25572_13396# cap_series_gyn a_25780_13880# vdd pmos_6p0 w=1.2u l=0.5u
X2307 a_16500_27132# cap_shunt_n a_16708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X2308 vdd a_18492_53687# a_18404_53784# vdd pmos_6p0 w=1.22u l=1u
X2309 a_13564_53687# a_13476_53784# vss vss nmos_6p0 w=0.82u l=1u
X2310 a_13460_26424# cap_shunt_n a_14392_26424# vss nmos_6p0 w=0.82u l=0.6u
X2311 a_1716_5180# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2312 a_1924_7970# cap_shunt_n a_1716_8316# vdd pmos_6p0 w=1.2u l=0.5u
X2313 vss cap_shunt_p a_4816_22020# vss nmos_6p0 w=0.82u l=0.6u
X2314 a_11572_5556# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2315 a_31808_29860# cap_shunt_p a_29700_29922# vss nmos_6p0 w=0.82u l=0.6u
X2316 a_21748_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2317 vdd tune_series_gygy[5] a_35692_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2318 a_3036_55688# a_2948_55732# vss vss nmos_6p0 w=0.82u l=1u
X2319 vss cap_shunt_n a_4032_7608# vss nmos_6p0 w=0.82u l=0.6u
X2320 a_1692_11784# a_1604_11828# vss vss nmos_6p0 w=0.82u l=1u
X2321 vdd tune_series_gy[5] a_24452_17724# vdd pmos_6p0 w=1.2u l=0.5u
X2322 a_25780_18584# cap_series_gyn a_26712_18584# vss nmos_6p0 w=0.82u l=0.6u
X2323 a_31808_26724# cap_shunt_p a_29700_26786# vss nmos_6p0 w=0.82u l=0.6u
X2324 vdd a_37420_16055# a_37332_16152# vdd pmos_6p0 w=1.22u l=1u
X2325 vdd tune_series_gygy[5] a_35692_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2326 a_12712_6040# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2327 vdd tune_shunt[3] a_32404_38108# vdd pmos_6p0 w=1.2u l=0.5u
X2328 vdd a_2140_27464# a_2052_27508# vdd pmos_6p0 w=1.22u l=1u
X2329 a_25780_15448# cap_series_gyp a_26712_15448# vss nmos_6p0 w=0.82u l=0.6u
X2330 a_14580_45240# cap_shunt_p a_14372_44756# vdd pmos_6p0 w=1.2u l=0.5u
X2331 a_6532_40052# cap_shunt_n a_6740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X2332 vdd a_24652_5512# a_24564_5556# vdd pmos_6p0 w=1.22u l=1u
X2333 a_6572_5556# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2334 a_23308_52119# a_23220_52216# vss vss nmos_6p0 w=0.82u l=1u
X2335 a_28484_33780# cap_shunt_p a_28692_34264# vdd pmos_6p0 w=1.2u l=0.5u
X2336 vdd a_37420_12919# a_37332_13016# vdd pmos_6p0 w=1.22u l=1u
X2337 a_3828_48376# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2338 a_34308_13020# cap_series_gygyp a_34516_12674# vdd pmos_6p0 w=1.2u l=0.5u
X2339 a_21540_5180# cap_series_gyp a_21748_4834# vdd pmos_6p0 w=1.2u l=0.5u
X2340 vdd a_33500_49416# a_33412_49460# vdd pmos_6p0 w=1.22u l=1u
X2341 a_28484_30644# cap_shunt_n a_28692_31128# vdd pmos_6p0 w=1.2u l=0.5u
X2342 a_17620_27508# cap_shunt_n a_17828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X2343 a_26768_4772# cap_series_gyp a_24660_4834# vss nmos_6p0 w=0.82u l=0.6u
X2344 a_17640_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2345 a_10988_54120# a_10900_54164# vss vss nmos_6p0 w=0.82u l=1u
X2346 vdd tune_series_gygy[3] a_35692_7124# vdd pmos_6p0 w=1.2u l=0.5u
X2347 a_36188_54120# a_36100_54164# vss vss nmos_6p0 w=0.82u l=1u
X2348 vss cap_shunt_p a_23072_22020# vss nmos_6p0 w=0.82u l=0.6u
X2349 vdd a_1692_53687# a_1604_53784# vdd pmos_6p0 w=1.22u l=1u
X2350 vss cap_shunt_p a_19936_48376# vss nmos_6p0 w=0.82u l=0.6u
X2351 a_10660_36194# cap_shunt_n a_11592_36132# vss nmos_6p0 w=0.82u l=0.6u
X2352 vdd a_20172_23895# a_20084_23992# vdd pmos_6p0 w=1.22u l=1u
X2353 a_36720_47893# cap_shunt_gyp a_36720_48438# vdd pmos_6p0 w=1.215u l=0.5u
X2354 vdd a_33500_46280# a_33412_46324# vdd pmos_6p0 w=1.22u l=1u
X2355 a_12788_18584# cap_shunt_p a_12580_18100# vdd pmos_6p0 w=1.2u l=0.5u
X2356 a_25780_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2357 a_2932_10744# cap_shunt_n a_2724_10260# vdd pmos_6p0 w=1.2u l=0.5u
X2358 a_3828_13880# cap_shunt_n a_3620_13396# vdd pmos_6p0 w=1.2u l=0.5u
X2359 a_17640_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2360 vdd a_25996_47848# a_25908_47892# vdd pmos_6p0 w=1.22u l=1u
X2361 a_25780_29560# cap_shunt_p a_25572_29076# vdd pmos_6p0 w=1.2u l=0.5u
X2362 vdd a_25548_55255# a_25460_55352# vdd pmos_6p0 w=1.22u l=1u
X2363 a_19836_50984# a_19748_51028# vss vss nmos_6p0 w=0.82u l=1u
X2364 vdd a_1692_50551# a_1604_50648# vdd pmos_6p0 w=1.22u l=1u
X2365 a_18612_4834# cap_series_gyp a_18404_5180# vdd pmos_6p0 w=1.2u l=0.5u
X2366 a_10680_8316# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X2367 vdd a_20172_20759# a_20084_20856# vdd pmos_6p0 w=1.22u l=1u
X2368 a_3828_42104# cap_shunt_p a_3620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X2369 a_13796_39330# cap_shunt_n a_13588_39676# vdd pmos_6p0 w=1.2u l=0.5u
X2370 vdd a_32604_18056# a_32516_18100# vdd pmos_6p0 w=1.22u l=1u
X2371 vdd tune_shunt[6] a_6532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X2372 a_16708_14242# cap_shunt_p a_17640_14180# vss nmos_6p0 w=0.82u l=0.6u
X2373 a_8064_38968# cap_shunt_n a_6740_38968# vss nmos_6p0 w=0.82u l=0.6u
X2374 a_28572_33303# a_28484_33400# vss vss nmos_6p0 w=0.82u l=1u
X2375 vdd a_25996_44712# a_25908_44756# vdd pmos_6p0 w=1.22u l=1u
X2376 vdd a_16028_32168# a_15940_32212# vdd pmos_6p0 w=1.22u l=1u
X2377 vdd a_25548_52119# a_25460_52216# vdd pmos_6p0 w=1.22u l=1u
X2378 a_30476_50984# a_30388_51028# vss vss nmos_6p0 w=0.82u l=1u
X2379 a_32404_25564# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2380 a_36296_21720# cap_series_gygyp a_35880_21236# vss nmos_6p0 w=0.82u l=0.6u
X2381 vdd a_18044_52552# a_17956_52596# vdd pmos_6p0 w=1.22u l=1u
X2382 vdd tune_shunt[7] a_13252_36916# vdd pmos_6p0 w=1.2u l=0.5u
X2383 a_32612_29922# cap_shunt_p a_32404_30268# vdd pmos_6p0 w=1.2u l=0.5u
X2384 a_37652_45540# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2385 vdd tune_shunt[6] a_3620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X2386 a_33500_38440# a_33412_38484# vss vss nmos_6p0 w=0.82u l=1u
X2387 a_23576_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X2388 a_22644_7608# cap_series_gyp a_22436_7124# vdd pmos_6p0 w=1.2u l=0.5u
X2389 a_7540_44380# cap_shunt_p a_7748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X2390 a_11668_40536# cap_shunt_n a_11460_40052# vdd pmos_6p0 w=1.2u l=0.5u
X2391 a_16028_27464# a_15940_27508# vss vss nmos_6p0 w=0.82u l=1u
X2392 a_20740_26424# cap_shunt_n a_20532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2393 a_37652_42404# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2394 a_25780_38968# cap_shunt_p a_25572_38484# vdd pmos_6p0 w=1.2u l=0.5u
X2395 vdd a_28348_21192# a_28260_21236# vdd pmos_6p0 w=1.22u l=1u
X2396 a_4424_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2397 vss tune_shunt[5] a_6740_53080# vss nmos_6p0 w=0.51u l=0.6u
X2398 vdd a_37868_5079# a_37780_5176# vdd pmos_6p0 w=1.22u l=1u
X2399 vdd tune_series_gygy[5] a_35692_16532# vdd pmos_6p0 w=1.2u l=0.5u
X2400 a_21748_17378# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2401 a_7540_41244# cap_shunt_n a_7748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X2402 a_16028_24328# a_15940_24372# vss vss nmos_6p0 w=0.82u l=1u
X2403 a_20740_23288# cap_shunt_p a_20532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2404 a_14692_9176# cap_series_gyn a_14484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X2405 a_16500_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2406 a_25780_35832# cap_shunt_p a_25572_35348# vdd pmos_6p0 w=1.2u l=0.5u
X2407 vdd tune_shunt[7] a_9220_20860# vdd pmos_6p0 w=1.2u l=0.5u
X2408 a_31808_17316# cap_series_gyp a_29700_17378# vss nmos_6p0 w=0.82u l=0.6u
X2409 a_15512_50244# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2410 a_4424_42404# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2411 vss tune_shunt[6] a_10548_38968# vss nmos_6p0 w=0.51u l=0.6u
X2412 vdd a_4492_3944# a_4404_3988# vdd pmos_6p0 w=1.22u l=1u
X2413 a_14468_3266# cap_series_gyn a_15400_3204# vss nmos_6p0 w=0.82u l=0.6u
X2414 a_13460_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2415 vss cap_shunt_p a_4704_49944# vss nmos_6p0 w=0.82u l=0.6u
X2416 a_13796_45602# cap_shunt_p a_13588_45948# vdd pmos_6p0 w=1.2u l=0.5u
X2417 a_6292_17378# cap_shunt_p a_6084_17724# vdd pmos_6p0 w=1.2u l=0.5u
X2418 a_5844_9176# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X2419 a_11592_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2420 a_14692_6040# cap_series_gyn a_14484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X2421 a_30924_52552# a_30836_52596# vss vss nmos_6p0 w=0.82u l=1u
X2422 a_12376_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2423 vss tune_shunt[7] a_13796_37762# vss nmos_6p0 w=0.51u l=0.6u
X2424 a_28484_24372# cap_shunt_p a_28692_24856# vdd pmos_6p0 w=1.2u l=0.5u
X2425 a_35292_3944# a_35204_3988# vss vss nmos_6p0 w=0.82u l=1u
X2426 a_25780_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2427 a_5152_35832# cap_shunt_n a_3828_35832# vss nmos_6p0 w=0.82u l=0.6u
X2428 a_25572_13396# cap_series_gyn a_25780_13880# vdd pmos_6p0 w=1.2u l=0.5u
X2429 a_30408_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2430 a_30688_45944# cap_shunt_gyn a_30708_45540# vss nmos_6p0 w=0.82u l=0.6u
X2431 a_15904_37700# cap_shunt_n a_13796_37762# vss nmos_6p0 w=0.82u l=0.6u
X2432 a_35628_34871# a_35540_34968# vss vss nmos_6p0 w=0.82u l=1u
X2433 a_13588_23996# cap_shunt_n a_13796_23650# vdd pmos_6p0 w=1.2u l=0.5u
X2434 vdd tune_series_gygy[5] a_35692_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2435 a_30632_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2436 vss tune_shunt[7] a_13796_34626# vss nmos_6p0 w=0.51u l=0.6u
X2437 a_25780_10744# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2438 vss tune_shunt[5] a_6292_51874# vss nmos_6p0 w=0.51u l=0.6u
X2439 a_25780_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2440 vdd a_25548_48983# a_25460_49080# vdd pmos_6p0 w=1.22u l=1u
X2441 a_23756_46280# a_23668_46324# vss vss nmos_6p0 w=0.82u l=1u
X2442 vdd a_1692_44279# a_1604_44376# vdd pmos_6p0 w=1.22u l=1u
X2443 vdd a_35292_19624# a_35204_19668# vdd pmos_6p0 w=1.22u l=1u
X2444 a_35628_31735# a_35540_31832# vss vss nmos_6p0 w=0.82u l=1u
X2445 vss cap_shunt_p a_18032_43972# vss nmos_6p0 w=0.82u l=0.6u
X2446 vdd tune_series_gygy[5] a_35692_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2447 vdd a_20172_14487# a_20084_14584# vdd pmos_6p0 w=1.22u l=1u
X2448 vss cap_series_gygyn a_32040_6340# vss nmos_6p0 w=0.82u l=0.6u
X2449 a_26376_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2450 a_25780_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2451 a_30476_44712# a_30388_44756# vss vss nmos_6p0 w=0.82u l=1u
X2452 a_2708_33058# cap_shunt_p a_4424_32996# vss nmos_6p0 w=0.82u l=0.6u
X2453 a_8860_9783# a_8772_9880# vss vss nmos_6p0 w=0.82u l=1u
X2454 a_28484_33780# cap_shunt_p a_28692_34264# vdd pmos_6p0 w=1.2u l=0.5u
X2455 a_19732_9176# cap_series_gyp a_19524_8692# vdd pmos_6p0 w=1.2u l=0.5u
X2456 a_14728_20452# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2457 vss cap_shunt_n a_18032_40836# vss nmos_6p0 w=0.82u l=0.6u
X2458 a_29624_32696# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2459 a_4940_7080# a_4852_7124# vss vss nmos_6p0 w=0.82u l=1u
X2460 vdd a_29244_43144# a_29156_43188# vdd pmos_6p0 w=1.22u l=1u
X2461 a_3828_32696# cap_shunt_p a_3620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X2462 vdd tune_shunt[7] a_6532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X2463 a_34308_13020# cap_series_gygyp a_34516_12674# vdd pmos_6p0 w=1.2u l=0.5u
X2464 a_26376_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2465 a_28572_23895# a_28484_23992# vss vss nmos_6p0 w=0.82u l=1u
X2466 a_36296_12312# cap_series_gygyp a_35880_11828# vss nmos_6p0 w=0.82u l=0.6u
X2467 a_28484_30644# cap_shunt_n a_28692_31128# vdd pmos_6p0 w=1.2u l=0.5u
X2468 vdd a_36076_30167# a_35988_30264# vdd pmos_6p0 w=1.22u l=1u
X2469 vdd tune_shunt[7] a_13252_27508# vdd pmos_6p0 w=1.2u l=0.5u
X2470 vss tune_series_gy[4] a_14692_9176# vss nmos_6p0 w=0.51u l=0.6u
X2471 vdd tune_shunt[7] a_16500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X2472 a_30364_52119# a_30276_52216# vss vss nmos_6p0 w=0.82u l=1u
X2473 vdd tune_shunt[7] a_3620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X2474 a_16708_44034# cap_shunt_p a_16500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X2475 a_36688_7608# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X2476 a_6956_6647# a_6868_6744# vss vss nmos_6p0 w=0.82u l=1u
X2477 vss tune_series_gy[4] a_18612_6402# vss nmos_6p0 w=0.51u l=0.6u
X2478 a_12788_18584# cap_shunt_p a_12580_18100# vdd pmos_6p0 w=1.2u l=0.5u
X2479 a_20740_17016# cap_shunt_p a_20532_16532# vdd pmos_6p0 w=1.2u l=0.5u
X2480 a_16500_36540# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2481 vdd tune_shunt[7] a_16500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X2482 a_25780_29560# cap_shunt_p a_25572_29076# vdd pmos_6p0 w=1.2u l=0.5u
X2483 a_9876_15448# cap_shunt_p a_9668_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2484 vdd a_31708_40008# a_31620_40052# vdd pmos_6p0 w=1.22u l=1u
X2485 vdd tune_shunt[7] a_12580_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2486 a_4424_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2487 a_16708_40898# cap_shunt_n a_16500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X2488 vdd a_3036_14920# a_2948_14964# vdd pmos_6p0 w=1.22u l=1u
X2489 a_20532_43188# cap_shunt_n a_20740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X2490 a_13796_39330# cap_shunt_n a_13588_39676# vdd pmos_6p0 w=1.2u l=0.5u
X2491 vdd tune_shunt[5] a_9668_51028# vdd pmos_6p0 w=1.2u l=0.5u
X2492 a_2500_47516# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2493 a_25780_34264# cap_shunt_p a_25572_33780# vdd pmos_6p0 w=1.2u l=0.5u
X2494 a_16500_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2495 a_14692_4472# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X2496 vdd tune_shunt[7] a_12580_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2497 a_9876_12312# cap_shunt_p a_9668_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2498 a_5152_29560# cap_shunt_n a_3828_29560# vss nmos_6p0 w=0.82u l=0.6u
X2499 vdd tune_series_gy[5] a_21540_13020# vdd pmos_6p0 w=1.2u l=0.5u
X2500 vss cap_series_gyp a_7176_7608# vss nmos_6p0 w=0.82u l=0.6u
X2501 a_9316_50306# cap_shunt_p a_10248_50244# vss nmos_6p0 w=0.82u l=0.6u
X2502 vss tune_shunt[7] a_12788_12312# vss nmos_6p0 w=0.51u l=0.6u
X2503 a_26892_50984# a_26804_51028# vss vss nmos_6p0 w=0.82u l=1u
X2504 a_33732_34264# cap_shunt_n a_35448_34264# vss nmos_6p0 w=0.82u l=0.6u
X2505 a_25780_31128# cap_shunt_p a_25572_30644# vdd pmos_6p0 w=1.2u l=0.5u
X2506 a_35628_28599# a_35540_28696# vss vss nmos_6p0 w=0.82u l=1u
X2507 vdd a_2140_47415# a_2052_47512# vdd pmos_6p0 w=1.22u l=1u
X2508 vss tune_shunt[7] a_13796_28354# vss nmos_6p0 w=0.51u l=0.6u
X2509 a_3620_25940# cap_shunt_p a_3828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X2510 a_3620_47892# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2511 a_5152_26424# cap_shunt_p a_3828_26424# vss nmos_6p0 w=0.82u l=0.6u
X2512 vdd tune_shunt[6] a_6196_47516# vdd pmos_6p0 w=1.2u l=0.5u
X2513 a_13796_20514# cap_shunt_n a_15512_20452# vss nmos_6p0 w=0.82u l=0.6u
X2514 vdd a_35740_53687# a_35652_53784# vdd pmos_6p0 w=1.22u l=1u
X2515 a_31708_32168# a_31620_32212# vss vss nmos_6p0 w=0.82u l=1u
X2516 a_33732_31128# cap_shunt_n a_35448_31128# vss nmos_6p0 w=0.82u l=0.6u
X2517 vdd tune_shunt[3] a_2724_8692# vdd pmos_6p0 w=1.2u l=0.5u
X2518 a_30812_53687# a_30724_53784# vss vss nmos_6p0 w=0.82u l=1u
X2519 vss tune_shunt[7] a_33732_27992# vss nmos_6p0 w=0.51u l=0.6u
X2520 a_13588_14588# cap_shunt_p a_13796_14242# vdd pmos_6p0 w=1.2u l=0.5u
X2521 a_23856_20452# cap_shunt_p a_21748_20514# vss nmos_6p0 w=0.82u l=0.6u
X2522 a_23868_50984# a_23780_51028# vss vss nmos_6p0 w=0.82u l=1u
X2523 a_2588_36872# a_2500_36916# vss vss nmos_6p0 w=0.82u l=1u
X2524 a_35628_25463# a_35540_25560# vss vss nmos_6p0 w=0.82u l=1u
X2525 vss tune_shunt[7] a_13796_25218# vss nmos_6p0 w=0.51u l=0.6u
X2526 a_3620_22804# cap_shunt_p a_3828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X2527 vdd tune_series_gygy[5] a_35692_16532# vdd pmos_6p0 w=1.2u l=0.5u
X2528 a_3620_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2529 a_10472_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2530 a_7224_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2531 a_25444_3266# cap_shunt_p a_25236_3612# vdd pmos_6p0 w=1.2u l=0.5u
X2532 vdd a_35740_50551# a_35652_50648# vdd pmos_6p0 w=1.22u l=1u
X2533 vss cap_shunt_p a_5936_43672# vss nmos_6p0 w=0.82u l=0.6u
X2534 a_31624_6748# cap_series_gygyn a_31436_6748# vdd pmos_6p0 w=1.2u l=0.5u
X2535 a_8176_53380# cap_shunt_n a_6852_53442# vss nmos_6p0 w=0.82u l=0.6u
X2536 a_30812_50551# a_30724_50648# vss vss nmos_6p0 w=0.82u l=1u
X2537 vdd tune_shunt[5] a_20532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X2538 a_14504_49944# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2539 a_14728_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2540 vss cap_shunt_n a_18032_34564# vss nmos_6p0 w=0.82u l=0.6u
X2541 vdd a_22076_52552# a_21988_52596# vdd pmos_6p0 w=1.22u l=1u
X2542 a_19724_45847# a_19636_45944# vss vss nmos_6p0 w=0.82u l=1u
X2543 a_26376_34564# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2544 vdd tune_series_gygy[5] a_34308_22428# vdd pmos_6p0 w=1.2u l=0.5u
X2545 a_1924_6402# cap_shunt_n a_1716_6748# vdd pmos_6p0 w=1.2u l=0.5u
X2546 a_25780_17016# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2547 a_6292_17378# cap_shunt_p a_6084_17724# vdd pmos_6p0 w=1.2u l=0.5u
X2548 a_13796_48738# cap_shunt_n a_14728_48676# vss nmos_6p0 w=0.82u l=0.6u
X2549 vss tune_shunt[5] a_21748_42466# vss nmos_6p0 w=0.51u l=0.6u
X2550 vss cap_shunt_n a_5936_40536# vss nmos_6p0 w=0.82u l=0.6u
X2551 a_2708_23650# cap_shunt_p a_4424_23588# vss nmos_6p0 w=0.82u l=0.6u
X2552 a_6292_50306# cap_shunt_p a_8008_50244# vss nmos_6p0 w=0.82u l=0.6u
X2553 a_28484_24372# cap_shunt_p a_28692_24856# vdd pmos_6p0 w=1.2u l=0.5u
X2554 vdd a_21516_53687# a_21428_53784# vdd pmos_6p0 w=1.22u l=1u
X2555 a_29624_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2556 vss tune_shunt[7] a_17828_21720# vss nmos_6p0 w=0.51u l=0.6u
X2557 vss cap_shunt_n a_18032_31428# vss nmos_6p0 w=0.82u l=0.6u
X2558 a_37080_24856# cap_series_gygyp a_35880_24372# vss nmos_6p0 w=0.82u l=0.6u
X2559 a_19724_42711# a_19636_42808# vss vss nmos_6p0 w=0.82u l=1u
X2560 a_26376_31428# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2561 a_8456_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2562 a_35692_19668# cap_series_gygyp a_35880_19668# vdd pmos_6p0 w=1.2u l=0.5u
X2563 a_17620_25940# cap_shunt_n a_17828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X2564 a_21056_7608# cap_series_gyp a_19732_7608# vss nmos_6p0 w=0.82u l=0.6u
X2565 a_31024_4772# cap_shunt_p a_29700_4834# vss nmos_6p0 w=0.82u l=0.6u
X2566 a_28484_8692# cap_series_gyn a_28692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X2567 vdd a_10316_53687# a_10228_53784# vdd pmos_6p0 w=1.22u l=1u
X2568 vdd a_21516_50551# a_21428_50648# vdd pmos_6p0 w=1.22u l=1u
X2569 a_22064_37400# cap_shunt_n a_20740_37400# vss nmos_6p0 w=0.82u l=0.6u
X2570 a_33732_34264# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2571 vss tune_shunt[7] a_6740_27992# vss nmos_6p0 w=0.51u l=0.6u
X2572 a_21748_17378# cap_shunt_p a_21540_17724# vdd pmos_6p0 w=1.2u l=0.5u
X2573 a_16708_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2574 vdd tune_shunt[7] a_16500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X2575 a_24660_22082# cap_shunt_p a_25592_22020# vss nmos_6p0 w=0.82u l=0.6u
X2576 a_18404_9884# cap_series_gyp a_18612_9538# vdd pmos_6p0 w=1.2u l=0.5u
X2577 a_30364_42711# a_30276_42808# vss vss nmos_6p0 w=0.82u l=1u
X2578 a_30428_21236# cap_series_gygyn a_30616_21236# vdd pmos_6p0 w=1.2u l=0.5u
X2579 vdd a_30924_55688# a_30836_55732# vdd pmos_6p0 w=1.22u l=1u
X2580 a_3380_18584# cap_shunt_p a_3172_18100# vdd pmos_6p0 w=1.2u l=0.5u
X2581 a_17620_22804# cap_shunt_n a_17828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X2582 vss cap_shunt_n a_4032_6340# vss nmos_6p0 w=0.82u l=0.6u
X2583 a_28484_5556# cap_shunt_n a_28692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X2584 a_2500_13020# cap_shunt_n a_2708_12674# vdd pmos_6p0 w=1.2u l=0.5u
X2585 a_19276_38007# a_19188_38104# vss vss nmos_6p0 w=0.82u l=1u
X2586 a_33732_31128# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2587 vss tune_shunt[7] a_6740_24856# vss nmos_6p0 w=0.51u l=0.6u
X2588 a_25572_7124# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2589 vdd a_36300_32168# a_36212_32212# vdd pmos_6p0 w=1.22u l=1u
X2590 vdd tune_shunt[7] a_16500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X2591 a_11800_7124# cap_series_gyp a_11824_7608# vss nmos_6p0 w=0.82u l=0.6u
X2592 a_18404_6748# cap_series_gyn a_18612_6402# vdd pmos_6p0 w=1.2u l=0.5u
X2593 a_34536_8316# cap_series_gygyp a_34348_8316# vdd pmos_6p0 w=1.2u l=0.5u
X2594 a_16500_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2595 a_15492_8316# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2596 a_12780_47415# a_12692_47512# vss vss nmos_6p0 w=0.82u l=1u
X2597 a_13460_32696# cap_shunt_n a_13252_32212# vdd pmos_6p0 w=1.2u l=0.5u
X2598 a_33500_41143# a_33412_41240# vss vss nmos_6p0 w=0.82u l=1u
X2599 vss cap_shunt_n a_23856_37700# vss nmos_6p0 w=0.82u l=0.6u
X2600 a_17828_21720# cap_shunt_p a_18760_21720# vss nmos_6p0 w=0.82u l=0.6u
X2601 vss cap_shunt_n a_8064_53080# vss nmos_6p0 w=0.82u l=0.6u
X2602 a_14372_46324# cap_shunt_p a_14580_46808# vdd pmos_6p0 w=1.2u l=0.5u
X2603 a_26892_44712# a_26804_44756# vss vss nmos_6p0 w=0.82u l=1u
X2604 vss cap_shunt_n a_4032_3204# vss nmos_6p0 w=0.82u l=0.6u
X2605 a_35880_24372# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2606 a_25780_24856# cap_shunt_p a_25572_24372# vdd pmos_6p0 w=1.2u l=0.5u
X2607 a_5636_11452# cap_shunt_n a_5844_11106# vdd pmos_6p0 w=1.2u l=0.5u
X2608 vss cap_shunt_n a_12992_43672# vss nmos_6p0 w=0.82u l=0.6u
X2609 a_2500_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2610 a_5636_11452# cap_shunt_n a_5844_11106# vdd pmos_6p0 w=1.2u l=0.5u
X2611 a_36300_27464# a_36212_27508# vss vss nmos_6p0 w=0.82u l=1u
X2612 vss tune_shunt[5] a_2708_18946# vss nmos_6p0 w=0.51u l=0.6u
X2613 a_29468_55255# a_29380_55352# vss vss nmos_6p0 w=0.82u l=1u
X2614 vdd tune_shunt[7] a_16500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X2615 a_13796_14242# cap_shunt_p a_15512_14180# vss nmos_6p0 w=0.82u l=0.6u
X2616 a_10452_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2617 a_23856_14180# cap_series_gyn a_21748_14242# vss nmos_6p0 w=0.82u l=0.6u
X2618 a_3484_55688# a_3396_55732# vss vss nmos_6p0 w=0.82u l=1u
X2619 a_13252_38484# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2620 a_24452_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2621 vdd a_20844_47848# a_20756_47892# vdd pmos_6p0 w=1.22u l=1u
X2622 vss cap_shunt_n a_12992_40536# vss nmos_6p0 w=0.82u l=0.6u
X2623 a_6532_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2624 a_25780_21720# cap_shunt_p a_25572_21236# vdd pmos_6p0 w=1.2u l=0.5u
X2625 a_3620_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2626 vdd a_2140_38007# a_2052_38104# vdd pmos_6p0 w=1.22u l=1u
X2627 a_37420_5079# a_37332_5176# vss vss nmos_6p0 w=0.82u l=1u
X2628 vdd a_13564_11351# a_13476_11448# vdd pmos_6p0 w=1.22u l=1u
X2629 vdd tune_series_gygy[5] a_34308_19292# vdd pmos_6p0 w=1.2u l=0.5u
X2630 a_20740_40536# cap_shunt_p a_20532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X2631 a_36188_53687# a_36100_53784# vss vss nmos_6p0 w=0.82u l=1u
X2632 a_3828_43672# cap_shunt_p a_3620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X2633 vdd tune_shunt[7] a_16500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X2634 a_31708_22760# a_31620_22804# vss vss nmos_6p0 w=0.82u l=1u
X2635 a_15120_43972# cap_shunt_n a_13796_44034# vss nmos_6p0 w=0.82u l=0.6u
X2636 vdd tune_shunt[6] a_20532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X2637 a_10452_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2638 a_9876_15448# cap_shunt_p a_9668_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2639 a_13252_35348# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2640 a_23856_11044# cap_series_gyn a_21748_11106# vss nmos_6p0 w=0.82u l=0.6u
X2641 a_36624_12612# cap_series_gygyp a_34516_12674# vss nmos_6p0 w=0.82u l=0.6u
X2642 vdd a_12220_52119# a_12132_52216# vdd pmos_6p0 w=1.22u l=1u
X2643 vss tune_shunt[4] a_21748_45602# vss nmos_6p0 w=0.51u l=0.6u
X2644 a_6740_37400# cap_shunt_n a_8456_37400# vss nmos_6p0 w=0.82u l=0.6u
X2645 vss cap_shunt_n a_18032_28292# vss nmos_6p0 w=0.82u l=0.6u
X2646 a_6620_54120# a_6532_54164# vss vss nmos_6p0 w=0.82u l=1u
X2647 a_17828_45240# cap_shunt_p a_19544_45240# vss nmos_6p0 w=0.82u l=0.6u
X2648 a_3620_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2649 a_2140_19191# a_2052_19288# vss vss nmos_6p0 w=0.82u l=1u
X2650 a_26376_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2651 a_21540_5180# cap_series_gyp a_21748_4834# vdd pmos_6p0 w=1.2u l=0.5u
X2652 vdd tune_series_gy[5] a_15532_11452# vdd pmos_6p0 w=1.2u l=0.5u
X2653 vdd tune_series_gygy[4] a_34308_16156# vdd pmos_6p0 w=1.2u l=0.5u
X2654 a_23756_52119# a_23668_52216# vss vss nmos_6p0 w=0.82u l=1u
X2655 vss cap_shunt_n a_5936_34264# vss nmos_6p0 w=0.82u l=0.6u
X2656 a_25780_34264# cap_shunt_p a_25572_33780# vdd pmos_6p0 w=1.2u l=0.5u
X2657 a_15120_40836# cap_shunt_n a_13796_40898# vss nmos_6p0 w=0.82u l=0.6u
X2658 vss tune_shunt[6] a_21748_36194# vss nmos_6p0 w=0.51u l=0.6u
X2659 vdd tune_shunt[6] a_20532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X2660 a_18612_11106# cap_series_gyn a_18404_11452# vdd pmos_6p0 w=1.2u l=0.5u
X2661 a_9876_12312# cap_shunt_p a_9668_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2662 a_10548_37400# cap_shunt_n a_10340_36916# vdd pmos_6p0 w=1.2u l=0.5u
X2663 a_22456_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2664 vss cap_shunt_n a_18032_25156# vss nmos_6p0 w=0.82u l=0.6u
X2665 a_29468_6647# a_29380_6744# vss vss nmos_6p0 w=0.82u l=1u
X2666 a_17828_42104# cap_shunt_n a_19544_42104# vss nmos_6p0 w=0.82u l=0.6u
X2667 a_2140_16055# a_2052_16152# vss vss nmos_6p0 w=0.82u l=1u
X2668 a_16688_45240# cap_shunt_p a_14580_45240# vss nmos_6p0 w=0.82u l=0.6u
X2669 a_27888_42104# cap_shunt_n a_25780_42104# vss nmos_6p0 w=0.82u l=0.6u
X2670 a_26376_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2671 a_37080_18584# cap_series_gygyn a_35880_18100# vss nmos_6p0 w=0.82u l=0.6u
X2672 a_19724_36439# a_19636_36536# vss vss nmos_6p0 w=0.82u l=1u
X2673 a_5636_8692# cap_shunt_p a_5844_9176# vdd pmos_6p0 w=1.2u l=0.5u
X2674 a_13796_39330# cap_shunt_n a_14728_39268# vss nmos_6p0 w=0.82u l=0.6u
X2675 vss cap_shunt_n a_5936_31128# vss nmos_6p0 w=0.82u l=0.6u
X2676 a_25780_31128# cap_shunt_p a_25572_30644# vdd pmos_6p0 w=1.2u l=0.5u
X2677 a_6292_49944# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2678 a_7672_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2679 vss tune_shunt[7] a_21748_33058# vss nmos_6p0 w=0.51u l=0.6u
X2680 vss tune_shunt[6] a_9316_50306# vss nmos_6p0 w=0.51u l=0.6u
X2681 vdd tune_shunt[7] a_16500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X2682 vdd tune_shunt[6] a_6196_47516# vdd pmos_6p0 w=1.2u l=0.5u
X2683 a_2140_52552# a_2052_52596# vss vss nmos_6p0 w=0.82u l=1u
X2684 a_16688_42104# cap_shunt_n a_14580_42104# vss nmos_6p0 w=0.82u l=0.6u
X2685 a_37080_15448# cap_series_gygyn a_35880_14964# vss nmos_6p0 w=0.82u l=0.6u
X2686 vdd a_32268_39575# a_32180_39672# vdd pmos_6p0 w=1.22u l=1u
X2687 vss tune_shunt[7] a_17828_35832# vss nmos_6p0 w=0.51u l=0.6u
X2688 vdd a_30924_49416# a_30836_49460# vdd pmos_6p0 w=1.22u l=1u
X2689 a_13460_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2690 vss cap_shunt_p a_27888_21720# vss nmos_6p0 w=0.82u l=0.6u
X2691 a_17620_16532# cap_shunt_p a_17828_17016# vdd pmos_6p0 w=1.2u l=0.5u
X2692 a_20740_20152# cap_shunt_p a_21672_20152# vss nmos_6p0 w=0.82u l=0.6u
X2693 vdd a_25996_55255# a_25908_55352# vdd pmos_6p0 w=1.22u l=1u
X2694 vss tune_shunt[5] a_6292_18584# vss nmos_6p0 w=0.51u l=0.6u
X2695 vdd tune_shunt[7] a_16500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X2696 a_17828_43672# cap_shunt_p a_17620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X2697 vdd a_30924_46280# a_30836_46324# vdd pmos_6p0 w=1.22u l=1u
X2698 a_13460_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2699 vdd a_16476_32168# a_16388_32212# vdd pmos_6p0 w=1.22u l=1u
X2700 a_29532_9884# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2701 vdd a_25996_52119# a_25908_52216# vdd pmos_6p0 w=1.22u l=1u
X2702 a_16924_32168# a_16836_32212# vss vss nmos_6p0 w=0.82u l=1u
X2703 a_10340_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2704 vss tune_shunt[7] a_6740_15448# vss nmos_6p0 w=0.51u l=0.6u
X2705 a_35880_18100# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2706 a_27228_20759# a_27140_20856# vss vss nmos_6p0 w=0.82u l=1u
X2707 a_35692_24372# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2708 a_6508_8215# a_6420_8312# vss vss nmos_6p0 w=0.82u l=1u
X2709 vdd a_18492_52552# a_18404_52596# vdd pmos_6p0 w=1.22u l=1u
X2710 a_13588_47516# cap_shunt_p a_13796_47170# vdd pmos_6p0 w=1.2u l=0.5u
X2711 vss tune_shunt[6] a_6740_38968# vss nmos_6p0 w=0.51u l=0.6u
X2712 a_24660_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2713 a_7768_8316# cap_series_gyn a_8576_7908# vss nmos_6p0 w=0.82u l=0.6u
X2714 a_10680_8316# cap_series_gyp a_10704_7908# vss nmos_6p0 w=0.82u l=0.6u
X2715 a_29468_48983# a_29380_49080# vss vss nmos_6p0 w=0.82u l=1u
X2716 vss tune_shunt[7] a_32612_26786# vss nmos_6p0 w=0.51u l=0.6u
X2717 vdd a_6060_31735# a_5972_31832# vdd pmos_6p0 w=1.22u l=1u
X2718 vss cap_series_gyp a_27888_9176# vss nmos_6p0 w=0.82u l=0.6u
X2719 a_6532_19668# cap_shunt_p a_6740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X2720 vss tune_shunt_gy[0] a_37632_33400# vss nmos_6p0 w=0.51u l=0.6u
X2721 a_35880_14964# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2722 a_35692_21236# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2723 a_23072_29860# cap_shunt_n a_21748_29922# vss nmos_6p0 w=0.82u l=0.6u
X2724 a_16476_27464# a_16388_27508# vss vss nmos_6p0 w=0.82u l=1u
X2725 a_1924_6040# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X2726 a_14692_9176# cap_series_gyn a_14484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X2727 vdd a_28796_21192# a_28708_21236# vdd pmos_6p0 w=1.22u l=1u
X2728 vdd tune_shunt[7] a_16500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X2729 a_27104_4472# cap_shunt_p a_25780_4472# vss nmos_6p0 w=0.82u l=0.6u
X2730 a_13796_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2731 a_10452_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2732 a_4032_4472# cap_shunt_p a_1924_4472# vss nmos_6p0 w=0.82u l=0.6u
X2733 a_30428_21236# cap_series_gygyn a_30616_21236# vdd pmos_6p0 w=1.2u l=0.5u
X2734 a_13252_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2735 vdd a_14908_53687# a_14820_53784# vdd pmos_6p0 w=1.22u l=1u
X2736 vss tune_shunt[6] a_21748_39330# vss nmos_6p0 w=0.51u l=0.6u
X2737 a_23072_26724# cap_shunt_n a_21748_26786# vss nmos_6p0 w=0.82u l=0.6u
X2738 a_16476_24328# a_16388_24372# vss vss nmos_6p0 w=0.82u l=1u
X2739 a_29492_17724# cap_series_gyp a_29700_17378# vdd pmos_6p0 w=1.2u l=0.5u
X2740 a_6740_48376# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X2741 a_3620_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2742 a_14692_6040# cap_series_gyn a_14484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X2743 a_11984_17016# cap_shunt_p a_9876_17016# vss nmos_6p0 w=0.82u l=0.6u
X2744 a_6740_26424# cap_shunt_n a_6532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2745 vdd tune_shunt[7] a_16500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X2746 a_11800_7124# cap_series_gyp a_11612_7124# vdd pmos_6p0 w=1.2u l=0.5u
X2747 a_30192_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2748 a_20740_46808# cap_shunt_p a_22456_46808# vss nmos_6p0 w=0.82u l=0.6u
X2749 a_15120_34564# cap_shunt_n a_13796_34626# vss nmos_6p0 w=0.82u l=0.6u
X2750 vdd tune_shunt[7] a_20532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X2751 a_13460_32696# cap_shunt_n a_13252_32212# vdd pmos_6p0 w=1.2u l=0.5u
X2752 vdd tune_shunt[7] a_13588_13020# vdd pmos_6p0 w=1.2u l=0.5u
X2753 vss tune_shunt[6] a_9316_47170# vss nmos_6p0 w=0.51u l=0.6u
X2754 vss cap_shunt_p a_35056_27992# vss nmos_6p0 w=0.82u l=0.6u
X2755 a_14372_46324# cap_shunt_p a_14580_46808# vdd pmos_6p0 w=1.2u l=0.5u
X2756 a_18816_32996# cap_shunt_n a_16708_33058# vss nmos_6p0 w=0.82u l=0.6u
X2757 a_35880_25940# cap_series_gygyp a_35692_25940# vdd pmos_6p0 w=1.2u l=0.5u
X2758 a_34396_19624# a_34308_19668# vss vss nmos_6p0 w=0.82u l=1u
X2759 a_36652_45540# cap_shunt_gyp a_36384_45540# vss nmos_6p0 w=0.82u l=0.6u
X2760 a_6740_23288# cap_shunt_p a_6532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2761 a_17416_9476# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2762 a_33544_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2763 a_7672_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2764 a_25780_24856# cap_shunt_p a_25572_24372# vdd pmos_6p0 w=1.2u l=0.5u
X2765 a_2708_48738# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2766 a_15120_31428# cap_shunt_n a_13796_31490# vss nmos_6p0 w=0.82u l=0.6u
X2767 a_4940_6647# a_4852_6744# vss vss nmos_6p0 w=0.82u l=1u
X2768 a_23464_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X2769 a_5612_30167# a_5524_30264# vss vss nmos_6p0 w=0.82u l=1u
X2770 a_22456_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2771 a_20328_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2772 vdd a_1692_52552# a_1604_52596# vdd pmos_6p0 w=1.22u l=1u
X2773 a_13796_34626# cap_shunt_n a_13588_34972# vdd pmos_6p0 w=1.2u l=0.5u
X2774 a_10548_27992# cap_shunt_n a_10340_27508# vdd pmos_6p0 w=1.2u l=0.5u
X2775 a_12580_13396# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2776 a_35880_22804# cap_series_gygyp a_35692_22804# vdd pmos_6p0 w=1.2u l=0.5u
X2777 a_1716_3988# cap_shunt_p a_1924_4472# vdd pmos_6p0 w=1.2u l=0.5u
X2778 vss tune_shunt[7] a_17828_29560# vss nmos_6p0 w=0.51u l=0.6u
X2779 a_13252_38484# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2780 a_28692_32696# cap_shunt_p a_28484_32212# vdd pmos_6p0 w=1.2u l=0.5u
X2781 a_32464_45302# cap_shunt_gyp a_32464_44757# vdd pmos_6p0 w=1.215u l=0.5u
X2782 a_36652_42404# cap_shunt_gyn a_36384_42404# vss nmos_6p0 w=0.82u l=0.6u
X2783 a_3620_40052# cap_shunt_n a_3828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X2784 a_7672_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2785 a_25780_21720# cap_shunt_p a_25572_21236# vdd pmos_6p0 w=1.2u l=0.5u
X2786 a_4940_3511# a_4852_3608# vss vss nmos_6p0 w=0.82u l=1u
X2787 vdd a_25548_54120# a_25460_54164# vdd pmos_6p0 w=1.22u l=1u
X2788 vdd a_25996_48983# a_25908_49080# vdd pmos_6p0 w=1.22u l=1u
X2789 vdd tune_shunt_gy[5] a_37444_49080# vdd pmos_6p0 w=1.215u l=0.5u
X2790 a_5612_27031# a_5524_27128# vss vss nmos_6p0 w=0.82u l=1u
X2791 vdd a_30812_6647# a_30724_6744# vdd pmos_6p0 w=1.22u l=1u
X2792 a_13796_31490# cap_shunt_n a_13588_31836# vdd pmos_6p0 w=1.2u l=0.5u
X2793 a_8344_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2794 vss tune_shunt[7] a_9876_20152# vss nmos_6p0 w=0.51u l=0.6u
X2795 vdd a_30812_20759# a_30724_20856# vdd pmos_6p0 w=1.22u l=1u
X2796 a_34308_13020# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2797 a_7748_29922# cap_shunt_n a_9464_29860# vss nmos_6p0 w=0.82u l=0.6u
X2798 vss tune_shunt[7] a_17828_26424# vss nmos_6p0 w=0.51u l=0.6u
X2799 a_9876_15448# cap_shunt_p a_9668_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2800 a_13252_35348# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2801 a_1716_5180# cap_shunt_p a_1924_4834# vdd pmos_6p0 w=1.2u l=0.5u
X2802 a_14784_21720# cap_shunt_n a_13460_21720# vss nmos_6p0 w=0.82u l=0.6u
X2803 vss cap_series_gyp a_27888_12312# vss nmos_6p0 w=0.82u l=0.6u
X2804 vss cap_series_gyn a_17024_4772# vss nmos_6p0 w=0.82u l=0.6u
X2805 vdd tune_shunt[5] a_2500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X2806 vdd a_25548_50984# a_25460_51028# vdd pmos_6p0 w=1.22u l=1u
X2807 a_34844_5512# a_34756_5556# vss vss nmos_6p0 w=0.82u l=1u
X2808 vdd tune_series_gy[5] a_15532_11452# vdd pmos_6p0 w=1.2u l=0.5u
X2809 a_27228_14487# a_27140_14584# vss vss nmos_6p0 w=0.82u l=1u
X2810 a_36160_44757# cap_shunt_gyn a_36160_45302# vdd pmos_6p0 w=1.215u l=0.5u
X2811 a_37080_6040# cap_series_gygyn a_35880_5556# vss nmos_6p0 w=0.82u l=0.6u
X2812 a_27104_13880# cap_series_gyn a_25780_13880# vss nmos_6p0 w=0.82u l=0.6u
X2813 a_7748_26786# cap_shunt_n a_9464_26724# vss nmos_6p0 w=0.82u l=0.6u
X2814 a_6060_5079# a_5972_5176# vss vss nmos_6p0 w=0.82u l=1u
X2815 a_9876_12312# cap_shunt_p a_9668_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2816 vdd a_29692_43144# a_29604_43188# vdd pmos_6p0 w=1.22u l=1u
X2817 a_13228_54120# a_13140_54164# vss vss nmos_6p0 w=0.82u l=1u
X2818 vdd a_6060_25463# a_5972_25560# vdd pmos_6p0 w=1.22u l=1u
X2819 a_16924_22760# a_16836_22804# vss vss nmos_6p0 w=0.82u l=1u
X2820 a_27228_11351# a_27140_11448# vss vss nmos_6p0 w=0.82u l=1u
X2821 a_27104_10744# cap_series_gyn a_25780_10744# vss nmos_6p0 w=0.82u l=0.6u
X2822 vdd tune_shunt[4] a_3620_13396# vdd pmos_6p0 w=1.2u l=0.5u
X2823 a_13588_38108# cap_shunt_n a_13796_37762# vdd pmos_6p0 w=1.2u l=0.5u
X2824 vdd tune_shunt[6] a_10452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X2825 a_21540_30268# cap_shunt_n a_21748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X2826 a_24660_17378# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2827 vdd a_28236_47848# a_28148_47892# vdd pmos_6p0 w=1.22u l=1u
X2828 a_20532_43188# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2829 a_7616_17316# cap_shunt_p a_6292_17378# vss nmos_6p0 w=0.82u l=0.6u
X2830 vdd tune_shunt[7] a_16500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X2831 a_13796_39330# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2832 a_21748_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2833 a_28692_6040# tune_shunt[0] vss vss nmos_6p0 w=0.51u l=0.6u
X2834 vdd a_24540_3511# a_24452_3608# vdd pmos_6p0 w=1.22u l=1u
X2835 vss cap_series_gyn a_26768_9476# vss nmos_6p0 w=0.82u l=0.6u
X2836 a_35880_13396# cap_series_gygyn a_36688_13880# vss nmos_6p0 w=0.82u l=0.6u
X2837 vdd a_28236_44712# a_28148_44756# vdd pmos_6p0 w=1.22u l=1u
X2838 a_10988_7080# a_10900_7124# vss vss nmos_6p0 w=0.82u l=1u
X2839 vdd a_31260_3944# a_31172_3988# vdd pmos_6p0 w=1.22u l=1u
X2840 vdd tune_shunt[7] a_16500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X2841 a_15120_28292# cap_shunt_n a_13796_28354# vss nmos_6p0 w=0.82u l=0.6u
X2842 vss tune_series_gy[4] a_32632_14588# vss nmos_6p0 w=0.51u l=0.6u
X2843 vdd a_4492_5079# a_4404_5176# vdd pmos_6p0 w=1.22u l=1u
X2844 vss tune_shunt[7] a_16708_37762# vss nmos_6p0 w=0.51u l=0.6u
X2845 a_23072_17316# cap_shunt_p a_21748_17378# vss nmos_6p0 w=0.82u l=0.6u
X2846 a_16016_7608# cap_series_gyp a_14692_7608# vss nmos_6p0 w=0.82u l=0.6u
X2847 a_25984_4772# cap_series_gyp a_24660_4834# vss nmos_6p0 w=0.82u l=0.6u
X2848 a_12264_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X2849 vss cap_series_gygyn a_37080_6040# vss nmos_6p0 w=0.82u l=0.6u
X2850 a_35880_10260# cap_series_gygyp a_36688_10744# vss nmos_6p0 w=0.82u l=0.6u
X2851 vdd a_2140_55688# a_2052_55732# vdd pmos_6p0 w=1.22u l=1u
X2852 a_25780_43672# cap_shunt_p a_26712_43672# vss nmos_6p0 w=0.82u l=0.6u
X2853 vdd tune_shunt[4] a_24452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X2854 a_36524_38007# a_36436_38104# vss vss nmos_6p0 w=0.82u l=1u
X2855 a_33524_35348# cap_shunt_n a_33732_35832# vdd pmos_6p0 w=1.2u l=0.5u
X2856 a_15120_25156# cap_shunt_n a_13796_25218# vss nmos_6p0 w=0.82u l=0.6u
X2857 vss tune_series_gy[3] a_32632_11452# vss nmos_6p0 w=0.51u l=0.6u
X2858 a_13588_47516# cap_shunt_p a_13796_47170# vdd pmos_6p0 w=1.2u l=0.5u
X2859 vss tune_shunt[7] a_16708_34626# vss nmos_6p0 w=0.51u l=0.6u
X2860 vdd tune_shunt[7] a_33524_27508# vdd pmos_6p0 w=1.2u l=0.5u
X2861 a_7176_6040# cap_series_gyp a_6760_5556# vss nmos_6p0 w=0.82u l=0.6u
X2862 a_18816_23588# cap_shunt_n a_16708_23650# vss nmos_6p0 w=0.82u l=0.6u
X2863 a_6628_12674# cap_shunt_p a_6420_13020# vdd pmos_6p0 w=1.2u l=0.5u
X2864 a_35880_16532# cap_series_gygyn a_35692_16532# vdd pmos_6p0 w=1.2u l=0.5u
X2865 a_21672_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2866 a_14580_43672# cap_shunt_n a_15512_43672# vss nmos_6p0 w=0.82u l=0.6u
X2867 a_25780_40536# cap_shunt_n a_26712_40536# vss nmos_6p0 w=0.82u l=0.6u
X2868 a_6760_3988# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X2869 a_7768_8316# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X2870 a_24452_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2871 a_5544_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2872 vss cap_shunt_p a_4032_20452# vss nmos_6p0 w=0.82u l=0.6u
X2873 a_31624_6748# cap_series_gygyn a_31436_6748# vdd pmos_6p0 w=1.2u l=0.5u
X2874 vdd a_1692_43144# a_1604_43188# vdd pmos_6p0 w=1.22u l=1u
X2875 a_13796_25218# cap_shunt_n a_13588_25564# vdd pmos_6p0 w=1.2u l=0.5u
X2876 a_18612_4834# cap_series_gyp a_19544_4772# vss nmos_6p0 w=0.82u l=0.6u
X2877 a_30428_21236# cap_series_gygyn a_30616_21236# vdd pmos_6p0 w=1.2u l=0.5u
X2878 a_14580_40536# cap_shunt_n a_15512_40536# vss nmos_6p0 w=0.82u l=0.6u
X2879 a_13252_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2880 a_16252_47848# a_16164_47892# vss vss nmos_6p0 w=0.82u l=1u
X2881 a_24428_47848# a_24340_47892# vss vss nmos_6p0 w=0.82u l=1u
X2882 vss tune_series_gygy[2] a_35880_5556# vss nmos_6p0 w=0.51u l=0.6u
X2883 a_7768_5180# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X2884 a_29492_17724# cap_series_gyp a_29700_17378# vdd pmos_6p0 w=1.2u l=0.5u
X2885 a_5612_17623# a_5524_17720# vss vss nmos_6p0 w=0.82u l=1u
X2886 a_27340_55255# a_27252_55352# vss vss nmos_6p0 w=0.82u l=1u
X2887 a_17640_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2888 a_13796_22082# cap_shunt_n a_13588_22428# vdd pmos_6p0 w=1.2u l=0.5u
X2889 a_17828_34264# cap_shunt_n a_17620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X2890 a_9316_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2891 a_18404_3988# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2892 vss tune_shunt[7] a_17828_17016# vss nmos_6p0 w=0.51u l=0.6u
X2893 vss cap_shunt_n a_19152_35832# vss nmos_6p0 w=0.82u l=0.6u
X2894 a_4032_32996# cap_shunt_p a_2708_33058# vss nmos_6p0 w=0.82u l=0.6u
X2895 a_21748_7970# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2896 a_32928_45944# cap_shunt_gyn a_32948_45540# vss nmos_6p0 w=0.82u l=0.6u
X2897 a_17620_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2898 vdd tune_shunt[3] a_2500_11452# vdd pmos_6p0 w=1.2u l=0.5u
X2899 vdd a_21964_53687# a_21876_53784# vdd pmos_6p0 w=1.22u l=1u
X2900 a_17640_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2901 a_17828_31128# cap_shunt_n a_17620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X2902 vss cap_series_gyn a_21840_13880# vss nmos_6p0 w=0.82u l=0.6u
X2903 a_10540_44712# a_10452_44756# vss vss nmos_6p0 w=0.82u l=1u
X2904 a_16500_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2905 vdd a_34396_25896# a_34308_25940# vdd pmos_6p0 w=1.22u l=1u
X2906 a_21748_4834# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X2907 a_28692_15448# cap_series_gyn a_28484_14964# vdd pmos_6p0 w=1.2u l=0.5u
X2908 a_15356_16488# a_15268_16532# vss vss nmos_6p0 w=0.82u l=1u
X2909 a_13796_34626# cap_shunt_n a_13588_34972# vdd pmos_6p0 w=1.2u l=0.5u
X2910 vdd tune_shunt[7] a_7540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X2911 a_35488_41621# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X2912 a_17620_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2913 a_2500_13020# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2914 vdd a_10764_53687# a_10676_53784# vdd pmos_6p0 w=1.22u l=1u
X2915 vdd a_21964_50551# a_21876_50648# vdd pmos_6p0 w=1.22u l=1u
X2916 a_10340_38484# cap_shunt_n a_10548_38968# vdd pmos_6p0 w=1.2u l=0.5u
X2917 a_21540_28700# cap_shunt_n a_21748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X2918 vss tune_series_gy[3] a_14692_4472# vss nmos_6p0 w=0.51u l=0.6u
X2919 vss cap_series_gyn a_21840_10744# vss nmos_6p0 w=0.82u l=0.6u
X2920 a_10808_13880# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2921 a_10540_41576# a_10452_41620# vss vss nmos_6p0 w=0.82u l=1u
X2922 vss cap_shunt_n a_8064_38968# vss nmos_6p0 w=0.82u l=0.6u
X2923 vdd a_34396_22760# a_34308_22804# vdd pmos_6p0 w=1.22u l=1u
X2924 vdd a_10540_3944# a_10452_3988# vdd pmos_6p0 w=1.22u l=1u
X2925 a_28692_12312# cap_series_gyn a_28484_11828# vdd pmos_6p0 w=1.2u l=0.5u
X2926 a_13796_31490# cap_shunt_n a_13588_31836# vdd pmos_6p0 w=1.2u l=0.5u
X2927 vdd a_27228_9783# a_27140_9880# vdd pmos_6p0 w=1.22u l=1u
X2928 vss tune_shunt[6] a_20740_37400# vss nmos_6p0 w=0.51u l=0.6u
X2929 vdd a_6060_12919# a_5972_13016# vdd pmos_6p0 w=1.22u l=1u
X2930 vss cap_shunt_p a_26768_32996# vss nmos_6p0 w=0.82u l=0.6u
X2931 vdd tune_shunt[7] a_9108_22428# vdd pmos_6p0 w=1.2u l=0.5u
X2932 a_21748_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2933 a_10340_35348# cap_shunt_n a_10548_35832# vdd pmos_6p0 w=1.2u l=0.5u
X2934 a_10808_10744# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2935 a_20532_18100# cap_shunt_p a_20740_18584# vdd pmos_6p0 w=1.2u l=0.5u
X2936 a_30800_38968# cap_shunt_n a_28692_38968# vss nmos_6p0 w=0.82u l=0.6u
X2937 vdd a_5500_11784# a_5412_11828# vdd pmos_6p0 w=1.22u l=1u
X2938 vdd a_2140_49416# a_2052_49460# vdd pmos_6p0 w=1.22u l=1u
X2939 a_28484_40052# cap_shunt_p a_28692_40536# vdd pmos_6p0 w=1.2u l=0.5u
X2940 vdd tune_shunt[6] a_24452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X2941 vdd tune_shunt[5] a_2500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X2942 a_33524_29076# cap_shunt_p a_33732_29560# vdd pmos_6p0 w=1.2u l=0.5u
X2943 vdd a_27228_6647# a_27140_6744# vdd pmos_6p0 w=1.22u l=1u
X2944 vss tune_shunt[7] a_16708_28354# vss nmos_6p0 w=0.51u l=0.6u
X2945 a_21748_42466# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X2946 a_32604_35304# a_32516_35348# vss vss nmos_6p0 w=0.82u l=1u
X2947 vdd tune_shunt[1] a_25572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X2948 vdd tune_shunt[6] a_24452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X2949 a_18404_13020# cap_series_gyn a_18612_12674# vdd pmos_6p0 w=1.2u l=0.5u
X2950 a_29532_16156# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2951 a_17828_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2952 vdd a_2140_46280# a_2052_46324# vdd pmos_6p0 w=1.22u l=1u
X2953 a_34144_45540# cap_shunt_gyn a_34144_45944# vdd pmos_6p0 w=1.215u l=0.5u
X2954 a_37632_41621# cap_shunt_gyp a_37652_42104# vss nmos_6p0 w=0.82u l=0.6u
X2955 a_25780_34264# cap_shunt_p a_26712_34264# vss nmos_6p0 w=0.82u l=0.6u
X2956 vdd tune_shunt[7] a_7540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X2957 a_9540_14242# cap_shunt_p a_9332_14588# vdd pmos_6p0 w=1.2u l=0.5u
X2958 a_35056_34264# cap_shunt_n a_33732_34264# vss nmos_6p0 w=0.82u l=0.6u
X2959 vdd a_6508_33303# a_6420_33400# vdd pmos_6p0 w=1.22u l=1u
X2960 a_13588_38108# cap_shunt_n a_13796_37762# vdd pmos_6p0 w=1.2u l=0.5u
X2961 vss cap_shunt_n a_4032_14180# vss nmos_6p0 w=0.82u l=0.6u
X2962 vss tune_shunt[7] a_16708_25218# vss nmos_6p0 w=0.51u l=0.6u
X2963 vdd a_35740_52552# a_35652_52596# vdd pmos_6p0 w=1.22u l=1u
X2964 a_6420_14588# cap_shunt_p a_6628_14242# vdd pmos_6p0 w=1.2u l=0.5u
X2965 a_13796_18946# cap_shunt_p a_13588_19292# vdd pmos_6p0 w=1.2u l=0.5u
X2966 vss tune_shunt[4] a_16708_48738# vss nmos_6p0 w=0.51u l=0.6u
X2967 a_20284_54120# a_20196_54164# vss vss nmos_6p0 w=0.82u l=1u
X2968 a_34144_42404# cap_shunt_gyn a_34144_42808# vdd pmos_6p0 w=1.215u l=0.5u
X2969 vss tune_shunt[5] a_24660_40898# vss nmos_6p0 w=0.51u l=0.6u
X2970 a_25780_31128# cap_shunt_p a_26712_31128# vss nmos_6p0 w=0.82u l=0.6u
X2971 a_6740_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2972 a_35056_31128# cap_shunt_n a_33732_31128# vss nmos_6p0 w=0.82u l=0.6u
X2973 a_24452_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2974 vss cap_shunt_n a_4032_11044# vss nmos_6p0 w=0.82u l=0.6u
X2975 a_27340_48983# a_27252_49080# vss vss nmos_6p0 w=0.82u l=1u
X2976 a_17620_46324# cap_shunt_n a_17828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X2977 vdd a_34844_24328# a_34756_24372# vdd pmos_6p0 w=1.22u l=1u
X2978 a_13796_15810# cap_shunt_p a_13588_16156# vdd pmos_6p0 w=1.2u l=0.5u
X2979 vdd a_32716_52552# a_32628_52596# vdd pmos_6p0 w=1.22u l=1u
X2980 a_36324_41621# cap_shunt_gyn a_36512_41621# vdd pmos_6p0 w=1.215u l=0.5u
X2981 a_33732_32696# cap_shunt_n a_33524_32212# vdd pmos_6p0 w=1.2u l=0.5u
X2982 vss cap_shunt_n a_19152_29560# vss nmos_6p0 w=0.82u l=0.6u
X2983 a_6740_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X2984 a_7540_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2985 a_12656_34264# cap_shunt_n a_10548_34264# vss nmos_6p0 w=0.82u l=0.6u
X2986 a_22436_10260# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X2987 a_19524_10260# cap_series_gyn a_19732_10744# vdd pmos_6p0 w=1.2u l=0.5u
X2988 a_30616_21236# cap_series_gygyn a_31424_21720# vss nmos_6p0 w=0.82u l=0.6u
X2989 a_29132_50984# a_29044_51028# vss vss nmos_6p0 w=0.82u l=1u
X2990 a_2140_38440# a_2052_38484# vss vss nmos_6p0 w=0.82u l=1u
X2991 vdd a_13340_52552# a_13252_52596# vdd pmos_6p0 w=1.22u l=1u
X2992 a_17640_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X2993 vss tune_shunt[5] a_3828_21720# vss nmos_6p0 w=0.51u l=0.6u
X2994 vdd a_34844_21192# a_34756_21236# vdd pmos_6p0 w=1.22u l=1u
X2995 a_7224_51512# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X2996 a_10660_44034# cap_shunt_n a_12376_43972# vss nmos_6p0 w=0.82u l=0.6u
X2997 a_17828_24856# cap_shunt_n a_17620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X2998 vss cap_shunt_n a_19152_26424# vss nmos_6p0 w=0.82u l=0.6u
X2999 a_35904_7608# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X3000 vdd a_32268_47848# a_32180_47892# vdd pmos_6p0 w=1.22u l=1u
X3001 a_12656_31128# cap_shunt_n a_10548_31128# vss nmos_6p0 w=0.82u l=0.6u
X3002 a_4032_23588# cap_shunt_p a_2708_23650# vss nmos_6p0 w=0.82u l=0.6u
X3003 a_7580_5180# cap_series_gyn a_7768_5180# vdd pmos_6p0 w=1.2u l=0.5u
X3004 vss cap_shunt_n a_13776_46808# vss nmos_6p0 w=0.82u l=0.6u
X3005 a_17620_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3006 a_37444_33781# cap_shunt_gyn a_37632_33781# vdd pmos_6p0 w=1.215u l=0.5u
X3007 a_17640_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3008 a_10660_40898# cap_shunt_n a_12376_40836# vss nmos_6p0 w=0.82u l=0.6u
X3009 a_10492_8316# cap_series_gyp a_10680_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3010 a_21748_12674# cap_series_gyn a_22680_12612# vss nmos_6p0 w=0.82u l=0.6u
X3011 a_21540_20860# cap_shunt_p a_21748_20514# vdd pmos_6p0 w=1.2u l=0.5u
X3012 a_17828_21720# cap_shunt_p a_17620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X3013 a_14692_4472# cap_series_gyp a_14484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3014 vdd a_34396_16488# a_34308_16532# vdd pmos_6p0 w=1.22u l=1u
X3015 a_13796_25218# cap_shunt_n a_13588_25564# vdd pmos_6p0 w=1.2u l=0.5u
X3016 vss tune_series_gy[5] a_21748_9538# vss nmos_6p0 w=0.51u l=0.6u
X3017 a_33024_47108# cap_shunt_gyn a_33024_47512# vdd pmos_6p0 w=1.215u l=0.5u
X3018 a_10340_29076# cap_shunt_n a_10548_29560# vdd pmos_6p0 w=1.2u l=0.5u
X3019 vdd a_12444_21192# a_12356_21236# vdd pmos_6p0 w=1.22u l=1u
X3020 a_13460_27992# cap_shunt_n a_15176_27992# vss nmos_6p0 w=0.82u l=0.6u
X3021 a_11648_12612# cap_shunt_p a_9540_12674# vss nmos_6p0 w=0.82u l=0.6u
X3022 a_29492_17724# cap_series_gyp a_29700_17378# vdd pmos_6p0 w=1.2u l=0.5u
X3023 vss cap_shunt_p a_8624_20452# vss nmos_6p0 w=0.82u l=0.6u
X3024 vss tune_series_gygy[5] a_30616_21236# vss nmos_6p0 w=0.51u l=0.6u
X3025 a_36384_47512# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X3026 vdd a_7404_55255# a_7316_55352# vdd pmos_6p0 w=1.22u l=1u
X3027 a_13796_22082# cap_shunt_n a_13588_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3028 a_35692_7124# cap_series_gygyp a_35880_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3029 a_6532_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3030 vss cap_shunt_p a_26768_23588# vss nmos_6p0 w=0.82u l=0.6u
X3031 a_27676_20759# a_27588_20856# vss vss nmos_6p0 w=0.82u l=1u
X3032 a_33500_54120# a_33412_54164# vss vss nmos_6p0 w=0.82u l=1u
X3033 a_21748_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3034 a_32604_29032# a_32516_29076# vss vss nmos_6p0 w=0.82u l=1u
X3035 a_13460_24856# cap_shunt_n a_15176_24856# vss nmos_6p0 w=0.82u l=0.6u
X3036 a_20740_20152# cap_shunt_p a_20532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X3037 vdd a_23420_54120# a_23332_54164# vdd pmos_6p0 w=1.22u l=1u
X3038 vdd a_31708_42711# a_31620_42808# vdd pmos_6p0 w=1.22u l=1u
X3039 vdd tune_shunt[3] a_2500_11452# vdd pmos_6p0 w=1.2u l=0.5u
X3040 a_7616_49944# cap_shunt_p a_6292_49944# vss nmos_6p0 w=0.82u l=0.6u
X3041 vdd tune_shunt[7] a_24452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X3042 a_20740_42104# cap_shunt_p a_20532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X3043 a_8576_6340# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X3044 a_31808_36132# cap_shunt_n a_29700_36194# vss nmos_6p0 w=0.82u l=0.6u
X3045 a_28692_15448# cap_series_gyn a_28484_14964# vdd pmos_6p0 w=1.2u l=0.5u
X3046 a_8008_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3047 a_16708_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3048 a_21748_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3049 a_32604_25896# a_32516_25940# vss vss nmos_6p0 w=0.82u l=1u
X3050 a_18404_5180# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3051 a_9668_13396# cap_shunt_p a_9876_13880# vdd pmos_6p0 w=1.2u l=0.5u
X3052 vdd a_23420_50984# a_23332_51028# vdd pmos_6p0 w=1.22u l=1u
X3053 vdd tune_shunt[6] a_14372_44756# vdd pmos_6p0 w=1.2u l=0.5u
X3054 a_10340_38484# cap_shunt_n a_10548_38968# vdd pmos_6p0 w=1.2u l=0.5u
X3055 vdd a_23308_14920# a_23220_14964# vdd pmos_6p0 w=1.22u l=1u
X3056 a_12580_49460# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3057 a_9540_9538# cap_shunt_p a_9332_9884# vdd pmos_6p0 w=1.2u l=0.5u
X3058 a_2708_9538# cap_shunt_n a_2500_9884# vdd pmos_6p0 w=1.2u l=0.5u
X3059 a_28692_12312# cap_series_gyn a_28484_11828# vdd pmos_6p0 w=1.2u l=0.5u
X3060 vss cap_shunt_p a_15120_18884# vss nmos_6p0 w=0.82u l=0.6u
X3061 a_7540_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3062 a_10340_35348# cap_shunt_n a_10548_35832# vdd pmos_6p0 w=1.2u l=0.5u
X3063 a_9428_20514# cap_shunt_p a_9220_20860# vdd pmos_6p0 w=1.2u l=0.5u
X3064 vss tune_shunt[7] a_10660_26786# vss nmos_6p0 w=0.51u l=0.6u
X3065 a_30028_49416# a_29940_49460# vss vss nmos_6p0 w=0.82u l=1u
X3066 a_29132_44712# a_29044_44756# vss vss nmos_6p0 w=0.82u l=1u
X3067 a_28484_40052# cap_shunt_p a_28692_40536# vdd pmos_6p0 w=1.2u l=0.5u
X3068 a_9668_16532# cap_shunt_p a_9876_17016# vdd pmos_6p0 w=1.2u l=0.5u
X3069 vss tune_shunt[6] a_25780_37400# vss nmos_6p0 w=0.51u l=0.6u
X3070 a_17640_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3071 a_6308_20860# cap_shunt_p a_6516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X3072 vss cap_shunt_p a_15120_15748# vss nmos_6p0 w=0.82u l=0.6u
X3073 a_16252_53687# a_16164_53784# vss vss nmos_6p0 w=0.82u l=1u
X3074 vdd a_22412_47415# a_22324_47512# vdd pmos_6p0 w=1.22u l=1u
X3075 vdd a_35292_38440# a_35204_38484# vdd pmos_6p0 w=1.22u l=1u
X3076 a_6740_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3077 a_7540_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3078 a_32612_29922# cap_shunt_p a_34328_29860# vss nmos_6p0 w=0.82u l=0.6u
X3079 vss tune_shunt[4] a_13796_50306# vss nmos_6p0 w=0.51u l=0.6u
X3080 a_30028_46280# a_29940_46324# vss vss nmos_6p0 w=0.82u l=1u
X3081 a_11780_6040# cap_series_gyn a_11572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X3082 a_33524_33780# cap_shunt_n a_33732_34264# vdd pmos_6p0 w=1.2u l=0.5u
X3083 a_18404_13020# cap_series_gyn a_18612_12674# vdd pmos_6p0 w=1.2u l=0.5u
X3084 a_29532_16156# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3085 a_17640_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3086 a_9540_14242# cap_shunt_p a_9332_14588# vdd pmos_6p0 w=1.2u l=0.5u
X3087 a_10660_34626# cap_shunt_n a_12376_34564# vss nmos_6p0 w=0.82u l=0.6u
X3088 vdd tune_series_gy[3] a_15492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X3089 vss cap_shunt_p a_19152_17016# vss nmos_6p0 w=0.82u l=0.6u
X3090 vdd a_20172_30167# a_20084_30264# vdd pmos_6p0 w=1.22u l=1u
X3091 a_32612_26786# cap_shunt_p a_34328_26724# vss nmos_6p0 w=0.82u l=0.6u
X3092 vdd a_8860_18056# a_8772_18100# vdd pmos_6p0 w=1.22u l=1u
X3093 a_13796_18946# cap_shunt_p a_13588_19292# vdd pmos_6p0 w=1.2u l=0.5u
X3094 a_13796_48738# cap_shunt_n a_13588_49084# vdd pmos_6p0 w=1.2u l=0.5u
X3095 vss tune_shunt[4] a_29700_23650# vss nmos_6p0 w=0.51u l=0.6u
X3096 a_33524_30644# cap_shunt_n a_33732_31128# vdd pmos_6p0 w=1.2u l=0.5u
X3097 a_6572_7124# cap_series_gyp a_6760_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3098 vdd a_25996_54120# a_25908_54164# vdd pmos_6p0 w=1.22u l=1u
X3099 a_8064_48376# cap_shunt_p a_6740_48376# vss nmos_6p0 w=0.82u l=0.6u
X3100 a_25780_42104# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3101 a_3932_55255# a_3844_55352# vss vss nmos_6p0 w=0.82u l=1u
X3102 a_10660_31490# cap_shunt_n a_12376_31428# vss nmos_6p0 w=0.82u l=0.6u
X3103 a_21540_11452# cap_series_gyn a_21748_11106# vdd pmos_6p0 w=1.2u l=0.5u
X3104 vss cap_shunt_n a_7952_3204# vss nmos_6p0 w=0.82u l=0.6u
X3105 vdd a_18156_50551# a_18068_50648# vdd pmos_6p0 w=1.22u l=1u
X3106 a_21636_6040# cap_series_gyp a_21428_5556# vdd pmos_6p0 w=1.2u l=0.5u
X3107 a_13796_15810# cap_shunt_p a_13588_16156# vdd pmos_6p0 w=1.2u l=0.5u
X3108 a_11592_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3109 a_17828_18584# cap_shunt_p a_17620_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3110 vdd tune_shunt[6] a_3620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X3111 vdd a_25996_50984# a_25908_51028# vdd pmos_6p0 w=1.22u l=1u
X3112 a_33500_47848# a_33412_47892# vss vss nmos_6p0 w=0.82u l=1u
X3113 a_19524_10260# cap_series_gyn a_19732_10744# vdd pmos_6p0 w=1.2u l=0.5u
X3114 a_27676_14487# a_27588_14584# vss vss nmos_6p0 w=0.82u l=1u
X3115 a_34516_18946# cap_series_gygyn a_35448_18884# vss nmos_6p0 w=0.82u l=0.6u
X3116 a_30528_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X3117 a_21748_42466# cap_shunt_n a_21540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X3118 a_13676_54120# a_13588_54164# vss vss nmos_6p0 w=0.82u l=1u
X3119 vss cap_shunt_n a_22064_37400# vss nmos_6p0 w=0.82u l=0.6u
X3120 vss tune_series_gy[1] a_10548_3266# vss nmos_6p0 w=0.51u l=0.6u
X3121 vdd a_4380_53687# a_4292_53784# vdd pmos_6p0 w=1.22u l=1u
X3122 a_27676_11351# a_27588_11448# vss vss nmos_6p0 w=0.82u l=1u
X3123 vdd a_3036_33736# a_2948_33780# vdd pmos_6p0 w=1.22u l=1u
X3124 a_34516_15810# cap_series_gygyn a_35448_15748# vss nmos_6p0 w=0.82u l=0.6u
X3125 a_24752_9176# cap_series_gyp a_22644_9176# vss nmos_6p0 w=0.82u l=0.6u
X3126 a_16028_33736# a_15940_33780# vss vss nmos_6p0 w=0.82u l=1u
X3127 a_20740_32696# cap_shunt_n a_20532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X3128 vdd a_28684_47848# a_28596_47892# vdd pmos_6p0 w=1.22u l=1u
X3129 a_13588_28700# cap_shunt_n a_13796_28354# vdd pmos_6p0 w=1.2u l=0.5u
X3130 vss tune_shunt[7] a_2708_23650# vss nmos_6p0 w=0.51u l=0.6u
X3131 vdd a_9644_3944# a_9556_3988# vdd pmos_6p0 w=1.22u l=1u
X3132 a_21540_20860# cap_shunt_p a_21748_20514# vdd pmos_6p0 w=1.2u l=0.5u
X3133 vdd a_28236_55255# a_28148_55352# vdd pmos_6p0 w=1.22u l=1u
X3134 vdd tune_shunt[6] a_17620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X3135 vss tune_shunt[7] a_10660_29922# vss nmos_6p0 w=0.51u l=0.6u
X3136 a_19732_12312# cap_series_gyn a_20664_12312# vss nmos_6p0 w=0.82u l=0.6u
X3137 vdd a_3036_30600# a_2948_30644# vdd pmos_6p0 w=1.22u l=1u
X3138 vss cap_series_gyn a_23632_4472# vss nmos_6p0 w=0.82u l=0.6u
X3139 a_32604_16488# a_32516_16532# vss vss nmos_6p0 w=0.82u l=1u
X3140 a_3828_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3141 a_10340_29076# cap_shunt_n a_10548_29560# vdd pmos_6p0 w=1.2u l=0.5u
X3142 a_24660_39330# cap_shunt_p a_24452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X3143 a_16028_30600# a_15940_30644# vss vss nmos_6p0 w=0.82u l=1u
X3144 a_3172_49460# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3145 vdd a_28684_44712# a_28596_44756# vdd pmos_6p0 w=1.22u l=1u
X3146 vss tune_shunt[5] a_2708_20514# vss nmos_6p0 w=0.51u l=0.6u
X3147 vdd a_28236_52119# a_28148_52216# vdd pmos_6p0 w=1.22u l=1u
X3148 vss tune_shunt[6] a_13796_47170# vss nmos_6p0 w=0.51u l=0.6u
X3149 a_5612_6647# a_5524_6744# vss vss nmos_6p0 w=0.82u l=1u
X3150 a_5152_45240# cap_shunt_p a_3828_45240# vss nmos_6p0 w=0.82u l=0.6u
X3151 a_20172_48983# a_20084_49080# vss vss nmos_6p0 w=0.82u l=1u
X3152 a_21540_45948# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3153 vdd tune_series_gy[5] a_22436_8692# vdd pmos_6p0 w=1.2u l=0.5u
X3154 vss cap_series_gyn a_16576_3204# vss nmos_6p0 w=0.82u l=0.6u
X3155 a_3620_19668# cap_shunt_p a_3828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X3156 a_10340_33780# cap_shunt_n a_10548_34264# vdd pmos_6p0 w=1.2u l=0.5u
X3157 a_34308_5180# cap_series_gygyp a_34516_4834# vdd pmos_6p0 w=1.2u l=0.5u
X3158 a_19936_27992# cap_shunt_n a_17828_27992# vss nmos_6p0 w=0.82u l=0.6u
X3159 a_7540_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3160 a_3620_41620# cap_shunt_p a_3828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X3161 vss tune_series_gygy[5] a_31624_20860# vss nmos_6p0 w=0.51u l=0.6u
X3162 vss tune_shunt[6] a_13796_44034# vss nmos_6p0 w=0.51u l=0.6u
X3163 a_25780_20152# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3164 a_5152_42104# cap_shunt_p a_3828_42104# vss nmos_6p0 w=0.82u l=0.6u
X3165 a_10492_8316# cap_series_gyp a_10680_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3166 a_11984_51512# cap_shunt_n a_9876_51512# vss nmos_6p0 w=0.82u l=0.6u
X3167 a_10660_28354# cap_shunt_n a_12376_28292# vss nmos_6p0 w=0.82u l=0.6u
X3168 a_9876_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3169 a_28692_27992# cap_shunt_p a_30408_27992# vss nmos_6p0 w=0.82u l=0.6u
X3170 a_10340_30644# cap_shunt_n a_10548_31128# vdd pmos_6p0 w=1.2u l=0.5u
X3171 a_13588_30268# cap_shunt_n a_13796_29922# vdd pmos_6p0 w=1.2u l=0.5u
X3172 a_19936_24856# cap_shunt_n a_17828_24856# vss nmos_6p0 w=0.82u l=0.6u
X3173 a_2140_44279# a_2052_44376# vss vss nmos_6p0 w=0.82u l=1u
X3174 vdd a_10092_7080# a_10004_7124# vdd pmos_6p0 w=1.22u l=1u
X3175 a_10660_25218# cap_shunt_n a_12376_25156# vss nmos_6p0 w=0.82u l=0.6u
X3176 a_14692_6040# cap_series_gyn a_16408_6040# vss nmos_6p0 w=0.82u l=0.6u
X3177 a_28692_24856# cap_shunt_p a_30408_24856# vss nmos_6p0 w=0.82u l=0.6u
X3178 vss cap_shunt_p a_5152_21720# vss nmos_6p0 w=0.82u l=0.6u
X3179 vdd a_34844_41143# a_34756_41240# vdd pmos_6p0 w=1.22u l=1u
X3180 a_33612_16055# a_33524_16152# vss vss nmos_6p0 w=0.82u l=1u
X3181 vdd a_16812_54120# a_16724_54164# vdd pmos_6p0 w=1.22u l=1u
X3182 vss tune_series_gy[5] a_29700_14242# vss nmos_6p0 w=0.51u l=0.6u
X3183 a_32464_46325# cap_shunt_gyn a_32464_46870# vdd pmos_6p0 w=1.215u l=0.5u
X3184 a_2140_41143# a_2052_41240# vss vss nmos_6p0 w=0.82u l=1u
X3185 a_24660_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3186 a_32444_11452# cap_series_gyp a_32632_11452# vdd pmos_6p0 w=1.2u l=0.5u
X3187 a_24876_47848# a_24788_47892# vss vss nmos_6p0 w=0.82u l=1u
X3188 a_29700_28354# cap_shunt_p a_29492_28700# vdd pmos_6p0 w=1.2u l=0.5u
X3189 a_9428_20514# cap_shunt_p a_9220_20860# vdd pmos_6p0 w=1.2u l=0.5u
X3190 a_24204_21192# a_24116_21236# vss vss nmos_6p0 w=0.82u l=1u
X3191 a_4816_47108# cap_shunt_p a_2708_47170# vss nmos_6p0 w=0.82u l=0.6u
X3192 a_7768_8316# cap_series_gyn a_7792_7908# vss nmos_6p0 w=0.82u l=0.6u
X3193 a_28484_40052# cap_shunt_p a_28692_40536# vdd pmos_6p0 w=1.2u l=0.5u
X3194 a_16708_37762# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3195 a_21748_36194# cap_shunt_n a_21540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X3196 vdd tune_shunt[6] a_16500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X3197 vss cap_shunt_n a_4816_29860# vss nmos_6p0 w=0.82u l=0.6u
X3198 a_11592_23588# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3199 vss tune_series_gy[4] a_29700_11106# vss nmos_6p0 w=0.51u l=0.6u
X3200 a_6308_20860# cap_shunt_p a_6516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X3201 a_26444_49416# a_26356_49460# vss vss nmos_6p0 w=0.82u l=1u
X3202 a_7748_23650# cap_shunt_p a_7540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X3203 vss tune_shunt[0] a_28692_6040# vss nmos_6p0 w=0.51u l=0.6u
X3204 a_16708_37762# cap_shunt_n a_18424_37700# vss nmos_6p0 w=0.82u l=0.6u
X3205 a_2856_4772# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3206 a_5096_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3207 a_26768_37700# cap_shunt_p a_24660_37762# vss nmos_6p0 w=0.82u l=0.6u
X3208 a_17620_41620# cap_shunt_n a_17828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X3209 a_16708_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3210 a_21748_33058# cap_shunt_n a_21540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X3211 a_24452_23996# cap_shunt_p a_24660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X3212 a_9204_51874# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3213 vss tune_shunt[6] a_6740_43672# vss nmos_6p0 w=0.51u l=0.6u
X3214 vss cap_shunt_p a_4816_26724# vss nmos_6p0 w=0.82u l=0.6u
X3215 vdd tune_shunt[6] a_16500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X3216 vss cap_shunt_n a_9856_39268# vss nmos_6p0 w=0.82u l=0.6u
X3217 vdd a_28236_48983# a_28148_49080# vdd pmos_6p0 w=1.22u l=1u
X3218 a_26444_46280# a_26356_46324# vss vss nmos_6p0 w=0.82u l=1u
X3219 vdd tune_series_gy[3] a_11612_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3220 a_34748_48376# cap_shunt_gyp a_34480_48438# vss nmos_6p0 w=0.82u l=0.6u
X3221 a_29700_34626# cap_shunt_p a_30632_34564# vss nmos_6p0 w=0.82u l=0.6u
X3222 vdd a_3036_24328# a_2948_24372# vdd pmos_6p0 w=1.22u l=1u
X3223 a_13796_48738# cap_shunt_n a_13588_49084# vdd pmos_6p0 w=1.2u l=0.5u
X3224 vdd a_38092_30600# a_38004_30644# vdd pmos_6p0 w=1.22u l=1u
X3225 a_20532_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3226 a_13564_55255# a_13476_55352# vss vss nmos_6p0 w=0.82u l=1u
X3227 a_6532_47892# cap_shunt_p a_6740_48376# vdd pmos_6p0 w=1.2u l=0.5u
X3228 a_1716_6748# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3229 vss tune_shunt[6] a_6740_40536# vss nmos_6p0 w=0.51u l=0.6u
X3230 a_35880_13396# cap_series_gygyn a_35692_13396# vdd pmos_6p0 w=1.2u l=0.5u
X3231 vss tune_shunt[4] a_2708_14242# vss nmos_6p0 w=0.51u l=0.6u
X3232 a_9876_21720# cap_shunt_p a_9668_21236# vdd pmos_6p0 w=1.2u l=0.5u
X3233 a_21540_11452# cap_series_gyn a_21748_11106# vdd pmos_6p0 w=1.2u l=0.5u
X3234 a_21748_9538# cap_series_gyp a_23464_9476# vss nmos_6p0 w=0.82u l=0.6u
X3235 a_21540_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3236 vss tune_shunt[6] a_2708_37762# vss nmos_6p0 w=0.51u l=0.6u
X3237 a_29700_31490# cap_shunt_p a_30632_31428# vss nmos_6p0 w=0.82u l=0.6u
X3238 a_34516_23650# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3239 vdd a_3036_21192# a_2948_21236# vdd pmos_6p0 w=1.22u l=1u
X3240 a_10660_4834# cap_series_gyp a_10452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X3241 a_20284_53687# a_20196_53784# vss vss nmos_6p0 w=0.82u l=1u
X3242 a_7616_51812# cap_shunt_p a_6292_51874# vss nmos_6p0 w=0.82u l=0.6u
X3243 a_6532_44756# cap_shunt_p a_6740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X3244 vss tune_series_gygy[3] a_34536_9884# vss nmos_6p0 w=0.51u l=0.6u
X3245 a_5948_11784# a_5860_11828# vss vss nmos_6p0 w=0.82u l=1u
X3246 a_25780_40536# cap_shunt_n a_25572_40052# vdd pmos_6p0 w=1.2u l=0.5u
X3247 vss tune_shunt[3] a_2708_11106# vss nmos_6p0 w=0.51u l=0.6u
X3248 a_20720_12612# cap_series_gyn a_18612_12674# vss nmos_6p0 w=0.82u l=0.6u
X3249 a_22680_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X3250 a_25780_4472# cap_shunt_p a_25572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3251 a_34308_17724# cap_series_gygyn a_34516_17378# vdd pmos_6p0 w=1.2u l=0.5u
X3252 a_20172_39575# a_20084_39672# vss vss nmos_6p0 w=0.82u l=1u
X3253 vss tune_shunt[6] a_2708_34626# vss nmos_6p0 w=0.51u l=0.6u
X3254 vss cap_shunt_n a_23072_29860# vss nmos_6p0 w=0.82u l=0.6u
X3255 a_34516_20514# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3256 a_21748_6402# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3257 vdd a_14012_8215# a_13924_8312# vdd pmos_6p0 w=1.22u l=1u
X3258 a_10340_24372# cap_shunt_n a_10548_24856# vdd pmos_6p0 w=1.2u l=0.5u
X3259 a_21540_9884# cap_series_gyp a_21748_9538# vdd pmos_6p0 w=1.2u l=0.5u
X3260 a_33052_52119# a_32964_52216# vss vss nmos_6p0 w=0.82u l=1u
X3261 a_19936_18584# cap_shunt_p a_17828_18584# vss nmos_6p0 w=0.82u l=0.6u
X3262 a_14580_40536# cap_shunt_n a_14372_40052# vdd pmos_6p0 w=1.2u l=0.5u
X3263 a_34536_8316# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X3264 vdd a_6956_33303# a_6868_33400# vdd pmos_6p0 w=1.22u l=1u
X3265 a_3620_32212# cap_shunt_p a_3828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X3266 vss cap_shunt_n a_23072_26724# vss nmos_6p0 w=0.82u l=0.6u
X3267 a_6532_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3268 a_21540_6748# cap_series_gyn a_21748_6402# vdd pmos_6p0 w=1.2u l=0.5u
X3269 vss cap_series_gygyp a_35736_6340# vss nmos_6p0 w=0.82u l=0.6u
X3270 a_35692_18100# cap_series_gygyn a_35880_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3271 a_28692_18584# cap_series_gyp a_30408_18584# vss nmos_6p0 w=0.82u l=0.6u
X3272 vss tune_shunt[4] a_33732_34264# vss nmos_6p0 w=0.51u l=0.6u
X3273 a_6572_3988# cap_series_gyp a_6760_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3274 a_19936_15448# cap_shunt_p a_17828_15448# vss nmos_6p0 w=0.82u l=0.6u
X3275 a_34516_15810# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3276 vss cap_shunt_p a_11984_17016# vss nmos_6p0 w=0.82u l=0.6u
X3277 vss cap_shunt_p a_8848_13880# vss nmos_6p0 w=0.82u l=0.6u
X3278 a_20740_15448# cap_series_gyn a_20532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X3279 vdd a_1692_18056# a_1604_18100# vdd pmos_6p0 w=1.22u l=1u
X3280 a_2140_34871# a_2052_34968# vss vss nmos_6p0 w=0.82u l=1u
X3281 a_18724_6040# cap_series_gyn a_19656_6040# vss nmos_6p0 w=0.82u l=0.6u
X3282 a_1716_8316# cap_shunt_n a_1924_7970# vdd pmos_6p0 w=1.2u l=0.5u
X3283 a_3640_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3284 a_11200_18584# cap_shunt_p a_9876_18584# vss nmos_6p0 w=0.82u l=0.6u
X3285 a_24660_39330# cap_shunt_p a_24452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X3286 a_28692_9176# cap_series_gyn a_28484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X3287 a_6532_11828# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3288 a_3172_49460# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3289 vss tune_shunt[7] a_10548_35832# vss nmos_6p0 w=0.51u l=0.6u
X3290 a_18612_9538# cap_series_gyp a_18404_9884# vdd pmos_6p0 w=1.2u l=0.5u
X3291 a_28692_15448# cap_series_gyn a_30408_15448# vss nmos_6p0 w=0.82u l=0.6u
X3292 a_37280_45302# cap_shunt_gyp a_37280_44757# vdd pmos_6p0 w=1.215u l=0.5u
X3293 vss tune_shunt[4] a_33732_31128# vss nmos_6p0 w=0.51u l=0.6u
X3294 a_16708_18946# cap_shunt_p a_17640_18884# vss nmos_6p0 w=0.82u l=0.6u
X3295 vdd a_35292_55255# a_35204_55352# vdd pmos_6p0 w=1.22u l=1u
X3296 a_2140_31735# a_2052_31832# vss vss nmos_6p0 w=0.82u l=1u
X3297 a_2932_12312# cap_shunt_n a_2724_11828# vdd pmos_6p0 w=1.2u l=0.5u
X3298 vss tune_series_gy[5] a_24660_12674# vss nmos_6p0 w=0.51u l=0.6u
X3299 vdd a_16028_36872# a_15940_36916# vdd pmos_6p0 w=1.22u l=1u
X3300 a_29580_50984# a_29492_51028# vss vss nmos_6p0 w=0.82u l=1u
X3301 a_11800_8692# cap_series_gyp a_11612_8692# vdd pmos_6p0 w=1.2u l=0.5u
X3302 a_11200_15448# cap_shunt_p a_9876_15448# vss nmos_6p0 w=0.82u l=0.6u
X3303 a_13788_52552# a_13700_52596# vss vss nmos_6p0 w=0.82u l=1u
X3304 vdd tune_shunt[5] a_29492_38108# vdd pmos_6p0 w=1.2u l=0.5u
X3305 a_28692_6040# cap_shunt_n a_28484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X3306 a_18612_6402# cap_series_gyn a_18404_6748# vdd pmos_6p0 w=1.2u l=0.5u
X3307 a_5612_52119# a_5524_52216# vss vss nmos_6p0 w=0.82u l=1u
X3308 a_16708_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3309 a_21748_26786# cap_shunt_n a_21540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X3310 a_16500_23996# cap_shunt_n a_16708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X3311 a_16708_15810# cap_shunt_p a_17640_15748# vss nmos_6p0 w=0.82u l=0.6u
X3312 a_23240_4472# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X3313 vdd a_35292_52119# a_35204_52216# vdd pmos_6p0 w=1.22u l=1u
X3314 a_22848_35832# cap_shunt_n a_20740_35832# vss nmos_6p0 w=0.82u l=0.6u
X3315 a_33500_53687# a_33412_53784# vss vss nmos_6p0 w=0.82u l=1u
X3316 a_29700_28354# cap_shunt_p a_30632_28292# vss nmos_6p0 w=0.82u l=0.6u
X3317 a_24660_20514# cap_shunt_p a_26376_20452# vss nmos_6p0 w=0.82u l=0.6u
X3318 vdd tune_shunt[7] a_25572_25940# vdd pmos_6p0 w=1.2u l=0.5u
X3319 a_11668_45240# cap_shunt_n a_11460_44756# vdd pmos_6p0 w=1.2u l=0.5u
X3320 a_17620_32212# cap_shunt_n a_17828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X3321 a_28124_6647# a_28036_6744# vss vss nmos_6p0 w=0.82u l=1u
X3322 vss tune_shunt[0] a_29700_4834# vss nmos_6p0 w=0.51u l=0.6u
X3323 a_24452_14588# cap_series_gyn a_24660_14242# vdd pmos_6p0 w=1.2u l=0.5u
X3324 vss tune_shunt[7] a_6740_34264# vss nmos_6p0 w=0.51u l=0.6u
X3325 a_16708_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3326 vss cap_shunt_p a_4816_17316# vss nmos_6p0 w=0.82u l=0.6u
X3327 a_10548_35832# cap_shunt_n a_11480_35832# vss nmos_6p0 w=0.82u l=0.6u
X3328 a_33500_50551# a_33412_50648# vss vss nmos_6p0 w=0.82u l=1u
X3329 a_9668_49460# cap_shunt_p a_9876_49944# vdd pmos_6p0 w=1.2u l=0.5u
X3330 a_29700_25218# cap_shunt_p a_30632_25156# vss nmos_6p0 w=0.82u l=0.6u
X3331 a_11480_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X3332 vss cap_series_gyn a_27104_13880# vss nmos_6p0 w=0.82u l=0.6u
X3333 vdd a_12892_21192# a_12804_21236# vdd pmos_6p0 w=1.22u l=1u
X3334 a_9668_49460# cap_shunt_p a_9876_49944# vdd pmos_6p0 w=1.2u l=0.5u
X3335 a_7540_45948# cap_shunt_p a_7748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X3336 vdd tune_shunt[7] a_25572_22804# vdd pmos_6p0 w=1.2u l=0.5u
X3337 a_6532_38484# cap_shunt_n a_6740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X3338 a_31436_6748# tune_series_gygy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3339 vss cap_series_gygyn a_36296_6040# vss nmos_6p0 w=0.82u l=0.6u
X3340 vss tune_series_gygy[5] a_30616_21236# vss nmos_6p0 w=0.51u l=0.6u
X3341 vss tune_shunt[7] a_6740_31128# vss nmos_6p0 w=0.51u l=0.6u
X3342 a_29700_28354# cap_shunt_p a_29492_28700# vdd pmos_6p0 w=1.2u l=0.5u
X3343 vdd a_7852_55255# a_7764_55352# vdd pmos_6p0 w=1.22u l=1u
X3344 a_24660_42466# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3345 vss tune_shunt[7] a_2708_28354# vss nmos_6p0 w=0.51u l=0.6u
X3346 vss cap_series_gyn a_27104_10744# vss nmos_6p0 w=0.82u l=0.6u
X3347 vdd a_24204_53687# a_24116_53784# vdd pmos_6p0 w=1.22u l=1u
X3348 vdd tune_shunt[6] a_16500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X3349 a_6532_35348# cap_shunt_n a_6740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X3350 a_10452_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3351 a_7748_23650# cap_shunt_p a_7540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X3352 a_7580_8316# cap_series_gyn a_7768_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3353 a_23072_45540# cap_shunt_p a_21748_45602# vss nmos_6p0 w=0.82u l=0.6u
X3354 vss cap_series_gygyn a_32040_20452# vss nmos_6p0 w=0.82u l=0.6u
X3355 a_29492_36540# cap_shunt_n a_29700_36194# vdd pmos_6p0 w=1.2u l=0.5u
X3356 vdd a_4828_55255# a_4740_55352# vdd pmos_6p0 w=1.22u l=1u
X3357 vdd a_24204_50551# a_24116_50648# vdd pmos_6p0 w=1.22u l=1u
X3358 a_11460_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3359 a_36300_33736# a_36212_33780# vss vss nmos_6p0 w=0.82u l=1u
X3360 vss tune_shunt[7] a_2708_25218# vss nmos_6p0 w=0.51u l=0.6u
X3361 vdd tune_shunt[6] a_16500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X3362 a_28484_25940# cap_shunt_p a_28692_26424# vdd pmos_6p0 w=1.2u l=0.5u
X3363 a_1716_3612# cap_shunt_n a_1924_3266# vdd pmos_6p0 w=1.2u l=0.5u
X3364 a_33052_42711# a_32964_42808# vss vss nmos_6p0 w=0.82u l=1u
X3365 a_10452_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3366 a_35692_10260# cap_series_gygyp a_35880_10260# vdd pmos_6p0 w=1.2u l=0.5u
X3367 a_30924_54120# a_30836_54164# vss vss nmos_6p0 w=0.82u l=1u
X3368 a_36624_22020# cap_series_gygyp a_34516_22082# vss nmos_6p0 w=0.82u l=0.6u
X3369 a_34144_47512# cap_shunt_gyp a_34144_47108# vdd pmos_6p0 w=1.215u l=0.5u
X3370 a_23072_42404# cap_shunt_n a_21748_42466# vss nmos_6p0 w=0.82u l=0.6u
X3371 a_29492_33404# cap_shunt_p a_29700_33058# vdd pmos_6p0 w=1.2u l=0.5u
X3372 a_2140_28599# a_2052_28696# vss vss nmos_6p0 w=0.82u l=1u
X3373 a_35880_25940# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3374 a_12608_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X3375 a_3640_14180# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3376 vdd a_4828_52119# a_4740_52216# vdd pmos_6p0 w=1.22u l=1u
X3377 vss cap_series_gyp a_17808_6340# vss nmos_6p0 w=0.82u l=0.6u
X3378 vdd a_23756_14920# a_23668_14964# vdd pmos_6p0 w=1.22u l=1u
X3379 vss tune_series_gy[5] a_24660_15810# vss nmos_6p0 w=0.51u l=0.6u
X3380 a_37548_43672# cap_shunt_gyp a_37280_43734# vss nmos_6p0 w=0.82u l=0.6u
X3381 a_36300_30600# a_36212_30644# vss vss nmos_6p0 w=0.82u l=1u
X3382 a_35880_13396# cap_series_gygyn a_35692_13396# vdd pmos_6p0 w=1.2u l=0.5u
X3383 vss cap_shunt_p a_23072_17316# vss nmos_6p0 w=0.82u l=0.6u
X3384 a_19836_49416# a_19748_49460# vss vss nmos_6p0 w=0.82u l=1u
X3385 a_6740_42104# cap_shunt_n a_6532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X3386 a_28484_22804# cap_shunt_p a_28692_23288# vdd pmos_6p0 w=1.2u l=0.5u
X3387 a_15120_50244# cap_shunt_p a_13796_50306# vss nmos_6p0 w=0.82u l=0.6u
X3388 vss tune_shunt[7] a_10548_29560# vss nmos_6p0 w=0.51u l=0.6u
X3389 a_22436_7124# cap_series_gyp a_22644_7608# vdd pmos_6p0 w=1.2u l=0.5u
X3390 a_25780_7608# cap_series_gyn a_25572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3391 a_9876_21720# cap_shunt_p a_9668_21236# vdd pmos_6p0 w=1.2u l=0.5u
X3392 vss tune_shunt[5] a_28692_32696# vss nmos_6p0 w=0.51u l=0.6u
X3393 a_15700_7970# cap_series_gyn a_15492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3394 vdd a_32716_9783# a_32628_9880# vdd pmos_6p0 w=1.22u l=1u
X3395 a_2140_25463# a_2052_25560# vss vss nmos_6p0 w=0.82u l=1u
X3396 a_3640_11044# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3397 vdd a_35628_14487# a_35540_14584# vdd pmos_6p0 w=1.22u l=1u
X3398 a_30476_49416# a_30388_49460# vss vss nmos_6p0 w=0.82u l=1u
X3399 a_29580_44712# a_29492_44756# vss vss nmos_6p0 w=0.82u l=1u
X3400 a_33524_33780# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3401 a_25780_40536# cap_shunt_n a_25572_40052# vdd pmos_6p0 w=1.2u l=0.5u
X3402 a_7672_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3403 vss tune_shunt[7] a_10548_26424# vss nmos_6p0 w=0.51u l=0.6u
X3404 a_5612_45847# a_5524_45944# vss vss nmos_6p0 w=0.82u l=1u
X3405 vss tune_shunt[6] a_7748_37762# vss nmos_6p0 w=0.51u l=0.6u
X3406 a_3828_37400# cap_shunt_n a_3620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X3407 vdd tune_shunt[6] a_6532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X3408 vss cap_series_gygyn a_32040_7908# vss nmos_6p0 w=0.82u l=0.6u
X3409 a_34308_17724# cap_series_gygyn a_34516_17378# vdd pmos_6p0 w=1.2u l=0.5u
X3410 a_31032_21720# cap_series_gygyn a_30616_21236# vss nmos_6p0 w=0.82u l=0.6u
X3411 vdd a_22860_47415# a_22772_47512# vdd pmos_6p0 w=1.22u l=1u
X3412 vdd tune_series_gy[3] a_15492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X3413 a_13796_50306# cap_shunt_p a_13588_50652# vdd pmos_6p0 w=1.2u l=0.5u
X3414 vdd a_16028_27464# a_15940_27508# vdd pmos_6p0 w=1.22u l=1u
X3415 vdd a_35628_11351# a_35540_11448# vdd pmos_6p0 w=1.22u l=1u
X3416 a_30476_46280# a_30388_46324# vss vss nmos_6p0 w=0.82u l=1u
X3417 vss tune_shunt[6] a_17828_45240# vss nmos_6p0 w=0.51u l=0.6u
X3418 a_33524_30644# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3419 a_22848_29560# cap_shunt_n a_20740_29560# vss nmos_6p0 w=0.82u l=0.6u
X3420 vdd tune_shunt[5] a_8996_52220# vdd pmos_6p0 w=1.2u l=0.5u
X3421 a_14580_40536# cap_shunt_n a_14372_40052# vdd pmos_6p0 w=1.2u l=0.5u
X3422 vdd a_36076_34871# a_35988_34968# vdd pmos_6p0 w=1.22u l=1u
X3423 a_24660_14242# cap_series_gyn a_26376_14180# vss nmos_6p0 w=0.82u l=0.6u
X3424 vdd a_23532_47848# a_23444_47892# vdd pmos_6p0 w=1.22u l=1u
X3425 a_7672_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3426 a_5612_42711# a_5524_42808# vss vss nmos_6p0 w=0.82u l=1u
X3427 vss tune_shunt[7] a_7748_34626# vss nmos_6p0 w=0.51u l=0.6u
X3428 a_7748_33058# cap_shunt_n a_8680_32996# vss nmos_6p0 w=0.82u l=0.6u
X3429 a_16500_14588# cap_shunt_p a_16708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X3430 vdd a_28348_19624# a_28260_19668# vdd pmos_6p0 w=1.22u l=1u
X3431 a_7748_45602# cap_shunt_p a_9464_45540# vss nmos_6p0 w=0.82u l=0.6u
X3432 vss tune_shunt[6] a_17828_42104# vss nmos_6p0 w=0.51u l=0.6u
X3433 a_10548_29560# cap_shunt_n a_11480_29560# vss nmos_6p0 w=0.82u l=0.6u
X3434 a_22848_26424# cap_shunt_n a_20740_26424# vss nmos_6p0 w=0.82u l=0.6u
X3435 vdd a_35292_7080# a_35204_7124# vdd pmos_6p0 w=1.22u l=1u
X3436 a_7540_39676# cap_shunt_n a_7748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X3437 a_24660_11106# cap_series_gyp a_26376_11044# vss nmos_6p0 w=0.82u l=0.6u
X3438 a_20740_15448# cap_series_gyn a_20532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X3439 vdd tune_series_gy[5] a_25572_16532# vdd pmos_6p0 w=1.2u l=0.5u
X3440 vdd a_19724_31735# a_19636_31832# vdd pmos_6p0 w=1.22u l=1u
X3441 a_6740_21720# cap_shunt_p a_7672_21720# vss nmos_6p0 w=0.82u l=0.6u
X3442 a_20832_6040# cap_series_gyn a_18724_6040# vss nmos_6p0 w=0.82u l=0.6u
X3443 a_26444_52119# a_26356_52216# vss vss nmos_6p0 w=0.82u l=1u
X3444 a_15512_48676# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3445 a_16708_45602# cap_shunt_p a_16500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X3446 a_25572_43188# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3447 a_6956_8215# a_6868_8312# vss vss nmos_6p0 w=0.82u l=1u
X3448 vss tune_shunt[6] a_6740_48376# vss nmos_6p0 w=0.51u l=0.6u
X3449 a_7748_42466# cap_shunt_n a_9464_42404# vss nmos_6p0 w=0.82u l=0.6u
X3450 a_24660_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3451 a_10548_26424# cap_shunt_n a_11480_26424# vss nmos_6p0 w=0.82u l=0.6u
X3452 vss tune_shunt[4] a_32612_36194# vss nmos_6p0 w=0.51u l=0.6u
X3453 vdd tune_shunt[2] a_1716_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3454 a_6760_3988# cap_series_gyp a_6572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3455 a_16500_17724# cap_shunt_p a_16708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X3456 a_36428_45240# cap_shunt_gyn a_36160_45302# vss nmos_6p0 w=0.82u l=0.6u
X3457 vdd a_6060_41143# a_5972_41240# vdd pmos_6p0 w=1.22u l=1u
X3458 a_6532_29076# cap_shunt_n a_6740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X3459 vdd tune_shunt[6] a_9108_50652# vdd pmos_6p0 w=1.2u l=0.5u
X3460 a_8680_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3461 a_14372_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3462 vdd tune_shunt[4] a_21540_17724# vdd pmos_6p0 w=1.2u l=0.5u
X3463 a_24660_33058# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3464 a_32268_23895# a_32180_23992# vss vss nmos_6p0 w=0.82u l=1u
X3465 a_35344_6340# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X3466 a_16500_23996# cap_shunt_n a_16708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X3467 a_20620_38007# a_20532_38104# vss vss nmos_6p0 w=0.82u l=1u
X3468 vss tune_shunt[4] a_32612_33058# vss nmos_6p0 w=0.51u l=0.6u
X3469 a_33500_5512# a_33412_5556# vss vss nmos_6p0 w=0.82u l=1u
X3470 a_9668_10260# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3471 a_30924_47848# a_30836_47892# vss vss nmos_6p0 w=0.82u l=1u
X3472 a_8680_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3473 a_16708_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3474 a_23072_36132# cap_shunt_n a_21748_36194# vss nmos_6p0 w=0.82u l=0.6u
X3475 vss tune_shunt[6] a_28692_35832# vss nmos_6p0 w=0.51u l=0.6u
X3476 a_16476_33736# a_16388_33780# vss vss nmos_6p0 w=0.82u l=1u
X3477 a_29492_27132# cap_shunt_p a_29700_26786# vdd pmos_6p0 w=1.2u l=0.5u
X3478 vss tune_series_gy[4] a_24660_9538# vss nmos_6p0 w=0.51u l=0.6u
X3479 a_31260_11784# a_31172_11828# vss vss nmos_6p0 w=0.82u l=1u
X3480 vss tune_shunt[5] a_6292_17016# vss nmos_6p0 w=0.51u l=0.6u
X3481 vdd a_28684_55255# a_28596_55352# vdd pmos_6p0 w=1.22u l=1u
X3482 a_11480_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3483 a_6292_18584# cap_shunt_p a_6084_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3484 a_28484_16532# cap_series_gyn a_28692_17016# vdd pmos_6p0 w=1.2u l=0.5u
X3485 a_5936_13880# cap_shunt_n a_3828_13880# vss nmos_6p0 w=0.82u l=0.6u
X3486 a_37868_12919# a_37780_13016# vss vss nmos_6p0 w=0.82u l=1u
X3487 a_31624_22428# cap_series_gygyn a_31436_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3488 a_16476_30600# a_16388_30644# vss vss nmos_6p0 w=0.82u l=1u
X3489 a_5636_11452# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3490 a_19544_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3491 a_19732_12312# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3492 a_35880_16532# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3493 vdd a_28684_52119# a_28596_52216# vdd pmos_6p0 w=1.22u l=1u
X3494 a_24660_7970# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3495 a_30812_55255# a_30724_55352# vss vss nmos_6p0 w=0.82u l=1u
X3496 a_6740_32696# cap_shunt_n a_6532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X3497 vdd a_12108_16055# a_12020_16152# vdd pmos_6p0 w=1.22u l=1u
X3498 a_14728_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3499 vss cap_series_gyn a_30800_9176# vss nmos_6p0 w=0.82u l=0.6u
X3500 vss tune_shunt[4] a_28692_23288# vss nmos_6p0 w=0.51u l=0.6u
X3501 a_11488_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X3502 a_10492_8316# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3503 a_13564_9783# a_13476_9880# vss vss nmos_6p0 w=0.82u l=1u
X3504 a_13796_44034# cap_shunt_n a_13588_44380# vdd pmos_6p0 w=1.2u l=0.5u
X3505 vss cap_shunt_n a_35056_34264# vss nmos_6p0 w=0.82u l=0.6u
X3506 a_8456_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3507 a_18612_9538# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3508 a_24660_4834# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X3509 vdd tune_shunt[7] a_9332_11452# vdd pmos_6p0 w=1.2u l=0.5u
X3510 vdd a_12108_12919# a_12020_13016# vdd pmos_6p0 w=1.22u l=1u
X3511 vdd a_36076_28599# a_35988_28696# vdd pmos_6p0 w=1.22u l=1u
X3512 a_14728_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3513 a_29492_36540# cap_shunt_n a_29700_36194# vdd pmos_6p0 w=1.2u l=0.5u
X3514 a_24660_29922# cap_shunt_n a_25592_29860# vss nmos_6p0 w=0.82u l=0.6u
X3515 vss tune_shunt[7] a_7748_28354# vss nmos_6p0 w=0.51u l=0.6u
X3516 a_3828_27992# cap_shunt_n a_3620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X3517 a_5612_36439# a_5524_36536# vss vss nmos_6p0 w=0.82u l=1u
X3518 a_21540_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3519 vdd tune_shunt[7] a_6532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X3520 a_13796_40898# cap_shunt_n a_13588_41244# vdd pmos_6p0 w=1.2u l=0.5u
X3521 vss cap_shunt_n a_35056_31128# vss nmos_6p0 w=0.82u l=0.6u
X3522 a_33936_29860# cap_shunt_p a_32612_29922# vss nmos_6p0 w=0.82u l=0.6u
X3523 a_8456_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3524 vdd tune_series_gy[4] a_14484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3525 vdd a_31260_53687# a_31172_53784# vdd pmos_6p0 w=1.22u l=1u
X3526 vdd a_19724_25463# a_19636_25560# vdd pmos_6p0 w=1.22u l=1u
X3527 a_2708_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3528 a_29492_33404# cap_shunt_p a_29700_33058# vdd pmos_6p0 w=1.2u l=0.5u
X3529 a_24660_26786# cap_shunt_p a_25592_26724# vss nmos_6p0 w=0.82u l=0.6u
X3530 vss tune_shunt[7] a_7748_25218# vss nmos_6p0 w=0.51u l=0.6u
X3531 a_7748_23650# cap_shunt_p a_8680_23588# vss nmos_6p0 w=0.82u l=0.6u
X3532 vdd a_31708_38440# a_31620_38484# vdd pmos_6p0 w=1.22u l=1u
X3533 a_21540_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3534 a_35040_45302# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3535 a_33936_26724# cap_shunt_p a_32612_26786# vss nmos_6p0 w=0.82u l=0.6u
X3536 a_16708_39330# cap_shunt_n a_16500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X3537 a_12788_17016# cap_shunt_p a_14504_17016# vss nmos_6p0 w=0.82u l=0.6u
X3538 a_7748_36194# cap_shunt_n a_9464_36132# vss nmos_6p0 w=0.82u l=0.6u
X3539 a_22848_17016# cap_shunt_p a_20740_17016# vss nmos_6p0 w=0.82u l=0.6u
X3540 a_9876_21720# cap_shunt_p a_9668_21236# vdd pmos_6p0 w=1.2u l=0.5u
X3541 vdd a_31260_50551# a_31172_50648# vdd pmos_6p0 w=1.22u l=1u
X3542 a_2500_17724# cap_shunt_p a_2708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X3543 a_6084_51028# cap_shunt_p a_6292_51512# vdd pmos_6p0 w=1.2u l=0.5u
X3544 a_28692_34264# cap_shunt_p a_28484_33780# vdd pmos_6p0 w=1.2u l=0.5u
X3545 a_2708_20514# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3546 vdd a_19724_22327# a_19636_22424# vdd pmos_6p0 w=1.22u l=1u
X3547 a_21748_12674# cap_series_gyn a_21540_13020# vdd pmos_6p0 w=1.2u l=0.5u
X3548 a_24652_21192# a_24564_21236# vss vss nmos_6p0 w=0.82u l=1u
X3549 a_17620_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3550 vdd a_31708_35304# a_31620_35348# vdd pmos_6p0 w=1.22u l=1u
X3551 a_6740_12312# cap_shunt_p a_7672_12312# vss nmos_6p0 w=0.82u l=0.6u
X3552 a_13460_37400# cap_shunt_n a_13252_36916# vdd pmos_6p0 w=1.2u l=0.5u
X3553 a_29700_11106# cap_series_gyp a_29492_11452# vdd pmos_6p0 w=1.2u l=0.5u
X3554 vss tune_shunt[7] a_6628_12674# vss nmos_6p0 w=0.51u l=0.6u
X3555 a_6084_19292# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3556 a_15512_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3557 a_27104_20152# cap_series_gyp a_25780_20152# vss nmos_6p0 w=0.82u l=0.6u
X3558 a_9316_48738# cap_shunt_p a_10248_48676# vss nmos_6p0 w=0.82u l=0.6u
X3559 vdd a_28348_45847# a_28260_45944# vdd pmos_6p0 w=1.22u l=1u
X3560 a_7792_6340# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X3561 a_8996_52220# cap_shunt_n a_9204_51874# vdd pmos_6p0 w=1.2u l=0.5u
X3562 a_26892_49416# a_26804_49460# vss vss nmos_6p0 w=0.82u l=1u
X3563 vdd a_34396_41576# a_34308_41620# vdd pmos_6p0 w=1.22u l=1u
X3564 vdd a_30364_22327# a_30276_22424# vdd pmos_6p0 w=1.22u l=1u
X3565 vss cap_shunt_n a_4032_7908# vss nmos_6p0 w=0.82u l=0.6u
X3566 a_1692_12919# a_1604_13016# vss vss nmos_6p0 w=0.82u l=1u
X3567 a_7540_34972# cap_shunt_n a_7748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X3568 a_28692_31128# cap_shunt_n a_28484_30644# vdd pmos_6p0 w=1.2u l=0.5u
X3569 a_13796_50306# cap_shunt_p a_13588_50652# vdd pmos_6p0 w=1.2u l=0.5u
X3570 vdd a_4380_52552# a_4292_52596# vdd pmos_6p0 w=1.22u l=1u
X3571 a_6532_47892# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3572 a_8680_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3573 a_6292_51874# cap_shunt_p a_6084_52220# vdd pmos_6p0 w=1.2u l=0.5u
X3574 a_6084_16156# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3575 vdd tune_shunt[5] a_8996_52220# vdd pmos_6p0 w=1.2u l=0.5u
X3576 vdd a_19276_17623# a_19188_17720# vdd pmos_6p0 w=1.22u l=1u
X3577 a_31624_19292# cap_series_gygyn a_31436_19292# vdd pmos_6p0 w=1.2u l=0.5u
X3578 a_6740_53080# cap_shunt_n a_6532_52596# vdd pmos_6p0 w=1.2u l=0.5u
X3579 vss tune_shunt[7] a_28692_29560# vss nmos_6p0 w=0.51u l=0.6u
X3580 a_26892_46280# a_26804_46324# vss vss nmos_6p0 w=0.82u l=1u
X3581 a_13796_18946# cap_shunt_p a_15512_18884# vss nmos_6p0 w=0.82u l=0.6u
X3582 vdd a_28236_54120# a_28148_54164# vdd pmos_6p0 w=1.22u l=1u
X3583 vdd a_28684_48983# a_28596_49080# vdd pmos_6p0 w=1.22u l=1u
X3584 a_7540_31836# cap_shunt_n a_7748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X3585 a_33948_13352# a_33860_13396# vss vss nmos_6p0 w=0.82u l=1u
X3586 a_16500_14588# cap_shunt_p a_16708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X3587 a_23856_18884# cap_shunt_p a_21748_18946# vss nmos_6p0 w=0.82u l=0.6u
X3588 a_23868_49416# a_23780_49460# vss vss nmos_6p0 w=0.82u l=1u
X3589 a_37280_43189# cap_shunt_gyp a_37280_43734# vdd pmos_6p0 w=1.215u l=0.5u
X3590 a_3620_14964# cap_shunt_p a_3828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X3591 a_6532_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3592 a_8680_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3593 vss tune_shunt[7] a_9876_21720# vss nmos_6p0 w=0.51u l=0.6u
X3594 vdd tune_shunt[7] a_17620_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3595 vss tune_shunt[5] a_16708_47170# vss nmos_6p0 w=0.51u l=0.6u
X3596 a_20740_45240# cap_shunt_n a_20532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X3597 vss tune_shunt[7] a_28692_26424# vss nmos_6p0 w=0.51u l=0.6u
X3598 a_13796_15810# cap_shunt_p a_15512_15748# vss nmos_6p0 w=0.82u l=0.6u
X3599 a_35880_19668# cap_series_gygyp a_36688_20152# vss nmos_6p0 w=0.82u l=0.6u
X3600 vdd a_28236_50984# a_28148_51028# vdd pmos_6p0 w=1.22u l=1u
X3601 a_30812_48983# a_30724_49080# vss vss nmos_6p0 w=0.82u l=1u
X3602 a_33948_10216# a_33860_10260# vss vss nmos_6p0 w=0.82u l=1u
X3603 vss tune_series_gy[5] a_22644_13880# vss nmos_6p0 w=0.51u l=0.6u
X3604 a_23856_15748# cap_series_gyn a_21748_15810# vss nmos_6p0 w=0.82u l=0.6u
X3605 a_12788_49944# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3606 a_3864_10744# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3607 a_34516_22082# cap_series_gygyp a_34308_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3608 a_28692_13880# cap_series_gyp a_29624_13880# vss nmos_6p0 w=0.82u l=0.6u
X3609 a_5388_5512# a_5300_5556# vss vss nmos_6p0 w=0.82u l=1u
X3610 vss tune_shunt[6] a_16708_44034# vss nmos_6p0 w=0.51u l=0.6u
X3611 a_21540_9884# cap_series_gyp a_21748_9538# vdd pmos_6p0 w=1.2u l=0.5u
X3612 a_10988_55255# a_10900_55352# vss vss nmos_6p0 w=0.82u l=1u
X3613 a_29492_11452# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3614 a_36188_55255# a_36100_55352# vss vss nmos_6p0 w=0.82u l=1u
X3615 vss cap_shunt_n a_5936_38968# vss nmos_6p0 w=0.82u l=0.6u
X3616 a_14692_10744# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3617 a_6292_48738# cap_shunt_p a_8008_48676# vss nmos_6p0 w=0.82u l=0.6u
X3618 vss tune_series_gy[5] a_22644_10744# vss nmos_6p0 w=0.51u l=0.6u
X3619 a_28692_10744# cap_series_gyp a_29624_10744# vss nmos_6p0 w=0.82u l=0.6u
X3620 a_19936_11044# cap_series_gyn a_18612_11106# vss nmos_6p0 w=0.82u l=0.6u
X3621 a_17828_46808# cap_shunt_n a_19544_46808# vss nmos_6p0 w=0.82u l=0.6u
X3622 vss cap_series_gyn a_30016_12312# vss nmos_6p0 w=0.82u l=0.6u
X3623 a_21540_6748# cap_series_gyn a_21748_6402# vdd pmos_6p0 w=1.2u l=0.5u
X3624 vss cap_shunt_n a_15120_43972# vss nmos_6p0 w=0.82u l=0.6u
X3625 a_19836_52119# a_19748_52216# vss vss nmos_6p0 w=0.82u l=1u
X3626 a_6740_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3627 a_20740_27992# cap_shunt_n a_21672_27992# vss nmos_6p0 w=0.82u l=0.6u
X3628 a_30588_41576# a_30500_41620# vss vss nmos_6p0 w=0.82u l=1u
X3629 a_29492_27132# cap_shunt_p a_29700_26786# vdd pmos_6p0 w=1.2u l=0.5u
X3630 a_29468_8215# a_29380_8312# vss vss nmos_6p0 w=0.82u l=1u
X3631 a_21540_25564# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3632 a_30428_19668# cap_series_gygyn a_30616_19668# vdd pmos_6p0 w=1.2u l=0.5u
X3633 a_16688_46808# cap_shunt_p a_14580_46808# vss nmos_6p0 w=0.82u l=0.6u
X3634 a_6292_18584# cap_shunt_p a_6084_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3635 a_9876_51512# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3636 vdd a_34844_40008# a_34756_40052# vdd pmos_6p0 w=1.22u l=1u
X3637 a_29492_23996# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3638 vss cap_series_gyn a_13104_6040# vss nmos_6p0 w=0.82u l=0.6u
X3639 a_8456_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3640 vss cap_shunt_n a_15120_40836# vss nmos_6p0 w=0.82u l=0.6u
X3641 a_13460_38968# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3642 vdd a_31260_44279# a_31172_44376# vdd pmos_6p0 w=1.22u l=1u
X3643 a_6740_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3644 a_20740_24856# cap_shunt_n a_21672_24856# vss nmos_6p0 w=0.82u l=0.6u
X3645 a_14908_6647# a_14820_6744# vss vss nmos_6p0 w=0.82u l=1u
X3646 vss cap_shunt_p a_19152_45240# vss nmos_6p0 w=0.82u l=0.6u
X3647 a_30920_12612# cap_series_gyn a_29720_13020# vss nmos_6p0 w=0.82u l=0.6u
X3648 a_2708_14242# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3649 vdd a_19724_16055# a_19636_16152# vdd pmos_6p0 w=1.22u l=1u
X3650 a_24660_17378# cap_series_gyp a_25592_17316# vss nmos_6p0 w=0.82u l=0.6u
X3651 a_2140_54120# a_2052_54164# vss vss nmos_6p0 w=0.82u l=1u
X3652 vdd a_31708_29032# a_31620_29076# vdd pmos_6p0 w=1.22u l=1u
X3653 vss tune_series_gygy[5] a_34516_23650# vss nmos_6p0 w=0.51u l=0.6u
X3654 a_21540_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3655 vdd tune_shunt[5] a_3172_51028# vdd pmos_6p0 w=1.2u l=0.5u
X3656 a_36384_47108# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3657 a_17828_40536# cap_shunt_n a_17620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X3658 a_19936_6340# cap_series_gyn a_18612_6402# vss nmos_6p0 w=0.82u l=0.6u
X3659 a_8748_55255# a_8660_55352# vss vss nmos_6p0 w=0.82u l=1u
X3660 vdd a_16476_36872# a_16388_36916# vdd pmos_6p0 w=1.22u l=1u
X3661 vss cap_shunt_n a_19152_42104# vss nmos_6p0 w=0.82u l=0.6u
X3662 a_10340_36916# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3663 a_28692_24856# cap_shunt_p a_28484_24372# vdd pmos_6p0 w=1.2u l=0.5u
X3664 a_2708_11106# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X3665 a_13796_44034# cap_shunt_n a_13588_44380# vdd pmos_6p0 w=1.2u l=0.5u
X3666 a_17620_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3667 vdd a_36300_27464# a_36212_27508# vdd pmos_6p0 w=1.22u l=1u
X3668 a_8680_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3669 vss tune_series_gygy[5] a_34516_20514# vss nmos_6p0 w=0.51u l=0.6u
X3670 a_16708_34626# cap_shunt_n a_16500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X3671 a_13460_27992# cap_shunt_n a_13252_27508# vdd pmos_6p0 w=1.2u l=0.5u
X3672 a_36232_23588# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X3673 vdd a_15804_49416# a_15716_49460# vdd pmos_6p0 w=1.22u l=1u
X3674 a_29492_36540# cap_shunt_n a_29700_36194# vdd pmos_6p0 w=1.2u l=0.5u
X3675 vss cap_shunt_p a_8064_48376# vss nmos_6p0 w=0.82u l=0.6u
X3676 a_18032_37700# cap_shunt_n a_16708_37762# vss nmos_6p0 w=0.82u l=0.6u
X3677 a_24452_28700# cap_shunt_n a_24660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X3678 a_7540_25564# cap_shunt_n a_7748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X3679 vdd a_27676_9783# a_27588_9880# vdd pmos_6p0 w=1.22u l=1u
X3680 a_13796_40898# cap_shunt_n a_13588_41244# vdd pmos_6p0 w=1.2u l=0.5u
X3681 a_4760_32696# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3682 vdd a_33948_3511# a_33860_3608# vdd pmos_6p0 w=1.22u l=1u
X3683 a_6532_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3684 vdd tune_series_gy[3] a_10492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3685 a_25780_20152# cap_series_gyp a_25572_19668# vdd pmos_6p0 w=1.2u l=0.5u
X3686 a_8680_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3687 a_11536_17316# cap_shunt_p a_9428_17378# vss nmos_6p0 w=0.82u l=0.6u
X3688 a_34516_18946# cap_series_gygyn a_34308_19292# vdd pmos_6p0 w=1.2u l=0.5u
X3689 a_5096_51512# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3690 a_16708_31490# cap_shunt_n a_16500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X3691 a_6740_43672# cap_shunt_p a_6532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X3692 a_20740_38968# cap_shunt_n a_20532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X3693 a_12788_15448# cap_shunt_p a_12580_14964# vdd pmos_6p0 w=1.2u l=0.5u
X3694 a_10808_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3695 a_29492_33404# cap_shunt_p a_29700_33058# vdd pmos_6p0 w=1.2u l=0.5u
X3696 vdd a_27676_6647# a_27588_6744# vdd pmos_6p0 w=1.22u l=1u
X3697 vss cap_series_gyn a_15792_3204# vss nmos_6p0 w=0.82u l=0.6u
X3698 vss cap_shunt_n a_18816_47108# vss nmos_6p0 w=0.82u l=0.6u
X3699 a_33292_43972# cap_shunt_gyn a_33024_43972# vss nmos_6p0 w=0.82u l=0.6u
X3700 a_6532_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3701 a_1924_7608# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X3702 vss tune_shunt[7] a_9876_12312# vss nmos_6p0 w=0.51u l=0.6u
X3703 a_34516_15810# cap_series_gygyn a_34308_16156# vdd pmos_6p0 w=1.2u l=0.5u
X3704 a_7748_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3705 a_6084_51028# cap_shunt_p a_6292_51512# vdd pmos_6p0 w=1.2u l=0.5u
X3706 a_2500_47516# cap_shunt_p a_2708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X3707 a_20740_35832# cap_shunt_n a_20532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X3708 a_28692_34264# cap_shunt_p a_28484_33780# vdd pmos_6p0 w=1.2u l=0.5u
X3709 a_7580_8316# cap_series_gyn a_7768_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3710 a_12788_12312# cap_shunt_p a_12580_11828# vdd pmos_6p0 w=1.2u l=0.5u
X3711 vss tune_series_gy[4] a_28692_17016# vss nmos_6p0 w=0.51u l=0.6u
X3712 a_21748_12674# cap_series_gyn a_21540_13020# vdd pmos_6p0 w=1.2u l=0.5u
X3713 a_18612_4472# cap_series_gyp a_18404_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3714 a_37444_33400# cap_shunt_gyp a_37632_33400# vdd pmos_6p0 w=1.215u l=0.5u
X3715 a_29700_11106# cap_series_gyp a_29492_11452# vdd pmos_6p0 w=1.2u l=0.5u
X3716 a_6084_19292# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3717 vdd a_24652_53687# a_24564_53784# vdd pmos_6p0 w=1.22u l=1u
X3718 a_13460_37400# cap_shunt_n a_13252_36916# vdd pmos_6p0 w=1.2u l=0.5u
X3719 vdd tune_shunt[7] a_13588_17724# vdd pmos_6p0 w=1.2u l=0.5u
X3720 vdd a_23308_33736# a_23220_33780# vdd pmos_6p0 w=1.22u l=1u
X3721 a_8996_52220# cap_shunt_n a_9204_51874# vdd pmos_6p0 w=1.2u l=0.5u
X3722 a_9108_47516# cap_shunt_p a_9316_47170# vdd pmos_6p0 w=1.2u l=0.5u
X3723 vdd a_16924_38440# a_16836_38484# vdd pmos_6p0 w=1.22u l=1u
X3724 a_25780_32696# cap_shunt_p a_27496_32696# vss nmos_6p0 w=0.82u l=0.6u
X3725 a_34396_24328# a_34308_24372# vss vss nmos_6p0 w=0.82u l=1u
X3726 vdd tune_shunt[7] a_6532_13396# vdd pmos_6p0 w=1.2u l=0.5u
X3727 a_28692_31128# cap_shunt_n a_28484_30644# vdd pmos_6p0 w=1.2u l=0.5u
X3728 vss cap_series_gyp a_23968_9176# vss nmos_6p0 w=0.82u l=0.6u
X3729 vdd a_34396_3944# a_34308_3988# vdd pmos_6p0 w=1.22u l=1u
X3730 a_3620_47892# cap_shunt_p a_3828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X3731 a_14692_6040# cap_series_gyn a_15624_6040# vss nmos_6p0 w=0.82u l=0.6u
X3732 a_6292_51874# cap_shunt_p a_6084_52220# vdd pmos_6p0 w=1.2u l=0.5u
X3733 a_15700_6402# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3734 a_6084_16156# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3735 vdd a_24652_50551# a_24564_50648# vdd pmos_6p0 w=1.22u l=1u
X3736 a_6404_47170# cap_shunt_p a_6196_47516# vdd pmos_6p0 w=1.2u l=0.5u
X3737 vss tune_shunt[6] a_9316_48738# vss nmos_6p0 w=0.51u l=0.6u
X3738 vdd a_23308_30600# a_23220_30644# vdd pmos_6p0 w=1.22u l=1u
X3739 a_21540_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3740 vdd a_16924_35304# a_16836_35348# vdd pmos_6p0 w=1.22u l=1u
X3741 a_28692_37400# cap_shunt_p a_28484_36916# vdd pmos_6p0 w=1.2u l=0.5u
X3742 a_3620_44756# cap_shunt_p a_3828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X3743 vss cap_shunt_n a_15120_34564# vss nmos_6p0 w=0.82u l=0.6u
X3744 a_30364_6647# a_30276_6744# vss vss nmos_6p0 w=0.82u l=1u
X3745 a_31624_6748# cap_series_gygyn a_32432_6340# vss nmos_6p0 w=0.82u l=0.6u
X3746 a_6740_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3747 a_4940_8215# a_4852_8312# vss vss nmos_6p0 w=0.82u l=1u
X3748 a_2724_8692# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3749 a_20740_18584# cap_shunt_p a_21672_18584# vss nmos_6p0 w=0.82u l=0.6u
X3750 vdd a_27228_38007# a_27140_38104# vdd pmos_6p0 w=1.22u l=1u
X3751 a_32156_36872# a_32068_36916# vss vss nmos_6p0 w=0.82u l=1u
X3752 vss tune_shunt[6] a_10660_42466# vss nmos_6p0 w=0.51u l=0.6u
X3753 a_2140_47848# a_2052_47892# vss vss nmos_6p0 w=0.82u l=1u
X3754 a_21748_39330# cap_shunt_p a_23464_39268# vss nmos_6p0 w=0.82u l=0.6u
X3755 a_21540_16156# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3756 a_34308_17724# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3757 a_9316_22082# cap_shunt_p a_9108_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3758 a_29492_14588# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3759 vss tune_shunt[5] a_6852_53442# vss nmos_6p0 w=0.51u l=0.6u
X3760 vss cap_shunt_n a_15120_31428# vss nmos_6p0 w=0.82u l=0.6u
X3761 a_34516_22082# cap_series_gygyp a_34308_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3762 vdd a_35292_54120# a_35204_54164# vdd pmos_6p0 w=1.22u l=1u
X3763 vss cap_shunt_n a_11984_51512# vss nmos_6p0 w=0.82u l=0.6u
X3764 a_6740_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3765 a_20740_15448# cap_series_gyn a_21672_15448# vss nmos_6p0 w=0.82u l=0.6u
X3766 a_31624_20860# cap_series_gygyn a_31436_20860# vdd pmos_6p0 w=1.2u l=0.5u
X3767 a_18424_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3768 vss cap_series_gyn a_11984_6340# vss nmos_6p0 w=0.82u l=0.6u
X3769 a_27228_19191# a_27140_19288# vss vss nmos_6p0 w=0.82u l=1u
X3770 vss tune_shunt[6] a_13796_40898# vss nmos_6p0 w=0.51u l=0.6u
X3771 a_2708_34626# cap_shunt_n a_2500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X3772 a_11460_43188# cap_shunt_n a_11668_43672# vdd pmos_6p0 w=1.2u l=0.5u
X3773 vdd a_9644_25896# a_9556_25940# vdd pmos_6p0 w=1.22u l=1u
X3774 a_1716_6748# cap_shunt_n a_1924_6402# vdd pmos_6p0 w=1.2u l=0.5u
X3775 a_32172_45540# cap_shunt_gyp a_31904_45540# vss nmos_6p0 w=0.82u l=0.6u
X3776 a_21748_22082# cap_shunt_p a_22680_22020# vss nmos_6p0 w=0.82u l=0.6u
X3777 vdd a_35292_50984# a_35204_51028# vdd pmos_6p0 w=1.22u l=1u
X3778 vdd a_16476_27464# a_16388_27508# vdd pmos_6p0 w=1.22u l=1u
X3779 vdd a_32268_54120# a_32180_54164# vdd pmos_6p0 w=1.22u l=1u
X3780 a_10340_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3781 a_34844_7080# a_34756_7124# vss vss nmos_6p0 w=0.82u l=1u
X3782 vdd tune_shunt[3] a_5636_9884# vdd pmos_6p0 w=1.2u l=0.5u
X3783 a_27228_16055# a_27140_16152# vss vss nmos_6p0 w=0.82u l=1u
X3784 a_37080_7608# cap_series_gygyp a_35880_7124# vss nmos_6p0 w=0.82u l=0.6u
X3785 a_18612_4472# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3786 a_35692_19668# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3787 vdd a_23980_47848# a_23892_47892# vdd pmos_6p0 w=1.22u l=1u
X3788 a_37444_40053# cap_shunt_gyn a_37632_40053# vdd pmos_6p0 w=1.215u l=0.5u
X3789 a_2708_31490# cap_shunt_p a_2500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X3790 a_16708_25218# cap_shunt_n a_16500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X3791 vdd a_9644_22760# a_9556_22804# vdd pmos_6p0 w=1.22u l=1u
X3792 a_24092_3511# a_24004_3608# vss vss nmos_6p0 w=0.82u l=1u
X3793 vdd a_28796_19624# a_28708_19668# vdd pmos_6p0 w=1.22u l=1u
X3794 vdd a_31708_55255# a_31620_55352# vdd pmos_6p0 w=1.22u l=1u
X3795 a_29492_27132# cap_shunt_p a_29700_26786# vdd pmos_6p0 w=1.2u l=0.5u
X3796 a_19732_7608# cap_series_gyp a_19524_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3797 a_1924_7608# cap_shunt_n a_1716_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3798 a_32716_12919# a_32628_13016# vss vss nmos_6p0 w=0.82u l=1u
X3799 vdd a_32268_50984# a_32180_51028# vdd pmos_6p0 w=1.22u l=1u
X3800 vss cap_shunt_p a_14896_48376# vss nmos_6p0 w=0.82u l=0.6u
X3801 vss cap_shunt_n a_12768_37700# vss nmos_6p0 w=0.82u l=0.6u
X3802 a_4760_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3803 a_34844_22760# a_34756_22804# vss vss nmos_6p0 w=0.82u l=1u
X3804 a_6292_18584# cap_shunt_p a_6084_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3805 a_30428_19668# cap_series_gygyn a_30616_19668# vdd pmos_6p0 w=1.2u l=0.5u
X3806 a_6532_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3807 vdd a_12332_55255# a_12244_55352# vdd pmos_6p0 w=1.22u l=1u
X3808 a_16708_22082# cap_shunt_n a_16500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3809 a_1924_4472# cap_shunt_p a_1716_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3810 a_13460_34264# cap_shunt_n a_15176_34264# vss nmos_6p0 w=0.82u l=0.6u
X3811 a_20740_29560# cap_shunt_n a_20532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X3812 vdd tune_series_gy[1] a_6572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3813 a_23576_12312# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X3814 vdd a_31708_52119# a_31620_52216# vdd pmos_6p0 w=1.22u l=1u
X3815 a_26892_52119# a_26804_52216# vss vss nmos_6p0 w=0.82u l=1u
X3816 a_3380_17016# cap_shunt_p a_5096_17016# vss nmos_6p0 w=0.82u l=0.6u
X3817 a_28692_7608# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X3818 a_16028_52552# a_15940_52596# vss vss nmos_6p0 w=0.82u l=1u
X3819 a_34144_48676# cap_shunt_gyn a_34144_49080# vdd pmos_6p0 w=1.215u l=0.5u
X3820 a_35880_25940# cap_series_gygyp a_35904_26424# vss nmos_6p0 w=0.82u l=0.6u
X3821 a_34348_8316# cap_series_gygyp a_34536_8316# vdd pmos_6p0 w=1.2u l=0.5u
X3822 a_34396_18056# a_34308_18100# vss vss nmos_6p0 w=0.82u l=1u
X3823 a_4312_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3824 vdd a_29468_19191# a_29380_19288# vdd pmos_6p0 w=1.22u l=1u
X3825 a_28692_24856# cap_shunt_p a_28484_24372# vdd pmos_6p0 w=1.2u l=0.5u
X3826 a_2500_38108# cap_shunt_n a_2708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X3827 a_13460_31128# cap_shunt_n a_15176_31128# vss nmos_6p0 w=0.82u l=0.6u
X3828 a_36308_39268# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X3829 a_7748_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3830 vss tune_shunt[7] a_13460_27992# vss nmos_6p0 w=0.51u l=0.6u
X3831 vdd a_4828_54120# a_4740_54164# vdd pmos_6p0 w=1.22u l=1u
X3832 a_13460_27992# cap_shunt_n a_13252_27508# vdd pmos_6p0 w=1.2u l=0.5u
X3833 a_16708_34626# cap_shunt_n a_16500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X3834 a_14392_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3835 a_21524_4472# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X3836 vss tune_series_gygy[5] a_35880_21236# vss nmos_6p0 w=0.51u l=0.6u
X3837 vdd a_23308_24328# a_23220_24372# vdd pmos_6p0 w=1.22u l=1u
X3838 a_25780_23288# cap_shunt_p a_27496_23288# vss nmos_6p0 w=0.82u l=0.6u
X3839 a_34396_14920# a_34308_14964# vss vss nmos_6p0 w=0.82u l=1u
X3840 vss tune_shunt[6] a_10660_45602# vss nmos_6p0 w=0.51u l=0.6u
X3841 a_13252_38484# cap_shunt_n a_13460_38968# vdd pmos_6p0 w=1.2u l=0.5u
X3842 vdd a_16924_29032# a_16836_29076# vdd pmos_6p0 w=1.22u l=1u
X3843 a_24452_28700# cap_shunt_n a_24660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X3844 vss cap_series_gygyp a_37080_7608# vss nmos_6p0 w=0.82u l=0.6u
X3845 a_7224_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3846 a_31648_20452# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X3847 a_3620_38484# cap_shunt_n a_3828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X3848 a_7748_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3849 vss cap_shunt_n a_15120_28292# vss nmos_6p0 w=0.82u l=0.6u
X3850 a_25780_20152# cap_series_gyp a_25572_19668# vdd pmos_6p0 w=1.2u l=0.5u
X3851 a_12668_52119# a_12580_52216# vss vss nmos_6p0 w=0.82u l=1u
X3852 vss tune_shunt[7] a_13460_24856# vss nmos_6p0 w=0.51u l=0.6u
X3853 a_34516_18946# cap_series_gygyn a_34308_19292# vdd pmos_6p0 w=1.2u l=0.5u
X3854 a_33052_55688# a_32964_55732# vss vss nmos_6p0 w=0.82u l=1u
X3855 vss tune_shunt[7] a_10660_36194# vss nmos_6p0 w=0.51u l=0.6u
X3856 a_16708_31490# cap_shunt_n a_16500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X3857 a_7176_7608# cap_series_gyp a_6760_7124# vss nmos_6p0 w=0.82u l=0.6u
X3858 vss tune_shunt[7] a_9876_18584# vss nmos_6p0 w=0.51u l=0.6u
X3859 vdd a_23308_21192# a_23220_21236# vdd pmos_6p0 w=1.22u l=1u
X3860 a_13252_35348# cap_shunt_n a_13460_35832# vdd pmos_6p0 w=1.2u l=0.5u
X3861 a_28692_27992# cap_shunt_p a_28484_27508# vdd pmos_6p0 w=1.2u l=0.5u
X3862 a_3620_35348# cap_shunt_n a_3828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X3863 vss cap_shunt_n a_15120_25156# vss nmos_6p0 w=0.82u l=0.6u
X3864 a_34516_15810# cap_series_gygyn a_34308_16156# vdd pmos_6p0 w=1.2u l=0.5u
X3865 a_19936_43672# cap_shunt_p a_17828_43672# vss nmos_6p0 w=0.82u l=0.6u
X3866 a_2500_47516# cap_shunt_p a_2708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X3867 vss tune_shunt[7] a_10660_33058# vss nmos_6p0 w=0.51u l=0.6u
X3868 vss tune_shunt[7] a_9876_15448# vss nmos_6p0 w=0.51u l=0.6u
X3869 vdd a_12556_16055# a_12468_16152# vdd pmos_6p0 w=1.22u l=1u
X3870 a_30028_55688# a_29940_55732# vss vss nmos_6p0 w=0.82u l=1u
X3871 vdd a_16252_13352# a_16164_13396# vdd pmos_6p0 w=1.22u l=1u
X3872 vss tune_series_gygy[3] a_35880_7124# vss nmos_6p0 w=0.51u l=0.6u
X3873 a_9108_47516# cap_shunt_p a_9316_47170# vdd pmos_6p0 w=1.2u l=0.5u
X3874 a_19936_40536# cap_shunt_n a_17828_40536# vss nmos_6p0 w=0.82u l=0.6u
X3875 a_18424_23588# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3876 a_32612_36194# cap_shunt_n a_34328_36132# vss nmos_6p0 w=0.82u l=0.6u
X3877 a_35692_7124# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3878 vdd a_12556_12919# a_12468_13016# vdd pmos_6p0 w=1.22u l=1u
X3879 a_2708_25218# cap_shunt_p a_2500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X3880 a_6292_51874# cap_shunt_p a_6084_52220# vdd pmos_6p0 w=1.2u l=0.5u
X3881 vss cap_shunt_n a_11872_35832# vss nmos_6p0 w=0.82u l=0.6u
X3882 a_16708_18946# cap_shunt_p a_16500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X3883 vdd tune_shunt[6] a_21540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X3884 vdd a_31708_48983# a_31620_49080# vdd pmos_6p0 w=1.22u l=1u
X3885 a_28692_40536# cap_shunt_p a_30408_40536# vss nmos_6p0 w=0.82u l=0.6u
X3886 a_2500_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3887 a_5612_55688# a_5524_55732# vss vss nmos_6p0 w=0.82u l=1u
X3888 a_16708_44034# cap_shunt_p a_17640_43972# vss nmos_6p0 w=0.82u l=0.6u
X3889 a_2708_22082# cap_shunt_p a_2500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3890 vdd a_12332_48983# a_12244_49080# vdd pmos_6p0 w=1.22u l=1u
X3891 a_10540_46280# a_10452_46324# vss vss nmos_6p0 w=0.82u l=1u
X3892 a_16708_15810# cap_shunt_p a_16500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X3893 vss cap_shunt_p a_4816_45540# vss nmos_6p0 w=0.82u l=0.6u
X3894 a_16708_40898# cap_shunt_n a_17640_40836# vss nmos_6p0 w=0.82u l=0.6u
X3895 a_2708_28354# cap_shunt_n a_2500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X3896 a_21748_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3897 a_28692_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3898 a_9316_22082# cap_shunt_p a_9108_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3899 a_25572_18100# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3900 a_31624_20860# cap_series_gygyn a_32432_20452# vss nmos_6p0 w=0.82u l=0.6u
X3901 a_31624_20860# cap_series_gygyn a_31436_20860# vdd pmos_6p0 w=1.2u l=0.5u
X3902 vdd a_25100_47415# a_25012_47512# vdd pmos_6p0 w=1.22u l=1u
X3903 a_1692_35304# a_1604_35348# vss vss nmos_6p0 w=0.82u l=1u
X3904 a_11984_29860# cap_shunt_n a_10660_29922# vss nmos_6p0 w=0.82u l=0.6u
X3905 a_16500_47516# cap_shunt_n a_16708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X3906 vdd a_28796_45847# a_28708_45944# vdd pmos_6p0 w=1.22u l=1u
X3907 a_6196_22428# cap_shunt_p a_6404_22082# vdd pmos_6p0 w=1.2u l=0.5u
X3908 a_5636_3612# cap_shunt_n a_5844_3266# vdd pmos_6p0 w=1.2u l=0.5u
X3909 vss cap_shunt_p a_4816_42404# vss nmos_6p0 w=0.82u l=0.6u
X3910 a_35880_16532# cap_series_gygyn a_35904_17016# vss nmos_6p0 w=0.82u l=0.6u
X3911 a_7748_37762# cap_shunt_n a_7540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X3912 a_9876_10744# cap_shunt_p a_9668_10260# vdd pmos_6p0 w=1.2u l=0.5u
X3913 vdd a_24204_43144# a_24116_43188# vdd pmos_6p0 w=1.22u l=1u
X3914 a_23464_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X3915 vdd a_33164_5079# a_33076_5176# vdd pmos_6p0 w=1.22u l=1u
X3916 vss tune_shunt[6] a_10660_39330# vss nmos_6p0 w=0.51u l=0.6u
X3917 a_25780_38968# cap_shunt_p a_26712_38968# vss nmos_6p0 w=0.82u l=0.6u
X3918 a_11984_26724# cap_shunt_n a_10660_26786# vss nmos_6p0 w=0.82u l=0.6u
X3919 a_8860_16488# a_8772_16532# vss vss nmos_6p0 w=0.82u l=1u
X3920 vdd a_3036_40008# a_2948_40052# vdd pmos_6p0 w=1.22u l=1u
X3921 a_7748_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3922 a_7336_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X3923 a_15492_5180# cap_series_gyn a_15700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X3924 a_3828_48376# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3925 vss tune_series_gy[4] a_24660_7970# vss nmos_6p0 w=0.51u l=0.6u
X3926 vss cap_shunt_p a_4032_18884# vss nmos_6p0 w=0.82u l=0.6u
X3927 a_3828_35832# cap_shunt_n a_5544_35832# vss nmos_6p0 w=0.82u l=0.6u
X3928 a_16708_25218# cap_shunt_n a_16500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X3929 vss tune_series_gygy[4] a_35880_11828# vss nmos_6p0 w=0.51u l=0.6u
X3930 vdd a_28684_54120# a_28596_54164# vdd pmos_6p0 w=1.22u l=1u
X3931 vdd a_37420_36439# a_37332_36536# vdd pmos_6p0 w=1.22u l=1u
X3932 a_14392_23288# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X3933 a_13252_29076# cap_shunt_n a_13460_29560# vdd pmos_6p0 w=1.2u l=0.5u
X3934 a_30428_19668# cap_series_gygyn a_30616_19668# vdd pmos_6p0 w=1.2u l=0.5u
X3935 a_3620_29076# cap_shunt_n a_3828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X3936 a_7748_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3937 vss tune_series_gy[5] a_18612_9538# vss nmos_6p0 w=0.51u l=0.6u
X3938 vss cap_shunt_p a_4032_15748# vss nmos_6p0 w=0.82u l=0.6u
X3939 a_16708_22082# cap_shunt_n a_16500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X3940 vss tune_series_gy[3] a_24660_4834# vss nmos_6p0 w=0.51u l=0.6u
X3941 vdd a_28684_50984# a_28596_51028# vdd pmos_6p0 w=1.22u l=1u
X3942 vss tune_shunt[5] a_6292_51512# vss nmos_6p0 w=0.51u l=0.6u
X3943 a_6084_16532# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3944 vss tune_shunt[5] a_2708_50306# vss nmos_6p0 w=0.51u l=0.6u
X3945 vss cap_shunt_gyn a_35532_48676# vss nmos_6p0 w=0.82u l=0.6u
X3946 vss cap_shunt_p a_23072_45540# vss nmos_6p0 w=0.82u l=0.6u
X3947 a_6532_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3948 a_12656_38968# cap_shunt_n a_10548_38968# vss nmos_6p0 w=0.82u l=0.6u
X3949 a_9668_13396# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3950 a_16364_54120# a_16276_54164# vss vss nmos_6p0 w=0.82u l=1u
X3951 a_11612_7124# cap_series_gyp a_11800_7124# vdd pmos_6p0 w=1.2u l=0.5u
X3952 a_19936_34264# cap_shunt_n a_17828_34264# vss nmos_6p0 w=0.82u l=0.6u
X3953 a_2500_38108# cap_shunt_n a_2708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X3954 a_20740_34264# cap_shunt_n a_20532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X3955 a_3036_32168# a_2948_32212# vss vss nmos_6p0 w=0.82u l=1u
X3956 a_2140_53687# a_2052_53784# vss vss nmos_6p0 w=0.82u l=1u
X3957 vdd a_31932_3511# a_31844_3608# vdd pmos_6p0 w=1.22u l=1u
X3958 a_2708_18946# cap_shunt_p a_2500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X3959 vss cap_shunt_n a_11872_29560# vss nmos_6p0 w=0.82u l=0.6u
X3960 vss cap_shunt_n a_23072_42404# vss nmos_6p0 w=0.82u l=0.6u
X3961 a_6532_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3962 a_28692_34264# cap_shunt_p a_30408_34264# vss nmos_6p0 w=0.82u l=0.6u
X3963 a_14012_5079# a_13924_5176# vss vss nmos_6p0 w=0.82u l=1u
X3964 a_22436_11828# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X3965 a_19524_11828# cap_series_gyn a_19732_12312# vdd pmos_6p0 w=1.2u l=0.5u
X3966 a_13252_38484# cap_shunt_n a_13460_38968# vdd pmos_6p0 w=1.2u l=0.5u
X3967 a_19936_31128# cap_shunt_n a_17828_31128# vss nmos_6p0 w=0.82u l=0.6u
X3968 a_24452_28700# cap_shunt_n a_24660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X3969 vss tune_shunt[7] a_24660_31490# vss nmos_6p0 w=0.51u l=0.6u
X3970 a_20740_31128# cap_shunt_n a_20532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X3971 a_2140_50551# a_2052_50648# vss vss nmos_6p0 w=0.82u l=1u
X3972 a_24660_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3973 a_2708_15810# cap_shunt_p a_2500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X3974 vss cap_shunt_n a_11872_26424# vss nmos_6p0 w=0.82u l=0.6u
X3975 a_1924_4472# cap_shunt_p a_1716_3988# vdd pmos_6p0 w=1.2u l=0.5u
X3976 a_28692_31128# cap_shunt_n a_30408_31128# vss nmos_6p0 w=0.82u l=0.6u
X3977 a_7580_6748# cap_series_gyp a_7768_6748# vdd pmos_6p0 w=1.2u l=0.5u
X3978 a_16708_47170# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X3979 a_13252_35348# cap_shunt_n a_13460_35832# vdd pmos_6p0 w=1.2u l=0.5u
X3980 a_16708_34626# cap_shunt_n a_17640_34564# vss nmos_6p0 w=0.82u l=0.6u
X3981 a_35880_18100# cap_series_gygyn a_35692_18100# vdd pmos_6p0 w=1.2u l=0.5u
X3982 a_2708_20514# cap_shunt_p a_2500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X3983 a_28484_38484# cap_shunt_n a_28692_38968# vdd pmos_6p0 w=1.2u l=0.5u
X3984 a_16016_10744# cap_series_gyn a_14692_10744# vss nmos_6p0 w=0.82u l=0.6u
X3985 a_1692_29032# a_1604_29076# vss vss nmos_6p0 w=0.82u l=1u
X3986 a_34560_6340# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X3987 a_22436_8692# cap_series_gyp a_22644_9176# vdd pmos_6p0 w=1.2u l=0.5u
X3988 a_10092_8648# a_10004_8692# vss vss nmos_6p0 w=0.82u l=1u
X3989 a_16708_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X3990 a_16708_31490# cap_shunt_n a_17640_31428# vss nmos_6p0 w=0.82u l=0.6u
X3991 a_21748_17378# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X3992 vss tune_shunt[5] a_6740_53080# vss nmos_6p0 w=0.51u l=0.6u
X3993 vss cap_shunt_n a_4816_36132# vss nmos_6p0 w=0.82u l=0.6u
X3994 a_33164_17623# a_33076_17720# vss vss nmos_6p0 w=0.82u l=1u
X3995 a_34516_20514# cap_series_gygyp a_34308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X3996 a_7748_29922# cap_shunt_n a_7540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X3997 a_9876_13880# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X3998 vss tune_shunt[6] a_11668_43672# vss nmos_6p0 w=0.51u l=0.6u
X3999 a_28484_35348# cap_shunt_p a_28692_35832# vdd pmos_6p0 w=1.2u l=0.5u
X4000 vdd tune_shunt[4] a_25572_41620# vdd pmos_6p0 w=1.2u l=0.5u
X4001 a_1692_25896# a_1604_25940# vss vss nmos_6p0 w=0.82u l=1u
X4002 a_4032_4772# cap_shunt_p a_1924_4834# vss nmos_6p0 w=0.82u l=0.6u
X4003 a_16500_38108# cap_shunt_n a_16708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X4004 a_24452_30268# cap_shunt_n a_24660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X4005 a_29700_33058# cap_shunt_p a_31416_32996# vss nmos_6p0 w=0.82u l=0.6u
X4006 a_3828_29560# cap_shunt_n a_5544_29560# vss nmos_6p0 w=0.82u l=0.6u
X4007 a_16708_18946# cap_shunt_p a_16500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X4008 a_15244_55688# a_15156_55732# vss vss nmos_6p0 w=0.82u l=1u
X4009 vdd tune_series_gygy[4] a_35692_36916# vdd pmos_6p0 w=1.2u l=0.5u
X4010 a_18404_9884# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4011 a_9876_10744# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4012 a_37632_41240# cap_shunt_gyp a_37444_41240# vdd pmos_6p0 w=1.215u l=0.5u
X4013 vss tune_shunt[6] a_11668_40536# vss nmos_6p0 w=0.51u l=0.6u
X4014 a_10340_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4015 vss tune_shunt[5] a_2708_47170# vss nmos_6p0 w=0.51u l=0.6u
X4016 vdd tune_shunt[6] a_14372_41620# vdd pmos_6p0 w=1.2u l=0.5u
X4017 a_16500_42812# cap_shunt_n a_16708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X4018 a_27496_37400# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4019 a_6084_50652# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4020 vss cap_shunt_gyp a_34412_47108# vss nmos_6p0 w=0.82u l=0.6u
X4021 a_3828_26424# cap_shunt_p a_5544_26424# vss nmos_6p0 w=0.82u l=0.6u
X4022 a_8576_7908# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4023 vdd tune_shunt[5] a_21540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X4024 vdd a_37420_27031# a_37332_27128# vdd pmos_6p0 w=1.22u l=1u
X4025 a_14484_7124# cap_series_gyp a_14692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X4026 a_16708_15810# cap_shunt_p a_16500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X4027 vdd tune_shunt_gy[6] a_30500_45944# vdd pmos_6p0 w=1.215u l=0.5u
X4028 a_18404_6748# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4029 a_32156_5512# a_32068_5556# vss vss nmos_6p0 w=0.82u l=1u
X4030 a_10704_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4031 a_6404_47170# cap_shunt_p a_7336_47108# vss nmos_6p0 w=0.82u l=0.6u
X4032 a_10340_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4033 a_27888_9176# cap_series_gyp a_25780_9176# vss nmos_6p0 w=0.82u l=0.6u
X4034 vss tune_shunt[6] a_2708_44034# vss nmos_6p0 w=0.51u l=0.6u
X4035 vdd a_14460_8215# a_14372_8312# vdd pmos_6p0 w=1.22u l=1u
X4036 a_9316_22082# cap_shunt_p a_9108_22428# vdd pmos_6p0 w=1.2u l=0.5u
X4037 a_29132_49416# a_29044_49460# vss vss nmos_6p0 w=0.82u l=1u
X4038 a_34536_8316# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X4039 a_11668_43672# cap_shunt_n a_12600_43672# vss nmos_6p0 w=0.82u l=0.6u
X4040 a_22644_13880# cap_series_gyn a_22436_13396# vdd pmos_6p0 w=1.2u l=0.5u
X4041 vss cap_shunt_p a_7616_17016# vss nmos_6p0 w=0.82u l=0.6u
X4042 a_7224_49944# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4043 a_38092_32168# a_38004_32212# vss vss nmos_6p0 w=0.82u l=1u
X4044 a_13588_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4045 vdd a_34844_19624# a_34756_19668# vdd pmos_6p0 w=1.22u l=1u
X4046 vss cap_shunt_n a_23072_36132# vss nmos_6p0 w=0.82u l=0.6u
X4047 vdd a_23756_33736# a_23668_33780# vdd pmos_6p0 w=1.22u l=1u
X4048 a_33732_27992# cap_shunt_p a_33524_27508# vdd pmos_6p0 w=1.2u l=0.5u
X4049 a_6532_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4050 a_14896_12312# cap_shunt_p a_12788_12312# vss nmos_6p0 w=0.82u l=0.6u
X4051 a_29132_46280# a_29044_46324# vss vss nmos_6p0 w=0.82u l=1u
X4052 vss cap_series_gygyp a_37080_37400# vss nmos_6p0 w=0.82u l=0.6u
X4053 a_11668_40536# cap_shunt_n a_12600_40536# vss nmos_6p0 w=0.82u l=0.6u
X4054 a_20740_24856# cap_shunt_n a_20532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X4055 a_3036_22760# a_2948_22804# vss vss nmos_6p0 w=0.82u l=1u
X4056 a_17828_20152# cap_shunt_p a_17620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X4057 a_16252_55255# a_16164_55352# vss vss nmos_6p0 w=0.82u l=1u
X4058 vdd a_23756_30600# a_23668_30644# vdd pmos_6p0 w=1.22u l=1u
X4059 vdd tune_series_gy[4] a_15492_9884# vdd pmos_6p0 w=1.2u l=0.5u
X4060 a_25780_4472# cap_shunt_p a_27496_4472# vss nmos_6p0 w=0.82u l=0.6u
X4061 a_6532_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4062 a_14728_43972# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4063 vdd a_20172_34871# a_20084_34968# vdd pmos_6p0 w=1.22u l=1u
X4064 a_9540_14242# cap_shunt_p a_10472_14180# vss nmos_6p0 w=0.82u l=0.6u
X4065 a_13252_29076# cap_shunt_n a_13460_29560# vdd pmos_6p0 w=1.2u l=0.5u
X4066 a_16708_28354# cap_shunt_n a_17640_28292# vss nmos_6p0 w=0.82u l=0.6u
X4067 vss tune_shunt[7] a_24660_22082# vss nmos_6p0 w=0.51u l=0.6u
X4068 vss cap_shunt_p a_8848_20152# vss nmos_6p0 w=0.82u l=0.6u
X4069 a_20740_21720# cap_shunt_p a_20532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X4070 a_34060_39575# a_33972_39672# vss vss nmos_6p0 w=0.82u l=1u
X4071 vdd a_27676_38007# a_27588_38104# vdd pmos_6p0 w=1.22u l=1u
X4072 a_28692_4472# cap_series_gyp a_28484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X4073 vdd a_35628_30167# a_35540_30264# vdd pmos_6p0 w=1.22u l=1u
X4074 vdd a_33948_8648# a_33860_8692# vdd pmos_6p0 w=1.22u l=1u
X4075 vdd tune_series_gy[4] a_15492_6748# vdd pmos_6p0 w=1.2u l=0.5u
X4076 a_14728_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4077 a_9540_11106# cap_shunt_p a_10472_11044# vss nmos_6p0 w=0.82u l=0.6u
X4078 a_37280_51574# cap_shunt_gyp a_37280_51029# vdd pmos_6p0 w=1.215u l=0.5u
X4079 vdd tune_series_gy[2] a_11572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X4080 a_34844_3511# a_34756_3608# vss vss nmos_6p0 w=0.82u l=1u
X4081 a_16708_25218# cap_shunt_n a_17640_25156# vss nmos_6p0 w=0.82u l=0.6u
X4082 a_6084_16532# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4083 vdd tune_shunt[1] a_1716_3612# vdd pmos_6p0 w=1.2u l=0.5u
X4084 a_27676_19191# a_27588_19288# vss vss nmos_6p0 w=0.82u l=1u
X4085 a_16632_6340# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4086 vdd a_33948_5512# a_33860_5556# vdd pmos_6p0 w=1.22u l=1u
X4087 a_2708_11106# cap_shunt_n a_2500_11452# vdd pmos_6p0 w=1.2u l=0.5u
X4088 a_22848_45240# cap_shunt_n a_20740_45240# vss nmos_6p0 w=0.82u l=0.6u
X4089 a_28484_29076# cap_shunt_p a_28692_29560# vdd pmos_6p0 w=1.2u l=0.5u
X4090 a_10452_28700# cap_shunt_n a_10660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X4091 a_29700_4834# cap_shunt_p a_29492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X4092 a_5844_9538# cap_shunt_p a_5636_9884# vdd pmos_6p0 w=1.2u l=0.5u
X4093 a_20740_34264# cap_shunt_n a_20532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X4094 a_28572_6647# a_28484_6744# vss vss nmos_6p0 w=0.82u l=1u
X4095 a_16500_30268# cap_shunt_n a_16708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X4096 a_7748_28354# cap_shunt_n a_7540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X4097 a_21636_6040# cap_series_gyp a_22568_6040# vss nmos_6p0 w=0.82u l=0.6u
X4098 a_19524_11828# cap_series_gyn a_19732_12312# vdd pmos_6p0 w=1.2u l=0.5u
X4099 a_27676_16055# a_27588_16152# vss vss nmos_6p0 w=0.82u l=1u
X4100 a_22848_42104# cap_shunt_p a_20740_42104# vss nmos_6p0 w=0.82u l=0.6u
X4101 vdd a_33500_13352# a_33412_13396# vdd pmos_6p0 w=1.22u l=1u
X4102 a_2500_42812# cap_shunt_p a_2708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X4103 a_1692_16488# a_1604_16532# vss vss nmos_6p0 w=0.82u l=1u
X4104 a_16028_38440# a_15940_38484# vss vss nmos_6p0 w=0.82u l=1u
X4105 a_16500_36540# cap_shunt_n a_16708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X4106 vdd tune_shunt[6] a_25572_32212# vdd pmos_6p0 w=1.2u l=0.5u
X4107 a_20740_31128# cap_shunt_n a_20532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X4108 a_20740_37400# cap_shunt_n a_20532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X4109 a_9316_48738# cap_shunt_p a_9108_49084# vdd pmos_6p0 w=1.2u l=0.5u
X4110 a_29700_23650# cap_shunt_p a_31416_23588# vss nmos_6p0 w=0.82u l=0.6u
X4111 vdd tune_shunt[6] a_21540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X4112 a_35692_8692# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4113 a_13460_35832# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4114 vss cap_series_gyp a_27104_20152# vss nmos_6p0 w=0.82u l=0.6u
X4115 vdd a_12780_55255# a_12692_55352# vdd pmos_6p0 w=1.22u l=1u
X4116 a_16500_33404# cap_shunt_n a_16708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X4117 a_12580_16532# cap_shunt_p a_12788_17016# vdd pmos_6p0 w=1.2u l=0.5u
X4118 a_2708_20514# cap_shunt_p a_2500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X4119 a_25572_10260# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4120 a_28484_38484# cap_shunt_n a_28692_38968# vdd pmos_6p0 w=1.2u l=0.5u
X4121 vdd tune_shunt[7] a_21540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X4122 a_25780_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4123 vdd a_23084_55688# a_22996_55732# vdd pmos_6p0 w=1.22u l=1u
X4124 a_16476_52552# a_16388_52596# vss vss nmos_6p0 w=0.82u l=1u
X4125 a_35692_5556# tune_series_gygy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4126 vss tune_shunt[7] a_33732_27992# vss nmos_6p0 w=0.51u l=0.6u
X4127 a_13796_44034# cap_shunt_n a_15512_43972# vss nmos_6p0 w=0.82u l=0.6u
X4128 a_13588_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4129 a_23856_43972# cap_shunt_n a_21748_44034# vss nmos_6p0 w=0.82u l=0.6u
X4130 a_34516_20514# cap_series_gygyp a_34308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X4131 a_13796_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4132 a_7748_29922# cap_shunt_n a_7540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X4133 vss tune_shunt[5] a_13796_48738# vss nmos_6p0 w=0.51u l=0.6u
X4134 a_28484_35348# cap_shunt_p a_28692_35832# vdd pmos_6p0 w=1.2u l=0.5u
X4135 a_25780_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4136 a_5612_8215# a_5524_8312# vss vss nmos_6p0 w=0.82u l=1u
X4137 a_26768_9476# cap_series_gyn a_24660_9538# vss nmos_6p0 w=0.82u l=0.6u
X4138 a_5152_46808# cap_shunt_p a_3828_46808# vss nmos_6p0 w=0.82u l=0.6u
X4139 vdd tune_series_gy[1] a_10340_3612# vdd pmos_6p0 w=1.2u l=0.5u
X4140 vss tune_series_gy[5] a_19732_9176# vss nmos_6p0 w=0.51u l=0.6u
X4141 a_13796_40898# cap_shunt_n a_15512_40836# vss nmos_6p0 w=0.82u l=0.6u
X4142 vdd a_23756_24328# a_23668_24372# vdd pmos_6p0 w=1.22u l=1u
X4143 a_25984_12612# cap_series_gyn a_24660_12674# vss nmos_6p0 w=0.82u l=0.6u
X4144 vdd a_21628_52552# a_21540_52596# vdd pmos_6p0 w=1.22u l=1u
X4145 a_23856_40836# cap_shunt_p a_21748_40898# vss nmos_6p0 w=0.82u l=0.6u
X4146 vss tune_shunt[7] a_9540_15810# vss nmos_6p0 w=0.51u l=0.6u
X4147 vss cap_shunt_n a_22848_32696# vss nmos_6p0 w=0.82u l=0.6u
X4148 a_28484_32212# cap_shunt_p a_28692_32696# vdd pmos_6p0 w=1.2u l=0.5u
X4149 a_9220_17724# cap_shunt_p a_9428_17378# vdd pmos_6p0 w=1.2u l=0.5u
X4150 vdd tune_series_gygy[4] a_35692_36916# vdd pmos_6p0 w=1.2u l=0.5u
X4151 vdd a_20172_28599# a_20084_28696# vdd pmos_6p0 w=1.22u l=1u
X4152 a_31436_8316# cap_series_gygyn a_31624_8316# vdd pmos_6p0 w=1.2u l=0.5u
X4153 a_18044_50984# a_17956_51028# vss vss nmos_6p0 w=0.82u l=1u
X4154 a_10660_42466# cap_shunt_n a_10452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X4155 a_2500_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4156 vdd tune_shunt[7] a_9220_19292# vdd pmos_6p0 w=1.2u l=0.5u
X4157 vdd a_23756_21192# a_23668_21236# vdd pmos_6p0 w=1.22u l=1u
X4158 a_6084_50652# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4159 a_14728_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4160 a_3828_46808# cap_shunt_p a_3620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X4161 vdd tune_shunt[6] a_6532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X4162 a_12600_45240# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4163 a_24660_4834# cap_series_gyp a_24452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X4164 a_24660_4834# cap_series_gyp a_26376_4772# vss nmos_6p0 w=0.82u l=0.6u
X4165 a_22436_10260# cap_series_gyp a_22644_10744# vdd pmos_6p0 w=1.2u l=0.5u
X4166 a_8456_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4167 a_14692_7608# cap_series_gyp a_16408_7608# vss nmos_6p0 w=0.82u l=0.6u
X4168 a_30476_55688# a_30388_55732# vss vss nmos_6p0 w=0.82u l=1u
X4169 a_36296_26424# cap_series_gygyp a_35880_25940# vss nmos_6p0 w=0.82u l=0.6u
X4170 vdd a_2140_23895# a_2052_23992# vdd pmos_6p0 w=1.22u l=1u
X4171 a_16708_20514# cap_shunt_p a_16500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X4172 a_14728_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4173 vss tune_shunt[6] a_7748_44034# vss nmos_6p0 w=0.51u l=0.6u
X4174 vdd tune_series_gy[2] a_7580_8316# vdd pmos_6p0 w=1.2u l=0.5u
X4175 vss tune_shunt[7] a_13796_15810# vss nmos_6p0 w=0.51u l=0.6u
X4176 a_12600_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4177 a_8456_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4178 vss cap_series_gyn a_20720_6340# vss nmos_6p0 w=0.82u l=0.6u
X4179 a_2588_13352# a_2500_13396# vss vss nmos_6p0 w=0.82u l=1u
X4180 a_2500_36540# cap_shunt_n a_2708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X4181 vdd a_2140_20759# a_2052_20856# vdd pmos_6p0 w=1.22u l=1u
X4182 a_20740_24856# cap_shunt_n a_20532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X4183 vss tune_shunt[1] a_5844_3266# vss nmos_6p0 w=0.51u l=0.6u
X4184 a_24660_42466# cap_shunt_n a_25592_42404# vss nmos_6p0 w=0.82u l=0.6u
X4185 vdd a_19724_41143# a_19636_41240# vdd pmos_6p0 w=1.22u l=1u
X4186 a_37652_47108# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4187 vdd tune_shunt[6] a_16500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X4188 a_7768_5180# cap_series_gyn a_7580_5180# vdd pmos_6p0 w=1.2u l=0.5u
X4189 vss tune_series_gy[3] a_28692_7608# vss nmos_6p0 w=0.51u l=0.6u
X4190 a_37632_45944# cap_shunt_gyn a_37652_45540# vss nmos_6p0 w=0.82u l=0.6u
X4191 vdd a_30364_41143# a_30276_41240# vdd pmos_6p0 w=1.22u l=1u
X4192 a_2500_33404# cap_shunt_p a_2708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X4193 a_13460_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4194 a_9332_13020# cap_shunt_p a_9540_12674# vdd pmos_6p0 w=1.2u l=0.5u
X4195 a_28484_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4196 a_20740_21720# cap_shunt_p a_20532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X4197 vdd a_12332_54120# a_12244_54164# vdd pmos_6p0 w=1.22u l=1u
X4198 vdd a_12780_48983# a_12692_49080# vdd pmos_6p0 w=1.22u l=1u
X4199 a_20740_27992# cap_shunt_n a_20532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X4200 a_16500_27132# cap_shunt_n a_16708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X4201 a_14484_3988# cap_series_gyp a_14692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X4202 a_16500_47516# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4203 vss tune_shunt[5] a_2708_18946# vss nmos_6p0 w=0.51u l=0.6u
X4204 a_20396_47848# a_20308_47892# vss vss nmos_6p0 w=0.82u l=1u
X4205 a_34664_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4206 a_4424_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4207 vdd tune_shunt[7] a_21540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X4208 a_13252_33780# cap_shunt_n a_13460_34264# vdd pmos_6p0 w=1.2u l=0.5u
X4209 a_13460_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4210 vdd a_37420_47848# a_37332_47892# vdd pmos_6p0 w=1.22u l=1u
X4211 a_37632_42808# cap_shunt_gyn a_37652_42404# vss nmos_6p0 w=0.82u l=0.6u
X4212 a_3172_16532# cap_shunt_p a_3380_17016# vdd pmos_6p0 w=1.2u l=0.5u
X4213 a_3620_33780# cap_shunt_n a_3828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X4214 a_2708_11106# cap_shunt_n a_2500_11452# vdd pmos_6p0 w=1.2u l=0.5u
X4215 vss tune_series_gygy[4] a_31624_19292# vss nmos_6p0 w=0.51u l=0.6u
X4216 a_35292_8648# a_35204_8692# vss vss nmos_6p0 w=0.82u l=1u
X4217 a_23308_47415# a_23220_47512# vss vss nmos_6p0 w=0.82u l=1u
X4218 vdd a_19276_33303# a_19188_33400# vdd pmos_6p0 w=1.22u l=1u
X4219 a_28484_29076# cap_shunt_p a_28692_29560# vdd pmos_6p0 w=1.2u l=0.5u
X4220 a_25780_18584# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X4221 a_11984_49944# cap_shunt_p a_9876_49944# vss nmos_6p0 w=0.82u l=0.6u
X4222 vdd a_24652_43144# a_24564_43188# vdd pmos_6p0 w=1.22u l=1u
X4223 a_13796_34626# cap_shunt_n a_15512_34564# vss nmos_6p0 w=0.82u l=0.6u
X4224 a_13252_30644# cap_shunt_n a_13460_31128# vdd pmos_6p0 w=1.2u l=0.5u
X4225 a_10660_6402# cap_series_gyn a_10452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X4226 a_20284_55255# a_20196_55352# vss vss nmos_6p0 w=0.82u l=1u
X4227 a_3380_51512# cap_shunt_n a_5096_51512# vss nmos_6p0 w=0.82u l=0.6u
X4228 a_16500_30268# cap_shunt_n a_16708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X4229 vdd a_32828_43144# a_32740_43188# vdd pmos_6p0 w=1.22u l=1u
X4230 a_23856_34564# cap_shunt_p a_21748_34626# vss nmos_6p0 w=0.82u l=0.6u
X4231 a_14012_11351# a_13924_11448# vss vss nmos_6p0 w=0.82u l=1u
X4232 a_14580_45240# cap_shunt_p a_14372_44756# vdd pmos_6p0 w=1.2u l=0.5u
X4233 a_3620_36916# cap_shunt_n a_3828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X4234 a_3620_30644# cap_shunt_n a_3828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X4235 vdd a_29468_53687# a_29380_53784# vdd pmos_6p0 w=1.22u l=1u
X4236 a_12264_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4237 a_37868_22327# a_37780_22424# vss vss nmos_6p0 w=0.82u l=1u
X4238 a_25780_15448# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4239 a_29244_41576# a_29156_41620# vss vss nmos_6p0 w=0.82u l=1u
X4240 vss cap_shunt_n a_33936_32996# vss nmos_6p0 w=0.82u l=0.6u
X4241 a_9072_37700# cap_shunt_n a_7748_37762# vss nmos_6p0 w=0.82u l=0.6u
X4242 a_10660_36194# cap_shunt_n a_10452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X4243 a_13796_31490# cap_shunt_n a_15512_31428# vss nmos_6p0 w=0.82u l=0.6u
X4244 a_5636_9884# cap_shunt_p a_5844_9538# vdd pmos_6p0 w=1.2u l=0.5u
X4245 a_12580_49460# cap_shunt_n a_12788_49944# vdd pmos_6p0 w=1.2u l=0.5u
X4246 a_23856_31428# cap_shunt_n a_21748_31490# vss nmos_6p0 w=0.82u l=0.6u
X4247 a_14728_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4248 vss cap_shunt_p a_22848_23288# vss nmos_6p0 w=0.82u l=0.6u
X4249 vss cap_series_gyn a_20720_12612# vss nmos_6p0 w=0.82u l=0.6u
X4250 a_16364_50551# a_16276_50648# vss vss nmos_6p0 w=0.82u l=1u
X4251 vdd tune_shunt[6] a_13588_42812# vdd pmos_6p0 w=1.2u l=0.5u
X4252 a_32612_28354# cap_shunt_p a_32404_28700# vdd pmos_6p0 w=1.2u l=0.5u
X4253 a_32444_11452# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4254 vdd a_20172_19191# a_20084_19288# vdd pmos_6p0 w=1.22u l=1u
X4255 a_5936_20152# cap_shunt_p a_3828_20152# vss nmos_6p0 w=0.82u l=0.6u
X4256 vdd a_29468_50551# a_29380_50648# vdd pmos_6p0 w=1.22u l=1u
X4257 vss cap_shunt_p a_18032_48676# vss nmos_6p0 w=0.82u l=0.6u
X4258 a_30016_37400# cap_shunt_p a_28692_37400# vss nmos_6p0 w=0.82u l=0.6u
X4259 a_3828_15448# cap_shunt_p a_3620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X4260 a_7224_51812# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4261 a_10660_33058# cap_shunt_n a_10452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X4262 a_2500_14588# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4263 vss cap_series_gygyp a_35736_7908# vss nmos_6p0 w=0.82u l=0.6u
X4264 a_28484_38484# cap_shunt_n a_28692_38968# vdd pmos_6p0 w=1.2u l=0.5u
X4265 a_14728_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4266 vss cap_shunt_p a_8736_14180# vss nmos_6p0 w=0.82u l=0.6u
X4267 a_6644_53788# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4268 vss tune_shunt[7] a_17828_35832# vss nmos_6p0 w=0.51u l=0.6u
X4269 a_21540_44380# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4270 a_8456_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4271 vdd tune_shunt[3] a_5636_10260# vdd pmos_6p0 w=1.2u l=0.5u
X4272 a_9316_50306# cap_shunt_p a_9108_50652# vdd pmos_6p0 w=1.2u l=0.5u
X4273 a_28012_3511# a_27924_3608# vss vss nmos_6p0 w=0.82u l=1u
X4274 vdd a_2140_14487# a_2052_14584# vdd pmos_6p0 w=1.22u l=1u
X4275 a_20740_43672# cap_shunt_n a_21672_43672# vss nmos_6p0 w=0.82u l=0.6u
X4276 a_28484_35348# cap_shunt_p a_28692_35832# vdd pmos_6p0 w=1.2u l=0.5u
X4277 a_36296_17016# cap_series_gygyn a_35880_16532# vss nmos_6p0 w=0.82u l=0.6u
X4278 a_2708_20514# cap_shunt_p a_3640_20452# vss nmos_6p0 w=0.82u l=0.6u
X4279 vdd tune_shunt[6] a_16500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X4280 a_24660_36194# cap_shunt_p a_25592_36132# vss nmos_6p0 w=0.82u l=0.6u
X4281 a_21540_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4282 a_33936_36132# cap_shunt_n a_32612_36194# vss nmos_6p0 w=0.82u l=0.6u
X4283 a_8456_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4284 a_11572_5556# cap_series_gyn a_11780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X4285 a_16708_48738# cap_shunt_p a_16500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X4286 vdd a_2140_11351# a_2052_11448# vdd pmos_6p0 w=1.22u l=1u
X4287 a_6740_13880# cap_shunt_p a_8456_13880# vss nmos_6p0 w=0.82u l=0.6u
X4288 a_20740_40536# cap_shunt_p a_21672_40536# vss nmos_6p0 w=0.82u l=0.6u
X4289 a_17620_36916# cap_shunt_n a_17828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X4290 a_2500_27132# cap_shunt_p a_2708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X4291 a_27228_44279# a_27140_44376# vss vss nmos_6p0 w=0.82u l=1u
X4292 a_11668_42104# cap_shunt_n a_11460_41620# vdd pmos_6p0 w=1.2u l=0.5u
X4293 vss tune_shunt[6] a_6740_38968# vss nmos_6p0 w=0.51u l=0.6u
X4294 a_32612_29922# cap_shunt_p a_32404_30268# vdd pmos_6p0 w=1.2u l=0.5u
X4295 a_10660_42466# cap_shunt_n a_10452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X4296 vdd tune_shunt[7] a_9220_19292# vdd pmos_6p0 w=1.2u l=0.5u
X4297 vdd tune_shunt[5] a_12580_19668# vdd pmos_6p0 w=1.2u l=0.5u
X4298 a_9876_20152# cap_shunt_p a_9668_19668# vdd pmos_6p0 w=1.2u l=0.5u
X4299 a_34664_29560# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4300 vdd tune_series_gy[0] a_28484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X4301 a_33500_55255# a_33412_55352# vss vss nmos_6p0 w=0.82u l=1u
X4302 vdd a_5612_31735# a_5524_31832# vdd pmos_6p0 w=1.22u l=1u
X4303 a_6760_7124# cap_series_gyp a_6572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X4304 a_17596_3944# a_17508_3988# vss vss nmos_6p0 w=0.82u l=1u
X4305 a_31416_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4306 a_17828_35832# cap_shunt_n a_18760_35832# vss nmos_6p0 w=0.82u l=0.6u
X4307 vdd a_3036_19624# a_2948_19668# vdd pmos_6p0 w=1.22u l=1u
X4308 a_1692_22327# a_1604_22424# vss vss nmos_6p0 w=0.82u l=1u
X4309 a_29624_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4310 a_28124_8215# a_28036_8312# vss vss nmos_6p0 w=0.82u l=1u
X4311 a_7540_44380# cap_shunt_p a_7748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X4312 a_27228_41143# a_27140_41240# vss vss nmos_6p0 w=0.82u l=1u
X4313 a_28692_40536# cap_shunt_p a_28484_40052# vdd pmos_6p0 w=1.2u l=0.5u
X4314 a_25780_38968# cap_shunt_p a_25572_38484# vdd pmos_6p0 w=1.2u l=0.5u
X4315 a_17828_15448# cap_shunt_p a_17620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X4316 a_16500_38108# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4317 a_14692_9176# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X4318 a_34516_18946# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4319 a_32040_20452# cap_series_gygyn a_31624_20860# vss nmos_6p0 w=0.82u l=0.6u
X4320 vdd a_17148_55255# a_17060_55352# vdd pmos_6p0 w=1.22u l=1u
X4321 a_13252_24372# cap_shunt_n a_13460_24856# vdd pmos_6p0 w=1.2u l=0.5u
X4322 vss tune_shunt[7] a_12788_17016# vss nmos_6p0 w=0.51u l=0.6u
X4323 a_9464_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4324 a_10660_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4325 a_13796_28354# cap_shunt_n a_15512_28292# vss nmos_6p0 w=0.82u l=0.6u
X4326 vss cap_series_gygyp a_36296_7608# vss nmos_6p0 w=0.82u l=0.6u
X4327 a_7540_41244# cap_shunt_n a_7748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X4328 a_23856_28292# cap_shunt_n a_21748_28354# vss nmos_6p0 w=0.82u l=0.6u
X4329 vdd a_6508_6647# a_6420_6744# vdd pmos_6p0 w=1.22u l=1u
X4330 a_18612_12674# cap_series_gyn a_18404_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4331 a_25780_35832# cap_shunt_p a_25572_35348# vdd pmos_6p0 w=1.2u l=0.5u
X4332 a_3620_24372# cap_shunt_p a_3828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X4333 vdd a_24204_18056# a_24116_18100# vdd pmos_6p0 w=1.22u l=1u
X4334 a_35600_49461# cap_shunt_gyp a_35600_50006# vdd pmos_6p0 w=1.215u l=0.5u
X4335 a_12264_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4336 a_6532_14964# cap_shunt_p a_6740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X4337 vdd a_17148_52119# a_17060_52216# vdd pmos_6p0 w=1.22u l=1u
X4338 a_22076_50984# a_21988_51028# vss vss nmos_6p0 w=0.82u l=1u
X4339 a_11460_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4340 a_13252_21236# cap_shunt_n a_13460_21720# vdd pmos_6p0 w=1.2u l=0.5u
X4341 a_15692_55688# a_15604_55732# vss vss nmos_6p0 w=0.82u l=1u
X4342 vdd tune_shunt[6] a_16500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X4343 a_13796_25218# cap_shunt_n a_15512_25156# vss nmos_6p0 w=0.82u l=0.6u
X4344 a_10452_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4345 a_23856_25156# cap_shunt_n a_21748_25218# vss nmos_6p0 w=0.82u l=0.6u
X4346 a_35692_14964# cap_series_gygyn a_35880_14964# vdd pmos_6p0 w=1.2u l=0.5u
X4347 a_33948_19624# a_33860_19668# vss vss nmos_6p0 w=0.82u l=1u
X4348 vdd tune_shunt[7] a_13588_36540# vdd pmos_6p0 w=1.2u l=0.5u
X4349 vdd a_5836_5512# a_5748_5556# vdd pmos_6p0 w=1.22u l=1u
X4350 a_3620_21236# cap_shunt_p a_3828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X4351 a_3620_27508# cap_shunt_n a_3828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X4352 a_35600_46325# cap_shunt_gyp a_35600_46870# vdd pmos_6p0 w=1.215u l=0.5u
X4353 vdd a_29468_44279# a_29380_44376# vdd pmos_6p0 w=1.22u l=1u
X4354 a_12264_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4355 a_9332_13020# cap_shunt_p a_9540_12674# vdd pmos_6p0 w=1.2u l=0.5u
X4356 a_3640_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4357 a_8860_50984# a_8772_51028# vss vss nmos_6p0 w=0.82u l=1u
X4358 a_6532_11828# cap_shunt_p a_6740_12312# vdd pmos_6p0 w=1.2u l=0.5u
X4359 a_3172_49460# cap_shunt_p a_3380_49944# vdd pmos_6p0 w=1.2u l=0.5u
X4360 a_10660_26786# cap_shunt_n a_10452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X4361 vss cap_shunt_p a_5936_48376# vss nmos_6p0 w=0.82u l=0.6u
X4362 a_13588_23996# cap_shunt_n a_13796_23650# vdd pmos_6p0 w=1.2u l=0.5u
X4363 a_35692_11828# cap_series_gygyp a_35880_11828# vdd pmos_6p0 w=1.2u l=0.5u
X4364 a_12668_55688# a_12580_55732# vss vss nmos_6p0 w=0.82u l=1u
X4365 vss cap_shunt_n a_18032_39268# vss nmos_6p0 w=0.82u l=0.6u
X4366 vdd tune_shunt[7] a_13588_33404# vdd pmos_6p0 w=1.2u l=0.5u
X4367 vss tune_shunt[7] a_17828_29560# vss nmos_6p0 w=0.51u l=0.6u
X4368 vdd tune_shunt[7] a_10452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X4369 a_34396_40008# a_34308_40052# vss vss nmos_6p0 w=0.82u l=1u
X4370 a_13252_33780# cap_shunt_n a_13460_34264# vdd pmos_6p0 w=1.2u l=0.5u
X4371 a_20328_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4372 a_3640_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4373 a_26108_45847# a_26020_45944# vss vss nmos_6p0 w=0.82u l=1u
X4374 a_26376_39268# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4375 vss cap_series_gyn a_17808_7908# vss nmos_6p0 w=0.82u l=0.6u
X4376 a_3172_16532# cap_shunt_p a_3380_17016# vdd pmos_6p0 w=1.2u l=0.5u
X4377 a_29580_49416# a_29492_49460# vss vss nmos_6p0 w=0.82u l=1u
X4378 a_6740_53080# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4379 vdd tune_series_gy[4] a_25572_8692# vdd pmos_6p0 w=1.2u l=0.5u
X4380 a_28484_29076# cap_shunt_p a_28692_29560# vdd pmos_6p0 w=1.2u l=0.5u
X4381 a_34516_4834# cap_series_gygyp a_34308_5180# vdd pmos_6p0 w=1.2u l=0.5u
X4382 a_34348_9884# cap_series_gygyn a_34536_9884# vdd pmos_6p0 w=1.2u l=0.5u
X4383 a_2708_14242# cap_shunt_n a_3640_14180# vss nmos_6p0 w=0.82u l=0.6u
X4384 vss tune_shunt[7] a_17828_26424# vss nmos_6p0 w=0.51u l=0.6u
X4385 vdd tune_series_gy[4] a_15492_9884# vdd pmos_6p0 w=1.2u l=0.5u
X4386 a_13252_30644# cap_shunt_n a_13460_31128# vdd pmos_6p0 w=1.2u l=0.5u
X4387 vss cap_series_gyp a_8968_6340# vss nmos_6p0 w=0.82u l=0.6u
X4388 vdd a_16924_50984# a_16836_51028# vdd pmos_6p0 w=1.22u l=1u
X4389 a_19724_47415# a_19636_47512# vss vss nmos_6p0 w=0.82u l=1u
X4390 a_29580_46280# a_29492_46324# vss vss nmos_6p0 w=0.82u l=1u
X4391 vss cap_shunt_p a_15120_50244# vss nmos_6p0 w=0.82u l=0.6u
X4392 a_14580_45240# cap_shunt_p a_14372_44756# vdd pmos_6p0 w=1.2u l=0.5u
X4393 vss cap_shunt_p a_27888_35832# vss nmos_6p0 w=0.82u l=0.6u
X4394 a_28692_4472# cap_series_gyp a_28484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X4395 a_24660_18946# cap_series_gyn a_26376_18884# vss nmos_6p0 w=0.82u l=0.6u
X4396 a_7672_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4397 a_20740_34264# cap_shunt_n a_21672_34264# vss nmos_6p0 w=0.82u l=0.6u
X4398 vdd tune_series_gy[3] a_25572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X4399 vdd tune_series_gy[4] a_15492_6748# vdd pmos_6p0 w=1.2u l=0.5u
X4400 a_34348_6748# cap_series_gygyp a_34536_6748# vdd pmos_6p0 w=1.2u l=0.5u
X4401 a_2708_11106# cap_shunt_n a_3640_11044# vss nmos_6p0 w=0.82u l=0.6u
X4402 a_22524_52552# a_22436_52596# vss vss nmos_6p0 w=0.82u l=1u
X4403 a_30364_47415# a_30276_47512# vss vss nmos_6p0 w=0.82u l=1u
X4404 a_36384_40836# cap_shunt_gyp a_36384_41240# vdd pmos_6p0 w=1.215u l=0.5u
X4405 a_10660_36194# cap_shunt_n a_10452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X4406 a_12580_49460# cap_shunt_n a_12788_49944# vdd pmos_6p0 w=1.2u l=0.5u
X4407 vss tune_shunt[5] a_17828_46808# vss nmos_6p0 w=0.51u l=0.6u
X4408 a_33500_48983# a_33412_49080# vss vss nmos_6p0 w=0.82u l=1u
X4409 a_29492_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4410 vdd a_5612_25463# a_5524_25560# vdd pmos_6p0 w=1.22u l=1u
X4411 a_15356_49416# a_15268_49460# vss vss nmos_6p0 w=0.82u l=1u
X4412 a_32444_11452# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4413 vss tune_series_gy[5] a_21748_12674# vss nmos_6p0 w=0.51u l=0.6u
X4414 a_24660_15810# cap_series_gyn a_26376_15748# vss nmos_6p0 w=0.82u l=0.6u
X4415 a_20740_31128# cap_shunt_n a_21672_31128# vss nmos_6p0 w=0.82u l=0.6u
X4416 a_17828_29560# cap_shunt_n a_18760_29560# vss nmos_6p0 w=0.82u l=0.6u
X4417 a_32612_28354# cap_shunt_p a_32404_28700# vdd pmos_6p0 w=1.2u l=0.5u
X4418 a_17620_27508# cap_shunt_n a_17828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X4419 a_1924_3266# cap_shunt_n a_1716_3612# vdd pmos_6p0 w=1.2u l=0.5u
X4420 a_27228_34871# a_27140_34968# vss vss nmos_6p0 w=0.82u l=1u
X4421 vss tune_series_gy[2] a_7768_6748# vss nmos_6p0 w=0.51u l=0.6u
X4422 a_10660_33058# cap_shunt_n a_10452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X4423 a_2708_50306# cap_shunt_n a_2500_50652# vdd pmos_6p0 w=1.2u l=0.5u
X4424 a_16708_44034# cap_shunt_p a_16500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X4425 vdd a_9644_41576# a_9556_41620# vdd pmos_6p0 w=1.22u l=1u
X4426 vdd a_5612_22327# a_5524_22424# vdd pmos_6p0 w=1.22u l=1u
X4427 a_21540_8316# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4428 a_17828_26424# cap_shunt_n a_18760_26424# vss nmos_6p0 w=0.82u l=0.6u
X4429 vdd a_6060_45847# a_5972_45944# vdd pmos_6p0 w=1.22u l=1u
X4430 a_2500_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4431 a_27228_31735# a_27140_31832# vss vss nmos_6p0 w=0.82u l=1u
X4432 a_19732_7608# cap_series_gyp a_20664_7608# vss nmos_6p0 w=0.82u l=0.6u
X4433 a_9316_50306# cap_shunt_p a_9108_50652# vdd pmos_6p0 w=1.2u l=0.5u
X4434 a_25780_29560# cap_shunt_p a_25572_29076# vdd pmos_6p0 w=1.2u l=0.5u
X4435 vss cap_series_gygyn a_32040_18884# vss nmos_6p0 w=0.82u l=0.6u
X4436 a_16708_40898# cap_shunt_n a_16500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X4437 a_1924_4472# cap_shunt_p a_3640_4472# vss nmos_6p0 w=0.82u l=0.6u
X4438 vdd tune_shunt[6] a_16500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X4439 a_9464_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4440 a_9668_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4441 vdd a_6060_42711# a_5972_42808# vdd pmos_6p0 w=1.22u l=1u
X4442 a_10452_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4443 a_32632_14588# cap_series_gyp a_32444_14588# vdd pmos_6p0 w=1.2u l=0.5u
X4444 a_20396_50551# a_20308_50648# vss vss nmos_6p0 w=0.82u l=1u
X4445 a_16476_38440# a_16388_38484# vss vss nmos_6p0 w=0.82u l=1u
X4446 a_31024_32996# cap_shunt_p a_29700_33058# vss nmos_6p0 w=0.82u l=0.6u
X4447 a_35344_7908# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X4448 a_21748_6402# cap_series_gyn a_22680_6340# vss nmos_6p0 w=0.82u l=0.6u
X4449 a_37420_9783# a_37332_9880# vss vss nmos_6p0 w=0.82u l=1u
X4450 a_18760_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4451 vss cap_shunt_n a_11984_29860# vss nmos_6p0 w=0.82u l=0.6u
X4452 a_33500_7080# a_33412_7124# vss vss nmos_6p0 w=0.82u l=1u
X4453 a_9668_11828# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4454 a_9876_20152# cap_shunt_p a_9668_19668# vdd pmos_6p0 w=1.2u l=0.5u
X4455 a_15120_48676# cap_shunt_n a_13796_48738# vss nmos_6p0 w=0.82u l=0.6u
X4456 a_36624_17316# cap_series_gygyn a_34516_17378# vss nmos_6p0 w=0.82u l=0.6u
X4457 vdd tune_shunt[7] a_13588_27132# vdd pmos_6p0 w=1.2u l=0.5u
X4458 vdd a_20620_17623# a_20532_17720# vdd pmos_6p0 w=1.22u l=1u
X4459 a_28692_40536# cap_shunt_p a_28484_40052# vdd pmos_6p0 w=1.2u l=0.5u
X4460 a_22848_3204# cap_series_gyp a_21524_3266# vss nmos_6p0 w=0.82u l=0.6u
X4461 a_6740_37400# cap_shunt_n a_6532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X4462 a_25780_38968# cap_shunt_p a_25572_38484# vdd pmos_6p0 w=1.2u l=0.5u
X4463 vss cap_shunt_n a_11984_26724# vss nmos_6p0 w=0.82u l=0.6u
X4464 vss cap_shunt_p a_4032_43972# vss nmos_6p0 w=0.82u l=0.6u
X4465 vss cap_shunt_n a_15568_37400# vss nmos_6p0 w=0.82u l=0.6u
X4466 a_13588_14588# cap_shunt_p a_13796_14242# vdd pmos_6p0 w=1.2u l=0.5u
X4467 a_19524_7124# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4468 a_15804_47848# a_15716_47892# vss vss nmos_6p0 w=0.82u l=1u
X4469 vdd a_23308_40008# a_23220_40052# vdd pmos_6p0 w=1.22u l=1u
X4470 a_13252_24372# cap_shunt_n a_13460_24856# vdd pmos_6p0 w=1.2u l=0.5u
X4471 a_1716_7124# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4472 a_35880_36916# cap_series_gygyp a_35692_36916# vdd pmos_6p0 w=1.2u l=0.5u
X4473 a_18612_12674# cap_series_gyn a_18404_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4474 vss cap_shunt_p a_27888_29560# vss nmos_6p0 w=0.82u l=0.6u
X4475 a_25780_35832# cap_shunt_p a_25572_35348# vdd pmos_6p0 w=1.2u l=0.5u
X4476 vss cap_shunt_p a_4032_40836# vss nmos_6p0 w=0.82u l=0.6u
X4477 vss cap_shunt_p a_7616_51512# vss nmos_6p0 w=0.82u l=0.6u
X4478 a_6532_14964# cap_shunt_p a_6740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X4479 vss tune_shunt[7] a_17828_17016# vss nmos_6p0 w=0.51u l=0.6u
X4480 a_13796_45602# cap_shunt_p a_13588_45948# vdd pmos_6p0 w=1.2u l=0.5u
X4481 vdd a_36524_33303# a_36436_33400# vdd pmos_6p0 w=1.22u l=1u
X4482 a_13252_21236# cap_shunt_n a_13460_21720# vdd pmos_6p0 w=1.2u l=0.5u
X4483 vss tune_shunt[6] a_25780_32696# vss nmos_6p0 w=0.51u l=0.6u
X4484 a_16576_3204# cap_series_gyn a_14468_3266# vss nmos_6p0 w=0.82u l=0.6u
X4485 a_13796_12674# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4486 a_6292_17378# cap_shunt_p a_6084_17724# vdd pmos_6p0 w=1.2u l=0.5u
X4487 a_14784_35832# cap_shunt_n a_13460_35832# vss nmos_6p0 w=0.82u l=0.6u
X4488 a_18492_50984# a_18404_51028# vss vss nmos_6p0 w=0.82u l=1u
X4489 vss cap_shunt_p a_27888_26424# vss nmos_6p0 w=0.82u l=0.6u
X4490 a_21524_4472# cap_series_gyn a_21316_3988# vdd pmos_6p0 w=1.2u l=0.5u
X4491 vdd tune_shunt[6] a_2500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X4492 a_12788_12312# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4493 a_25572_13396# cap_series_gyn a_25780_13880# vdd pmos_6p0 w=1.2u l=0.5u
X4494 a_25572_43188# cap_shunt_p a_25780_43672# vdd pmos_6p0 w=1.2u l=0.5u
X4495 a_27228_28599# a_27140_28696# vss vss nmos_6p0 w=0.82u l=1u
X4496 a_6532_11828# cap_shunt_p a_6740_12312# vdd pmos_6p0 w=1.2u l=0.5u
X4497 a_19732_13880# cap_series_gyn a_19524_13396# vdd pmos_6p0 w=1.2u l=0.5u
X4498 vdd a_31260_18056# a_31172_18100# vdd pmos_6p0 w=1.22u l=1u
X4499 a_3172_49460# cap_shunt_p a_3380_49944# vdd pmos_6p0 w=1.2u l=0.5u
X4500 vdd a_33948_25896# a_33860_25940# vdd pmos_6p0 w=1.22u l=1u
X4501 a_2708_44034# cap_shunt_p a_2500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X4502 a_27104_27992# cap_shunt_p a_25780_27992# vss nmos_6p0 w=0.82u l=0.6u
X4503 a_10660_26786# cap_shunt_n a_10452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X4504 a_13588_23996# cap_shunt_n a_13796_23650# vdd pmos_6p0 w=1.2u l=0.5u
X4505 vss cap_series_gyp a_31024_14180# vss nmos_6p0 w=0.82u l=0.6u
X4506 vdd a_5612_16055# a_5524_16152# vdd pmos_6p0 w=1.22u l=1u
X4507 a_23308_32168# a_23220_32212# vss vss nmos_6p0 w=0.82u l=1u
X4508 vdd a_27340_53687# a_27252_53784# vdd pmos_6p0 w=1.22u l=1u
X4509 a_22412_53687# a_22324_53784# vss vss nmos_6p0 w=0.82u l=1u
X4510 vdd a_6060_39575# a_5972_39672# vdd pmos_6p0 w=1.22u l=1u
X4511 vdd tune_shunt[7] a_2500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X4512 a_18724_6040# cap_series_gyn a_18516_5556# vdd pmos_6p0 w=1.2u l=0.5u
X4513 a_21748_17378# cap_shunt_p a_21540_17724# vdd pmos_6p0 w=1.2u l=0.5u
X4514 a_14372_43188# cap_shunt_n a_14580_43672# vdd pmos_6p0 w=1.2u l=0.5u
X4515 a_2500_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4516 a_27228_25463# a_27140_25560# vss vss nmos_6p0 w=0.82u l=1u
X4517 a_16408_6040# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4518 a_27104_24856# cap_shunt_p a_25780_24856# vss nmos_6p0 w=0.82u l=0.6u
X4519 vdd a_33948_22760# a_33860_22804# vdd pmos_6p0 w=1.22u l=1u
X4520 a_2708_40898# cap_shunt_p a_2500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X4521 vss tune_shunt[6] a_20740_37400# vss nmos_6p0 w=0.51u l=0.6u
X4522 vdd a_9644_32168# a_9556_32212# vdd pmos_6p0 w=1.22u l=1u
X4523 vss cap_series_gyp a_31024_11044# vss nmos_6p0 w=0.82u l=0.6u
X4524 vdd a_5612_12919# a_5524_13016# vdd pmos_6p0 w=1.22u l=1u
X4525 a_11780_6040# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X4526 a_11612_8692# cap_series_gyp a_11800_8692# vdd pmos_6p0 w=1.2u l=0.5u
X4527 a_17828_17016# cap_shunt_p a_18760_17016# vss nmos_6p0 w=0.82u l=0.6u
X4528 a_11212_53687# a_11124_53784# vss vss nmos_6p0 w=0.82u l=1u
X4529 vdd a_27340_50551# a_27252_50648# vdd pmos_6p0 w=1.22u l=1u
X4530 a_22412_50551# a_22324_50648# vss vss nmos_6p0 w=0.82u l=1u
X4531 vdd a_6060_36439# a_5972_36536# vdd pmos_6p0 w=1.22u l=1u
X4532 a_2500_13020# cap_shunt_n a_2708_12674# vdd pmos_6p0 w=1.2u l=0.5u
X4533 a_2500_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4534 a_19152_32696# cap_shunt_n a_17828_32696# vss nmos_6p0 w=0.82u l=0.6u
X4535 a_7792_7908# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4536 a_27104_9176# cap_series_gyp a_25780_9176# vss nmos_6p0 w=0.82u l=0.6u
X4537 a_2932_9176# cap_shunt_n a_3864_9176# vss nmos_6p0 w=0.82u l=0.6u
X4538 vss cap_series_gyn a_16016_10744# vss nmos_6p0 w=0.82u l=0.6u
X4539 a_21748_42466# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4540 a_9644_27464# a_9556_27508# vss vss nmos_6p0 w=0.82u l=1u
X4541 vdd a_11996_17623# a_11908_17720# vdd pmos_6p0 w=1.22u l=1u
X4542 a_17828_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4543 vdd a_12780_54120# a_12692_54164# vdd pmos_6p0 w=1.22u l=1u
X4544 a_18940_52552# a_18852_52596# vss vss nmos_6p0 w=0.82u l=1u
X4545 a_31024_23588# cap_shunt_p a_29700_23650# vss nmos_6p0 w=0.82u l=0.6u
X4546 a_24660_7970# cap_series_gyp a_24452_8316# vdd pmos_6p0 w=1.2u l=0.5u
X4547 a_11984_45540# cap_shunt_n a_10660_45602# vss nmos_6p0 w=0.82u l=0.6u
X4548 a_35880_24372# cap_series_gygyp a_36688_24856# vss nmos_6p0 w=0.82u l=0.6u
X4549 a_1692_50984# a_1604_51028# vss vss nmos_6p0 w=0.82u l=1u
X4550 a_15120_39268# cap_shunt_n a_13796_39330# vss nmos_6p0 w=0.82u l=0.6u
X4551 a_16708_44034# cap_shunt_p a_16500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X4552 a_9644_24328# a_9556_24372# vss vss nmos_6p0 w=0.82u l=1u
X4553 vdd a_37420_55255# a_37332_55352# vdd pmos_6p0 w=1.22u l=1u
X4554 vss tune_shunt[4] a_16708_48738# vss nmos_6p0 w=0.51u l=0.6u
X4555 a_21524_4472# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X4556 a_12788_18584# cap_shunt_p a_12580_18100# vdd pmos_6p0 w=1.2u l=0.5u
X4557 a_11984_42404# cap_shunt_n a_10660_42466# vss nmos_6p0 w=0.82u l=0.6u
X4558 a_23756_47415# a_23668_47512# vss vss nmos_6p0 w=0.82u l=1u
X4559 a_11572_3988# cap_series_gyp a_11780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X4560 a_9316_50306# cap_shunt_p a_9108_50652# vdd pmos_6p0 w=1.2u l=0.5u
X4561 a_7748_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4562 a_25780_29560# cap_shunt_p a_25572_29076# vdd pmos_6p0 w=1.2u l=0.5u
X4563 a_6740_27992# cap_shunt_n a_6532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X4564 vdd tune_shunt[7] a_12580_14964# vdd pmos_6p0 w=1.2u l=0.5u
X4565 a_13796_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4566 a_24452_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4567 vss tune_shunt[7] a_13460_34264# vss nmos_6p0 w=0.51u l=0.6u
X4568 a_25780_4472# cap_shunt_p a_26712_4472# vss nmos_6p0 w=0.82u l=0.6u
X4569 vss cap_shunt_n a_4032_34564# vss nmos_6p0 w=0.82u l=0.6u
X4570 a_5388_7080# a_5300_7124# vss vss nmos_6p0 w=0.82u l=1u
X4571 a_23464_9476# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4572 vdd a_37420_52119# a_37332_52216# vdd pmos_6p0 w=1.22u l=1u
X4573 a_16708_40898# cap_shunt_n a_16500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X4574 a_13796_39330# cap_shunt_n a_13588_39676# vdd pmos_6p0 w=1.2u l=0.5u
X4575 a_14460_11351# a_14372_11448# vss vss nmos_6p0 w=0.82u l=1u
X4576 vdd a_11324_55688# a_11236_55732# vdd pmos_6p0 w=1.22u l=1u
X4577 a_14784_29560# cap_shunt_n a_13460_29560# vss nmos_6p0 w=0.82u l=0.6u
X4578 a_36652_47108# cap_shunt_gyp a_36384_47108# vss nmos_6p0 w=0.82u l=0.6u
X4579 vdd tune_shunt[7] a_12580_11828# vdd pmos_6p0 w=1.2u l=0.5u
X4580 a_32632_14588# cap_series_gyp a_32444_14588# vdd pmos_6p0 w=1.2u l=0.5u
X4581 a_29692_41576# a_29604_41620# vss vss nmos_6p0 w=0.82u l=1u
X4582 a_24452_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4583 vss tune_shunt[7] a_13460_31128# vss nmos_6p0 w=0.51u l=0.6u
X4584 vss tune_shunt[5] a_3828_21720# vss nmos_6p0 w=0.51u l=0.6u
X4585 a_1924_3266# cap_shunt_n a_1716_3612# vdd pmos_6p0 w=1.2u l=0.5u
X4586 vss cap_shunt_p a_4032_31428# vss nmos_6p0 w=0.82u l=0.6u
X4587 vss cap_shunt_gyp a_36652_45540# vss nmos_6p0 w=0.82u l=0.6u
X4588 a_17828_48376# cap_shunt_p a_17620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X4589 a_18516_5556# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4590 a_9876_20152# cap_shunt_p a_9668_19668# vdd pmos_6p0 w=1.2u l=0.5u
X4591 a_14784_26424# cap_shunt_n a_13460_26424# vss nmos_6p0 w=0.82u l=0.6u
X4592 vss tune_shunt[7] a_25780_23288# vss nmos_6p0 w=0.51u l=0.6u
X4593 a_3620_25940# cap_shunt_p a_3828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X4594 a_24660_12674# cap_series_gyn a_24452_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4595 vss cap_series_gyp a_27888_17016# vss nmos_6p0 w=0.82u l=0.6u
X4596 a_2708_18946# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4597 vss cap_series_gyn a_17024_9476# vss nmos_6p0 w=0.82u l=0.6u
X4598 vdd tune_shunt[7] a_2500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X4599 a_25572_7124# cap_series_gyn a_25780_7608# vdd pmos_6p0 w=1.2u l=0.5u
X4600 vss cap_series_gyp a_23072_4772# vss nmos_6p0 w=0.82u l=0.6u
X4601 a_3248_4472# cap_shunt_p a_1924_4472# vss nmos_6p0 w=0.82u l=0.6u
X4602 vss cap_shunt_gyn a_36652_42404# vss nmos_6p0 w=0.82u l=0.6u
X4603 vdd tune_series_gygy[3] a_34348_8316# vdd pmos_6p0 w=1.2u l=0.5u
X4604 vdd a_33948_16488# a_33860_16532# vdd pmos_6p0 w=1.22u l=1u
X4605 a_27104_18584# cap_series_gyn a_25780_18584# vss nmos_6p0 w=0.82u l=0.6u
X4606 a_17828_45240# cap_shunt_p a_17620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X4607 a_15492_8316# cap_series_gyn a_15700_7970# vdd pmos_6p0 w=1.2u l=0.5u
X4608 a_21740_55688# a_21652_55732# vss vss nmos_6p0 w=0.82u l=1u
X4609 a_11200_53080# cap_shunt_n a_9876_53080# vss nmos_6p0 w=0.82u l=0.6u
X4610 a_14908_8215# a_14820_8312# vss vss nmos_6p0 w=0.82u l=1u
X4611 a_13588_14588# cap_shunt_p a_13796_14242# vdd pmos_6p0 w=1.2u l=0.5u
X4612 vss cap_shunt_n a_19152_46808# vss nmos_6p0 w=0.82u l=0.6u
X4613 a_3620_22804# cap_shunt_p a_3828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X4614 a_23308_22760# a_23220_22804# vss vss nmos_6p0 w=0.82u l=1u
X4615 vdd a_7516_54120# a_7428_54164# vdd pmos_6p0 w=1.22u l=1u
X4616 a_19656_6040# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4617 a_17620_36916# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4618 a_2500_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4619 vdd tune_shunt[5] a_2500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X4620 vdd tune_shunt[7] a_32404_30268# vdd pmos_6p0 w=1.2u l=0.5u
X4621 a_15492_5180# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4622 a_27104_15448# cap_series_gyp a_25780_15448# vss nmos_6p0 w=0.82u l=0.6u
X4623 a_19936_7908# cap_series_gyp a_18612_7970# vss nmos_6p0 w=0.82u l=0.6u
X4624 vss cap_series_gyn a_30920_12612# vss nmos_6p0 w=0.82u l=0.6u
X4625 a_20740_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4626 a_15356_52119# a_15268_52216# vss vss nmos_6p0 w=0.82u l=1u
X4627 a_3828_21720# cap_shunt_p a_4760_21720# vss nmos_6p0 w=0.82u l=0.6u
X4628 vdd a_34396_36872# a_34308_36916# vdd pmos_6p0 w=1.22u l=1u
X4629 a_6532_14964# cap_shunt_p a_6740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X4630 a_13796_45602# cap_shunt_p a_13588_45948# vdd pmos_6p0 w=1.2u l=0.5u
X4631 vdd a_6060_27031# a_5972_27128# vdd pmos_6p0 w=1.22u l=1u
X4632 a_19152_23288# cap_shunt_n a_17828_23288# vss nmos_6p0 w=0.82u l=0.6u
X4633 a_21748_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4634 vss cap_shunt_p a_30800_37400# vss nmos_6p0 w=0.82u l=0.6u
X4635 a_27676_44279# a_27588_44376# vss vss nmos_6p0 w=0.82u l=1u
X4636 a_6196_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4637 vdd tune_shunt[6] a_2500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X4638 a_1692_44712# a_1604_44756# vss vss nmos_6p0 w=0.82u l=1u
X4639 a_25572_43188# cap_shunt_p a_25780_43672# vdd pmos_6p0 w=1.2u l=0.5u
X4640 a_6532_11828# cap_shunt_p a_6740_12312# vdd pmos_6p0 w=1.2u l=0.5u
X4641 a_35880_18100# cap_series_gygyn a_36688_18584# vss nmos_6p0 w=0.82u l=0.6u
X4642 vss tune_shunt[3] a_2708_9538# vss nmos_6p0 w=0.51u l=0.6u
X4643 a_21748_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4644 a_27676_41143# a_27588_41240# vss vss nmos_6p0 w=0.82u l=1u
X4645 a_23464_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4646 a_25984_9476# cap_series_gyn a_24660_9538# vss nmos_6p0 w=0.82u l=0.6u
X4647 vdd tune_shunt[7] a_2500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X4648 a_21748_17378# cap_shunt_p a_21540_17724# vdd pmos_6p0 w=1.2u l=0.5u
X4649 vdd a_22524_49416# a_22436_49460# vdd pmos_6p0 w=1.22u l=1u
X4650 a_14372_43188# cap_shunt_n a_14580_43672# vdd pmos_6p0 w=1.2u l=0.5u
X4651 a_1692_41576# a_1604_41620# vss vss nmos_6p0 w=0.82u l=1u
X4652 a_11984_36132# cap_shunt_n a_10660_36194# vss nmos_6p0 w=0.82u l=0.6u
X4653 a_17828_35832# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4654 a_35880_14964# cap_series_gygyn a_36688_15448# vss nmos_6p0 w=0.82u l=0.6u
X4655 vdd a_17596_55255# a_17508_55352# vdd pmos_6p0 w=1.22u l=1u
X4656 vss cap_shunt_n a_4032_28292# vss nmos_6p0 w=0.82u l=0.6u
X4657 a_3828_45240# cap_shunt_p a_5544_45240# vss nmos_6p0 w=0.82u l=0.6u
X4658 a_3380_18584# cap_shunt_p a_3172_18100# vdd pmos_6p0 w=1.2u l=0.5u
X4659 a_14260_3612# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4660 a_36296_6040# cap_series_gygyn a_35880_5556# vss nmos_6p0 w=0.82u l=0.6u
X4661 vdd a_32604_10216# a_32516_10260# vdd pmos_6p0 w=1.22u l=1u
X4662 vdd a_24652_18056# a_24564_18100# vdd pmos_6p0 w=1.22u l=1u
X4663 a_8300_55688# a_8212_55732# vss vss nmos_6p0 w=0.82u l=1u
X4664 vdd a_17596_52119# a_17508_52216# vdd pmos_6p0 w=1.22u l=1u
X4665 a_13000_7608# cap_series_gyp a_11800_7124# vss nmos_6p0 w=0.82u l=0.6u
X4666 a_35880_3988# tune_series_gygy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X4667 vss cap_shunt_p a_4032_25156# vss nmos_6p0 w=0.82u l=0.6u
X4668 a_24452_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4669 a_3828_42104# cap_shunt_p a_5544_42104# vss nmos_6p0 w=0.82u l=0.6u
X4670 a_15804_53687# a_15716_53784# vss vss nmos_6p0 w=0.82u l=1u
X4671 vdd a_34844_38440# a_34756_38484# vdd pmos_6p0 w=1.22u l=1u
X4672 a_18612_9538# cap_series_gyp a_19544_9476# vss nmos_6p0 w=0.82u l=0.6u
X4673 vdd a_30812_19191# a_30724_19288# vdd pmos_6p0 w=1.22u l=1u
X4674 a_9876_49944# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4675 a_6740_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4676 a_14692_7608# cap_series_gyp a_15624_7608# vss nmos_6p0 w=0.82u l=0.6u
X4677 a_24660_4834# cap_series_gyp a_25592_4772# vss nmos_6p0 w=0.82u l=0.6u
X4678 a_18724_6040# cap_series_gyn a_18516_5556# vdd pmos_6p0 w=1.2u l=0.5u
X4679 a_5636_11452# cap_shunt_n a_5844_11106# vdd pmos_6p0 w=1.2u l=0.5u
X4680 a_9428_20514# cap_shunt_p a_11144_20452# vss nmos_6p0 w=0.82u l=0.6u
X4681 a_24452_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4682 vdd tune_shunt[5] a_2500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X4683 vss tune_shunt[2] a_1924_7970# vss nmos_6p0 w=0.51u l=0.6u
X4684 a_17640_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4685 vss tune_shunt[6] a_3828_35832# vss nmos_6p0 w=0.51u l=0.6u
X4686 a_37420_23895# a_37332_23992# vss vss nmos_6p0 w=0.82u l=1u
X4687 a_17828_38968# cap_shunt_n a_17620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X4688 a_10452_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4689 a_21748_29922# cap_shunt_n a_22680_29860# vss nmos_6p0 w=0.82u l=0.6u
X4690 a_31624_8316# cap_series_gygyn a_32432_7908# vss nmos_6p0 w=0.82u l=0.6u
X4691 a_30364_8215# a_30276_8312# vss vss nmos_6p0 w=0.82u l=1u
X4692 a_26556_45847# a_26468_45944# vss vss nmos_6p0 w=0.82u l=1u
X4693 a_6532_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4694 a_14460_5079# a_14372_5176# vss vss nmos_6p0 w=0.82u l=1u
X4695 vss cap_shunt_n a_12656_27992# vss nmos_6p0 w=0.82u l=0.6u
X4696 vss cap_series_gyn a_25984_12612# vss nmos_6p0 w=0.82u l=0.6u
X4697 vdd tune_shunt[7] a_2500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X4698 a_17808_6340# cap_series_gyp a_15700_6402# vss nmos_6p0 w=0.82u l=0.6u
X4699 vss tune_shunt[2] a_1924_4834# vss nmos_6p0 w=0.51u l=0.6u
X4700 vss tune_series_gygy[5] a_34516_18946# vss nmos_6p0 w=0.51u l=0.6u
X4701 a_20740_40536# cap_shunt_p a_20532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X4702 vdd a_2140_13352# a_2052_13396# vdd pmos_6p0 w=1.22u l=1u
X4703 vdd a_17708_50551# a_17620_50648# vdd pmos_6p0 w=1.22u l=1u
X4704 a_3828_43672# cap_shunt_p a_3620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X4705 a_17828_35832# cap_shunt_n a_17620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X4706 a_10452_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4707 a_21540_34972# cap_shunt_p a_21748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X4708 a_21748_26786# cap_shunt_n a_22680_26724# vss nmos_6p0 w=0.82u l=0.6u
X4709 a_21748_9538# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4710 a_13796_39330# cap_shunt_n a_13588_39676# vdd pmos_6p0 w=1.2u l=0.5u
X4711 a_17620_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4712 vss cap_shunt_n a_12656_24856# vss nmos_6p0 w=0.82u l=0.6u
X4713 a_5096_49944# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4714 vdd a_33612_23895# a_33524_23992# vdd pmos_6p0 w=1.22u l=1u
X4715 vss tune_shunt[7] a_13460_21720# vss nmos_6p0 w=0.51u l=0.6u
X4716 vss cap_series_gyp a_13000_7608# vss nmos_6p0 w=0.82u l=0.6u
X4717 a_21540_31836# cap_shunt_n a_21748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X4718 vss tune_series_gy[4] a_14692_9176# vss nmos_6p0 w=0.51u l=0.6u
X4719 a_10808_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4720 a_22972_52552# a_22884_52596# vss vss nmos_6p0 w=0.82u l=1u
X4721 a_14484_7124# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4722 vss tune_series_gy[5] a_25780_13880# vss nmos_6p0 w=0.51u l=0.6u
X4723 vdd a_3932_53687# a_3844_53784# vdd pmos_6p0 w=1.22u l=1u
X4724 a_27676_34871# a_27588_34968# vss vss nmos_6p0 w=0.82u l=1u
X4725 a_24660_12674# cap_series_gyn a_24452_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4726 a_13460_38968# cap_shunt_n a_15176_38968# vss nmos_6p0 w=0.82u l=0.6u
X4727 a_10808_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4728 a_6084_19292# cap_shunt_p a_6292_18946# vdd pmos_6p0 w=1.2u l=0.5u
X4729 a_35740_50984# a_35652_51028# vss vss nmos_6p0 w=0.82u l=1u
X4730 a_22680_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4731 vdd tune_shunt[7] a_2500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X4732 a_17828_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4733 vss tune_series_gy[4] a_25780_10744# vss nmos_6p0 w=0.51u l=0.6u
X4734 a_31904_45540# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4735 a_27676_31735# a_27588_31832# vss vss nmos_6p0 w=0.82u l=1u
X4736 vdd a_32604_8648# a_32516_8692# vdd pmos_6p0 w=1.22u l=1u
X4737 a_6084_16156# cap_shunt_p a_6292_15810# vdd pmos_6p0 w=1.2u l=0.5u
X4738 a_9876_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4739 vdd tune_shunt[5] a_2500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X4740 a_14692_4472# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X4741 vdd tune_shunt[6] a_24452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X4742 a_17828_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4743 a_32716_50984# a_32628_51028# vss vss nmos_6p0 w=0.82u l=1u
X4744 vdd a_6508_38007# a_6420_38104# vdd pmos_6p0 w=1.22u l=1u
X4745 a_33500_3511# a_33412_3608# vss vss nmos_6p0 w=0.82u l=1u
X4746 a_24452_19292# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4747 a_4816_32996# cap_shunt_p a_2708_33058# vss nmos_6p0 w=0.82u l=0.6u
X4748 vdd a_32604_5512# a_32516_5556# vdd pmos_6p0 w=1.22u l=1u
X4749 vss cap_shunt_p a_31808_29860# vss nmos_6p0 w=0.82u l=0.6u
X4750 a_13340_50984# a_13252_51028# vss vss nmos_6p0 w=0.82u l=1u
X4751 a_10340_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4752 vdd tune_shunt[7] a_20532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X4753 a_18404_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4754 vss cap_shunt_p a_8400_18584# vss nmos_6p0 w=0.82u l=0.6u
X4755 a_6196_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4756 a_24452_16156# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4757 a_25780_43672# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X4758 a_25572_43188# cap_shunt_p a_25780_43672# vdd pmos_6p0 w=1.2u l=0.5u
X4759 vss tune_shunt[7] a_3828_29560# vss nmos_6p0 w=0.51u l=0.6u
X4760 vss cap_shunt_p a_31808_26724# vss nmos_6p0 w=0.82u l=0.6u
X4761 vdd a_18940_7080# a_18852_7124# vdd pmos_6p0 w=1.22u l=1u
X4762 a_11880_7908# cap_series_gyp a_10680_8316# vss nmos_6p0 w=0.82u l=0.6u
X4763 vdd tune_shunt[7] a_20532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X4764 vss cap_shunt_p a_11984_49944# vss nmos_6p0 w=0.82u l=0.6u
X4765 a_19524_7124# cap_series_gyp a_19732_7608# vdd pmos_6p0 w=1.2u l=0.5u
X4766 a_5844_11106# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X4767 a_29532_13020# cap_series_gyn a_29720_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4768 a_29132_55688# a_29044_55732# vss vss nmos_6p0 w=0.82u l=1u
X4769 a_14580_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4770 a_25780_40536# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4771 a_17640_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4772 vss tune_shunt[7] a_3828_26424# vss nmos_6p0 w=0.51u l=0.6u
X4773 a_10452_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4774 a_17828_29560# cap_shunt_n a_17620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X4775 vdd a_23756_40008# a_23668_40052# vdd pmos_6p0 w=1.22u l=1u
X4776 vdd a_18940_49416# a_18852_49460# vdd pmos_6p0 w=1.22u l=1u
X4777 vss cap_shunt_n a_9072_37700# vss nmos_6p0 w=0.82u l=0.6u
X4778 a_35880_8692# cap_series_gygyn a_35692_8692# vdd pmos_6p0 w=1.2u l=0.5u
X4779 vdd a_20172_44279# a_20084_44376# vdd pmos_6p0 w=1.22u l=1u
X4780 vss tune_shunt[5] a_29700_37762# vss nmos_6p0 w=0.51u l=0.6u
X4781 a_14580_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4782 a_37444_38485# cap_shunt_gyp a_37632_38485# vdd pmos_6p0 w=1.215u l=0.5u
X4783 a_25236_3612# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4784 a_26108_55688# a_26020_55732# vss vss nmos_6p0 w=0.82u l=1u
X4785 a_6740_26424# cap_shunt_n a_6532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X4786 a_34980_44376# cap_shunt_gyn a_35168_44376# vdd pmos_6p0 w=1.215u l=0.5u
X4787 a_21540_25564# cap_shunt_n a_21748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X4788 a_21748_17378# cap_shunt_p a_22680_17316# vss nmos_6p0 w=0.82u l=0.6u
X4789 vdd tune_shunt[7] a_13588_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4790 a_26712_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4791 a_28124_38007# a_28036_38104# vss vss nmos_6p0 w=0.82u l=1u
X4792 a_35880_5556# cap_series_gygyn a_35692_5556# vdd pmos_6p0 w=1.2u l=0.5u
X4793 a_14728_50244# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4794 vss tune_shunt[6] a_29700_34626# vss nmos_6p0 w=0.51u l=0.6u
X4795 a_27676_28599# a_27588_28696# vss vss nmos_6p0 w=0.82u l=1u
X4796 a_6740_23288# cap_shunt_p a_6532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X4797 vss tune_series_gygy[2] a_34536_6748# vss nmos_6p0 w=0.51u l=0.6u
X4798 vdd tune_series_gy[2] a_14260_3612# vdd pmos_6p0 w=1.2u l=0.5u
X4799 a_5636_11452# cap_shunt_n a_5844_11106# vdd pmos_6p0 w=1.2u l=0.5u
X4800 a_21540_22428# cap_shunt_p a_21748_22082# vdd pmos_6p0 w=1.2u l=0.5u
X4801 a_16700_13352# a_16612_13396# vss vss nmos_6p0 w=0.82u l=1u
X4802 a_31904_45944# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X4803 vdd tune_shunt[5] a_2500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X4804 a_12580_13396# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4805 a_23756_32168# a_23668_32212# vss vss nmos_6p0 w=0.82u l=1u
X4806 a_22860_53687# a_22772_53784# vss vss nmos_6p0 w=0.82u l=1u
X4807 a_9876_48376# cap_shunt_p a_9668_47892# vdd pmos_6p0 w=1.2u l=0.5u
X4808 vdd tune_shunt[6] a_12580_47892# vdd pmos_6p0 w=1.2u l=0.5u
X4809 vdd a_37644_30600# a_37556_30644# vdd pmos_6p0 w=1.22u l=1u
X4810 a_21540_28700# cap_shunt_n a_21748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X4811 a_27676_25463# a_27588_25560# vss vss nmos_6p0 w=0.82u l=1u
X4812 a_15904_20452# cap_shunt_n a_13796_20514# vss nmos_6p0 w=0.82u l=0.6u
X4813 vdd a_3036_47848# a_2948_47892# vdd pmos_6p0 w=1.22u l=1u
X4814 vdd tune_shunt[7] a_2500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X4815 a_28692_4472# cap_series_gyp a_30408_4472# vss nmos_6p0 w=0.82u l=0.6u
X4816 a_20740_40536# cap_shunt_p a_20532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X4817 vss cap_series_gygyp a_36296_21720# vss nmos_6p0 w=0.82u l=0.6u
X4818 a_36720_50006# cap_shunt_gyp a_36720_49461# vdd pmos_6p0 w=1.215u l=0.5u
X4819 a_20740_46808# cap_shunt_p a_20532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X4820 a_9876_15448# cap_shunt_p a_9668_14964# vdd pmos_6p0 w=1.2u l=0.5u
X4821 a_11660_53687# a_11572_53784# vss vss nmos_6p0 w=0.82u l=1u
X4822 a_22860_50551# a_22772_50648# vss vss nmos_6p0 w=0.82u l=1u
X4823 vss tune_shunt[6] a_2708_37762# vss nmos_6p0 w=0.51u l=0.6u
X4824 a_21540_34972# cap_shunt_p a_21748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X4825 vss tune_series_gy[2] a_11780_6040# vss nmos_6p0 w=0.51u l=0.6u
X4826 a_25572_8692# cap_series_gyp a_25780_9176# vdd pmos_6p0 w=1.2u l=0.5u
X4827 a_31648_18884# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X4828 vdd a_3036_44712# a_2948_44756# vdd pmos_6p0 w=1.22u l=1u
X4829 a_15492_9884# cap_series_gyn a_15700_9538# vdd pmos_6p0 w=1.2u l=0.5u
X4830 a_17828_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4831 a_36720_46870# cap_shunt_gyp a_36720_46325# vdd pmos_6p0 w=1.215u l=0.5u
X4832 vdd tune_shunt[4] a_29492_23996# vdd pmos_6p0 w=1.2u l=0.5u
X4833 a_9876_12312# cap_shunt_p a_9668_11828# vdd pmos_6p0 w=1.2u l=0.5u
X4834 a_35292_36872# a_35204_36916# vss vss nmos_6p0 w=0.82u l=1u
X4835 vss tune_shunt[6] a_2708_34626# vss nmos_6p0 w=0.51u l=0.6u
X4836 a_21540_31836# cap_shunt_n a_21748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X4837 vdd a_23308_19624# a_23220_19668# vdd pmos_6p0 w=1.22u l=1u
X4838 vdd a_13564_53687# a_13476_53784# vdd pmos_6p0 w=1.22u l=1u
X4839 a_4816_23588# cap_shunt_p a_2708_23650# vss nmos_6p0 w=0.82u l=0.6u
X4840 a_32604_52119# a_32516_52216# vss vss nmos_6p0 w=0.82u l=1u
X4841 a_25572_5556# cap_series_gyp a_25780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X4842 a_19544_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4843 a_15492_6748# cap_series_gyp a_15700_6402# vdd pmos_6p0 w=1.2u l=0.5u
X4844 a_28692_18584# cap_series_gyp a_28484_18100# vdd pmos_6p0 w=1.2u l=0.5u
X4845 a_11424_47108# cap_shunt_p a_9316_47170# vss nmos_6p0 w=0.82u l=0.6u
X4846 a_30708_45540# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4847 vdd tune_shunt[4] a_3620_13396# vdd pmos_6p0 w=1.2u l=0.5u
X4848 vdd tune_shunt[4] a_20532_16532# vdd pmos_6p0 w=1.2u l=0.5u
X4849 a_25780_34264# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4850 a_6084_19292# cap_shunt_p a_6292_18946# vdd pmos_6p0 w=1.2u l=0.5u
X4851 a_20532_43188# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4852 vss cap_series_gyp a_8184_6340# vss nmos_6p0 w=0.82u l=0.6u
X4853 a_9332_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4854 vss tune_shunt[4] a_33732_34264# vss nmos_6p0 w=0.51u l=0.6u
X4855 vss cap_series_gyp a_31808_17316# vss nmos_6p0 w=0.82u l=0.6u
X4856 a_13796_50306# cap_shunt_p a_15512_50244# vss nmos_6p0 w=0.82u l=0.6u
X4857 a_25984_22020# cap_shunt_p a_24660_22082# vss nmos_6p0 w=0.82u l=0.6u
X4858 a_19936_38968# cap_shunt_n a_17828_38968# vss nmos_6p0 w=0.82u l=0.6u
X4859 a_7540_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4860 a_21748_7970# cap_series_gyp a_21540_8316# vdd pmos_6p0 w=1.2u l=0.5u
X4861 a_34480_47893# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X4862 a_3640_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4863 a_20740_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X4864 a_25780_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X4865 a_6760_5556# cap_series_gyp a_6572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X4866 a_6084_16156# cap_shunt_p a_6292_15810# vdd pmos_6p0 w=1.2u l=0.5u
X4867 a_3828_34264# cap_shunt_n a_3620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X4868 a_9420_53687# a_9332_53784# vss vss nmos_6p0 w=0.82u l=1u
X4869 a_10660_39330# cap_shunt_n a_12376_39268# vss nmos_6p0 w=0.82u l=0.6u
X4870 vss tune_shunt[4] a_33732_31128# vss nmos_6p0 w=0.51u l=0.6u
X4871 a_28692_38968# cap_shunt_n a_30408_38968# vss nmos_6p0 w=0.82u l=0.6u
X4872 vss cap_shunt_n a_5152_35832# vss nmos_6p0 w=0.82u l=0.6u
X4873 a_16528_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4874 a_21540_19292# cap_shunt_p a_21748_18946# vdd pmos_6p0 w=1.2u l=0.5u
X4875 vdd a_34844_55255# a_34756_55352# vdd pmos_6p0 w=1.22u l=1u
X4876 vdd a_11772_55688# a_11684_55732# vdd pmos_6p0 w=1.22u l=1u
X4877 a_3620_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4878 vss cap_shunt_n a_15904_37700# vss nmos_6p0 w=0.82u l=0.6u
X4879 vss tune_shunt[7] a_29700_28354# vss nmos_6p0 w=0.51u l=0.6u
X4880 a_2140_55255# a_2052_55352# vss vss nmos_6p0 w=0.82u l=1u
X4881 a_3640_40836# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4882 a_33524_35348# cap_shunt_n a_33732_35832# vdd pmos_6p0 w=1.2u l=0.5u
X4883 a_3828_31128# cap_shunt_n a_3620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X4884 a_8456_53080# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4885 a_24204_35304# a_24116_35348# vss vss nmos_6p0 w=0.82u l=1u
X4886 a_35692_7124# cap_series_gygyp a_35880_7124# vdd pmos_6p0 w=1.2u l=0.5u
X4887 a_2500_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4888 a_21540_16156# cap_series_gyn a_21748_15810# vdd pmos_6p0 w=1.2u l=0.5u
X4889 vdd a_34844_52119# a_34756_52216# vdd pmos_6p0 w=1.22u l=1u
X4890 a_26712_12312# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4891 a_13384_43672# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4892 a_3620_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4893 a_6628_12674# cap_shunt_p a_6420_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4894 a_8400_17016# cap_shunt_p a_6292_17016# vss nmos_6p0 w=0.82u l=0.6u
X4895 a_28484_18100# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4896 a_25572_18100# cap_series_gyn a_25780_18584# vdd pmos_6p0 w=1.2u l=0.5u
X4897 vss tune_shunt[7] a_29700_25218# vss nmos_6p0 w=0.51u l=0.6u
X4898 a_31624_19292# cap_series_gygyn a_32432_18884# vss nmos_6p0 w=0.82u l=0.6u
X4899 vdd tune_series_gygy[5] a_31436_20860# vdd pmos_6p0 w=1.2u l=0.5u
X4900 vdd a_27340_52552# a_27252_52596# vdd pmos_6p0 w=1.22u l=1u
X4901 vss tune_series_gy[5] a_22644_9176# vss nmos_6p0 w=0.51u l=0.6u
X4902 a_15904_14180# cap_shunt_p a_13796_14242# vss nmos_6p0 w=0.82u l=0.6u
X4903 a_16500_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4904 a_24660_44034# cap_shunt_p a_26376_43972# vss nmos_6p0 w=0.82u l=0.6u
X4905 a_29532_13020# cap_series_gyn a_29720_13020# vdd pmos_6p0 w=1.2u l=0.5u
X4906 a_24452_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4907 vdd a_2140_30167# a_2052_30264# vdd pmos_6p0 w=1.22u l=1u
X4908 a_30632_14180# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4909 a_16708_48738# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X4910 a_13384_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4911 a_15492_5180# cap_series_gyn a_15700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X4912 vdd a_7964_54120# a_7876_54164# vdd pmos_6p0 w=1.22u l=1u
X4913 a_23756_22760# a_23668_22804# vss vss nmos_6p0 w=0.82u l=1u
X4914 vdd a_24316_52552# a_24228_52596# vdd pmos_6p0 w=1.22u l=1u
X4915 a_10340_3612# cap_series_gyn a_10548_3266# vdd pmos_6p0 w=1.2u l=0.5u
X4916 a_24660_40898# cap_shunt_n a_26376_40836# vss nmos_6p0 w=0.82u l=0.6u
X4917 vdd a_3036_38440# a_2948_38484# vdd pmos_6p0 w=1.22u l=1u
X4918 a_34560_7908# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X4919 a_2588_19624# a_2500_19668# vss vss nmos_6p0 w=0.82u l=1u
X4920 a_30632_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X4921 a_8848_37400# cap_shunt_n a_6740_37400# vss nmos_6p0 w=0.82u l=0.6u
X4922 a_6740_26424# cap_shunt_n a_6532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X4923 vss cap_series_gygyp a_36296_12312# vss nmos_6p0 w=0.82u l=0.6u
X4924 vdd a_9532_55688# a_9444_55732# vdd pmos_6p0 w=1.22u l=1u
X4925 a_17828_34264# cap_shunt_n a_17620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X4926 vss tune_shunt[7] a_2708_28354# vss nmos_6p0 w=0.51u l=0.6u
X4927 a_21540_25564# cap_shunt_n a_21748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X4928 a_9108_47516# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4929 a_37632_45944# cap_shunt_gyn a_37444_45944# vdd pmos_6p0 w=1.215u l=0.5u
X4930 vdd a_3036_35304# a_2948_35348# vdd pmos_6p0 w=1.22u l=1u
X4931 a_3828_21720# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X4932 a_17620_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4933 a_6740_23288# cap_shunt_p a_6532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X4934 a_1716_7124# cap_shunt_n a_1924_7608# vdd pmos_6p0 w=1.2u l=0.5u
X4935 a_9428_18946# cap_shunt_p a_9220_19292# vdd pmos_6p0 w=1.2u l=0.5u
X4936 a_17828_31128# cap_shunt_n a_17620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X4937 vss tune_shunt[7] a_2708_25218# vss nmos_6p0 w=0.51u l=0.6u
X4938 a_21540_22428# cap_shunt_p a_21748_22082# vdd pmos_6p0 w=1.2u l=0.5u
X4939 a_15624_10744# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X4940 vdd tune_series_gy[5] a_29492_14588# vdd pmos_6p0 w=1.2u l=0.5u
X4941 vdd a_6508_55688# a_6420_55732# vdd pmos_6p0 w=1.22u l=1u
X4942 vss tune_shunt[5] a_6292_49944# vss nmos_6p0 w=0.51u l=0.6u
X4943 a_37632_42808# cap_shunt_gyn a_37444_42808# vdd pmos_6p0 w=1.215u l=0.5u
X4944 a_6532_33780# cap_shunt_n a_6740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X4945 vdd tune_shunt[7] a_7540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X4946 vss tune_shunt[5] a_2708_48738# vss nmos_6p0 w=0.51u l=0.6u
X4947 a_32604_42711# a_32516_42808# vss vss nmos_6p0 w=0.82u l=1u
X4948 vdd a_32380_41576# a_32292_41620# vdd pmos_6p0 w=1.22u l=1u
X4949 a_35180_38007# a_35092_38104# vss vss nmos_6p0 w=0.82u l=1u
X4950 a_17620_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4951 a_9876_48376# cap_shunt_p a_9668_47892# vdd pmos_6p0 w=1.2u l=0.5u
X4952 a_10340_38484# cap_shunt_n a_10548_38968# vdd pmos_6p0 w=1.2u l=0.5u
X4953 vdd a_22972_49416# a_22884_49460# vdd pmos_6p0 w=1.22u l=1u
X4954 a_3620_46324# cap_shunt_p a_3828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X4955 a_3620_40052# cap_shunt_n a_3828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X4956 a_14484_8692# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4957 vss cap_shunt_p a_19936_21720# vss nmos_6p0 w=0.82u l=0.6u
X4958 a_32156_7080# a_32068_7124# vss vss nmos_6p0 w=0.82u l=1u
X4959 a_6532_30644# cap_shunt_n a_6740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X4960 a_22064_20152# cap_shunt_p a_20740_20152# vss nmos_6p0 w=0.82u l=0.6u
X4961 vss cap_shunt_n a_5152_29560# vss nmos_6p0 w=0.82u l=0.6u
X4962 a_15792_3204# cap_series_gyn a_14468_3266# vss nmos_6p0 w=0.82u l=0.6u
X4963 a_34308_13020# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4964 a_10340_35348# cap_shunt_n a_10548_35832# vdd pmos_6p0 w=1.2u l=0.5u
X4965 vdd tune_series_gy[4] a_29492_17724# vdd pmos_6p0 w=1.2u l=0.5u
X4966 vss cap_shunt_n a_8848_27992# vss nmos_6p0 w=0.82u l=0.6u
X4967 a_14484_5556# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4968 a_2140_48983# a_2052_49080# vss vss nmos_6p0 w=0.82u l=1u
X4969 a_3640_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X4970 a_33524_29076# cap_shunt_p a_33732_29560# vdd pmos_6p0 w=1.2u l=0.5u
X4971 a_3828_24856# cap_shunt_p a_3620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X4972 a_19276_20759# a_19188_20856# vss vss nmos_6p0 w=0.82u l=1u
X4973 vdd a_33052_41143# a_32964_41240# vdd pmos_6p0 w=1.22u l=1u
X4974 vdd tune_shunt[5] a_32404_34972# vdd pmos_6p0 w=1.2u l=0.5u
X4975 a_24204_29032# a_24116_29076# vss vss nmos_6p0 w=0.82u l=1u
X4976 vdd a_15020_54120# a_14932_54164# vdd pmos_6p0 w=1.22u l=1u
X4977 vss cap_shunt_p a_5152_26424# vss nmos_6p0 w=0.82u l=0.6u
X4978 a_23084_47848# a_22996_47892# vss vss nmos_6p0 w=0.82u l=1u
X4979 vdd tune_shunt[7] a_9668_16532# vdd pmos_6p0 w=1.2u l=0.5u
X4980 vss tune_shunt[6] a_17828_45240# vss nmos_6p0 w=0.51u l=0.6u
X4981 vss tune_shunt[7] a_24660_26786# vss nmos_6p0 w=0.51u l=0.6u
X4982 vss cap_shunt_p a_8848_24856# vss nmos_6p0 w=0.82u l=0.6u
X4983 a_3640_31428# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X4984 vss cap_shunt_p a_23856_20452# vss nmos_6p0 w=0.82u l=0.6u
X4985 vdd a_35628_34871# a_35540_34968# vdd pmos_6p0 w=1.22u l=1u
X4986 a_11612_8692# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X4987 a_3828_21720# cap_shunt_p a_3620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X4988 a_28460_3511# a_28372_3608# vss vss nmos_6p0 w=0.82u l=1u
X4989 vdd tune_shunt[4] a_32404_31836# vdd pmos_6p0 w=1.2u l=0.5u
X4990 a_24204_25896# a_24116_25940# vss vss nmos_6p0 w=0.82u l=1u
X4991 a_9540_15810# cap_shunt_p a_10472_15748# vss nmos_6p0 w=0.82u l=0.6u
X4992 a_4492_5512# a_4404_5556# vss vss nmos_6p0 w=0.82u l=1u
X4993 a_19732_12312# cap_series_gyn a_21448_12312# vss nmos_6p0 w=0.82u l=0.6u
X4994 vss cap_shunt_n a_8176_53380# vss nmos_6p0 w=0.82u l=0.6u
X4995 vss tune_shunt[6] a_17828_42104# vss nmos_6p0 w=0.51u l=0.6u
X4996 a_12788_49944# cap_shunt_n a_14504_49944# vss nmos_6p0 w=0.82u l=0.6u
X4997 vdd tune_shunt[4] a_16500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X4998 a_24752_13880# cap_series_gyn a_22644_13880# vss nmos_6p0 w=0.82u l=0.6u
X4999 a_14580_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5000 vdd tune_shunt[6] a_11460_41620# vdd pmos_6p0 w=1.2u l=0.5u
X5001 a_24660_34626# cap_shunt_p a_26376_34564# vss nmos_6p0 w=0.82u l=0.6u
X5002 a_24452_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5003 vdd tune_shunt[6] a_10452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X5004 vss tune_shunt[7] a_21748_31490# vss nmos_6p0 w=0.51u l=0.6u
X5005 vss cap_shunt_p a_31808_4772# vss nmos_6p0 w=0.82u l=0.6u
X5006 a_17620_46324# cap_shunt_n a_17828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X5007 vss cap_series_gyp a_21840_7608# vss nmos_6p0 w=0.82u l=0.6u
X5008 vss tune_shunt[6] a_6740_48376# vss nmos_6p0 w=0.51u l=0.6u
X5009 a_21748_37762# cap_shunt_n a_21540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X5010 a_24752_10744# cap_series_gyp a_22644_10744# vss nmos_6p0 w=0.82u l=0.6u
X5011 a_14580_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5012 a_16632_7908# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X5013 a_21540_19292# cap_shunt_p a_21748_18946# vdd pmos_6p0 w=1.2u l=0.5u
X5014 a_22848_46808# cap_shunt_p a_20740_46808# vss nmos_6p0 w=0.82u l=0.6u
X5015 a_7540_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5016 a_14484_7124# cap_series_gyp a_14692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X5017 vdd a_5612_41143# a_5524_41240# vdd pmos_6p0 w=1.22u l=1u
X5018 a_37632_39672# cap_shunt_gyp a_37444_39672# vdd pmos_6p0 w=1.215u l=0.5u
X5019 a_29700_39330# cap_shunt_p a_30632_39268# vss nmos_6p0 w=0.82u l=0.6u
X5020 a_24660_31490# cap_shunt_p a_26376_31428# vss nmos_6p0 w=0.82u l=0.6u
X5021 vss cap_shunt_p a_27104_27992# vss nmos_6p0 w=0.82u l=0.6u
X5022 a_22436_10260# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5023 a_19052_50551# a_18964_50648# vss vss nmos_6p0 w=0.82u l=1u
X5024 a_17828_45240# cap_shunt_p a_18760_45240# vss nmos_6p0 w=0.82u l=0.6u
X5025 vdd tune_shunt[6] a_25572_36916# vdd pmos_6p0 w=1.2u l=0.5u
X5026 vdd a_3036_29032# a_2948_29076# vdd pmos_6p0 w=1.22u l=1u
X5027 a_6740_20152# cap_shunt_p a_8456_20152# vss nmos_6p0 w=0.82u l=0.6u
X5028 a_21748_42466# cap_shunt_n a_21540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X5029 vdd a_38092_35304# a_38004_35348# vdd pmos_6p0 w=1.22u l=1u
X5030 a_35448_27992# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5031 a_28572_8215# a_28484_8312# vss vss nmos_6p0 w=0.82u l=1u
X5032 a_25592_32996# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5033 a_17828_24856# cap_shunt_n a_17620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X5034 a_21540_16156# cap_series_gyn a_21748_15810# vdd pmos_6p0 w=1.2u l=0.5u
X5035 a_2708_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5036 vss cap_shunt_p a_27104_24856# vss nmos_6p0 w=0.82u l=0.6u
X5037 a_28692_6040# tune_shunt[0] vss vss nmos_6p0 w=0.51u l=0.6u
X5038 a_25572_18100# cap_series_gyn a_25780_18584# vdd pmos_6p0 w=1.2u l=0.5u
X5039 a_17828_42104# cap_shunt_n a_18760_42104# vss nmos_6p0 w=0.82u l=0.6u
X5040 vdd a_34508_39575# a_34420_39672# vdd pmos_6p0 w=1.22u l=1u
X5041 a_17620_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5042 vdd a_6956_6647# a_6868_6744# vdd pmos_6p0 w=1.22u l=1u
X5043 a_18612_6402# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5044 vdd tune_series_gygy[5] a_31436_20860# vdd pmos_6p0 w=1.2u l=0.5u
X5045 a_25572_14964# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5046 vdd a_8412_10216# a_8324_10260# vdd pmos_6p0 w=1.22u l=1u
X5047 a_17828_21720# cap_shunt_p a_17620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X5048 a_22680_9476# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5049 a_6532_24372# cap_shunt_p a_6740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X5050 a_29700_23650# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5051 vdd a_17596_54120# a_17508_54164# vdd pmos_6p0 w=1.22u l=1u
X5052 a_31260_35304# a_31172_35348# vss vss nmos_6p0 w=0.82u l=1u
X5053 a_10340_29076# cap_shunt_n a_10548_29560# vdd pmos_6p0 w=1.2u l=0.5u
X5054 a_35692_24372# cap_series_gygyp a_35880_24372# vdd pmos_6p0 w=1.2u l=0.5u
X5055 a_5844_3266# cap_shunt_n a_5636_3612# vdd pmos_6p0 w=1.2u l=0.5u
X5056 a_25572_11828# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5057 a_9856_29860# cap_shunt_n a_7748_29922# vss nmos_6p0 w=0.82u l=0.6u
X5058 a_29492_17724# cap_series_gyp a_29700_17378# vdd pmos_6p0 w=1.2u l=0.5u
X5059 a_34396_52552# a_34308_52596# vss vss nmos_6p0 w=0.82u l=1u
X5060 vdd a_6956_38007# a_6868_38104# vdd pmos_6p0 w=1.22u l=1u
X5061 a_3640_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5062 vdd a_19164_55688# a_19076_55732# vdd pmos_6p0 w=1.22u l=1u
X5063 vdd a_17596_50984# a_17508_51028# vdd pmos_6p0 w=1.22u l=1u
X5064 a_33920_43734# cap_shunt_gyn a_33920_43189# vdd pmos_6p0 w=1.215u l=0.5u
X5065 vss tune_shunt[7] a_24660_29922# vss nmos_6p0 w=0.51u l=0.6u
X5066 a_19276_14487# a_19188_14584# vss vss nmos_6p0 w=0.82u l=1u
X5067 a_6532_21236# cap_shunt_p a_6740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X5068 a_6532_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5069 a_28484_36916# cap_shunt_p a_28692_37400# vdd pmos_6p0 w=1.2u l=0.5u
X5070 vss cap_shunt_n a_11984_45540# vss nmos_6p0 w=0.82u l=0.6u
X5071 vdd a_2588_25896# a_2500_25940# vdd pmos_6p0 w=1.22u l=1u
X5072 a_15700_4834# cap_series_gyn a_15492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X5073 a_35692_21236# cap_series_gygyp a_35880_21236# vdd pmos_6p0 w=1.2u l=0.5u
X5074 a_9856_26724# cap_shunt_n a_7748_26786# vss nmos_6p0 w=0.82u l=0.6u
X5075 a_34536_9884# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X5076 a_21524_3266# cap_series_gyp a_21316_3612# vdd pmos_6p0 w=1.2u l=0.5u
X5077 vss cap_series_gyn a_23856_14180# vss nmos_6p0 w=0.82u l=0.6u
X5078 a_20740_20152# cap_shunt_p a_20532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X5079 a_2140_39575# a_2052_39672# vss vss nmos_6p0 w=0.82u l=1u
X5080 vdd a_20620_33303# a_20532_33400# vdd pmos_6p0 w=1.22u l=1u
X5081 vdd a_35628_28599# a_35540_28696# vdd pmos_6p0 w=1.22u l=1u
X5082 a_3640_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5083 vdd a_31372_52552# a_31284_52596# vdd pmos_6p0 w=1.22u l=1u
X5084 vdd a_27788_47415# a_27700_47512# vdd pmos_6p0 w=1.22u l=1u
X5085 vdd tune_shunt[4] a_32404_25564# vdd pmos_6p0 w=1.2u l=0.5u
X5086 a_9428_18946# cap_shunt_p a_9220_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5087 vss cap_shunt_n a_11984_42404# vss nmos_6p0 w=0.82u l=0.6u
X5088 a_13588_30268# cap_shunt_n a_13796_29922# vdd pmos_6p0 w=1.2u l=0.5u
X5089 vdd a_2588_22760# a_2500_22804# vdd pmos_6p0 w=1.22u l=1u
X5090 a_6084_16532# cap_shunt_p a_6292_17016# vdd pmos_6p0 w=1.2u l=0.5u
X5091 a_6532_33780# cap_shunt_n a_6740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X5092 a_9668_13396# cap_shunt_p a_9876_13880# vdd pmos_6p0 w=1.2u l=0.5u
X5093 vss cap_shunt_p a_8848_15448# vss nmos_6p0 w=0.82u l=0.6u
X5094 a_10752_20452# cap_shunt_p a_9428_20514# vss nmos_6p0 w=0.82u l=0.6u
X5095 vdd a_30812_53687# a_30724_53784# vdd pmos_6p0 w=1.22u l=1u
X5096 vss tune_shunt[5] a_9876_53080# vss nmos_6p0 w=0.51u l=0.6u
X5097 vdd tune_shunt[7] a_10452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X5098 a_24660_9538# cap_series_gyn a_24452_9884# vdd pmos_6p0 w=1.2u l=0.5u
X5099 vss cap_series_gyn a_23856_11044# vss nmos_6p0 w=0.82u l=0.6u
X5100 a_9668_13396# cap_shunt_p a_9876_13880# vdd pmos_6p0 w=1.2u l=0.5u
X5101 vss tune_series_gy[5] a_24660_17378# vss nmos_6p0 w=0.51u l=0.6u
X5102 a_9876_48376# cap_shunt_p a_9668_47892# vdd pmos_6p0 w=1.2u l=0.5u
X5103 a_13796_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5104 a_29580_55688# a_29492_55732# vss vss nmos_6p0 w=0.82u l=1u
X5105 a_24204_16488# a_24116_16532# vss vss nmos_6p0 w=0.82u l=1u
X5106 a_24660_28354# cap_shunt_n a_26376_28292# vss nmos_6p0 w=0.82u l=0.6u
X5107 vdd tune_shunt[7] a_10452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X5108 a_6532_30644# cap_shunt_n a_6740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X5109 vdd a_30812_50551# a_30724_50648# vdd pmos_6p0 w=1.22u l=1u
X5110 a_12600_46808# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5111 a_24660_6402# cap_series_gyn a_24452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X5112 a_22436_11828# cap_series_gyn a_22644_12312# vdd pmos_6p0 w=1.2u l=0.5u
X5113 a_20740_32696# cap_shunt_n a_22456_32696# vss nmos_6p0 w=0.82u l=0.6u
X5114 a_7540_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5115 a_32632_14588# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5116 a_26556_55688# a_26468_55732# vss vss nmos_6p0 w=0.82u l=1u
X5117 vss cap_shunt_p a_16688_45240# vss nmos_6p0 w=0.82u l=0.6u
X5118 vss cap_shunt_n a_27888_42104# vss nmos_6p0 w=0.82u l=0.6u
X5119 a_24660_25218# cap_shunt_p a_26376_25156# vss nmos_6p0 w=0.82u l=0.6u
X5120 vss tune_shunt[7] a_21748_22082# vss nmos_6p0 w=0.51u l=0.6u
X5121 vdd a_13564_5079# a_13476_5176# vdd pmos_6p0 w=1.22u l=1u
X5122 vdd a_19724_45847# a_19636_45944# vdd pmos_6p0 w=1.22u l=1u
X5123 vdd tune_shunt[7] a_10452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X5124 vdd a_38092_29032# a_38004_29076# vdd pmos_6p0 w=1.22u l=1u
X5125 a_18724_6040# cap_series_gyn a_20440_6040# vss nmos_6p0 w=0.82u l=0.6u
X5126 vss tune_shunt[7] a_6628_12674# vss nmos_6p0 w=0.51u l=0.6u
X5127 vdd tune_shunt[5] a_2500_50652# vdd pmos_6p0 w=1.2u l=0.5u
X5128 a_21748_36194# cap_shunt_n a_21540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X5129 a_6740_35832# cap_shunt_n a_7672_35832# vss nmos_6p0 w=0.82u l=0.6u
X5130 a_28572_38007# a_28484_38104# vss vss nmos_6p0 w=0.82u l=1u
X5131 a_29700_34626# cap_shunt_p a_29492_34972# vdd pmos_6p0 w=1.2u l=0.5u
X5132 a_6308_20860# cap_shunt_p a_6516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X5133 a_27104_43672# cap_shunt_p a_25780_43672# vss nmos_6p0 w=0.82u l=0.6u
X5134 vdd a_33948_41576# a_33860_41620# vdd pmos_6p0 w=1.22u l=1u
X5135 vss cap_series_gygyp a_36624_23588# vss nmos_6p0 w=0.82u l=0.6u
X5136 a_7540_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5137 vss cap_series_gyp a_20720_7908# vss nmos_6p0 w=0.82u l=0.6u
X5138 vdd a_3932_52552# a_3844_52596# vdd pmos_6p0 w=1.22u l=1u
X5139 a_32632_11452# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X5140 vss cap_shunt_n a_16688_42104# vss nmos_6p0 w=0.82u l=0.6u
X5141 vdd tune_shunt[7] a_25572_27508# vdd pmos_6p0 w=1.2u l=0.5u
X5142 vss cap_series_gyn a_27104_18584# vss nmos_6p0 w=0.82u l=0.6u
X5143 vdd a_19724_42711# a_19636_42808# vdd pmos_6p0 w=1.22u l=1u
X5144 vdd a_6060_55255# a_5972_55352# vdd pmos_6p0 w=1.22u l=1u
X5145 a_37084_40008# a_36996_40052# vss vss nmos_6p0 w=0.82u l=1u
X5146 a_21748_33058# cap_shunt_n a_21540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X5147 a_7768_6748# cap_series_gyp a_7580_6748# vdd pmos_6p0 w=1.2u l=0.5u
X5148 a_29700_31490# cap_shunt_p a_29492_31836# vdd pmos_6p0 w=1.2u l=0.5u
X5149 a_15904_43672# cap_shunt_n a_14580_43672# vss nmos_6p0 w=0.82u l=0.6u
X5150 vdd tune_shunt[6] a_3620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X5151 a_27104_40536# cap_shunt_n a_25780_40536# vss nmos_6p0 w=0.82u l=0.6u
X5152 a_25592_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5153 a_31260_29032# a_31172_29076# vss vss nmos_6p0 w=0.82u l=1u
X5154 a_8860_17623# a_8772_17720# vss vss nmos_6p0 w=0.82u l=1u
X5155 vdd a_30364_42711# a_30276_42808# vdd pmos_6p0 w=1.22u l=1u
X5156 vss cap_series_gyp a_27104_15448# vss nmos_6p0 w=0.82u l=0.6u
X5157 vdd tune_shunt[4] a_16500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X5158 a_17620_43188# cap_shunt_p a_17828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X5159 a_22644_9176# cap_series_gyp a_22436_8692# vdd pmos_6p0 w=1.2u l=0.5u
X5160 vdd a_3036_55255# a_2948_55352# vdd pmos_6p0 w=1.22u l=1u
X5161 a_37868_30167# a_37780_30264# vss vss nmos_6p0 w=0.82u l=1u
X5162 vdd tune_shunt[6] a_11460_41620# vdd pmos_6p0 w=1.2u l=0.5u
X5163 a_15904_40536# cap_shunt_n a_14580_40536# vss nmos_6p0 w=0.82u l=0.6u
X5164 a_16708_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5165 a_31436_8316# cap_series_gygyn a_31624_8316# vdd pmos_6p0 w=1.2u l=0.5u
X5166 a_29700_14242# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5167 a_31260_25896# a_31172_25940# vss vss nmos_6p0 w=0.82u l=1u
X5168 a_10340_25940# cap_shunt_n a_10548_26424# vdd pmos_6p0 w=1.2u l=0.5u
X5169 vdd tune_shunt[2] a_1716_5180# vdd pmos_6p0 w=1.2u l=0.5u
X5170 a_1716_8316# cap_shunt_n a_1924_7970# vdd pmos_6p0 w=1.2u l=0.5u
X5171 a_9668_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5172 a_6060_33303# a_5972_33400# vss vss nmos_6p0 w=0.82u l=1u
X5173 a_5936_27992# cap_shunt_n a_3828_27992# vss nmos_6p0 w=0.82u l=0.6u
X5174 vdd tune_series_gy[5] a_19524_7124# vdd pmos_6p0 w=1.2u l=0.5u
X5175 vdd a_3036_52119# a_2948_52216# vdd pmos_6p0 w=1.22u l=1u
X5176 a_9644_43144# a_9556_43188# vss vss nmos_6p0 w=0.82u l=1u
X5177 a_37868_27031# a_37780_27128# vss vss nmos_6p0 w=0.82u l=1u
X5178 a_18044_49416# a_17956_49460# vss vss nmos_6p0 w=0.82u l=1u
X5179 a_29492_38108# cap_shunt_n a_29700_37762# vdd pmos_6p0 w=1.2u l=0.5u
X5180 a_19544_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5181 a_29700_11106# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5182 a_6084_50652# cap_shunt_p a_6292_50306# vdd pmos_6p0 w=1.2u l=0.5u
X5183 a_21748_42466# cap_shunt_n a_21540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X5184 a_29492_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5185 a_29492_5180# tune_shunt[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5186 vdd a_23756_19624# a_23668_19668# vdd pmos_6p0 w=1.22u l=1u
X5187 a_6740_46808# cap_shunt_p a_6532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X5188 a_28484_27508# cap_shunt_p a_28692_27992# vdd pmos_6p0 w=1.2u l=0.5u
X5189 vss cap_shunt_n a_11984_36132# vss nmos_6p0 w=0.82u l=0.6u
X5190 a_5936_24856# cap_shunt_p a_3828_24856# vss nmos_6p0 w=0.82u l=0.6u
X5191 a_10340_22804# cap_shunt_n a_10548_23288# vdd pmos_6p0 w=1.2u l=0.5u
X5192 vss cap_series_gyn a_23856_6340# vss nmos_6p0 w=0.82u l=0.6u
X5193 a_9644_40008# a_9556_40052# vss vss nmos_6p0 w=0.82u l=1u
X5194 vdd a_2588_16488# a_2500_16532# vdd pmos_6p0 w=1.22u l=1u
X5195 vss cap_shunt_p a_30016_35832# vss nmos_6p0 w=0.82u l=0.6u
X5196 a_25572_18100# cap_series_gyn a_25780_18584# vdd pmos_6p0 w=1.2u l=0.5u
X5197 a_34308_23996# cap_series_gygyp a_34516_23650# vdd pmos_6p0 w=1.2u l=0.5u
X5198 a_29492_31836# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5199 a_21448_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5200 vdd a_18044_10216# a_17956_10260# vdd pmos_6p0 w=1.22u l=1u
X5201 a_34144_45540# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5202 a_21748_7970# cap_series_gyp a_21540_8316# vdd pmos_6p0 w=1.2u l=0.5u
X5203 a_13588_28700# cap_shunt_n a_13796_28354# vdd pmos_6p0 w=1.2u l=0.5u
X5204 a_21540_20860# cap_shunt_p a_21748_20514# vdd pmos_6p0 w=1.2u l=0.5u
X5205 vss cap_shunt_n a_4032_50244# vss nmos_6p0 w=0.82u l=0.6u
X5206 vdd tune_shunt[6] a_17620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X5207 vdd a_36188_53687# a_36100_53784# vdd pmos_6p0 w=1.22u l=1u
X5208 a_6532_24372# cap_shunt_p a_6740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X5209 vdd a_30812_44279# a_30724_44376# vdd pmos_6p0 w=1.22u l=1u
X5210 a_8456_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5211 a_13796_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5212 a_34144_42404# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5213 a_33524_35348# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5214 vss cap_shunt_n a_18816_32996# vss nmos_6p0 w=0.82u l=0.6u
X5215 vss cap_series_gyp a_12216_7608# vss nmos_6p0 w=0.82u l=0.6u
X5216 vdd a_1692_9783# a_1604_9880# vdd pmos_6p0 w=1.22u l=1u
X5217 vdd a_19724_39575# a_19636_39672# vdd pmos_6p0 w=1.22u l=1u
X5218 a_2708_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5219 vdd tune_shunt[7] a_10452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X5220 a_5612_47415# a_5524_47512# vss vss nmos_6p0 w=0.82u l=1u
X5221 vdd tune_shunt[6] a_2500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X5222 a_29744_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X5223 a_21540_45948# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5224 a_6740_29560# cap_shunt_n a_7672_29560# vss nmos_6p0 w=0.82u l=0.6u
X5225 a_6532_21236# cap_shunt_p a_6740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X5226 a_2708_37762# cap_shunt_n a_4424_37700# vss nmos_6p0 w=0.82u l=0.6u
X5227 a_20740_23288# cap_shunt_p a_22456_23288# vss nmos_6p0 w=0.82u l=0.6u
X5228 vdd a_29468_6647# a_29380_6744# vdd pmos_6p0 w=1.22u l=1u
X5229 a_1692_30167# a_1604_30264# vss vss nmos_6p0 w=0.82u l=1u
X5230 a_7540_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5231 a_3620_41620# cap_shunt_p a_3828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X5232 vdd tune_shunt[3] a_5636_8692# vdd pmos_6p0 w=1.2u l=0.5u
X5233 a_29624_37400# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5234 vdd a_19724_36439# a_19636_36536# vdd pmos_6p0 w=1.22u l=1u
X5235 a_2708_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5236 a_20740_20152# cap_shunt_p a_20532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X5237 vdd tune_shunt[6] a_2500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X5238 a_24652_35304# a_24564_35348# vss vss nmos_6p0 w=0.82u l=1u
X5239 vss tune_shunt[7] a_29700_29922# vss nmos_6p0 w=0.51u l=0.6u
X5240 a_21748_26786# cap_shunt_n a_21540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X5241 a_6740_26424# cap_shunt_n a_7672_26424# vss nmos_6p0 w=0.82u l=0.6u
X5242 a_29700_25218# cap_shunt_p a_29492_25564# vdd pmos_6p0 w=1.2u l=0.5u
X5243 a_27104_34264# cap_shunt_p a_25780_34264# vss nmos_6p0 w=0.82u l=0.6u
X5244 a_1692_27031# a_1604_27128# vss vss nmos_6p0 w=0.82u l=1u
X5245 a_6084_16532# cap_shunt_p a_6292_17016# vdd pmos_6p0 w=1.2u l=0.5u
X5246 vdd a_34396_55688# a_34308_55732# vdd pmos_6p0 w=1.22u l=1u
X5247 a_6532_33780# cap_shunt_n a_6740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X5248 a_13588_30268# cap_shunt_n a_13796_29922# vdd pmos_6p0 w=1.2u l=0.5u
X5249 a_27788_52552# a_27700_52596# vss vss nmos_6p0 w=0.82u l=1u
X5250 vss cap_shunt_n a_14784_21720# vss nmos_6p0 w=0.82u l=0.6u
X5251 vss tune_shunt[6] a_16708_40898# vss nmos_6p0 w=0.51u l=0.6u
X5252 a_11572_3988# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5253 a_35880_3988# cap_series_gygyp a_35692_3988# vdd pmos_6p0 w=1.2u l=0.5u
X5254 a_27104_31128# cap_shunt_p a_25780_31128# vss nmos_6p0 w=0.82u l=0.6u
X5255 vdd a_27228_23895# a_27140_23992# vdd pmos_6p0 w=1.22u l=1u
X5256 a_3380_49944# cap_shunt_p a_5096_49944# vss nmos_6p0 w=0.82u l=0.6u
X5257 a_6532_30644# cap_shunt_n a_6740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X5258 a_7540_45948# cap_shunt_p a_7748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X5259 a_29492_5180# cap_shunt_p a_29700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X5260 vdd a_24764_52552# a_24676_52596# vdd pmos_6p0 w=1.22u l=1u
X5261 a_10548_35832# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5262 a_28692_32696# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5263 a_14484_10260# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5264 vdd a_27228_20759# a_27140_20856# vdd pmos_6p0 w=1.22u l=1u
X5265 a_19544_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5266 a_31816_21720# cap_series_gygyn a_30616_21236# vss nmos_6p0 w=0.82u l=0.6u
X5267 vdd a_9980_55688# a_9892_55732# vdd pmos_6p0 w=1.22u l=1u
X5268 vdd tune_shunt[5] a_2500_50652# vdd pmos_6p0 w=1.2u l=0.5u
X5269 a_21748_36194# cap_shunt_n a_21540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X5270 a_31260_16488# a_31172_16532# vss vss nmos_6p0 w=0.82u l=1u
X5271 a_29700_34626# cap_shunt_p a_29492_34972# vdd pmos_6p0 w=1.2u l=0.5u
X5272 a_33948_24328# a_33860_24372# vss vss nmos_6p0 w=0.82u l=1u
X5273 a_23968_7608# cap_series_gyp a_22644_7608# vss nmos_6p0 w=0.82u l=0.6u
X5274 a_6308_20860# cap_shunt_p a_6516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X5275 a_12768_43972# cap_shunt_n a_10660_44034# vss nmos_6p0 w=0.82u l=0.6u
X5276 a_28692_27992# cap_shunt_p a_29624_27992# vss nmos_6p0 w=0.82u l=0.6u
X5277 a_6060_23895# a_5972_23992# vss vss nmos_6p0 w=0.82u l=1u
X5278 a_37868_17623# a_37780_17720# vss vss nmos_6p0 w=0.82u l=1u
X5279 a_9644_33736# a_9556_33780# vss vss nmos_6p0 w=0.82u l=1u
X5280 vss cap_shunt_p a_30016_29560# vss nmos_6p0 w=0.82u l=0.6u
X5281 vss cap_shunt_p a_7616_17316# vss nmos_6p0 w=0.82u l=0.6u
X5282 a_9668_52596# cap_shunt_n a_9876_53080# vdd pmos_6p0 w=1.2u l=0.5u
X5283 a_19544_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5284 a_29492_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5285 a_25100_53687# a_25012_53784# vss vss nmos_6p0 w=0.82u l=1u
X5286 a_21748_33058# cap_shunt_n a_21540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X5287 vss cap_series_gygyp a_34952_6340# vss nmos_6p0 w=0.82u l=0.6u
X5288 vdd a_6956_55688# a_6868_55732# vdd pmos_6p0 w=1.22u l=1u
X5289 a_29700_31490# cap_shunt_p a_29492_31836# vdd pmos_6p0 w=1.2u l=0.5u
X5290 a_28484_7124# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5291 a_13796_12674# cap_shunt_p a_14728_12612# vss nmos_6p0 w=0.82u l=0.6u
X5292 a_5936_15448# cap_shunt_p a_3828_15448# vss nmos_6p0 w=0.82u l=0.6u
X5293 a_24452_44380# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5294 a_28692_24856# cap_shunt_p a_29624_24856# vss nmos_6p0 w=0.82u l=0.6u
X5295 a_5844_10744# cap_shunt_p a_5636_10260# vdd pmos_6p0 w=1.2u l=0.5u
X5296 a_12768_40836# cap_shunt_n a_10660_40898# vss nmos_6p0 w=0.82u l=0.6u
X5297 a_9644_30600# a_9556_30644# vss vss nmos_6p0 w=0.82u l=1u
X5298 vss cap_shunt_p a_30016_26424# vss nmos_6p0 w=0.82u l=0.6u
X5299 a_18404_8316# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5300 a_20532_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5301 a_13796_48738# cap_shunt_n a_13588_49084# vdd pmos_6p0 w=1.2u l=0.5u
X5302 a_25100_50551# a_25012_50648# vss vss nmos_6p0 w=0.82u l=1u
X5303 a_31708_36872# a_31620_36916# vss vss nmos_6p0 w=0.82u l=1u
X5304 a_33524_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5305 a_24660_9538# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5306 a_6508_44279# a_6420_44376# vss vss nmos_6p0 w=0.82u l=1u
X5307 a_21540_11452# cap_series_gyn a_21748_11106# vdd pmos_6p0 w=1.2u l=0.5u
X5308 vdd tune_shunt[7] a_9332_16156# vdd pmos_6p0 w=1.2u l=0.5u
X5309 a_2708_18946# cap_shunt_p a_3640_18884# vss nmos_6p0 w=0.82u l=0.6u
X5310 a_24452_41244# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5311 vdd a_17596_7080# a_17508_7124# vdd pmos_6p0 w=1.22u l=1u
X5312 a_21540_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5313 a_15568_27992# cap_shunt_n a_13460_27992# vss nmos_6p0 w=0.82u l=0.6u
X5314 a_20328_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5315 a_4648_9176# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5316 vdd a_34844_54120# a_34756_54164# vdd pmos_6p0 w=1.22u l=1u
X5317 a_29384_3612# cap_series_gyn a_29196_3612# vdd pmos_6p0 w=1.2u l=0.5u
X5318 vss tune_shunt[7] a_20740_20152# vss nmos_6p0 w=0.51u l=0.6u
X5319 a_7068_54120# a_6980_54164# vss vss nmos_6p0 w=0.82u l=1u
X5320 a_20740_38968# cap_shunt_n a_21672_38968# vss nmos_6p0 w=0.82u l=0.6u
X5321 vss cap_shunt_n a_18816_23588# vss nmos_6p0 w=0.82u l=0.6u
X5322 a_6508_41143# a_6420_41240# vss vss nmos_6p0 w=0.82u l=1u
X5323 a_2708_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5324 a_2708_15810# cap_shunt_p a_3640_15748# vss nmos_6p0 w=0.82u l=0.6u
X5325 a_29492_38108# cap_shunt_n a_29700_37762# vdd pmos_6p0 w=1.2u l=0.5u
X5326 a_24652_29032# a_24564_29076# vss vss nmos_6p0 w=0.82u l=1u
X5327 a_2500_23996# cap_shunt_p a_2708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X5328 a_6084_50652# cap_shunt_p a_6292_50306# vdd pmos_6p0 w=1.2u l=0.5u
X5329 a_36384_45540# cap_shunt_gyp a_36384_45944# vdd pmos_6p0 w=1.215u l=0.5u
X5330 a_15568_24856# cap_shunt_n a_13460_24856# vss nmos_6p0 w=0.82u l=0.6u
X5331 a_14468_3266# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X5332 vss cap_series_gyn a_8968_7908# vss nmos_6p0 w=0.82u l=0.6u
X5333 vss cap_series_gyp a_11096_7908# vss nmos_6p0 w=0.82u l=0.6u
X5334 vdd a_34844_50984# a_34756_51028# vdd pmos_6p0 w=1.22u l=1u
X5335 a_33920_44757# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X5336 vdd a_4940_6647# a_4852_6744# vdd pmos_6p0 w=1.22u l=1u
X5337 a_18180_3612# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5338 a_36524_14487# a_36436_14584# vss vss nmos_6p0 w=0.82u l=1u
X5339 a_21748_45602# cap_shunt_p a_22680_45540# vss nmos_6p0 w=0.82u l=0.6u
X5340 vdd a_34396_49416# a_34308_49460# vdd pmos_6p0 w=1.22u l=1u
X5341 a_28692_38968# cap_shunt_n a_28484_38484# vdd pmos_6p0 w=1.2u l=0.5u
X5342 a_3620_32212# cap_shunt_p a_3828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X5343 a_2708_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5344 vdd a_19724_27031# a_19636_27128# vdd pmos_6p0 w=1.22u l=1u
X5345 a_24652_25896# a_24564_25940# vss vss nmos_6p0 w=0.82u l=1u
X5346 a_34308_23996# cap_series_gygyp a_34516_23650# vdd pmos_6p0 w=1.2u l=0.5u
X5347 a_22524_54120# a_22436_54164# vss vss nmos_6p0 w=0.82u l=1u
X5348 a_17620_46324# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5349 a_36384_42404# cap_shunt_gyn a_36384_42808# vdd pmos_6p0 w=1.215u l=0.5u
X5350 a_29700_4834# tune_shunt[0] vss vss nmos_6p0 w=0.51u l=0.6u
X5351 vdd tune_shunt[6] a_9108_49084# vdd pmos_6p0 w=1.2u l=0.5u
X5352 vdd a_25212_55688# a_25124_55732# vdd pmos_6p0 w=1.22u l=1u
X5353 a_26444_47415# a_26356_47512# vss vss nmos_6p0 w=0.82u l=1u
X5354 a_24452_5180# cap_series_gyp a_24660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X5355 vdd a_4940_3511# a_4852_3608# vdd pmos_6p0 w=1.22u l=1u
X5356 a_27496_4472# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5357 a_36524_11351# a_36436_11448# vss vss nmos_6p0 w=0.82u l=1u
X5358 a_32040_18884# cap_series_gygyn a_31624_19292# vss nmos_6p0 w=0.82u l=0.6u
X5359 a_21748_42466# cap_shunt_n a_22680_42404# vss nmos_6p0 w=0.82u l=0.6u
X5360 vdd a_15356_14920# a_15268_14964# vdd pmos_6p0 w=1.22u l=1u
X5361 a_1692_17623# a_1604_17720# vss vss nmos_6p0 w=0.82u l=1u
X5362 a_8400_51512# cap_shunt_p a_6292_51512# vss nmos_6p0 w=0.82u l=0.6u
X5363 a_7540_39676# cap_shunt_n a_7748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X5364 a_28692_35832# cap_shunt_p a_28484_35348# vdd pmos_6p0 w=1.2u l=0.5u
X5365 a_6532_24372# cap_shunt_p a_6740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X5366 a_10548_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5367 vdd a_12444_50984# a_12356_51028# vdd pmos_6p0 w=1.22u l=1u
X5368 a_8680_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5369 a_16708_45602# cap_shunt_p a_16500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X5370 a_22076_49416# a_21988_49460# vss vss nmos_6p0 w=0.82u l=1u
X5371 vdd a_15356_11784# a_15268_11828# vdd pmos_6p0 w=1.22u l=1u
X5372 a_32156_13352# a_32068_13396# vss vss nmos_6p0 w=0.82u l=1u
X5373 vdd a_27228_14487# a_27140_14584# vdd pmos_6p0 w=1.22u l=1u
X5374 vdd tune_shunt[6] a_2500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X5375 a_10660_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5376 a_6740_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5377 a_6532_21236# cap_shunt_p a_6740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X5378 vss tune_series_gy[1] a_10548_3266# vss nmos_6p0 w=0.51u l=0.6u
X5379 a_33948_18056# a_33860_18100# vss vss nmos_6p0 w=0.82u l=1u
X5380 a_35448_20452# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X5381 vss cap_shunt_gyn a_36428_43672# vss nmos_6p0 w=0.82u l=0.6u
X5382 a_10548_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5383 a_3620_19668# cap_shunt_p a_3828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X5384 a_28484_7124# cap_series_gyp a_28692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X5385 a_7580_5180# cap_series_gyn a_7768_5180# vdd pmos_6p0 w=1.2u l=0.5u
X5386 a_7748_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5387 a_28692_23288# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5388 a_8860_49416# a_8772_49460# vss vss nmos_6p0 w=0.82u l=1u
X5389 vss cap_shunt_p a_7728_22020# vss nmos_6p0 w=0.82u l=0.6u
X5390 a_32156_10216# a_32068_10260# vss vss nmos_6p0 w=0.82u l=1u
X5391 vdd a_27228_11351# a_27140_11448# vdd pmos_6p0 w=1.22u l=1u
X5392 vdd tune_shunt[6] a_2500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X5393 a_21748_26786# cap_shunt_n a_21540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X5394 vss tune_series_gygy[5] a_35880_21236# vss nmos_6p0 w=0.51u l=0.6u
X5395 a_17828_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5396 a_9876_13880# cap_shunt_p a_10808_13880# vss nmos_6p0 w=0.82u l=0.6u
X5397 a_37444_47512# cap_shunt_gyp a_37632_47512# vdd pmos_6p0 w=1.215u l=0.5u
X5398 a_29700_25218# cap_shunt_p a_29492_25564# vdd pmos_6p0 w=1.2u l=0.5u
X5399 a_22568_6040# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5400 a_33948_14920# a_33860_14964# vss vss nmos_6p0 w=0.82u l=1u
X5401 vdd tune_shunt[7] a_21540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X5402 a_28692_18584# cap_series_gyp a_29624_18584# vss nmos_6p0 w=0.82u l=0.6u
X5403 vdd a_34956_39575# a_34868_39672# vdd pmos_6p0 w=1.22u l=1u
X5404 a_34396_38440# a_34308_38484# vss vss nmos_6p0 w=0.82u l=1u
X5405 a_12768_34564# cap_shunt_n a_10660_34626# vss nmos_6p0 w=0.82u l=0.6u
X5406 a_7748_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5407 a_35264_47108# cap_shunt_gyn a_35264_47512# vdd pmos_6p0 w=1.215u l=0.5u
X5408 a_21748_7970# cap_series_gyp a_22680_7908# vss nmos_6p0 w=0.82u l=0.6u
X5409 vdd a_8860_10216# a_8772_10260# vdd pmos_6p0 w=1.22u l=1u
X5410 a_19544_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5411 a_18516_5556# cap_series_gyn a_18724_6040# vdd pmos_6p0 w=1.2u l=0.5u
X5412 a_16920_11044# cap_series_gyp a_15720_11452# vss nmos_6p0 w=0.82u l=0.6u
X5413 a_17828_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5414 a_9876_10744# cap_shunt_p a_10808_10744# vss nmos_6p0 w=0.82u l=0.6u
X5415 a_28692_15448# cap_series_gyn a_29624_15448# vss nmos_6p0 w=0.82u l=0.6u
X5416 vdd a_23308_44712# a_23220_44756# vdd pmos_6p0 w=1.22u l=1u
X5417 a_12768_31428# cap_shunt_n a_10660_31490# vss nmos_6p0 w=0.82u l=0.6u
X5418 a_9668_49460# cap_shunt_p a_9876_49944# vdd pmos_6p0 w=1.2u l=0.5u
X5419 a_35904_23288# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X5420 vss cap_series_gyn a_30016_17016# vss nmos_6p0 w=0.82u l=0.6u
X5421 a_18044_52119# a_17956_52216# vss vss nmos_6p0 w=0.82u l=1u
X5422 vss cap_shunt_n a_15120_48676# vss nmos_6p0 w=0.82u l=0.6u
X5423 a_6740_48376# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5424 a_29916_20759# a_29828_20856# vss vss nmos_6p0 w=0.82u l=1u
X5425 vdd tune_shunt[6] a_20532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X5426 a_6508_34871# a_6420_34968# vss vss nmos_6p0 w=0.82u l=1u
X5427 vss tune_shunt[2] a_1924_7970# vss nmos_6p0 w=0.51u l=0.6u
X5428 vdd a_15804_13352# a_15716_13396# vdd pmos_6p0 w=1.22u l=1u
X5429 vss tune_shunt[6] a_3828_45240# vss nmos_6p0 w=0.51u l=0.6u
X5430 a_10452_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5431 a_7748_23650# cap_shunt_p a_7540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X5432 vss tune_series_gy[1] a_6760_3988# vss nmos_6p0 w=0.51u l=0.6u
X5433 a_30016_4472# cap_series_gyp a_28692_4472# vss nmos_6p0 w=0.82u l=0.6u
X5434 a_22456_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5435 a_32404_36540# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5436 a_6508_31735# a_6420_31832# vss vss nmos_6p0 w=0.82u l=1u
X5437 a_2500_14588# cap_shunt_n a_2708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X5438 vdd a_16588_55688# a_16500_55732# vdd pmos_6p0 w=1.22u l=1u
X5439 vss cap_shunt_p a_25984_22020# vss nmos_6p0 w=0.82u l=0.6u
X5440 a_11460_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5441 a_31260_5512# a_31172_5556# vss vss nmos_6p0 w=0.82u l=1u
X5442 vss tune_shunt[2] a_1924_4834# vss nmos_6p0 w=0.51u l=0.6u
X5443 a_6644_53788# cap_shunt_n a_6852_53442# vdd pmos_6p0 w=1.2u l=0.5u
X5444 vss cap_shunt_gyp a_35308_45240# vss nmos_6p0 w=0.82u l=0.6u
X5445 vss tune_shunt[6] a_3828_42104# vss nmos_6p0 w=0.51u l=0.6u
X5446 a_10452_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5447 a_21540_44380# cap_shunt_n a_21748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X5448 a_21748_36194# cap_shunt_n a_22680_36132# vss nmos_6p0 w=0.82u l=0.6u
X5449 a_34516_20514# cap_series_gygyp a_36232_20452# vss nmos_6p0 w=0.82u l=0.6u
X5450 a_13588_20860# cap_shunt_n a_13796_20514# vdd pmos_6p0 w=1.2u l=0.5u
X5451 a_5844_10744# cap_shunt_p a_5636_10260# vdd pmos_6p0 w=1.2u l=0.5u
X5452 a_32404_33404# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5453 a_28692_29560# cap_shunt_p a_28484_29076# vdd pmos_6p0 w=1.2u l=0.5u
X5454 a_13796_48738# cap_shunt_n a_13588_49084# vdd pmos_6p0 w=1.2u l=0.5u
X5455 vss cap_shunt_n a_12656_34264# vss nmos_6p0 w=0.82u l=0.6u
X5456 a_21056_12312# cap_series_gyn a_19732_12312# vss nmos_6p0 w=0.82u l=0.6u
X5457 a_24652_16488# a_24564_16532# vss vss nmos_6p0 w=0.82u l=1u
X5458 a_2708_45602# cap_shunt_p a_2500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X5459 a_6740_42104# cap_shunt_n a_6532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X5460 a_16708_39330# cap_shunt_n a_16500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X5461 vdd a_9644_36872# a_9556_36916# vdd pmos_6p0 w=1.22u l=1u
X5462 a_21540_41244# cap_shunt_p a_21748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X5463 a_22412_55255# a_22324_55352# vss vss nmos_6p0 w=0.82u l=1u
X5464 a_2500_17724# cap_shunt_p a_2708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X5465 a_16408_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5466 a_26376_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5467 vdd tune_series_gy[5] a_24452_13020# vdd pmos_6p0 w=1.2u l=0.5u
X5468 a_33524_33780# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5469 vss cap_shunt_n a_12656_31128# vss nmos_6p0 w=0.82u l=0.6u
X5470 a_29492_38108# cap_shunt_n a_29700_37762# vdd pmos_6p0 w=1.2u l=0.5u
X5471 a_2500_23996# cap_shunt_p a_2708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X5472 a_12788_20152# cap_shunt_p a_12580_19668# vdd pmos_6p0 w=1.2u l=0.5u
X5473 a_16924_36872# a_16836_36916# vss vss nmos_6p0 w=0.82u l=1u
X5474 a_11872_32696# cap_shunt_n a_10548_32696# vss nmos_6p0 w=0.82u l=0.6u
X5475 a_6740_12312# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5476 vss tune_series_gy[4] a_25780_20152# vss nmos_6p0 w=0.51u l=0.6u
X5477 vss tune_shunt_gy[1] a_37632_40053# vss nmos_6p0 w=0.51u l=0.6u
X5478 a_33524_30644# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5479 a_12768_28292# cap_shunt_n a_10660_28354# vss nmos_6p0 w=0.82u l=0.6u
X5480 a_2708_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5481 vss tune_shunt[7] a_9876_17016# vss nmos_6p0 w=0.51u l=0.6u
X5482 a_7748_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5483 a_28692_38968# cap_shunt_n a_28484_38484# vdd pmos_6p0 w=1.2u l=0.5u
X5484 a_35692_25940# cap_series_gygyp a_35880_25940# vdd pmos_6p0 w=1.2u l=0.5u
X5485 a_6572_7124# cap_series_gyp a_6760_7124# vdd pmos_6p0 w=1.2u l=0.5u
X5486 vss tune_series_gygy[4] a_35880_11828# vss nmos_6p0 w=0.51u l=0.6u
X5487 a_12768_25156# cap_shunt_n a_10660_25218# vss nmos_6p0 w=0.82u l=0.6u
X5488 vdd tune_series_gy[5] a_21540_14588# vdd pmos_6p0 w=1.2u l=0.5u
X5489 a_18940_54120# a_18852_54164# vss vss nmos_6p0 w=0.82u l=1u
X5490 vdd a_23308_38440# a_23220_38484# vdd pmos_6p0 w=1.22u l=1u
X5491 a_7748_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5492 a_5544_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5493 a_28692_35832# cap_shunt_p a_28484_35348# vdd pmos_6p0 w=1.2u l=0.5u
X5494 a_35692_22804# cap_series_gygyp a_35880_22804# vdd pmos_6p0 w=1.2u l=0.5u
X5495 vdd a_3484_55255# a_3396_55352# vdd pmos_6p0 w=1.22u l=1u
X5496 vss tune_shunt[3] a_5844_9538# vss nmos_6p0 w=0.51u l=0.6u
X5497 vss cap_shunt_gyn a_33292_43972# vss nmos_6p0 w=0.82u l=0.6u
X5498 vss tune_shunt[7] a_13460_38968# vss nmos_6p0 w=0.51u l=0.6u
X5499 a_37868_49416# a_37780_49460# vss vss nmos_6p0 w=0.82u l=1u
X5500 a_16708_45602# cap_shunt_p a_16500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X5501 a_6508_28599# a_6420_28696# vss vss nmos_6p0 w=0.82u l=1u
X5502 vss tune_shunt[5] a_2708_50306# vss nmos_6p0 w=0.51u l=0.6u
X5503 vss cap_shunt_p a_7616_49944# vss nmos_6p0 w=0.82u l=0.6u
X5504 vdd a_27788_49416# a_27700_49460# vdd pmos_6p0 w=1.22u l=1u
X5505 vdd a_23308_35304# a_23220_35348# vdd pmos_6p0 w=1.22u l=1u
X5506 a_15916_54120# a_15828_54164# vss vss nmos_6p0 w=0.82u l=1u
X5507 vdd a_3484_52119# a_3396_52216# vdd pmos_6p0 w=1.22u l=1u
X5508 vss cap_shunt_n a_31808_36132# vss nmos_6p0 w=0.82u l=0.6u
X5509 vss cap_shunt_n a_15120_39268# vss nmos_6p0 w=0.82u l=0.6u
X5510 a_28692_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5511 a_18492_49416# a_18404_49460# vss vss nmos_6p0 w=0.82u l=1u
X5512 vdd tune_shunt[7] a_20532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X5513 a_37868_46280# a_37780_46324# vss vss nmos_6p0 w=0.82u l=1u
X5514 a_6508_25463# a_6420_25560# vss vss nmos_6p0 w=0.82u l=1u
X5515 vdd a_27788_46280# a_27700_46324# vdd pmos_6p0 w=1.22u l=1u
X5516 a_18816_37700# cap_shunt_n a_16708_37762# vss nmos_6p0 w=0.82u l=0.6u
X5517 a_6628_12674# cap_shunt_p a_8344_12612# vss nmos_6p0 w=0.82u l=0.6u
X5518 a_16500_23996# cap_shunt_n a_16708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X5519 a_10540_5512# a_10452_5556# vss vss nmos_6p0 w=0.82u l=1u
X5520 a_33544_37700# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5521 a_28692_10744# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5522 a_24660_17378# cap_series_gyp a_24452_17724# vdd pmos_6p0 w=1.2u l=0.5u
X5523 vdd a_18492_10216# a_18404_10260# vdd pmos_6p0 w=1.22u l=1u
X5524 vss cap_shunt_p a_22064_20152# vss nmos_6p0 w=0.82u l=0.6u
X5525 a_32404_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5526 vdd tune_shunt[7] a_25572_25940# vdd pmos_6p0 w=1.2u l=0.5u
X5527 a_12580_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5528 a_2708_39330# cap_shunt_n a_2500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X5529 a_20740_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5530 vss tune_shunt_gy[2] a_36512_41621# vss nmos_6p0 w=0.51u l=0.6u
X5531 a_22412_48983# a_22324_49080# vss vss nmos_6p0 w=0.82u l=1u
X5532 a_31624_22428# cap_series_gygyn a_31436_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5533 a_35840_27992# cap_shunt_p a_33732_27992# vss nmos_6p0 w=0.82u l=0.6u
X5534 a_3620_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5535 vdd tune_shunt[7] a_25572_22804# vdd pmos_6p0 w=1.2u l=0.5u
X5536 a_25572_8692# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5537 a_18940_8648# a_18852_8692# vss vss nmos_6p0 w=0.82u l=1u
X5538 a_34536_9884# cap_series_gygyn a_34348_9884# vdd pmos_6p0 w=1.2u l=0.5u
X5539 a_15492_9884# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5540 a_20740_24856# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5541 a_6740_32696# cap_shunt_n a_6532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X5542 vdd a_9644_27464# a_9556_27508# vdd pmos_6p0 w=1.22u l=1u
X5543 a_17820_55688# a_17732_55732# vss vss nmos_6p0 w=0.82u l=1u
X5544 a_32716_17623# a_32628_17720# vss vss nmos_6p0 w=0.82u l=1u
X5545 a_25572_5556# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5546 vss cap_shunt_gyp a_32172_45540# vss nmos_6p0 w=0.82u l=0.6u
X5547 a_15492_6748# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5548 a_34536_6748# cap_series_gygyp a_34348_6748# vdd pmos_6p0 w=1.2u l=0.5u
X5549 a_23464_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5550 a_1692_49416# a_1604_49460# vss vss nmos_6p0 w=0.82u l=1u
X5551 a_2500_14588# cap_shunt_n a_2708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X5552 a_16700_19624# a_16612_19668# vss vss nmos_6p0 w=0.82u l=1u
X5553 a_11872_23288# cap_shunt_n a_10548_23288# vss nmos_6p0 w=0.82u l=0.6u
X5554 vdd tune_series_gygy[0] a_35692_3988# vdd pmos_6p0 w=1.2u l=0.5u
X5555 a_11572_3988# cap_series_gyp a_11780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X5556 vss tune_shunt[5] a_2708_47170# vss nmos_6p0 w=0.51u l=0.6u
X5557 a_21540_44380# cap_shunt_n a_21748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X5558 a_23464_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5559 a_35692_10260# cap_series_gygyp a_35880_10260# vdd pmos_6p0 w=1.2u l=0.5u
X5560 a_10660_33058# cap_shunt_n a_11592_32996# vss nmos_6p0 w=0.82u l=0.6u
X5561 a_5844_10744# cap_shunt_p a_5636_10260# vdd pmos_6p0 w=1.2u l=0.5u
X5562 a_35692_16532# cap_series_gygyn a_35880_16532# vdd pmos_6p0 w=1.2u l=0.5u
X5563 a_1692_46280# a_1604_46324# vss vss nmos_6p0 w=0.82u l=1u
X5564 a_28692_29560# cap_shunt_p a_28484_29076# vdd pmos_6p0 w=1.2u l=0.5u
X5565 vdd a_1692_10216# a_1604_10260# vdd pmos_6p0 w=1.22u l=1u
X5566 a_12788_15448# cap_shunt_p a_12580_14964# vdd pmos_6p0 w=1.2u l=0.5u
X5567 a_17620_18100# cap_shunt_p a_17828_18584# vdd pmos_6p0 w=1.2u l=0.5u
X5568 vdd a_3036_54120# a_2948_54164# vdd pmos_6p0 w=1.22u l=1u
X5569 vdd a_27676_23895# a_27588_23992# vdd pmos_6p0 w=1.22u l=1u
X5570 vdd a_33164_16055# a_33076_16152# vdd pmos_6p0 w=1.22u l=1u
X5571 a_6308_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5572 a_6740_42104# cap_shunt_n a_6532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X5573 a_16708_39330# cap_shunt_n a_16500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X5574 vss tune_series_gygy[5] a_35880_25940# vss nmos_6p0 w=0.51u l=0.6u
X5575 a_9876_21720# cap_shunt_p a_9668_21236# vdd pmos_6p0 w=1.2u l=0.5u
X5576 a_9876_51512# cap_shunt_n a_9668_51028# vdd pmos_6p0 w=1.2u l=0.5u
X5577 vss tune_shunt[6] a_2708_44034# vss nmos_6p0 w=0.51u l=0.6u
X5578 a_21540_41244# cap_shunt_p a_21748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X5579 vdd a_23308_29032# a_23220_29076# vdd pmos_6p0 w=1.22u l=1u
X5580 a_33024_44376# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X5581 a_10548_35832# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5582 vdd a_32604_14920# a_32516_14964# vdd pmos_6p0 w=1.22u l=1u
X5583 a_12788_12312# cap_shunt_p a_12580_11828# vdd pmos_6p0 w=1.2u l=0.5u
X5584 a_17620_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5585 vdd a_37196_32168# a_37108_32212# vdd pmos_6p0 w=1.22u l=1u
X5586 a_29700_11106# cap_series_gyp a_29492_11452# vdd pmos_6p0 w=1.2u l=0.5u
X5587 vdd a_33164_12919# a_33076_13016# vdd pmos_6p0 w=1.22u l=1u
X5588 a_24660_12674# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5589 vdd a_27676_20759# a_27588_20856# vdd pmos_6p0 w=1.22u l=1u
X5590 a_37644_32168# a_37556_32212# vss vss nmos_6p0 w=0.82u l=1u
X5591 a_16252_11784# a_16164_11828# vss vss nmos_6p0 w=0.82u l=1u
X5592 a_3828_46808# cap_shunt_p a_5544_46808# vss nmos_6p0 w=0.82u l=0.6u
X5593 vdd tune_shunt[7] a_29492_30268# vdd pmos_6p0 w=1.2u l=0.5u
X5594 a_34396_41143# a_34308_41240# vss vss nmos_6p0 w=0.82u l=1u
X5595 a_36296_7608# cap_series_gygyp a_35880_7124# vss nmos_6p0 w=0.82u l=0.6u
X5596 vdd a_32604_11784# a_32516_11828# vdd pmos_6p0 w=1.22u l=1u
X5597 a_6532_47892# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5598 a_20720_6340# cap_series_gyn a_18612_6402# vss nmos_6p0 w=0.82u l=0.6u
X5599 vdd tune_shunt[5] a_29492_36540# vdd pmos_6p0 w=1.2u l=0.5u
X5600 a_31624_19292# cap_series_gygyn a_31436_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5601 a_19936_48376# cap_shunt_p a_17828_48376# vss nmos_6p0 w=0.82u l=0.6u
X5602 a_16708_20514# cap_shunt_p a_18424_20452# vss nmos_6p0 w=0.82u l=0.6u
X5603 a_15804_55255# a_15716_55352# vss vss nmos_6p0 w=0.82u l=1u
X5604 vss tune_series_gygy[0] a_31624_6748# vss nmos_6p0 w=0.51u l=0.6u
X5605 a_26768_20452# cap_shunt_p a_24660_20514# vss nmos_6p0 w=0.82u l=0.6u
X5606 a_37196_27464# a_37108_27508# vss vss nmos_6p0 w=0.82u l=1u
X5607 a_2500_9884# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5608 a_16500_14588# cap_shunt_p a_16708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X5609 vdd a_36188_52552# a_36100_52596# vdd pmos_6p0 w=1.22u l=1u
X5610 vss cap_shunt_p a_5152_45240# vss nmos_6p0 w=0.82u l=0.6u
X5611 a_6532_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5612 a_15176_21720# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5613 a_29384_3612# cap_series_gyn a_29196_3612# vdd pmos_6p0 w=1.2u l=0.5u
X5614 vdd tune_shunt[7] a_17620_18100# vdd pmos_6p0 w=1.2u l=0.5u
X5615 a_33612_39575# a_33524_39672# vss vss nmos_6p0 w=0.82u l=1u
X5616 vdd tune_shunt[5] a_29492_33404# vdd pmos_6p0 w=1.2u l=0.5u
X5617 a_10340_3612# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5618 vss cap_shunt_p a_8848_43672# vss nmos_6p0 w=0.82u l=0.6u
X5619 vdd tune_series_gy[5] a_25572_16532# vdd pmos_6p0 w=1.2u l=0.5u
X5620 a_20740_45240# cap_shunt_n a_20532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X5621 vdd a_1692_8648# a_1604_8692# vdd pmos_6p0 w=1.22u l=1u
X5622 a_3640_50244# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5623 a_6956_44279# a_6868_44376# vss vss nmos_6p0 w=0.82u l=1u
X5624 a_27496_13880# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X5625 a_3828_40536# cap_shunt_n a_3620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X5626 a_20740_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5627 a_11200_48376# cap_shunt_p a_9876_48376# vss nmos_6p0 w=0.82u l=0.6u
X5628 a_24204_44712# a_24116_44756# vss vss nmos_6p0 w=0.82u l=1u
X5629 vss cap_shunt_p a_5152_42104# vss nmos_6p0 w=0.82u l=0.6u
X5630 a_16708_48738# cap_shunt_p a_17640_48676# vss nmos_6p0 w=0.82u l=0.6u
X5631 vss cap_shunt_n a_8848_40536# vss nmos_6p0 w=0.82u l=0.6u
X5632 a_3620_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5633 a_17808_7908# cap_series_gyn a_15700_7970# vss nmos_6p0 w=0.82u l=0.6u
X5634 vdd a_16252_53687# a_16164_53784# vdd pmos_6p0 w=1.22u l=1u
X5635 vss tune_shunt[4] a_24660_42466# vss nmos_6p0 w=0.51u l=0.6u
X5636 a_6956_41143# a_6868_41240# vss vss nmos_6p0 w=0.82u l=1u
X5637 a_2708_34626# cap_shunt_n a_2500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X5638 a_27496_10744# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X5639 a_20740_15448# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5640 a_11460_43188# cap_shunt_n a_11668_43672# vdd pmos_6p0 w=1.2u l=0.5u
X5641 a_24204_41576# a_24116_41620# vss vss nmos_6p0 w=0.82u l=1u
X5642 a_4032_37700# cap_shunt_n a_2708_37762# vss nmos_6p0 w=0.82u l=0.6u
X5643 a_2708_31490# cap_shunt_p a_2500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X5644 a_24660_17378# cap_series_gyp a_24452_17724# vdd pmos_6p0 w=1.2u l=0.5u
X5645 a_22972_54120# a_22884_54164# vss vss nmos_6p0 w=0.82u l=1u
X5646 a_1924_4834# cap_shunt_p a_3640_4772# vss nmos_6p0 w=0.82u l=0.6u
X5647 vss cap_series_gygyn a_37080_13880# vss nmos_6p0 w=0.82u l=0.6u
X5648 vdd a_25660_55688# a_25572_55732# vdd pmos_6p0 w=1.22u l=1u
X5649 a_26892_47415# a_26804_47512# vss vss nmos_6p0 w=0.82u l=1u
X5650 vss tune_shunt[7] a_16708_15810# vss nmos_6p0 w=0.51u l=0.6u
X5651 a_6292_18584# cap_shunt_p a_6084_18100# vdd pmos_6p0 w=1.2u l=0.5u
X5652 vss cap_shunt_p a_4816_47108# vss nmos_6p0 w=0.82u l=0.6u
X5653 a_23464_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5654 a_10660_23650# cap_shunt_n a_11592_23588# vss nmos_6p0 w=0.82u l=0.6u
X5655 a_10548_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5656 a_31624_22428# cap_series_gygyn a_31436_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5657 vss cap_series_gygyp a_37080_10744# vss nmos_6p0 w=0.82u l=0.6u
X5658 vdd a_12892_50984# a_12804_51028# vdd pmos_6p0 w=1.22u l=1u
X5659 vss cap_shunt_p a_27104_43672# vss nmos_6p0 w=0.82u l=0.6u
X5660 a_15532_11452# cap_series_gyp a_15720_11452# vdd pmos_6p0 w=1.2u l=0.5u
X5661 vdd a_27676_14487# a_27588_14584# vdd pmos_6p0 w=1.22u l=1u
X5662 vdd a_22636_55688# a_22548_55732# vdd pmos_6p0 w=1.22u l=1u
X5663 vss cap_shunt_p a_26768_37700# vss nmos_6p0 w=0.82u l=0.6u
X5664 a_25572_33780# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5665 a_6740_32696# cap_shunt_n a_6532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X5666 a_21540_5180# cap_series_gyp a_21748_4834# vdd pmos_6p0 w=1.2u l=0.5u
X5667 vss tune_series_gygy[5] a_35880_16532# vss nmos_6p0 w=0.51u l=0.6u
X5668 a_17828_40536# cap_shunt_n a_17620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X5669 vdd a_37980_44712# a_37892_44756# vdd pmos_6p0 w=1.22u l=1u
X5670 a_10340_36916# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5671 a_10548_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5672 vss cap_shunt_n a_27104_40536# vss nmos_6p0 w=0.82u l=0.6u
X5673 a_20664_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5674 a_30632_4772# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5675 a_17620_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5676 vdd a_27676_11351# a_27588_11448# vdd pmos_6p0 w=1.22u l=1u
X5677 a_9428_18946# cap_shunt_p a_11144_18884# vss nmos_6p0 w=0.82u l=0.6u
X5678 a_6292_18946# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5679 a_25572_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5680 a_18404_5180# cap_series_gyp a_18612_4834# vdd pmos_6p0 w=1.2u l=0.5u
X5681 vss tune_series_gy[4] a_24660_9538# vss nmos_6p0 w=0.51u l=0.6u
X5682 a_16708_14242# cap_shunt_p a_18424_14180# vss nmos_6p0 w=0.82u l=0.6u
X5683 a_29492_36540# cap_shunt_n a_29700_36194# vdd pmos_6p0 w=1.2u l=0.5u
X5684 a_10452_34972# cap_shunt_n a_10660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X5685 a_26768_14180# cap_series_gyn a_24660_14242# vss nmos_6p0 w=0.82u l=0.6u
X5686 a_6532_40052# cap_shunt_n a_6740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X5687 a_37652_32996# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5688 vdd a_23308_55255# a_23220_55352# vdd pmos_6p0 w=1.22u l=1u
X5689 vdd a_11884_47415# a_11796_47512# vdd pmos_6p0 w=1.22u l=1u
X5690 a_6532_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5691 vdd tune_shunt[7] a_29492_27132# vdd pmos_6p0 w=1.2u l=0.5u
X5692 vss cap_shunt_p a_7616_51812# vss nmos_6p0 w=0.82u l=0.6u
X5693 a_37868_52119# a_37780_52216# vss vss nmos_6p0 w=0.82u l=1u
X5694 a_9856_45540# cap_shunt_p a_7748_45602# vss nmos_6p0 w=0.82u l=0.6u
X5695 a_20740_38968# cap_shunt_n a_20532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X5696 a_29492_33404# cap_shunt_p a_29700_33058# vdd pmos_6p0 w=1.2u l=0.5u
X5697 a_10452_31836# cap_shunt_n a_10660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X5698 a_12788_15448# cap_shunt_p a_12580_14964# vdd pmos_6p0 w=1.2u l=0.5u
X5699 a_26768_11044# cap_series_gyp a_24660_11106# vss nmos_6p0 w=0.82u l=0.6u
X5700 vdd a_10988_43144# a_10900_43188# vdd pmos_6p0 w=1.22u l=1u
X5701 a_31624_22428# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5702 vdd a_23756_44712# a_23668_44756# vdd pmos_6p0 w=1.22u l=1u
X5703 vdd a_23308_52119# a_23220_52216# vdd pmos_6p0 w=1.22u l=1u
X5704 a_18492_52119# a_18404_52216# vss vss nmos_6p0 w=0.82u l=1u
X5705 a_6532_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5706 a_4424_32996# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5707 vdd a_5612_6647# a_5524_6744# vdd pmos_6p0 w=1.22u l=1u
X5708 a_11780_4472# cap_series_gyp a_11572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X5709 a_14012_9783# a_13924_9880# vss vss nmos_6p0 w=0.82u l=1u
X5710 a_8064_21720# cap_shunt_p a_6740_21720# vss nmos_6p0 w=0.82u l=0.6u
X5711 a_9876_51512# cap_shunt_n a_9668_51028# vdd pmos_6p0 w=1.2u l=0.5u
X5712 vdd a_2588_41576# a_2500_41620# vdd pmos_6p0 w=1.22u l=1u
X5713 a_32380_43144# a_32292_43188# vss vss nmos_6p0 w=0.82u l=1u
X5714 a_9856_42404# cap_shunt_n a_7748_42466# vss nmos_6p0 w=0.82u l=0.6u
X5715 vss tune_shunt[6] a_24660_36194# vss nmos_6p0 w=0.51u l=0.6u
X5716 a_20740_35832# cap_shunt_n a_20532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X5717 vss cap_shunt_n a_8848_34264# vss nmos_6p0 w=0.82u l=0.6u
X5718 a_12788_12312# cap_shunt_p a_12580_11828# vdd pmos_6p0 w=1.2u l=0.5u
X5719 vdd tune_series_gy[4] a_32444_14588# vdd pmos_6p0 w=1.2u l=0.5u
X5720 a_6956_34871# a_6868_34968# vss vss nmos_6p0 w=0.82u l=1u
X5721 a_21748_12674# cap_series_gyn a_21540_13020# vdd pmos_6p0 w=1.2u l=0.5u
X5722 a_29700_11106# cap_series_gyp a_29492_11452# vdd pmos_6p0 w=1.2u l=0.5u
X5723 vdd tune_shunt[7] a_13588_17724# vdd pmos_6p0 w=1.2u l=0.5u
X5724 a_9644_5512# a_9556_5556# vss vss nmos_6p0 w=0.82u l=1u
X5725 vss tune_series_gy[4] a_29720_16156# vss nmos_6p0 w=0.51u l=0.6u
X5726 vdd a_4940_5512# a_4852_5556# vdd pmos_6p0 w=1.22u l=1u
X5727 a_33500_21192# a_33412_21236# vss vss nmos_6p0 w=0.82u l=1u
X5728 a_16708_39330# cap_shunt_n a_17640_39268# vss nmos_6p0 w=0.82u l=0.6u
X5729 vss tune_shunt[6] a_24660_33058# vss nmos_6p0 w=0.51u l=0.6u
X5730 vss cap_shunt_n a_8848_31128# vss nmos_6p0 w=0.82u l=0.6u
X5731 a_6956_31735# a_6868_31832# vss vss nmos_6p0 w=0.82u l=1u
X5732 a_2708_25218# cap_shunt_p a_2500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X5733 a_6292_51874# cap_shunt_p a_6084_52220# vdd pmos_6p0 w=1.2u l=0.5u
X5734 a_6404_47170# cap_shunt_p a_6196_47516# vdd pmos_6p0 w=1.2u l=0.5u
X5735 vdd tune_shunt[6] a_9108_47516# vdd pmos_6p0 w=1.2u l=0.5u
X5736 a_36384_47512# cap_shunt_gyp a_36384_47108# vdd pmos_6p0 w=1.215u l=0.5u
X5737 a_31624_19292# cap_series_gygyn a_31436_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5738 a_16800_6040# cap_series_gyn a_14692_6040# vss nmos_6p0 w=0.82u l=0.6u
X5739 a_14692_9176# cap_series_gyn a_14484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X5740 vdd a_28124_17623# a_28036_17720# vdd pmos_6p0 w=1.22u l=1u
X5741 a_2708_22082# cap_shunt_p a_2500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5742 a_9876_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5743 a_6292_17378# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5744 a_37632_49080# cap_shunt_gyn a_37444_49080# vdd pmos_6p0 w=1.215u l=0.5u
X5745 a_32716_49416# a_32628_49460# vss vss nmos_6p0 w=0.82u l=1u
X5746 a_20740_45240# cap_shunt_n a_20532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X5747 a_4032_9476# cap_shunt_n a_2708_9538# vss nmos_6p0 w=0.82u l=0.6u
X5748 vss cap_shunt_gyp a_32732_45240# vss nmos_6p0 w=0.82u l=0.6u
X5749 a_22860_55255# a_22772_55352# vss vss nmos_6p0 w=0.82u l=1u
X5750 a_14692_6040# cap_series_gyn a_14484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X5751 vss tune_series_gy[5] a_19732_12312# vss nmos_6p0 w=0.51u l=0.6u
X5752 a_18940_53687# a_18852_53784# vss vss nmos_6p0 w=0.82u l=1u
X5753 a_34516_22082# cap_series_gygyp a_34308_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5754 a_9876_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5755 vss tune_shunt[5] a_12788_49944# vss nmos_6p0 w=0.51u l=0.6u
X5756 a_31624_20860# cap_series_gygyn a_31436_20860# vdd pmos_6p0 w=1.2u l=0.5u
X5757 a_1692_52119# a_1604_52216# vss vss nmos_6p0 w=0.82u l=1u
X5758 vdd tune_shunt[6] a_14372_46324# vdd pmos_6p0 w=1.2u l=0.5u
X5759 vss cap_shunt_p a_27104_34264# vss nmos_6p0 w=0.82u l=0.6u
X5760 a_10248_50244# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5761 a_16500_47516# cap_shunt_n a_16708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X5762 a_6196_22428# cap_shunt_p a_6404_22082# vdd pmos_6p0 w=1.2u l=0.5u
X5763 a_2708_34626# cap_shunt_n a_2500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X5764 a_35448_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5765 a_25572_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5766 a_10340_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5767 a_13588_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5768 vss cap_shunt_p a_27104_31128# vss nmos_6p0 w=0.82u l=0.6u
X5769 a_25984_29860# cap_shunt_n a_24660_29922# vss nmos_6p0 w=0.82u l=0.6u
X5770 vdd a_13340_10216# a_13252_10260# vdd pmos_6p0 w=1.22u l=1u
X5771 vdd a_23308_48983# a_23220_49080# vdd pmos_6p0 w=1.22u l=1u
X5772 a_2708_31490# cap_shunt_p a_2500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X5773 a_35448_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5774 a_18388_3266# cap_series_gyn a_18180_3612# vdd pmos_6p0 w=1.2u l=0.5u
X5775 a_25572_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5776 a_25780_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5777 a_10452_25564# cap_shunt_n a_10660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X5778 a_16708_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5779 a_29492_27132# cap_shunt_p a_29700_26786# vdd pmos_6p0 w=1.2u l=0.5u
X5780 a_9668_18100# cap_shunt_p a_9876_18584# vdd pmos_6p0 w=1.2u l=0.5u
X5781 a_3864_9176# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5782 a_9332_14588# cap_shunt_p a_9540_14242# vdd pmos_6p0 w=1.2u l=0.5u
X5783 vss tune_shunt[6] a_24660_39330# vss nmos_6p0 w=0.51u l=0.6u
X5784 vdd a_23756_38440# a_23668_38484# vdd pmos_6p0 w=1.22u l=1u
X5785 a_13588_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5786 a_25984_26724# cap_shunt_p a_24660_26786# vss nmos_6p0 w=0.82u l=0.6u
X5787 a_6532_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5788 a_10452_5180# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5789 a_5936_43672# cap_shunt_p a_3828_43672# vss nmos_6p0 w=0.82u l=0.6u
X5790 a_34536_9884# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X5791 a_6628_14242# cap_shunt_p a_6420_14588# vdd pmos_6p0 w=1.2u l=0.5u
X5792 vdd a_16700_16488# a_16612_16532# vdd pmos_6p0 w=1.22u l=1u
X5793 a_14896_17016# cap_shunt_p a_12788_17016# vss nmos_6p0 w=0.82u l=0.6u
X5794 a_9856_36132# cap_shunt_n a_7748_36194# vss nmos_6p0 w=0.82u l=0.6u
X5795 vdd a_20284_53687# a_20196_53784# vdd pmos_6p0 w=1.22u l=1u
X5796 a_20740_29560# cap_shunt_n a_20532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X5797 a_25572_3988# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5798 vss cap_series_gyn a_8184_7908# vss nmos_6p0 w=0.82u l=0.6u
X5799 a_15532_11452# cap_series_gyp a_15720_11452# vdd pmos_6p0 w=1.2u l=0.5u
X5800 a_6956_28599# a_6868_28696# vss vss nmos_6p0 w=0.82u l=1u
X5801 a_37868_6647# a_37780_6744# vss vss nmos_6p0 w=0.82u l=1u
X5802 a_13796_12674# cap_shunt_p a_13588_13020# vdd pmos_6p0 w=1.2u l=0.5u
X5803 vdd a_23756_35304# a_23668_35348# vdd pmos_6p0 w=1.22u l=1u
X5804 a_16500_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5805 a_10660_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5806 a_25780_9176# cap_series_gyp a_27496_9176# vss nmos_6p0 w=0.82u l=0.6u
X5807 a_8064_12312# cap_shunt_p a_6740_12312# vss nmos_6p0 w=0.82u l=0.6u
X5808 a_14728_48676# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5809 a_5936_40536# cap_shunt_n a_3828_40536# vss nmos_6p0 w=0.82u l=0.6u
X5810 a_4424_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5811 vss tune_series_gy[4] a_21748_6402# vss nmos_6p0 w=0.51u l=0.6u
X5812 vdd a_2588_32168# a_2500_32212# vdd pmos_6p0 w=1.22u l=1u
X5813 a_3248_4772# cap_shunt_p a_1924_4834# vss nmos_6p0 w=0.82u l=0.6u
X5814 a_6956_25463# a_6868_25560# vss vss nmos_6p0 w=0.82u l=1u
X5815 a_37868_3511# a_37780_3608# vss vss nmos_6p0 w=0.82u l=1u
X5816 a_2708_18946# cap_shunt_p a_2500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5817 a_26712_4472# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5818 a_19732_10744# cap_series_gyn a_19524_10260# vdd pmos_6p0 w=1.2u l=0.5u
X5819 a_16708_34626# cap_shunt_n a_16500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X5820 a_3640_4472# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5821 a_2708_44034# cap_shunt_p a_3640_43972# vss nmos_6p0 w=0.82u l=0.6u
X5822 a_10452_34972# cap_shunt_n a_10660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X5823 a_33500_11784# a_33412_11828# vss vss nmos_6p0 w=0.82u l=1u
X5824 a_6532_40052# cap_shunt_n a_6740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X5825 vss tune_shunt[7] a_13796_29922# vss nmos_6p0 w=0.51u l=0.6u
X5826 vdd tune_shunt[2] a_1716_8316# vdd pmos_6p0 w=1.2u l=0.5u
X5827 a_15904_18884# cap_shunt_p a_13796_18946# vss nmos_6p0 w=0.82u l=0.6u
X5828 a_2708_15810# cap_shunt_p a_2500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X5829 a_34516_18946# cap_series_gygyn a_34308_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5830 a_20620_20759# a_20532_20856# vss vss nmos_6p0 w=0.82u l=1u
X5831 a_9316_50306# cap_shunt_p a_11032_50244# vss nmos_6p0 w=0.82u l=0.6u
X5832 a_2588_27464# a_2500_27508# vss vss nmos_6p0 w=0.82u l=1u
X5833 vdd a_2140_34871# a_2052_34968# vdd pmos_6p0 w=1.22u l=1u
X5834 a_16708_31490# cap_shunt_n a_16500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X5835 a_15700_6402# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X5836 a_25572_8692# cap_series_gyp a_25780_9176# vdd pmos_6p0 w=1.2u l=0.5u
X5837 a_20740_38968# cap_shunt_n a_20532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X5838 a_10452_31836# cap_shunt_n a_10660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X5839 a_2708_40898# cap_shunt_p a_3640_40836# vss nmos_6p0 w=0.82u l=0.6u
X5840 a_6404_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5841 a_15492_9884# cap_series_gyn a_15700_9538# vdd pmos_6p0 w=1.2u l=0.5u
X5842 a_35840_20452# cap_series_gygyp a_34516_20514# vss nmos_6p0 w=0.82u l=0.6u
X5843 a_37084_52552# a_36996_52596# vss vss nmos_6p0 w=0.82u l=1u
X5844 a_6740_45240# cap_shunt_p a_7672_45240# vss nmos_6p0 w=0.82u l=0.6u
X5845 vss tune_shunt[7] a_9540_15810# vss nmos_6p0 w=0.51u l=0.6u
X5846 a_22860_48983# a_22772_49080# vss vss nmos_6p0 w=0.82u l=1u
X5847 a_15904_15748# cap_shunt_p a_13796_15810# vss nmos_6p0 w=0.82u l=0.6u
X5848 a_34516_15810# cap_series_gygyn a_34308_16156# vdd pmos_6p0 w=1.2u l=0.5u
X5849 a_9876_51512# cap_shunt_n a_9668_51028# vdd pmos_6p0 w=1.2u l=0.5u
X5850 a_2588_24328# a_2500_24372# vss vss nmos_6p0 w=0.82u l=1u
X5851 vdd a_30364_55255# a_30276_55352# vdd pmos_6p0 w=1.22u l=1u
X5852 a_36988_49944# cap_shunt_gyp a_36720_50006# vss nmos_6p0 w=0.82u l=0.6u
X5853 a_2500_47516# cap_shunt_p a_2708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X5854 a_1692_45847# a_1604_45944# vss vss nmos_6p0 w=0.82u l=1u
X5855 a_25572_5556# cap_series_gyp a_25780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X5856 a_30016_13880# cap_series_gyp a_28692_13880# vss nmos_6p0 w=0.82u l=0.6u
X5857 a_2708_50306# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5858 a_20740_35832# cap_shunt_n a_20532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X5859 a_11592_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5860 vss tune_shunt[7] a_7748_23650# vss nmos_6p0 w=0.51u l=0.6u
X5861 a_15492_6748# cap_series_gyp a_15700_6402# vdd pmos_6p0 w=1.2u l=0.5u
X5862 a_6740_42104# cap_shunt_n a_7672_42104# vss nmos_6p0 w=0.82u l=0.6u
X5863 a_6084_49084# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5864 vss tune_series_gy[4] a_14692_10744# vss nmos_6p0 w=0.51u l=0.6u
X5865 a_17708_12919# a_17620_13016# vss vss nmos_6p0 w=0.82u l=1u
X5866 vdd a_28124_9783# a_28036_9880# vdd pmos_6p0 w=1.22u l=1u
X5867 vdd a_30364_52119# a_30276_52216# vdd pmos_6p0 w=1.22u l=1u
X5868 a_36988_46808# cap_shunt_gyp a_36720_46870# vss nmos_6p0 w=0.82u l=0.6u
X5869 a_1692_42711# a_1604_42808# vss vss nmos_6p0 w=0.82u l=1u
X5870 a_30016_10744# cap_series_gyp a_28692_10744# vss nmos_6p0 w=0.82u l=0.6u
X5871 vdd tune_shunt[7] a_6532_13396# vdd pmos_6p0 w=1.2u l=0.5u
X5872 a_3828_13880# cap_shunt_n a_3620_13396# vdd pmos_6p0 w=1.2u l=0.5u
X5873 a_30408_12312# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X5874 vdd a_33500_53687# a_33412_53784# vdd pmos_6p0 w=1.22u l=1u
X5875 a_16500_38108# cap_shunt_n a_16708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X5876 a_19724_33303# a_19636_33400# vss vss nmos_6p0 w=0.82u l=1u
X5877 a_3620_47892# cap_shunt_p a_3828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X5878 a_2708_25218# cap_shunt_p a_2500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X5879 a_21628_50984# a_21540_51028# vss vss nmos_6p0 w=0.82u l=1u
X5880 a_6404_47170# cap_shunt_p a_6196_47516# vdd pmos_6p0 w=1.2u l=0.5u
X5881 a_20532_43188# cap_shunt_n a_20740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X5882 vdd tune_shunt[6] a_21540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X5883 vdd a_19276_47415# a_19188_47512# vdd pmos_6p0 w=1.22u l=1u
X5884 a_16708_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5885 vdd a_28124_6647# a_28036_6744# vdd pmos_6p0 w=1.22u l=1u
X5886 a_22064_27992# cap_shunt_n a_20740_27992# vss nmos_6p0 w=0.82u l=0.6u
X5887 a_13796_48738# cap_shunt_n a_15512_48676# vss nmos_6p0 w=0.82u l=0.6u
X5888 a_13588_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5889 vdd a_33500_50551# a_33412_50648# vdd pmos_6p0 w=1.22u l=1u
X5890 a_31624_6748# cap_series_gygyn a_31436_6748# vdd pmos_6p0 w=1.2u l=0.5u
X5891 vdd a_3484_54120# a_3396_54164# vdd pmos_6p0 w=1.22u l=1u
X5892 vss tune_shunt[5] a_9876_51512# vss nmos_6p0 w=0.51u l=0.6u
X5893 a_3620_44756# cap_shunt_p a_3828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X5894 a_2708_22082# cap_shunt_p a_2500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5895 a_37868_36439# a_37780_36536# vss vss nmos_6p0 w=0.82u l=1u
X5896 a_19544_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5897 a_22064_24856# cap_shunt_n a_20740_24856# vss nmos_6p0 w=0.82u l=0.6u
X5898 a_13588_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5899 a_9540_12674# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X5900 a_34308_17724# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5901 vdd a_23756_29032# a_23668_29076# vdd pmos_6p0 w=1.22u l=1u
X5902 a_25984_17316# cap_series_gyp a_24660_17378# vss nmos_6p0 w=0.82u l=0.6u
X5903 a_33948_40008# a_33860_40052# vss vss nmos_6p0 w=0.82u l=1u
X5904 a_10340_32212# cap_shunt_n a_10548_32696# vdd pmos_6p0 w=1.2u l=0.5u
X5905 a_5936_34264# cap_shunt_n a_3828_34264# vss nmos_6p0 w=0.82u l=0.6u
X5906 a_34516_22082# cap_series_gygyp a_34308_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5907 vdd tune_shunt[5] a_6532_52596# vdd pmos_6p0 w=1.2u l=0.5u
X5908 vdd tune_series_gy[4] a_18404_5180# vdd pmos_6p0 w=1.2u l=0.5u
X5909 a_19544_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5910 a_6196_22428# cap_shunt_p a_6404_22082# vdd pmos_6p0 w=1.2u l=0.5u
X5911 a_16500_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5912 a_11668_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5913 a_14728_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5914 a_5936_31128# cap_shunt_n a_3828_31128# vss nmos_6p0 w=0.82u l=0.6u
X5915 a_28692_40536# cap_shunt_p a_29624_40536# vss nmos_6p0 w=0.82u l=0.6u
X5916 a_11996_20759# a_11908_20856# vss vss nmos_6p0 w=0.82u l=1u
X5917 a_24452_20860# cap_shunt_p a_24660_20514# vdd pmos_6p0 w=1.2u l=0.5u
X5918 a_8456_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X5919 vdd a_33052_42711# a_32964_42808# vdd pmos_6p0 w=1.22u l=1u
X5920 a_24660_9538# cap_series_gyn a_26376_9476# vss nmos_6p0 w=0.82u l=0.6u
X5921 a_9540_11106# cap_shunt_p a_9332_11452# vdd pmos_6p0 w=1.2u l=0.5u
X5922 a_7952_12612# cap_shunt_p a_6628_12674# vss nmos_6p0 w=0.82u l=0.6u
X5923 a_19732_9176# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5924 a_20620_14487# a_20532_14584# vss vss nmos_6p0 w=0.82u l=1u
X5925 a_11668_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5926 vdd a_2140_28599# a_2052_28696# vdd pmos_6p0 w=1.22u l=1u
X5927 a_16708_25218# cap_shunt_n a_16500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X5928 a_10452_25564# cap_shunt_n a_10660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X5929 a_30428_21236# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5930 vdd a_19724_48983# a_19636_49080# vdd pmos_6p0 w=1.22u l=1u
X5931 a_2708_47170# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X5932 vss tune_shunt[5] a_17828_46808# vss nmos_6p0 w=0.51u l=0.6u
X5933 a_2708_34626# cap_shunt_n a_3640_34564# vss nmos_6p0 w=0.82u l=0.6u
X5934 vdd tune_series_gy[4] a_22436_7124# vdd pmos_6p0 w=1.2u l=0.5u
X5935 a_25592_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X5936 vdd tune_series_gygy[1] a_31436_8316# vdd pmos_6p0 w=1.2u l=0.5u
X5937 a_2588_18056# a_2500_18100# vss vss nmos_6p0 w=0.82u l=1u
X5938 a_6740_27992# cap_shunt_n a_8456_27992# vss nmos_6p0 w=0.82u l=0.6u
X5939 a_16708_22082# cap_shunt_n a_16500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X5940 vdd a_30364_48983# a_30276_49080# vdd pmos_6p0 w=1.22u l=1u
X5941 a_4492_7080# a_4404_7124# vss vss nmos_6p0 w=0.82u l=1u
X5942 a_24652_44712# a_24564_44756# vss vss nmos_6p0 w=0.82u l=1u
X5943 a_2708_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5944 a_2708_31490# cap_shunt_p a_3640_31428# vss nmos_6p0 w=0.82u l=0.6u
X5945 a_20740_29560# cap_shunt_n a_20532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X5946 vss tune_shunt[4] a_29700_39330# vss nmos_6p0 w=0.51u l=0.6u
X5947 a_13796_12674# cap_shunt_p a_13588_13020# vdd pmos_6p0 w=1.2u l=0.5u
X5948 a_14580_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5949 a_13900_3511# a_13812_3608# vss vss nmos_6p0 w=0.82u l=1u
X5950 vdd a_5612_45847# a_5524_45944# vdd pmos_6p0 w=1.22u l=1u
X5951 a_2588_14920# a_2500_14964# vss vss nmos_6p0 w=0.82u l=1u
X5952 a_35740_52119# a_35652_52216# vss vss nmos_6p0 w=0.82u l=1u
X5953 a_1692_36439# a_1604_36536# vss vss nmos_6p0 w=0.82u l=1u
X5954 a_17828_32696# cap_shunt_n a_19544_32696# vss nmos_6p0 w=0.82u l=0.6u
X5955 a_6740_24856# cap_shunt_p a_8456_24856# vss nmos_6p0 w=0.82u l=0.6u
X5956 a_2500_38108# cap_shunt_n a_2708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X5957 a_27888_32696# cap_shunt_p a_25780_32696# vss nmos_6p0 w=0.82u l=0.6u
X5958 a_24652_41576# a_24564_41620# vss vss nmos_6p0 w=0.82u l=1u
X5959 a_2708_18946# cap_shunt_p a_2500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5960 a_32828_41576# a_32740_41620# vss vss nmos_6p0 w=0.82u l=1u
X5961 a_7748_28354# cap_shunt_n a_7540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X5962 a_19732_10744# cap_series_gyn a_19524_10260# vdd pmos_6p0 w=1.2u l=0.5u
X5963 a_12580_13396# cap_shunt_p a_12788_13880# vdd pmos_6p0 w=1.2u l=0.5u
X5964 a_10808_53080# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X5965 vdd a_5612_42711# a_5524_42808# vdd pmos_6p0 w=1.22u l=1u
X5966 a_10452_34972# cap_shunt_n a_10660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X5967 a_22436_11828# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5968 vss cap_series_gyn a_21056_12312# vss nmos_6p0 w=0.82u l=0.6u
X5969 a_12788_48376# cap_shunt_p a_12580_47892# vdd pmos_6p0 w=1.2u l=0.5u
X5970 a_17828_46808# cap_shunt_n a_18760_46808# vss nmos_6p0 w=0.82u l=0.6u
X5971 a_13252_38484# cap_shunt_n a_13460_38968# vdd pmos_6p0 w=1.2u l=0.5u
X5972 a_37632_47512# cap_shunt_gyp a_37652_47108# vss nmos_6p0 w=0.82u l=0.6u
X5973 a_2500_42812# cap_shunt_p a_2708_42466# vdd pmos_6p0 w=1.2u l=0.5u
X5974 a_6532_40052# cap_shunt_n a_6740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X5975 a_24452_28700# cap_shunt_n a_24660_28354# vdd pmos_6p0 w=1.2u l=0.5u
X5976 a_13588_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5977 a_3620_38484# cap_shunt_n a_3828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X5978 a_19724_23895# a_19636_23992# vss vss nmos_6p0 w=0.82u l=1u
X5979 a_5844_3266# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X5980 a_2708_15810# cap_shunt_p a_2500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X5981 a_34516_18946# cap_series_gygyn a_34308_19292# vdd pmos_6p0 w=1.2u l=0.5u
X5982 vdd a_31036_43144# a_30948_43188# vdd pmos_6p0 w=1.22u l=1u
X5983 vdd a_19276_38007# a_19188_38104# vdd pmos_6p0 w=1.22u l=1u
X5984 a_10452_31836# cap_shunt_n a_10660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X5985 vdd a_27228_30167# a_27140_30264# vdd pmos_6p0 w=1.22u l=1u
X5986 a_28692_7608# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X5987 a_22064_18584# cap_shunt_p a_20740_18584# vss nmos_6p0 w=0.82u l=0.6u
X5988 a_13252_35348# cap_shunt_n a_13460_35832# vdd pmos_6p0 w=1.2u l=0.5u
X5989 a_21516_52119# a_21428_52216# vss vss nmos_6p0 w=0.82u l=1u
X5990 a_10660_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X5991 a_13796_39330# cap_shunt_n a_15512_39268# vss nmos_6p0 w=0.82u l=0.6u
X5992 vss cap_series_gyn a_20496_3204# vss nmos_6p0 w=0.82u l=0.6u
X5993 a_13588_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X5994 vss cap_shunt_p a_8400_18884# vss nmos_6p0 w=0.82u l=0.6u
X5995 a_23856_39268# cap_shunt_p a_21748_39330# vss nmos_6p0 w=0.82u l=0.6u
X5996 a_35880_18100# cap_series_gygyn a_35692_18100# vdd pmos_6p0 w=1.2u l=0.5u
X5997 a_3620_35348# cap_shunt_n a_3828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X5998 a_34516_15810# cap_series_gygyn a_34308_16156# vdd pmos_6p0 w=1.2u l=0.5u
X5999 a_12580_16532# cap_shunt_p a_12788_17016# vdd pmos_6p0 w=1.2u l=0.5u
X6000 a_22064_15448# cap_series_gyn a_20740_15448# vss nmos_6p0 w=0.82u l=0.6u
X6001 a_19276_19191# a_19188_19288# vss vss nmos_6p0 w=0.82u l=1u
X6002 a_25780_9176# cap_series_gyp a_25572_8692# vdd pmos_6p0 w=1.2u l=0.5u
X6003 vss cap_shunt_p a_8400_15748# vss nmos_6p0 w=0.82u l=0.6u
X6004 a_6084_49084# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6005 a_34348_9884# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6006 a_15700_9538# cap_series_gyn a_15492_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6007 vdd tune_shunt[6] a_13588_47516# vdd pmos_6p0 w=1.2u l=0.5u
X6008 a_13796_22082# cap_shunt_n a_14728_22020# vss nmos_6p0 w=0.82u l=0.6u
X6009 a_28692_34264# cap_shunt_p a_29624_34264# vss nmos_6p0 w=0.82u l=0.6u
X6010 vss cap_shunt_p a_23856_18884# vss nmos_6p0 w=0.82u l=0.6u
X6011 a_34396_54120# a_34308_54164# vss vss nmos_6p0 w=0.82u l=1u
X6012 vdd tune_shunt[6] a_6532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X6013 a_19276_16055# a_19188_16152# vss vss nmos_6p0 w=0.82u l=1u
X6014 a_3828_20152# cap_shunt_p a_3620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X6015 a_10660_37762# cap_shunt_n a_10452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X6016 a_25780_6040# cap_series_gyp a_25572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X6017 a_6404_47170# cap_shunt_p a_6196_47516# vdd pmos_6p0 w=1.2u l=0.5u
X6018 a_20532_43188# cap_shunt_n a_20740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X6019 a_15700_6402# cap_series_gyp a_15492_6748# vdd pmos_6p0 w=1.2u l=0.5u
X6020 a_34348_6748# tune_series_gygy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6021 a_16708_18946# cap_shunt_p a_16500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X6022 a_2708_28354# cap_shunt_n a_3640_28292# vss nmos_6p0 w=0.82u l=0.6u
X6023 vdd a_37420_5079# a_37332_5176# vdd pmos_6p0 w=1.22u l=1u
X6024 vdd a_23756_55255# a_23668_55352# vdd pmos_6p0 w=1.22u l=1u
X6025 a_28692_31128# cap_shunt_n a_29624_31128# vss nmos_6p0 w=0.82u l=0.6u
X6026 a_2932_10744# cap_shunt_n a_3864_10744# vss nmos_6p0 w=0.82u l=0.6u
X6027 vss cap_series_gyn a_23856_15748# vss nmos_6p0 w=0.82u l=0.6u
X6028 a_18032_20452# cap_shunt_p a_16708_20514# vss nmos_6p0 w=0.82u l=0.6u
X6029 a_24452_11452# cap_series_gyp a_24660_11106# vdd pmos_6p0 w=1.2u l=0.5u
X6030 a_16708_15810# cap_shunt_p a_16500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X6031 vdd a_2140_19191# a_2052_19288# vdd pmos_6p0 w=1.22u l=1u
X6032 a_2708_25218# cap_shunt_p a_3640_25156# vss nmos_6p0 w=0.82u l=0.6u
X6033 a_31624_22428# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6034 vdd a_23756_52119# a_23668_52216# vdd pmos_6p0 w=1.22u l=1u
X6035 a_14468_3266# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X6036 a_15568_34264# cap_shunt_n a_13460_34264# vss nmos_6p0 w=0.82u l=0.6u
X6037 a_22436_10260# cap_series_gyp a_22644_10744# vdd pmos_6p0 w=1.2u l=0.5u
X6038 a_6572_5556# cap_series_gyp a_6760_5556# vdd pmos_6p0 w=1.2u l=0.5u
X6039 a_5488_17016# cap_shunt_p a_3380_17016# vss nmos_6p0 w=0.82u l=0.6u
X6040 vdd a_5612_39575# a_5524_39672# vdd pmos_6p0 w=1.22u l=1u
X6041 a_24660_42466# cap_shunt_n a_24452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X6042 vss tune_shunt[7] a_21748_26786# vss nmos_6p0 w=0.51u l=0.6u
X6043 vss tune_shunt[7] a_6740_21720# vss nmos_6p0 w=0.51u l=0.6u
X6044 a_11668_46808# cap_shunt_n a_11460_46324# vdd pmos_6p0 w=1.2u l=0.5u
X6045 a_2500_30268# cap_shunt_n a_2708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X6046 vdd tune_series_gy[4] a_18516_5556# vdd pmos_6p0 w=1.2u l=0.5u
X6047 a_15568_31128# cap_shunt_n a_13460_31128# vss nmos_6p0 w=0.82u l=0.6u
X6048 vdd a_5612_36439# a_5524_36536# vdd pmos_6p0 w=1.22u l=1u
X6049 vss cap_shunt_p a_31024_34564# vss nmos_6p0 w=0.82u l=0.6u
X6050 vss cap_shunt_p a_16688_46808# vss nmos_6p0 w=0.82u l=0.6u
X6051 a_17596_8648# a_17508_8692# vss vss nmos_6p0 w=0.82u l=1u
X6052 a_6740_15448# cap_shunt_p a_8456_15448# vss nmos_6p0 w=0.82u l=0.6u
X6053 a_2500_36540# cap_shunt_n a_2708_36194# vdd pmos_6p0 w=1.2u l=0.5u
X6054 a_17828_23288# cap_shunt_n a_19544_23288# vss nmos_6p0 w=0.82u l=0.6u
X6055 a_35880_7124# cap_series_gygyp a_35692_7124# vdd pmos_6p0 w=1.2u l=0.5u
X6056 a_29624_9176# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X6057 a_16500_28700# cap_shunt_n a_16708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X6058 a_27888_23288# cap_shunt_p a_25780_23288# vss nmos_6p0 w=0.82u l=0.6u
X6059 a_24452_20860# cap_shunt_p a_24660_20514# vdd pmos_6p0 w=1.2u l=0.5u
X6060 a_28692_7608# cap_series_gyp a_28484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X6061 a_17828_20152# cap_shunt_p a_17620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X6062 a_18612_7970# cap_series_gyp a_18404_8316# vdd pmos_6p0 w=1.2u l=0.5u
X6063 vss cap_shunt_p a_31024_31428# vss nmos_6p0 w=0.82u l=0.6u
X6064 a_10452_25564# cap_shunt_n a_10660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X6065 a_30428_21236# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6066 a_13252_29076# cap_shunt_n a_13460_29560# vdd pmos_6p0 w=1.2u l=0.5u
X6067 vdd a_28572_17623# a_28484_17720# vdd pmos_6p0 w=1.22u l=1u
X6068 a_10660_36194# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6069 a_2500_33404# cap_shunt_p a_2708_33058# vdd pmos_6p0 w=1.2u l=0.5u
X6070 vdd a_10988_8648# a_10900_8692# vdd pmos_6p0 w=1.22u l=1u
X6071 a_3620_29076# cap_shunt_n a_3828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X6072 a_2708_9538# cap_shunt_n a_2500_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6073 vdd a_37532_54120# a_37444_54164# vdd pmos_6p0 w=1.22u l=1u
X6074 a_35040_43189# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X6075 vdd tune_series_gy[4] a_18404_5180# vdd pmos_6p0 w=1.2u l=0.5u
X6076 a_6532_19668# cap_shunt_p a_6740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X6077 a_10548_3266# cap_series_gyn a_10340_3612# vdd pmos_6p0 w=1.2u l=0.5u
X6078 a_10660_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6079 vdd a_10988_5512# a_10900_5556# vdd pmos_6p0 w=1.22u l=1u
X6080 vdd a_13900_55688# a_13812_55732# vdd pmos_6p0 w=1.22u l=1u
X6081 a_17620_25940# cap_shunt_n a_17828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X6082 a_35692_19668# cap_series_gygyp a_35880_19668# vdd pmos_6p0 w=1.2u l=0.5u
X6083 a_7748_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6084 a_18388_3266# cap_series_gyn a_18180_3612# vdd pmos_6p0 w=1.2u l=0.5u
X6085 a_30408_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6086 vdd tune_series_gy[0] a_29196_3612# vdd pmos_6p0 w=1.2u l=0.5u
X6087 vdd tune_shunt[2] a_1716_6748# vdd pmos_6p0 w=1.2u l=0.5u
X6088 a_9332_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6089 a_7748_28354# cap_shunt_n a_7540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X6090 a_9876_20152# cap_shunt_p a_10808_20152# vss nmos_6p0 w=0.82u l=0.6u
X6091 vdd a_10092_41576# a_10004_41620# vdd pmos_6p0 w=1.22u l=1u
X6092 a_12580_13396# cap_shunt_p a_12788_13880# vdd pmos_6p0 w=1.2u l=0.5u
X6093 vdd tune_shunt[7] a_13588_38108# vdd pmos_6p0 w=1.2u l=0.5u
X6094 vdd tune_shunt[7] a_21540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X6095 a_17620_22804# cap_shunt_n a_17828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X6096 a_23744_6040# cap_series_gyp a_21636_6040# vss nmos_6p0 w=0.82u l=0.6u
X6097 a_10752_18884# cap_shunt_p a_9428_18946# vss nmos_6p0 w=0.82u l=0.6u
X6098 vdd a_23756_48983# a_23668_49080# vdd pmos_6p0 w=1.22u l=1u
X6099 a_13252_38484# cap_shunt_n a_13460_38968# vdd pmos_6p0 w=1.2u l=0.5u
X6100 a_29720_13020# cap_series_gyn a_29532_13020# vdd pmos_6p0 w=1.2u l=0.5u
X6101 a_18032_14180# cap_shunt_p a_16708_14242# vss nmos_6p0 w=0.82u l=0.6u
X6102 a_9316_48738# cap_shunt_p a_9108_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6103 vss cap_series_gyp a_23856_7908# vss nmos_6p0 w=0.82u l=0.6u
X6104 vdd a_15132_50984# a_15044_51028# vdd pmos_6p0 w=1.22u l=1u
X6105 a_36384_48676# cap_shunt_gyn a_36384_49080# vdd pmos_6p0 w=1.215u l=0.5u
X6106 vss tune_shunt[6] a_9876_48376# vss nmos_6p0 w=0.51u l=0.6u
X6107 a_13252_35348# cap_shunt_n a_13460_35832# vdd pmos_6p0 w=1.2u l=0.5u
X6108 a_13796_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6109 vdd a_18044_11784# a_17956_11828# vdd pmos_6p0 w=1.22u l=1u
X6110 a_35880_18100# cap_series_gygyn a_35692_18100# vdd pmos_6p0 w=1.2u l=0.5u
X6111 a_24660_36194# cap_shunt_p a_24452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X6112 a_25572_10260# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6113 a_2708_20514# cap_shunt_p a_2500_20860# vdd pmos_6p0 w=1.2u l=0.5u
X6114 a_9668_52596# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6115 a_20532_14964# cap_series_gyn a_20740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X6116 vss tune_shunt[6] a_28692_37400# vss nmos_6p0 w=0.51u l=0.6u
X6117 a_32612_34626# cap_shunt_n a_32404_34972# vdd pmos_6p0 w=1.2u l=0.5u
X6118 a_8400_17316# cap_shunt_p a_6292_17378# vss nmos_6p0 w=0.82u l=0.6u
X6119 a_8184_6340# cap_series_gyp a_7768_6748# vss nmos_6p0 w=0.82u l=0.6u
X6120 a_24660_33058# cap_shunt_p a_24452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X6121 vss cap_shunt_p a_31024_28292# vss nmos_6p0 w=0.82u l=0.6u
X6122 a_21428_5556# cap_series_gyp a_21636_6040# vdd pmos_6p0 w=1.2u l=0.5u
X6123 a_15512_12612# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6124 a_7748_29922# cap_shunt_n a_7540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X6125 vss tune_shunt[7] a_6740_12312# vss nmos_6p0 w=0.51u l=0.6u
X6126 vss tune_shunt[4] a_21748_17378# vss nmos_6p0 w=0.51u l=0.6u
X6127 vdd tune_shunt[6] a_2500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X6128 a_32612_31490# cap_shunt_n a_32404_31836# vdd pmos_6p0 w=1.2u l=0.5u
X6129 vdd tune_shunt[4] a_25572_41620# vdd pmos_6p0 w=1.2u l=0.5u
X6130 a_27228_39575# a_27140_39672# vss vss nmos_6p0 w=0.82u l=1u
X6131 a_37084_38440# a_36996_38484# vss vss nmos_6p0 w=0.82u l=1u
X6132 vss tune_shunt[7] a_10660_31490# vss nmos_6p0 w=0.51u l=0.6u
X6133 a_1924_7970# cap_shunt_n a_1716_8316# vdd pmos_6p0 w=1.2u l=0.5u
X6134 a_14908_52119# a_14820_52216# vss vss nmos_6p0 w=0.82u l=1u
X6135 vdd a_33948_36872# a_33860_36916# vdd pmos_6p0 w=1.22u l=1u
X6136 a_29468_22327# a_29380_22424# vss vss nmos_6p0 w=0.82u l=1u
X6137 vdd a_14908_9783# a_14820_9880# vdd pmos_6p0 w=1.22u l=1u
X6138 a_27104_38968# cap_shunt_p a_25780_38968# vss nmos_6p0 w=0.82u l=0.6u
X6139 a_10660_37762# cap_shunt_n a_10452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X6140 a_20740_43672# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6141 a_20532_43188# cap_shunt_n a_20740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X6142 a_16708_48738# cap_shunt_p a_16500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6143 vdd a_9644_46280# a_9556_46324# vdd pmos_6p0 w=1.22u l=1u
X6144 vdd a_5612_27031# a_5524_27128# vdd pmos_6p0 w=1.22u l=1u
X6145 vss cap_shunt_p a_31024_25156# vss nmos_6p0 w=0.82u l=0.6u
X6146 a_7748_37762# cap_shunt_n a_8680_37700# vss nmos_6p0 w=0.82u l=0.6u
X6147 a_11668_42104# cap_shunt_n a_11460_41620# vdd pmos_6p0 w=1.2u l=0.5u
X6148 a_2500_27132# cap_shunt_p a_2708_26786# vdd pmos_6p0 w=1.2u l=0.5u
X6149 a_2500_47516# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6150 a_24452_11452# cap_series_gyp a_24660_11106# vdd pmos_6p0 w=1.2u l=0.5u
X6151 a_10660_42466# cap_shunt_n a_10452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X6152 vdd a_14908_6647# a_14820_6744# vdd pmos_6p0 w=1.22u l=1u
X6153 a_28692_13880# cap_series_gyp a_28484_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6154 a_20740_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6155 vdd a_10540_40008# a_10452_40052# vdd pmos_6p0 w=1.22u l=1u
X6156 a_27788_54120# a_27700_54164# vss vss nmos_6p0 w=0.82u l=1u
X6157 a_7540_42812# cap_shunt_n a_7748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X6158 a_22436_10260# cap_series_gyp a_22644_10744# vdd pmos_6p0 w=1.2u l=0.5u
X6159 a_9668_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6160 vdd a_6060_5079# a_5972_5176# vdd pmos_6p0 w=1.22u l=1u
X6161 a_29196_3612# cap_series_gyn a_29384_3612# vdd pmos_6p0 w=1.2u l=0.5u
X6162 vdd tune_series_gy[5] a_19524_8692# vdd pmos_6p0 w=1.2u l=0.5u
X6163 a_23464_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6164 a_24660_42466# cap_shunt_n a_24452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X6165 a_17828_35832# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6166 a_7768_6748# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X6167 a_6292_51874# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6168 a_2500_30268# cap_shunt_n a_2708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X6169 a_21672_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6170 a_9644_38440# a_9556_38484# vss vss nmos_6p0 w=0.82u l=1u
X6171 a_17620_16532# cap_shunt_p a_17828_17016# vdd pmos_6p0 w=1.2u l=0.5u
X6172 a_23464_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6173 vdd a_32604_33736# a_32516_33780# vdd pmos_6p0 w=1.22u l=1u
X6174 a_16500_28700# cap_shunt_n a_16708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X6175 a_24452_20860# cap_shunt_p a_24660_20514# vdd pmos_6p0 w=1.2u l=0.5u
X6176 a_17828_43672# cap_shunt_p a_17620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X6177 a_24660_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6178 a_13796_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6179 a_22644_12312# cap_series_gyn a_23576_12312# vss nmos_6p0 w=0.82u l=0.6u
X6180 vss cap_shunt_p a_4032_48676# vss nmos_6p0 w=0.82u l=0.6u
X6181 a_13252_29076# cap_shunt_n a_13460_29560# vdd pmos_6p0 w=1.2u l=0.5u
X6182 a_25100_55255# a_25012_55352# vss vss nmos_6p0 w=0.82u l=1u
X6183 a_6084_49460# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6184 vdd a_32604_30600# a_32516_30644# vdd pmos_6p0 w=1.22u l=1u
X6185 vss tune_shunt[7] a_20740_27992# vss nmos_6p0 w=0.51u l=0.6u
X6186 vdd tune_series_gy[5] a_22436_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6187 vss cap_series_gygyp a_34952_7908# vss nmos_6p0 w=0.82u l=0.6u
X6188 a_35880_10260# cap_series_gygyp a_35692_10260# vdd pmos_6p0 w=1.2u l=0.5u
X6189 vss cap_series_gyp a_30800_13880# vss nmos_6p0 w=0.82u l=0.6u
X6190 a_3380_18584# cap_shunt_p a_4312_18584# vss nmos_6p0 w=0.82u l=0.6u
X6191 vdd a_20284_52552# a_20196_52596# vdd pmos_6p0 w=1.22u l=1u
X6192 vss tune_shunt[6] a_3828_35832# vss nmos_6p0 w=0.51u l=0.6u
X6193 vdd tune_shunt[7] a_9332_13020# vdd pmos_6p0 w=1.2u l=0.5u
X6194 a_37868_55688# a_37780_55732# vss vss nmos_6p0 w=0.82u l=1u
X6195 a_5636_3612# cap_shunt_n a_5844_3266# vdd pmos_6p0 w=1.2u l=0.5u
X6196 a_6532_19668# cap_shunt_p a_6740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X6197 a_31424_21720# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X6198 vdd a_36524_38007# a_36436_38104# vdd pmos_6p0 w=1.22u l=1u
X6199 a_8512_22020# cap_shunt_p a_6404_22082# vss nmos_6p0 w=0.82u l=0.6u
X6200 vdd tune_shunt[7] a_9668_16532# vdd pmos_6p0 w=1.2u l=0.5u
X6201 a_35692_3988# cap_series_gygyp a_35880_3988# vdd pmos_6p0 w=1.2u l=0.5u
X6202 a_13460_32696# cap_shunt_n a_14392_32696# vss nmos_6p0 w=0.82u l=0.6u
X6203 vss tune_shunt[5] a_20740_24856# vss nmos_6p0 w=0.51u l=0.6u
X6204 a_11592_13880# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6205 a_13796_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6206 a_24360_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6207 vss cap_series_gyp a_30800_10744# vss nmos_6p0 w=0.82u l=0.6u
X6208 a_2708_11106# cap_shunt_n a_2500_11452# vdd pmos_6p0 w=1.2u l=0.5u
X6209 a_24660_26786# cap_shunt_p a_24452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X6210 a_21524_3266# cap_series_gyp a_22456_3204# vss nmos_6p0 w=0.82u l=0.6u
X6211 vdd a_32156_25896# a_32068_25940# vdd pmos_6p0 w=1.22u l=1u
X6212 a_4492_6647# a_4404_6744# vss vss nmos_6p0 w=0.82u l=1u
X6213 a_12788_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6214 vdd tune_shunt[6] a_2500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X6215 a_32612_25218# cap_shunt_p a_32404_25564# vdd pmos_6p0 w=1.2u l=0.5u
X6216 vss tune_series_gy[4] a_15700_6402# vss nmos_6p0 w=0.51u l=0.6u
X6217 a_11668_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6218 vdd tune_shunt[7] a_24452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X6219 a_16500_30268# cap_shunt_n a_16708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X6220 vdd a_6508_23895# a_6420_23992# vdd pmos_6p0 w=1.22u l=1u
X6221 a_2708_48738# cap_shunt_p a_2500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6222 vdd tune_shunt[7] a_28484_25940# vdd pmos_6p0 w=1.2u l=0.5u
X6223 a_11592_10744# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6224 a_3620_36916# cap_shunt_n a_3828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X6225 a_31808_32996# cap_shunt_p a_29700_33058# vss nmos_6p0 w=0.82u l=0.6u
X6226 vdd a_32156_22760# a_32068_22804# vdd pmos_6p0 w=1.22u l=1u
X6227 a_4492_3511# a_4404_3608# vss vss nmos_6p0 w=0.82u l=1u
X6228 vdd a_30364_6647# a_30276_6744# vdd pmos_6p0 w=1.22u l=1u
X6229 vss cap_shunt_p a_8064_21720# vss nmos_6p0 w=0.82u l=0.6u
X6230 a_11668_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6231 vdd tune_shunt[6] a_25572_32212# vdd pmos_6p0 w=1.2u l=0.5u
X6232 a_9316_48738# cap_shunt_p a_9108_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6233 a_10660_36194# cap_shunt_n a_10452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X6234 a_24452_9884# cap_series_gyn a_24660_9538# vdd pmos_6p0 w=1.2u l=0.5u
X6235 a_20740_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6236 vdd tune_shunt[4] a_28484_22804# vdd pmos_6p0 w=1.2u l=0.5u
X6237 vdd tune_shunt[6] a_13588_42812# vdd pmos_6p0 w=1.2u l=0.5u
X6238 a_3828_35832# cap_shunt_n a_4760_35832# vss nmos_6p0 w=0.82u l=0.6u
X6239 a_27788_47848# a_27700_47892# vss vss nmos_6p0 w=0.82u l=1u
X6240 a_32612_28354# cap_shunt_p a_32404_28700# vdd pmos_6p0 w=1.2u l=0.5u
X6241 a_14468_3266# cap_series_gyn a_16184_3204# vss nmos_6p0 w=0.82u l=0.6u
X6242 a_8624_20452# cap_shunt_p a_6516_20514# vss nmos_6p0 w=0.82u l=0.6u
X6243 a_10640_50244# cap_shunt_p a_9316_50306# vss nmos_6p0 w=0.82u l=0.6u
X6244 a_7540_36540# cap_shunt_n a_7748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X6245 a_2500_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6246 a_35840_34264# cap_shunt_n a_33732_34264# vss nmos_6p0 w=0.82u l=0.6u
X6247 a_34396_5512# a_34308_5556# vss vss nmos_6p0 w=0.82u l=1u
X6248 a_3828_15448# cap_shunt_p a_3620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X6249 a_10660_33058# cap_shunt_n a_10452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X6250 a_17828_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6251 a_24452_6748# cap_series_gyn a_24660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X6252 a_2708_50306# cap_shunt_n a_2500_50652# vdd pmos_6p0 w=1.2u l=0.5u
X6253 a_24660_36194# cap_shunt_p a_24452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X6254 a_20740_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6255 vdd tune_series_gy[5] a_19524_10260# vdd pmos_6p0 w=1.2u l=0.5u
X6256 a_6644_53788# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6257 a_2708_9538# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X6258 a_7540_33404# cap_shunt_n a_7748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X6259 a_8008_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6260 a_31904_45540# cap_shunt_gyp a_31904_45944# vdd pmos_6p0 w=1.215u l=0.5u
X6261 a_35840_31128# cap_shunt_n a_33732_31128# vss nmos_6p0 w=0.82u l=0.6u
X6262 a_13588_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6263 a_14260_3612# cap_series_gyn a_14468_3266# vdd pmos_6p0 w=1.2u l=0.5u
X6264 a_17828_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6265 a_35264_45944# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X6266 a_23464_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6267 a_24660_33058# cap_shunt_p a_24452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X6268 vss cap_series_gyn a_16016_6040# vss nmos_6p0 w=0.82u l=0.6u
X6269 vdd a_33500_52552# a_33412_52596# vdd pmos_6p0 w=1.22u l=1u
X6270 vdd tune_shunt[6] a_2500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X6271 a_31808_4772# cap_shunt_p a_29700_4834# vss nmos_6p0 w=0.82u l=0.6u
X6272 a_1692_55688# a_1604_55732# vss vss nmos_6p0 w=0.82u l=1u
X6273 vdd a_29916_47415# a_29828_47512# vdd pmos_6p0 w=1.22u l=1u
X6274 a_1924_4472# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X6275 a_32612_34626# cap_shunt_n a_33544_34564# vss nmos_6p0 w=0.82u l=0.6u
X6276 vdd a_24092_3511# a_24004_3608# vdd pmos_6p0 w=1.22u l=1u
X6277 a_7580_6748# cap_series_gyp a_7768_6748# vdd pmos_6p0 w=1.2u l=0.5u
X6278 vss cap_series_gyn a_19936_12612# vss nmos_6p0 w=0.82u l=0.6u
X6279 a_20532_18100# cap_shunt_p a_20740_18584# vdd pmos_6p0 w=1.2u l=0.5u
X6280 a_16708_48738# cap_shunt_p a_16500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6281 a_34396_53687# a_34308_53784# vss vss nmos_6p0 w=0.82u l=1u
X6282 a_35264_42808# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X6283 vdd a_32604_24328# a_32516_24372# vdd pmos_6p0 w=1.22u l=1u
X6284 a_10864_14180# cap_shunt_p a_9540_14242# vss nmos_6p0 w=0.82u l=0.6u
X6285 a_25100_48983# a_25012_49080# vss vss nmos_6p0 w=0.82u l=1u
X6286 a_17828_46808# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6287 a_11668_42104# cap_shunt_n a_11460_41620# vdd pmos_6p0 w=1.2u l=0.5u
X6288 a_29700_23650# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X6289 a_6572_3988# cap_series_gyp a_6760_3988# vdd pmos_6p0 w=1.2u l=0.5u
X6290 a_24452_11452# cap_series_gyp a_24660_11106# vdd pmos_6p0 w=1.2u l=0.5u
X6291 a_10660_42466# cap_shunt_n a_10452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X6292 vdd a_31484_43144# a_31396_43188# vdd pmos_6p0 w=1.22u l=1u
X6293 a_32612_31490# cap_shunt_n a_33544_31428# vss nmos_6p0 w=0.82u l=0.6u
X6294 vdd a_27676_30167# a_27588_30264# vdd pmos_6p0 w=1.22u l=1u
X6295 vss tune_shunt[7] a_3828_29560# vss nmos_6p0 w=0.51u l=0.6u
X6296 a_24660_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6297 vdd tune_shunt[5] a_12580_19668# vdd pmos_6p0 w=1.2u l=0.5u
X6298 vss cap_shunt_n a_4032_39268# vss nmos_6p0 w=0.82u l=0.6u
X6299 a_24452_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6300 a_25780_9176# cap_series_gyp a_26712_9176# vss nmos_6p0 w=0.82u l=0.6u
X6301 a_21964_52119# a_21876_52216# vss vss nmos_6p0 w=0.82u l=1u
X6302 vdd tune_series_gygy[5] a_34308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X6303 a_34396_50551# a_34308_50648# vss vss nmos_6p0 w=0.82u l=1u
X6304 a_7540_42812# cap_shunt_n a_7748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X6305 a_2140_21192# a_2052_21236# vss vss nmos_6p0 w=0.82u l=1u
X6306 a_10864_11044# cap_shunt_p a_9540_11106# vss nmos_6p0 w=0.82u l=0.6u
X6307 a_21748_12674# cap_series_gyn a_23464_12612# vss nmos_6p0 w=0.82u l=0.6u
X6308 vss tune_shunt[7] a_20740_18584# vss nmos_6p0 w=0.51u l=0.6u
X6309 a_22436_10260# cap_series_gyp a_22644_10744# vdd pmos_6p0 w=1.2u l=0.5u
X6310 a_5844_11106# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X6311 a_17828_15448# cap_shunt_p a_17620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X6312 vss tune_shunt[7] a_3828_26424# vss nmos_6p0 w=0.51u l=0.6u
X6313 a_1716_5180# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6314 vss cap_shunt_n a_25984_29860# vss nmos_6p0 w=0.82u l=0.6u
X6315 a_1924_7970# cap_shunt_n a_1716_8316# vdd pmos_6p0 w=1.2u l=0.5u
X6316 vdd a_30028_47848# a_29940_47892# vdd pmos_6p0 w=1.22u l=1u
X6317 a_34328_29860# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6318 vss cap_series_gyp a_16920_11044# vss nmos_6p0 w=0.82u l=0.6u
X6319 a_13460_23288# cap_shunt_n a_14392_23288# vss nmos_6p0 w=0.82u l=0.6u
X6320 vss tune_series_gy[5] a_20740_15448# vss nmos_6p0 w=0.51u l=0.6u
X6321 a_6760_3988# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X6322 vdd a_33612_9783# a_33524_9880# vdd pmos_6p0 w=1.22u l=1u
X6323 vdd a_32156_16488# a_32068_16532# vdd pmos_6p0 w=1.22u l=1u
X6324 vss cap_shunt_p a_25984_26724# vss nmos_6p0 w=0.82u l=0.6u
X6325 vss cap_shunt_n a_8848_53080# vss nmos_6p0 w=0.82u l=0.6u
X6326 a_11460_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6327 vdd a_30028_44712# a_29940_44756# vdd pmos_6p0 w=1.22u l=1u
X6328 a_34328_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6329 vdd tune_series_gy[5] a_24452_14588# vdd pmos_6p0 w=1.2u l=0.5u
X6330 vss tune_shunt[6] a_3828_46808# vss nmos_6p0 w=0.51u l=0.6u
X6331 vss cap_series_gyp a_23072_9476# vss nmos_6p0 w=0.82u l=0.6u
X6332 vss cap_shunt_gyp a_36652_47108# vss nmos_6p0 w=0.82u l=0.6u
X6333 a_10452_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6334 vdd tune_series_gy[4] a_28484_16532# vdd pmos_6p0 w=1.2u l=0.5u
X6335 a_3828_29560# cap_shunt_n a_4760_29560# vss nmos_6p0 w=0.82u l=0.6u
X6336 vdd tune_shunt[7] a_13588_36540# vdd pmos_6p0 w=1.2u l=0.5u
X6337 a_3620_27508# cap_shunt_n a_3828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X6338 a_31808_23588# cap_shunt_p a_29700_23650# vss nmos_6p0 w=0.82u l=0.6u
X6339 a_21540_8316# cap_series_gyp a_21748_7970# vdd pmos_6p0 w=1.2u l=0.5u
X6340 a_8400_49944# cap_shunt_p a_6292_49944# vss nmos_6p0 w=0.82u l=0.6u
X6341 a_34144_47512# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X6342 a_34480_46870# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6343 a_9332_13020# cap_shunt_p a_9540_12674# vdd pmos_6p0 w=1.2u l=0.5u
X6344 vdd tune_shunt_gy[2] a_36324_41621# vdd pmos_6p0 w=1.215u l=0.5u
X6345 vss cap_shunt_n a_12656_38968# vss nmos_6p0 w=0.82u l=0.6u
X6346 a_6084_49460# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6347 a_31260_7080# a_31172_7124# vss vss nmos_6p0 w=0.82u l=1u
X6348 a_6572_5556# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6349 a_2932_10744# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X6350 vss cap_shunt_p a_8064_12312# vss nmos_6p0 w=0.82u l=0.6u
X6351 vdd tune_series_gy[5] a_22436_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6352 vss tune_shunt[7] a_13460_35832# vss nmos_6p0 w=0.51u l=0.6u
X6353 a_29492_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6354 a_10660_26786# cap_shunt_n a_10452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X6355 a_2708_44034# cap_shunt_p a_2500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X6356 a_37196_30600# a_37108_30644# vss vss nmos_6p0 w=0.82u l=1u
X6357 vss cap_series_gyn a_20832_6040# vss nmos_6p0 w=0.82u l=0.6u
X6358 a_27496_20152# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6359 a_21540_45948# cap_shunt_p a_21748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X6360 a_3828_26424# cap_shunt_p a_4760_26424# vss nmos_6p0 w=0.82u l=0.6u
X6361 vdd tune_shunt[7] a_13588_33404# vdd pmos_6p0 w=1.2u l=0.5u
X6362 a_21540_5180# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6363 a_6532_19668# cap_shunt_p a_6740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X6364 a_10660_4834# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X6365 a_30800_12312# cap_series_gyn a_28692_12312# vss nmos_6p0 w=0.82u l=0.6u
X6366 a_35448_18884# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X6367 vss tune_shunt[7] a_25780_27992# vss nmos_6p0 w=0.51u l=0.6u
X6368 a_7540_27132# cap_shunt_n a_7748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X6369 vdd tune_series_gy[5] a_24452_17724# vdd pmos_6p0 w=1.2u l=0.5u
X6370 a_15904_43972# cap_shunt_n a_13796_44034# vss nmos_6p0 w=0.82u l=0.6u
X6371 a_2708_40898# cap_shunt_p a_2500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X6372 a_24660_26786# cap_shunt_p a_24452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X6373 a_7540_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6374 vss tune_shunt[6] a_13796_40898# vss nmos_6p0 w=0.51u l=0.6u
X6375 vdd tune_shunt[6] a_2500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X6376 vdd tune_shunt_gy[0] a_37444_33781# vdd pmos_6p0 w=1.215u l=0.5u
X6377 a_34536_6748# cap_series_gygyp a_35344_6340# vss nmos_6p0 w=0.82u l=0.6u
X6378 a_5636_8692# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6379 a_35448_15748# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X6380 a_32612_28354# cap_shunt_p a_33544_28292# vss nmos_6p0 w=0.82u l=0.6u
X6381 vss tune_shunt[7] a_25780_24856# vss nmos_6p0 w=0.51u l=0.6u
X6382 vdd tune_shunt[7] a_28484_25940# vdd pmos_6p0 w=1.2u l=0.5u
X6383 a_15904_40836# cap_shunt_n a_13796_40898# vss nmos_6p0 w=0.82u l=0.6u
X6384 vdd a_28124_33303# a_28036_33400# vdd pmos_6p0 w=1.22u l=1u
X6385 a_9540_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6386 a_17828_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6387 a_2708_9538# cap_shunt_n a_2500_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6388 a_34844_36872# a_34756_36916# vss vss nmos_6p0 w=0.82u l=1u
X6389 vdd a_10092_3944# a_10004_3988# vdd pmos_6p0 w=1.22u l=1u
X6390 vss cap_series_gygyp a_37080_20152# vss nmos_6p0 w=0.82u l=0.6u
X6391 a_4760_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6392 a_25780_32696# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6393 a_4256_10744# cap_shunt_n a_2932_10744# vss nmos_6p0 w=0.82u l=0.6u
X6394 a_9316_48738# cap_shunt_p a_9108_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6395 a_10660_36194# cap_shunt_n a_10452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X6396 a_32612_25218# cap_shunt_p a_33544_25156# vss nmos_6p0 w=0.82u l=0.6u
X6397 a_12580_49460# cap_shunt_n a_12788_49944# vdd pmos_6p0 w=1.2u l=0.5u
X6398 vdd tune_shunt[4] a_28484_22804# vdd pmos_6p0 w=1.2u l=0.5u
X6399 vdd a_37980_54120# a_37892_54164# vdd pmos_6p0 w=1.22u l=1u
X6400 a_7540_36540# cap_shunt_n a_7748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X6401 a_29916_19191# a_29828_19288# vss vss nmos_6p0 w=0.82u l=1u
X6402 a_29700_14242# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6403 a_14012_53687# a_13924_53784# vss vss nmos_6p0 w=0.82u l=1u
X6404 a_10660_33058# cap_shunt_n a_10452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X6405 a_2708_50306# cap_shunt_n a_2500_50652# vdd pmos_6p0 w=1.2u l=0.5u
X6406 a_25572_40052# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6407 a_35880_8692# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X6408 a_29532_9884# cap_series_gyn a_29720_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6409 a_10452_44380# cap_shunt_n a_10660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X6410 vdd a_37980_50984# a_37892_51028# vdd pmos_6p0 w=1.22u l=1u
X6411 a_7540_33404# cap_shunt_n a_7748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X6412 a_13588_50652# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6413 a_24660_9538# cap_series_gyn a_25592_9476# vss nmos_6p0 w=0.82u l=0.6u
X6414 a_2932_10744# cap_shunt_n a_2724_10260# vdd pmos_6p0 w=1.2u l=0.5u
X6415 a_2140_11784# a_2052_11828# vss vss nmos_6p0 w=0.82u l=1u
X6416 vdd tune_shunt[6] a_20532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X6417 a_32404_36540# cap_shunt_n a_32612_36194# vdd pmos_6p0 w=1.2u l=0.5u
X6418 vss cap_shunt_n a_22064_27992# vss nmos_6p0 w=0.82u l=0.6u
X6419 a_29700_11106# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X6420 a_14372_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6421 a_21840_7608# cap_series_gyp a_19732_7608# vss nmos_6p0 w=0.82u l=0.6u
X6422 vss tune_shunt[7] a_3380_17016# vss nmos_6p0 w=0.51u l=0.6u
X6423 a_25780_37400# cap_shunt_p a_27496_37400# vss nmos_6p0 w=0.82u l=0.6u
X6424 a_10452_41244# cap_shunt_n a_10660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X6425 a_10452_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6426 a_25984_42404# cap_shunt_n a_24660_42466# vss nmos_6p0 w=0.82u l=0.6u
X6427 a_32404_33404# cap_shunt_n a_32612_33058# vdd pmos_6p0 w=1.2u l=0.5u
X6428 vss cap_shunt_n a_22064_24856# vss nmos_6p0 w=0.82u l=0.6u
X6429 a_14460_9783# a_14372_9880# vss vss nmos_6p0 w=0.82u l=1u
X6430 a_20532_18100# cap_shunt_p a_20740_18584# vdd pmos_6p0 w=1.2u l=0.5u
X6431 a_34516_18946# cap_series_gygyn a_36232_18884# vss nmos_6p0 w=0.82u l=0.6u
X6432 a_31248_44757# cap_shunt_gyn a_31268_45240# vss nmos_6p0 w=0.82u l=0.6u
X6433 a_32632_14588# cap_series_gyp a_32444_14588# vdd pmos_6p0 w=1.2u l=0.5u
X6434 vdd tune_series_gygy[4] a_35692_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6435 vss cap_series_gyp a_25984_17316# vss nmos_6p0 w=0.82u l=0.6u
X6436 a_10540_7080# a_10452_7124# vss vss nmos_6p0 w=0.82u l=1u
X6437 vss tune_series_gygy[0] a_35880_3988# vss nmos_6p0 w=0.51u l=0.6u
X6438 a_20532_14964# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6439 vss tune_shunt[7] a_13460_29560# vss nmos_6p0 w=0.51u l=0.6u
X6440 vdd a_15580_50984# a_15492_51028# vdd pmos_6p0 w=1.22u l=1u
X6441 a_21540_39676# cap_shunt_p a_21748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X6442 a_23856_6340# cap_series_gyn a_21748_6402# vss nmos_6p0 w=0.82u l=0.6u
X6443 a_35292_13352# a_35204_13396# vss vss nmos_6p0 w=0.82u l=1u
X6444 a_26712_35832# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6445 vdd tune_shunt[7] a_13588_27132# vdd pmos_6p0 w=1.2u l=0.5u
X6446 vdd a_18492_11784# a_18404_11828# vdd pmos_6p0 w=1.22u l=1u
X6447 a_34516_15810# cap_series_gygyn a_36232_15748# vss nmos_6p0 w=0.82u l=0.6u
X6448 a_33524_33780# cap_shunt_n a_33732_34264# vdd pmos_6p0 w=1.2u l=0.5u
X6449 a_21180_52552# a_21092_52596# vss vss nmos_6p0 w=0.82u l=1u
X6450 vss tune_shunt[7] a_13460_26424# vss nmos_6p0 w=0.51u l=0.6u
X6451 vss cap_shunt_p a_14896_12312# vss nmos_6p0 w=0.82u l=0.6u
X6452 a_11436_54120# a_11348_54164# vss vss nmos_6p0 w=0.82u l=1u
X6453 a_6740_37400# cap_shunt_n a_6532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X6454 a_35292_10216# a_35204_10260# vss vss nmos_6p0 w=0.82u l=1u
X6455 vdd a_2140_53687# a_2052_53784# vdd pmos_6p0 w=1.22u l=1u
X6456 a_18424_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6457 vss cap_shunt_p a_7952_12612# vss nmos_6p0 w=0.82u l=0.6u
X6458 a_27788_53687# a_27700_53784# vss vss nmos_6p0 w=0.82u l=1u
X6459 a_5152_32696# cap_shunt_p a_3828_32696# vss nmos_6p0 w=0.82u l=0.6u
X6460 a_14112_13880# cap_shunt_p a_12788_13880# vss nmos_6p0 w=0.82u l=0.6u
X6461 a_33524_30644# cap_shunt_n a_33732_31128# vdd pmos_6p0 w=1.2u l=0.5u
X6462 vss tune_series_gy[4] a_25780_18584# vss nmos_6p0 w=0.51u l=0.6u
X6463 vss tune_shunt[6] a_13796_45602# vss nmos_6p0 w=0.51u l=0.6u
X6464 a_5488_51512# cap_shunt_n a_3380_51512# vss nmos_6p0 w=0.82u l=0.6u
X6465 vdd a_26444_47848# a_26356_47892# vdd pmos_6p0 w=1.22u l=1u
X6466 a_27676_39575# a_27588_39672# vss vss nmos_6p0 w=0.82u l=1u
X6467 a_15904_34564# cap_shunt_n a_13796_34626# vss nmos_6p0 w=0.82u l=0.6u
X6468 a_12216_7608# cap_series_gyp a_11800_7124# vss nmos_6p0 w=0.82u l=0.6u
X6469 a_15700_6402# cap_series_gyp a_17416_6340# vss nmos_6p0 w=0.82u l=0.6u
X6470 a_2588_43144# a_2500_43188# vss vss nmos_6p0 w=0.82u l=1u
X6471 a_35740_55688# a_35652_55732# vss vss nmos_6p0 w=0.82u l=1u
X6472 vdd a_2140_50551# a_2052_50648# vdd pmos_6p0 w=1.22u l=1u
X6473 vss cap_shunt_p a_35840_27992# vss nmos_6p0 w=0.82u l=0.6u
X6474 a_27788_50551# a_27700_50648# vss vss nmos_6p0 w=0.82u l=1u
X6475 a_30632_34564# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6476 vss tune_series_gy[5] a_25780_15448# vss nmos_6p0 w=0.51u l=0.6u
X6477 a_18044_3944# a_17956_3988# vss vss nmos_6p0 w=0.82u l=1u
X6478 a_3828_21720# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6479 a_35692_14964# cap_series_gygyn a_35880_14964# vdd pmos_6p0 w=1.2u l=0.5u
X6480 vdd tune_series_gy[4] a_28484_16532# vdd pmos_6p0 w=1.2u l=0.5u
X6481 vdd a_26444_44712# a_26356_44756# vdd pmos_6p0 w=1.22u l=1u
X6482 a_15904_31428# cap_shunt_n a_13796_31490# vss nmos_6p0 w=0.82u l=0.6u
X6483 a_2588_40008# a_2500_40052# vss vss nmos_6p0 w=0.82u l=1u
X6484 vdd a_1692_14920# a_1604_14964# vdd pmos_6p0 w=1.22u l=1u
X6485 a_3172_49460# cap_shunt_p a_3380_49944# vdd pmos_6p0 w=1.2u l=0.5u
X6486 a_30632_31428# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6487 a_14692_9176# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X6488 a_10660_26786# cap_shunt_n a_10452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X6489 a_25780_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6490 a_2708_44034# cap_shunt_p a_2500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X6491 vss tune_shunt[5] a_2708_48738# vss nmos_6p0 w=0.51u l=0.6u
X6492 a_21540_45948# cap_shunt_p a_21748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X6493 vdd a_31932_41576# a_31844_41620# vdd pmos_6p0 w=1.22u l=1u
X6494 a_35692_11828# cap_series_gygyp a_35880_11828# vdd pmos_6p0 w=1.2u l=0.5u
X6495 vdd a_18940_13352# a_18852_13396# vdd pmos_6p0 w=1.22u l=1u
X6496 a_7540_27132# cap_shunt_n a_7748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X6497 vdd a_1692_11784# a_1604_11828# vdd pmos_6p0 w=1.22u l=1u
X6498 a_13588_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6499 a_2708_40898# cap_shunt_p a_2500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X6500 vdd tune_series_gy[1] a_6572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X6501 a_22064_43672# cap_shunt_n a_20740_43672# vss nmos_6p0 w=0.82u l=0.6u
X6502 a_21748_23650# cap_shunt_p a_21540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X6503 a_13588_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6504 a_25984_36132# cap_shunt_p a_24660_36194# vss nmos_6p0 w=0.82u l=0.6u
X6505 a_25780_26424# cap_shunt_p a_25572_25940# vdd pmos_6p0 w=1.2u l=0.5u
X6506 vdd tune_shunt[7] a_20532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X6507 a_32404_27132# cap_shunt_p a_32612_26786# vdd pmos_6p0 w=1.2u l=0.5u
X6508 vss cap_shunt_p a_22064_18584# vss nmos_6p0 w=0.82u l=0.6u
X6509 vdd a_32604_41143# a_32516_41240# vdd pmos_6p0 w=1.22u l=1u
X6510 a_14392_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6511 a_20440_6040# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X6512 a_18388_3266# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X6513 a_8848_13880# cap_shunt_p a_6740_13880# vss nmos_6p0 w=0.82u l=0.6u
X6514 a_3828_48376# cap_shunt_p a_3620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X6515 a_19276_44279# a_19188_44376# vss vss nmos_6p0 w=0.82u l=1u
X6516 a_22064_40536# cap_shunt_p a_20740_40536# vss nmos_6p0 w=0.82u l=0.6u
X6517 a_22636_47848# a_22548_47892# vss vss nmos_6p0 w=0.82u l=1u
X6518 a_20720_7908# cap_series_gyp a_18612_7970# vss nmos_6p0 w=0.82u l=0.6u
X6519 a_26712_29560# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6520 a_25780_23288# cap_shunt_p a_25572_22804# vdd pmos_6p0 w=1.2u l=0.5u
X6521 a_5040_9176# cap_shunt_n a_2932_9176# vss nmos_6p0 w=0.82u l=0.6u
X6522 vss cap_series_gyn a_22064_15448# vss nmos_6p0 w=0.82u l=0.6u
X6523 a_19524_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6524 vdd tune_shunt[5] a_6084_51028# vdd pmos_6p0 w=1.2u l=0.5u
X6525 vss cap_shunt_n a_23856_43972# vss nmos_6p0 w=0.82u l=0.6u
X6526 vdd a_35180_33303# a_35092_33400# vdd pmos_6p0 w=1.22u l=1u
X6527 a_4380_52119# a_4292_52216# vss vss nmos_6p0 w=0.82u l=1u
X6528 a_3828_45240# cap_shunt_p a_3620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X6529 a_19276_41143# a_19188_41240# vss vss nmos_6p0 w=0.82u l=1u
X6530 vss cap_shunt_p a_5152_46808# vss nmos_6p0 w=0.82u l=0.6u
X6531 a_16500_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6532 a_26712_26424# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6533 a_16708_44034# cap_shunt_p a_16500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X6534 a_22644_7608# cap_series_gyp a_24360_7608# vss nmos_6p0 w=0.82u l=0.6u
X6535 vss cap_series_gyn a_19936_6340# vss nmos_6p0 w=0.82u l=0.6u
X6536 a_18404_5180# cap_series_gyp a_18612_4834# vdd pmos_6p0 w=1.2u l=0.5u
X6537 a_10452_44380# cap_shunt_n a_10660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X6538 a_3620_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6539 vss cap_shunt_p a_23856_40836# vss nmos_6p0 w=0.82u l=0.6u
X6540 vss tune_shunt[7] a_13796_39330# vss nmos_6p0 w=0.51u l=0.6u
X6541 a_32404_36540# cap_shunt_n a_32612_36194# vdd pmos_6p0 w=1.2u l=0.5u
X6542 a_15904_28292# cap_shunt_n a_13796_28354# vss nmos_6p0 w=0.82u l=0.6u
X6543 a_24204_46280# a_24116_46324# vss vss nmos_6p0 w=0.82u l=1u
X6544 a_24452_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6545 a_6740_27992# cap_shunt_n a_6532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X6546 vdd a_16252_18056# a_16164_18100# vdd pmos_6p0 w=1.22u l=1u
X6547 a_16700_18056# a_16612_18100# vss vss nmos_6p0 w=0.82u l=1u
X6548 a_11460_40052# cap_shunt_n a_11668_40536# vdd pmos_6p0 w=1.2u l=0.5u
X6549 a_8400_51812# cap_shunt_p a_6292_51874# vss nmos_6p0 w=0.82u l=0.6u
X6550 vdd a_2140_44279# a_2052_44376# vdd pmos_6p0 w=1.22u l=1u
X6551 a_16708_40898# cap_shunt_n a_16500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X6552 a_30632_28292# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6553 vdd a_6956_23895# a_6868_23992# vdd pmos_6p0 w=1.22u l=1u
X6554 a_20104_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X6555 a_2708_50306# cap_shunt_n a_3640_50244# vss nmos_6p0 w=0.82u l=0.6u
X6556 a_10452_41244# cap_shunt_n a_10660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X6557 vdd tune_shunt[7] a_32404_28700# vdd pmos_6p0 w=1.2u l=0.5u
X6558 a_5152_23288# cap_shunt_p a_3828_23288# vss nmos_6p0 w=0.82u l=0.6u
X6559 a_11800_8692# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X6560 a_18604_50551# a_18516_50648# vss vss nmos_6p0 w=0.82u l=1u
X6561 vdd a_37644_35304# a_37556_35348# vdd pmos_6p0 w=1.22u l=1u
X6562 a_32404_33404# cap_shunt_n a_32612_33058# vdd pmos_6p0 w=1.2u l=0.5u
X6563 a_15904_25156# cap_shunt_n a_13796_25218# vss nmos_6p0 w=0.82u l=0.6u
X6564 a_20532_18100# cap_shunt_p a_20740_18584# vdd pmos_6p0 w=1.2u l=0.5u
X6565 a_24452_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6566 a_25444_3266# cap_shunt_p a_25236_3612# vdd pmos_6p0 w=1.2u l=0.5u
X6567 a_19524_8692# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6568 a_32632_14588# cap_series_gyp a_32444_14588# vdd pmos_6p0 w=1.2u l=0.5u
X6569 a_6740_43672# cap_shunt_p a_8456_43672# vss nmos_6p0 w=0.82u l=0.6u
X6570 a_2588_33736# a_2500_33780# vss vss nmos_6p0 w=0.82u l=1u
X6571 vdd tune_series_gygy[4] a_35692_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6572 a_16700_14920# a_16612_14964# vss vss nmos_6p0 w=0.82u l=1u
X6573 a_30632_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6574 a_28692_9176# cap_series_gyn a_30408_9176# vss nmos_6p0 w=0.82u l=0.6u
X6575 a_10660_4834# cap_series_gyp a_10452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X6576 vss cap_series_gygyp a_36296_26424# vss nmos_6p0 w=0.82u l=0.6u
X6577 a_9876_20152# cap_shunt_p a_9668_19668# vdd pmos_6p0 w=1.2u l=0.5u
X6578 a_17828_48376# cap_shunt_p a_17620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X6579 a_21540_39676# cap_shunt_p a_21748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X6580 vdd a_28572_9783# a_28484_9880# vdd pmos_6p0 w=1.22u l=1u
X6581 vdd a_34844_3511# a_34756_3608# vdd pmos_6p0 w=1.22u l=1u
X6582 a_25780_4472# cap_shunt_p a_25572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X6583 a_24660_12674# cap_series_gyn a_24452_13020# vdd pmos_6p0 w=1.2u l=0.5u
X6584 a_6740_40536# cap_shunt_n a_8456_40536# vss nmos_6p0 w=0.82u l=0.6u
X6585 a_3828_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6586 a_33524_33780# cap_shunt_n a_33732_34264# vdd pmos_6p0 w=1.2u l=0.5u
X6587 a_2588_30600# a_2500_30644# vss vss nmos_6p0 w=0.82u l=1u
X6588 a_14260_3612# cap_series_gyn a_14468_3266# vdd pmos_6p0 w=1.2u l=0.5u
X6589 a_20172_22327# a_20084_22424# vss vss nmos_6p0 w=0.82u l=1u
X6590 a_6740_37400# cap_shunt_n a_6532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X6591 a_21540_9884# cap_series_gyp a_21748_9538# vdd pmos_6p0 w=1.2u l=0.5u
X6592 a_17828_45240# cap_shunt_p a_17620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X6593 vdd a_28572_6647# a_28484_6744# vdd pmos_6p0 w=1.22u l=1u
X6594 a_6532_47892# cap_shunt_p a_6740_48376# vdd pmos_6p0 w=1.2u l=0.5u
X6595 a_22960_6040# cap_series_gyp a_21636_6040# vss nmos_6p0 w=0.82u l=0.6u
X6596 a_33524_30644# cap_shunt_n a_33732_31128# vdd pmos_6p0 w=1.2u l=0.5u
X6597 a_17620_36916# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6598 a_28484_8692# cap_series_gyn a_28692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X6599 vdd a_37196_27464# a_37108_27508# vdd pmos_6p0 w=1.22u l=1u
X6600 a_35692_25940# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6601 a_33948_52552# a_33860_52596# vss vss nmos_6p0 w=0.82u l=1u
X6602 a_18404_9884# cap_series_gyp a_18612_9538# vdd pmos_6p0 w=1.2u l=0.5u
X6603 a_16708_18946# cap_shunt_p a_18424_18884# vss nmos_6p0 w=0.82u l=0.6u
X6604 vdd a_18716_55688# a_18628_55732# vdd pmos_6p0 w=1.22u l=1u
X6605 vss cap_shunt_n a_19936_35832# vss nmos_6p0 w=0.82u l=0.6u
X6606 a_21540_6748# cap_series_gyn a_21748_6402# vdd pmos_6p0 w=1.2u l=0.5u
X6607 a_26768_18884# cap_series_gyn a_24660_18946# vss nmos_6p0 w=0.82u l=0.6u
X6608 a_6532_44756# cap_shunt_p a_6740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X6609 a_21748_14242# cap_series_gyn a_21540_14588# vdd pmos_6p0 w=1.2u l=0.5u
X6610 a_33732_35832# cap_shunt_n a_34664_35832# vss nmos_6p0 w=0.82u l=0.6u
X6611 a_22064_34264# cap_shunt_n a_20740_34264# vss nmos_6p0 w=0.82u l=0.6u
X6612 a_11780_6040# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X6613 a_35880_8692# cap_series_gygyn a_35692_8692# vdd pmos_6p0 w=1.2u l=0.5u
X6614 a_17828_18584# cap_shunt_p a_17620_18100# vdd pmos_6p0 w=1.2u l=0.5u
X6615 vss tune_shunt[7] a_9316_22082# vss nmos_6p0 w=0.51u l=0.6u
X6616 a_28484_5556# cap_shunt_n a_28692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X6617 a_25780_17016# cap_series_gyp a_25572_16532# vdd pmos_6p0 w=1.2u l=0.5u
X6618 a_35692_22804# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6619 a_18404_6748# cap_series_gyn a_18612_6402# vdd pmos_6p0 w=1.2u l=0.5u
X6620 a_16708_15810# cap_shunt_p a_18424_15748# vss nmos_6p0 w=0.82u l=0.6u
X6621 vdd a_30924_52552# a_30836_52596# vdd pmos_6p0 w=1.22u l=1u
X6622 vdd a_35292_3944# a_35204_3988# vdd pmos_6p0 w=1.22u l=1u
X6623 a_3640_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6624 a_6776_10744# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6625 a_26768_15748# cap_series_gyn a_24660_15810# vss nmos_6p0 w=0.82u l=0.6u
X6626 a_3172_49460# cap_shunt_p a_3380_49944# vdd pmos_6p0 w=1.2u l=0.5u
X6627 a_3828_38968# cap_shunt_n a_3620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X6628 a_19276_34871# a_19188_34968# vss vss nmos_6p0 w=0.82u l=1u
X6629 vdd a_33052_55255# a_32964_55352# vdd pmos_6p0 w=1.22u l=1u
X6630 a_22064_31128# cap_shunt_n a_20740_31128# vss nmos_6p0 w=0.82u l=0.6u
X6631 a_35880_5556# cap_series_gygyn a_35692_5556# vdd pmos_6p0 w=1.2u l=0.5u
X6632 a_27340_50984# a_27252_51028# vss vss nmos_6p0 w=0.82u l=1u
X6633 vdd tune_series_gy[5] a_18404_13020# vdd pmos_6p0 w=1.2u l=0.5u
X6634 vss cap_shunt_n a_8848_38968# vss nmos_6p0 w=0.82u l=0.6u
X6635 vss cap_shunt_p a_23856_34564# vss nmos_6p0 w=0.82u l=0.6u
X6636 a_21748_17378# cap_shunt_p a_21540_17724# vdd pmos_6p0 w=1.2u l=0.5u
X6637 a_14372_43188# cap_shunt_n a_14580_43672# vdd pmos_6p0 w=1.2u l=0.5u
X6638 a_3828_35832# cap_shunt_n a_3620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X6639 a_19276_31735# a_19188_31832# vss vss nmos_6p0 w=0.82u l=1u
X6640 vdd a_33052_52119# a_32964_52216# vdd pmos_6p0 w=1.22u l=1u
X6641 vdd a_30476_47848# a_30388_47892# vdd pmos_6p0 w=1.22u l=1u
X6642 a_10548_35832# cap_shunt_n a_12264_35832# vss nmos_6p0 w=0.82u l=0.6u
X6643 vdd a_37868_31735# a_37780_31832# vdd pmos_6p0 w=1.22u l=1u
X6644 a_9668_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6645 vss cap_series_gyp a_22960_6040# vss nmos_6p0 w=0.82u l=0.6u
X6646 a_26712_17016# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6647 a_24316_50984# a_24228_51028# vss vss nmos_6p0 w=0.82u l=1u
X6648 a_3036_36872# a_2948_36916# vss vss nmos_6p0 w=0.82u l=1u
X6649 a_3620_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6650 vss cap_shunt_n a_23856_31428# vss nmos_6p0 w=0.82u l=0.6u
X6651 a_25780_26424# cap_shunt_p a_25572_25940# vdd pmos_6p0 w=1.2u l=0.5u
X6652 vdd a_30476_44712# a_30388_44756# vdd pmos_6p0 w=1.22u l=1u
X6653 vdd a_37644_29032# a_37556_29076# vdd pmos_6p0 w=1.22u l=1u
X6654 a_32404_27132# cap_shunt_p a_32612_26786# vdd pmos_6p0 w=1.2u l=0.5u
X6655 a_24452_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6656 a_9644_7080# a_9556_7124# vss vss nmos_6p0 w=0.82u l=1u
X6657 a_24660_6402# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X6658 a_5844_9176# cap_shunt_p a_7560_9176# vss nmos_6p0 w=0.82u l=0.6u
X6659 vdd a_6172_54120# a_6084_54164# vdd pmos_6p0 w=1.22u l=1u
X6660 a_23072_32996# cap_shunt_n a_21748_33058# vss nmos_6p0 w=0.82u l=0.6u
X6661 a_29492_23996# cap_shunt_p a_29700_23650# vdd pmos_6p0 w=1.2u l=0.5u
X6662 a_3620_13396# cap_shunt_n a_3828_13880# vdd pmos_6p0 w=1.2u l=0.5u
X6663 vdd tune_series_gygy[5] a_31436_22428# vdd pmos_6p0 w=1.2u l=0.5u
X6664 a_25780_23288# cap_shunt_p a_25572_22804# vdd pmos_6p0 w=1.2u l=0.5u
X6665 vdd a_5612_55255# a_5524_55352# vdd pmos_6p0 w=1.22u l=1u
X6666 a_36636_40008# a_36548_40052# vss vss nmos_6p0 w=0.82u l=1u
X6667 a_12376_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6668 a_24452_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6669 a_16800_7608# cap_series_gyp a_14692_7608# vss nmos_6p0 w=0.82u l=0.6u
X6670 vss tune_shunt[5] a_21748_42466# vss nmos_6p0 w=0.51u l=0.6u
X6671 a_6740_34264# cap_shunt_n a_8456_34264# vss nmos_6p0 w=0.82u l=0.6u
X6672 a_3828_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6673 vdd tune_shunt[5] a_6084_51028# vdd pmos_6p0 w=1.2u l=0.5u
X6674 a_1924_6040# cap_shunt_p a_1716_5556# vdd pmos_6p0 w=1.2u l=0.5u
X6675 a_21540_13020# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6676 vss cap_series_gygyn a_36296_17016# vss nmos_6p0 w=0.82u l=0.6u
X6677 a_17828_38968# cap_shunt_n a_17620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X6678 vdd a_5612_52119# a_5524_52216# vdd pmos_6p0 w=1.22u l=1u
X6679 a_10452_44380# cap_shunt_n a_10660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X6680 vss cap_shunt_p a_27104_38968# vss nmos_6p0 w=0.82u l=0.6u
X6681 a_12376_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6682 a_22644_9176# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6683 a_6740_31128# cap_shunt_n a_8456_31128# vss nmos_6p0 w=0.82u l=0.6u
X6684 a_3828_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6685 a_9668_47892# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6686 vss cap_shunt_gyn a_32732_46808# vss nmos_6p0 w=0.82u l=0.6u
X6687 a_17828_35832# cap_shunt_n a_17620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X6688 vss cap_shunt_n a_19936_29560# vss nmos_6p0 w=0.82u l=0.6u
X6689 a_6740_27992# cap_shunt_n a_6532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X6690 a_34308_5180# tune_series_gygy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6691 a_18940_55255# a_18852_55352# vss vss nmos_6p0 w=0.82u l=1u
X6692 a_11460_40052# cap_shunt_n a_11668_40536# vdd pmos_6p0 w=1.2u l=0.5u
X6693 a_29700_37762# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6694 a_7672_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6695 a_6532_38484# cap_shunt_n a_6740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X6696 a_10452_41244# cap_shunt_n a_10660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X6697 a_5612_33303# a_5524_33400# vss vss nmos_6p0 w=0.82u l=1u
X6698 a_33732_29560# cap_shunt_p a_34664_29560# vss nmos_6p0 w=0.82u l=0.6u
X6699 vdd a_21180_49416# a_21092_49460# vdd pmos_6p0 w=1.22u l=1u
X6700 vdd a_28572_33303# a_28484_33400# vdd pmos_6p0 w=1.22u l=1u
X6701 a_17620_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6702 a_9428_20514# cap_shunt_p a_9220_20860# vdd pmos_6p0 w=1.2u l=0.5u
X6703 a_8008_51512# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6704 a_35692_16532# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6705 a_29700_37762# cap_shunt_n a_31416_37700# vss nmos_6p0 w=0.82u l=0.6u
X6706 vss tune_shunt[7] a_17828_32696# vss nmos_6p0 w=0.51u l=0.6u
X6707 vdd tune_series_gy[3] a_14484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X6708 vdd a_8860_16055# a_8772_16152# vdd pmos_6p0 w=1.22u l=1u
X6709 vdd a_1692_31735# a_1604_31832# vdd pmos_6p0 w=1.22u l=1u
X6710 vss cap_shunt_n a_19936_26424# vss nmos_6p0 w=0.82u l=0.6u
X6711 a_18612_11106# cap_series_gyn a_18404_11452# vdd pmos_6p0 w=1.2u l=0.5u
X6712 a_6532_35348# cap_shunt_n a_6740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X6713 a_29700_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6714 a_19544_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X6715 vdd a_33052_48983# a_32964_49080# vdd pmos_6p0 w=1.22u l=1u
X6716 a_19276_28599# a_19188_28696# vss vss nmos_6p0 w=0.82u l=1u
X6717 vdd a_31260_10216# a_31172_10260# vdd pmos_6p0 w=1.22u l=1u
X6718 a_29532_9884# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6719 a_27340_44712# a_27252_44756# vss vss nmos_6p0 w=0.82u l=1u
X6720 a_7748_33058# cap_shunt_n a_9464_32996# vss nmos_6p0 w=0.82u l=0.6u
X6721 a_17620_41620# cap_shunt_n a_17828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X6722 a_24660_12674# cap_series_gyn a_24452_13020# vdd pmos_6p0 w=1.2u l=0.5u
X6723 a_3640_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6724 vss cap_shunt_n a_23856_28292# vss nmos_6p0 w=0.82u l=0.6u
X6725 a_31416_14180# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6726 a_14460_53687# a_14372_53784# vss vss nmos_6p0 w=0.82u l=1u
X6727 vdd a_20620_47415# a_20532_47512# vdd pmos_6p0 w=1.22u l=1u
X6728 a_13796_17378# cap_shunt_p a_13588_17724# vdd pmos_6p0 w=1.2u l=0.5u
X6729 a_10548_29560# cap_shunt_n a_12264_29560# vss nmos_6p0 w=0.82u l=0.6u
X6730 a_3828_29560# cap_shunt_n a_3620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X6731 a_19276_25463# a_19188_25560# vss vss nmos_6p0 w=0.82u l=1u
X6732 vdd a_37868_25463# a_37780_25560# vdd pmos_6p0 w=1.22u l=1u
X6733 a_10452_6748# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6734 vdd a_2588_36872# a_2500_36916# vdd pmos_6p0 w=1.22u l=1u
X6735 a_8412_3511# a_8324_3608# vss vss nmos_6p0 w=0.82u l=1u
X6736 a_6532_47892# cap_shunt_p a_6740_48376# vdd pmos_6p0 w=1.2u l=0.5u
X6737 vss cap_shunt_n a_23856_25156# vss nmos_6p0 w=0.82u l=0.6u
X6738 a_31416_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6739 a_37868_8215# a_37780_8312# vss vss nmos_6p0 w=0.82u l=1u
X6740 vdd a_14012_11351# a_13924_11448# vdd pmos_6p0 w=1.22u l=1u
X6741 vdd tune_series_gygy[4] a_31436_19292# vdd pmos_6p0 w=1.2u l=0.5u
X6742 a_10548_26424# cap_shunt_n a_12264_26424# vss nmos_6p0 w=0.82u l=0.6u
X6743 vdd a_37868_22327# a_37780_22424# vdd pmos_6p0 w=1.22u l=1u
X6744 a_24452_19292# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6745 a_20532_33780# cap_shunt_n a_20740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X6746 vdd a_36972_55688# a_36884_55732# vdd pmos_6p0 w=1.22u l=1u
X6747 a_6532_44756# cap_shunt_p a_6740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X6748 a_11480_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6749 a_25780_17016# cap_series_gyp a_25572_16532# vdd pmos_6p0 w=1.2u l=0.5u
X6750 a_24204_52119# a_24116_52216# vss vss nmos_6p0 w=0.82u l=1u
X6751 vdd a_16364_50551# a_16276_50648# vdd pmos_6p0 w=1.22u l=1u
X6752 a_13796_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6753 a_19732_12312# cap_series_gyn a_19524_11828# vdd pmos_6p0 w=1.2u l=0.5u
X6754 vdd a_5612_48983# a_5524_49080# vdd pmos_6p0 w=1.22u l=1u
X6755 vdd tune_shunt[6] a_11460_46324# vdd pmos_6p0 w=1.2u l=0.5u
X6756 a_24660_39330# cap_shunt_p a_26376_39268# vss nmos_6p0 w=0.82u l=0.6u
X6757 a_16408_10744# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X6758 vdd tune_shunt[7] a_17620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X6759 a_24452_16156# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6760 vss tune_shunt[6] a_21748_36194# vss nmos_6p0 w=0.51u l=0.6u
X6761 a_23072_23588# cap_shunt_p a_21748_23650# vss nmos_6p0 w=0.82u l=0.6u
X6762 a_11800_7124# cap_series_gyp a_11612_7124# vdd pmos_6p0 w=1.2u l=0.5u
X6763 a_20532_30644# cap_shunt_n a_20740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X6764 a_29492_14588# cap_series_gyp a_29700_14242# vdd pmos_6p0 w=1.2u l=0.5u
X6765 a_25572_43188# cap_shunt_p a_25780_43672# vdd pmos_6p0 w=1.2u l=0.5u
X6766 a_11480_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6767 vdd a_33948_55688# a_33860_55732# vdd pmos_6p0 w=1.22u l=1u
X6768 a_18760_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6769 vss cap_shunt_gyn a_34748_46808# vss nmos_6p0 w=0.82u l=0.6u
X6770 a_18612_12674# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6771 a_10248_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6772 vss tune_shunt[6] a_16708_40898# vss nmos_6p0 w=0.51u l=0.6u
X6773 vss tune_shunt[7] a_21748_33058# vss nmos_6p0 w=0.51u l=0.6u
X6774 a_11884_54120# a_11796_54164# vss vss nmos_6p0 w=0.82u l=1u
X6775 vdd a_28012_3511# a_27924_3608# vdd pmos_6p0 w=1.22u l=1u
X6776 a_37084_54120# a_36996_54164# vss vss nmos_6p0 w=0.82u l=1u
X6777 a_6740_46808# cap_shunt_p a_7672_46808# vss nmos_6p0 w=0.82u l=0.6u
X6778 a_14372_43188# cap_shunt_n a_14580_43672# vdd pmos_6p0 w=1.2u l=0.5u
X6779 a_33920_43734# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6780 a_37280_44757# tune_shunt_gy[3] vdd vdd pmos_6p0 w=1.215u l=0.5u
X6781 a_17828_29560# cap_shunt_n a_17620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X6782 vss tune_shunt[7] a_13796_15810# vss nmos_6p0 w=0.51u l=0.6u
X6783 vdd a_26892_47848# a_26804_47892# vdd pmos_6p0 w=1.22u l=1u
X6784 vss cap_series_gygyp a_35840_20452# vss nmos_6p0 w=0.82u l=0.6u
X6785 vdd a_26444_55255# a_26356_55352# vdd pmos_6p0 w=1.22u l=1u
X6786 a_25572_19668# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6787 vdd a_1692_25463# a_1604_25560# vdd pmos_6p0 w=1.22u l=1u
X6788 a_29700_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6789 a_29492_23996# cap_shunt_p a_29700_23650# vdd pmos_6p0 w=1.2u l=0.5u
X6790 a_7672_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6791 vdd a_33500_18056# a_33412_18100# vdd pmos_6p0 w=1.22u l=1u
X6792 a_6532_29076# cap_shunt_n a_6740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X6793 a_5612_23895# a_5524_23992# vss vss nmos_6p0 w=0.82u l=1u
X6794 a_1716_5180# cap_shunt_p a_1924_4834# vdd pmos_6p0 w=1.2u l=0.5u
X6795 vdd a_26892_44712# a_26804_44756# vdd pmos_6p0 w=1.22u l=1u
X6796 vdd a_26444_52119# a_26356_52216# vdd pmos_6p0 w=1.22u l=1u
X6797 a_31372_50984# a_31284_51028# vss vss nmos_6p0 w=0.82u l=1u
X6798 vdd tune_series_gygy[5] a_31436_22428# vdd pmos_6p0 w=1.2u l=0.5u
X6799 vss tune_shunt[7] a_17828_23288# vss nmos_6p0 w=0.51u l=0.6u
X6800 vdd a_1692_22327# a_1604_22424# vdd pmos_6p0 w=1.22u l=1u
X6801 a_34720_29860# cap_shunt_p a_32612_29922# vss nmos_6p0 w=0.82u l=0.6u
X6802 a_29624_13880# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6803 vss cap_shunt_p a_19936_17016# vss nmos_6p0 w=0.82u l=0.6u
X6804 a_6292_17016# cap_shunt_p a_8008_17016# vss nmos_6p0 w=0.82u l=0.6u
X6805 a_3380_51512# cap_shunt_n a_3172_51028# vdd pmos_6p0 w=1.2u l=0.5u
X6806 a_29700_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6807 a_10340_36916# cap_shunt_n a_10548_37400# vdd pmos_6p0 w=1.2u l=0.5u
X6808 vdd tune_shunt[6] a_12580_47892# vdd pmos_6p0 w=1.2u l=0.5u
X6809 a_5936_38968# cap_shunt_n a_3828_38968# vss nmos_6p0 w=0.82u l=0.6u
X6810 a_9644_54120# a_9556_54164# vss vss nmos_6p0 w=0.82u l=1u
X6811 a_17620_32212# cap_shunt_n a_17828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X6812 a_7748_23650# cap_shunt_p a_9464_23588# vss nmos_6p0 w=0.82u l=0.6u
X6813 a_34720_26724# cap_shunt_p a_32612_26786# vss nmos_6p0 w=0.82u l=0.6u
X6814 vdd tune_series_gy[5] a_18404_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6815 a_29624_10744# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X6816 a_19544_46808# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6817 vdd a_20620_38007# a_20532_38104# vdd pmos_6p0 w=1.22u l=1u
X6818 vdd tune_shunt[7] a_7540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X6819 a_21748_4834# cap_series_gyp a_21540_5180# vdd pmos_6p0 w=1.2u l=0.5u
X6820 vdd a_29244_21192# a_29156_21236# vdd pmos_6p0 w=1.22u l=1u
X6821 vdd a_37868_16055# a_37780_16152# vdd pmos_6p0 w=1.22u l=1u
X6822 a_21540_34972# cap_shunt_p a_21748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X6823 a_13796_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6824 vdd a_2588_27464# a_2500_27508# vdd pmos_6p0 w=1.22u l=1u
X6825 vss tune_shunt[7] a_20740_20152# vss nmos_6p0 w=0.51u l=0.6u
X6826 a_6532_38484# cap_shunt_n a_6740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X6827 vdd tune_series_gy[4] a_18404_6748# vdd pmos_6p0 w=1.2u l=0.5u
X6828 vdd tune_shunt[7] a_7540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X6829 a_20620_19191# a_20532_19288# vss vss nmos_6p0 w=0.82u l=1u
X6830 vss tune_shunt[5] a_20740_43672# vss nmos_6p0 w=0.51u l=0.6u
X6831 a_13796_36194# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6832 a_9316_48738# cap_shunt_p a_11032_48676# vss nmos_6p0 w=0.82u l=0.6u
X6833 vss cap_shunt_n a_22848_37400# vss nmos_6p0 w=0.82u l=0.6u
X6834 vdd a_37868_12919# a_37780_13016# vdd pmos_6p0 w=1.22u l=1u
X6835 a_21540_31836# cap_shunt_n a_21748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X6836 vss tune_shunt[5] a_3380_51512# vss nmos_6p0 w=0.51u l=0.6u
X6837 a_20532_24372# cap_shunt_n a_20740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X6838 a_35840_18884# cap_series_gygyn a_34516_18946# vss nmos_6p0 w=0.82u l=0.6u
X6839 a_6532_35348# cap_shunt_n a_6740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X6840 vdd a_32268_9783# a_32180_9880# vdd pmos_6p0 w=1.22u l=1u
X6841 vdd a_33948_49416# a_33860_49460# vdd pmos_6p0 w=1.22u l=1u
X6842 a_10092_43144# a_10004_43188# vss vss nmos_6p0 w=0.82u l=1u
X6843 vss tune_shunt[6] a_20740_40536# vss nmos_6p0 w=0.51u l=0.6u
X6844 a_13796_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6845 a_2500_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6846 a_20620_16055# a_20532_16152# vss vss nmos_6p0 w=0.82u l=1u
X6847 a_31820_52552# a_31732_52596# vss vss nmos_6p0 w=0.82u l=1u
X6848 vdd a_26108_45847# a_26020_45944# vdd pmos_6p0 w=1.22u l=1u
X6849 a_15512_22020# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X6850 a_2708_48738# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6851 vdd tune_shunt[6] a_10452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X6852 a_35840_15748# cap_series_gygyn a_34516_15810# vss nmos_6p0 w=0.82u l=0.6u
X6853 a_6084_19292# cap_shunt_p a_6292_18946# vdd pmos_6p0 w=1.2u l=0.5u
X6854 a_20532_21236# cap_shunt_p a_20740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X6855 a_13796_17378# cap_shunt_p a_13588_17724# vdd pmos_6p0 w=1.2u l=0.5u
X6856 a_29700_39330# cap_shunt_p a_29492_39676# vdd pmos_6p0 w=1.2u l=0.5u
X6857 vdd a_2140_52552# a_2052_52596# vdd pmos_6p0 w=1.22u l=1u
X6858 a_35264_48676# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6859 a_36524_34871# a_36436_34968# vss vss nmos_6p0 w=0.82u l=1u
X6860 a_6740_13880# cap_shunt_p a_6532_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6861 a_10092_40008# a_10004_40052# vss vss nmos_6p0 w=0.82u l=1u
X6862 a_7540_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6863 a_6532_47892# cap_shunt_p a_6740_48376# vdd pmos_6p0 w=1.2u l=0.5u
X6864 vdd tune_series_gy[3] a_29532_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6865 a_24652_46280# a_24564_46324# vss vss nmos_6p0 w=0.82u l=1u
X6866 vss cap_shunt_n a_14784_35832# vss nmos_6p0 w=0.82u l=0.6u
X6867 a_6084_16156# cap_shunt_p a_6292_15810# vdd pmos_6p0 w=1.2u l=0.5u
X6868 vdd a_26444_48983# a_26356_49080# vdd pmos_6p0 w=1.22u l=1u
X6869 a_21748_37762# cap_shunt_n a_21540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X6870 a_35880_13396# cap_series_gygyn a_35692_13396# vdd pmos_6p0 w=1.2u l=0.5u
X6871 a_31708_13352# a_31620_13396# vss vss nmos_6p0 w=0.82u l=1u
X6872 vdd tune_series_gygy[4] a_31436_19292# vdd pmos_6p0 w=1.2u l=0.5u
X6873 a_21628_49416# a_21540_49460# vss vss nmos_6p0 w=0.82u l=1u
X6874 a_3828_34264# cap_shunt_n a_3620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X6875 a_36524_31735# a_36436_31832# vss vss nmos_6p0 w=0.82u l=1u
X6876 a_13252_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6877 a_3620_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6878 a_6532_44756# cap_shunt_p a_6740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X6879 a_36076_30167# a_35988_30264# vss vss nmos_6p0 w=0.82u l=1u
X6880 vdd tune_shunt[4] a_24452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X6881 a_31708_10216# a_31620_10260# vss vss nmos_6p0 w=0.82u l=1u
X6882 vss tune_shunt[6] a_9876_49944# vss nmos_6p0 w=0.51u l=0.6u
X6883 a_3828_31128# cap_shunt_n a_3620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X6884 vdd tune_shunt[7] a_20532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X6885 a_19732_12312# cap_series_gyn a_19524_11828# vdd pmos_6p0 w=1.2u l=0.5u
X6886 vdd a_1692_16055# a_1604_16152# vdd pmos_6p0 w=1.22u l=1u
X6887 vdd tune_shunt[6] a_11460_46324# vdd pmos_6p0 w=1.2u l=0.5u
X6888 a_13252_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6889 a_17828_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6890 vdd a_27228_34871# a_27140_34968# vdd pmos_6p0 w=1.22u l=1u
X6891 a_14484_8692# cap_series_gyn a_14692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X6892 a_3620_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6893 a_29492_14588# cap_series_gyp a_29700_14242# vdd pmos_6p0 w=1.2u l=0.5u
X6894 a_36076_27031# a_35988_27128# vss vss nmos_6p0 w=0.82u l=1u
X6895 a_28484_18100# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6896 a_6516_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6897 a_33948_38440# a_33860_38484# vss vss nmos_6p0 w=0.82u l=1u
X6898 a_13796_29922# cap_shunt_n a_14728_29860# vss nmos_6p0 w=0.82u l=0.6u
X6899 vss tune_shunt[7] a_21748_23650# vss nmos_6p0 w=0.51u l=0.6u
X6900 vdd tune_shunt[7] a_20532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X6901 vss cap_shunt_p a_5936_21720# vss nmos_6p0 w=0.82u l=0.6u
X6902 vss cap_shunt_n a_19152_32696# vss nmos_6p0 w=0.82u l=0.6u
X6903 a_29532_13020# cap_series_gyn a_29720_13020# vdd pmos_6p0 w=1.2u l=0.5u
X6904 vdd a_1692_12919# a_1604_13016# vdd pmos_6p0 w=1.22u l=1u
X6905 a_17828_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6906 a_14484_5556# cap_series_gyn a_14692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X6907 a_31260_52119# a_31172_52216# vss vss nmos_6p0 w=0.82u l=1u
X6908 a_29492_39676# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6909 a_22644_13880# cap_series_gyn a_24360_13880# vss nmos_6p0 w=0.82u l=0.6u
X6910 vss cap_series_gyn a_30136_15748# vss nmos_6p0 w=0.82u l=0.6u
X6911 a_26376_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X6912 a_13796_39330# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6913 a_10340_27508# cap_shunt_n a_10548_27992# vdd pmos_6p0 w=1.2u l=0.5u
X6914 a_13796_26786# cap_shunt_n a_14728_26724# vss nmos_6p0 w=0.82u l=0.6u
X6915 a_28692_38968# cap_shunt_n a_29624_38968# vss nmos_6p0 w=0.82u l=0.6u
X6916 vss tune_shunt[7] a_21748_20514# vss nmos_6p0 w=0.51u l=0.6u
X6917 a_11996_19191# a_11908_19288# vss vss nmos_6p0 w=0.82u l=1u
X6918 vdd tune_shunt[7] a_7540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X6919 a_22644_10744# cap_series_gyp a_24360_10744# vss nmos_6p0 w=0.82u l=0.6u
X6920 vdd a_20396_50551# a_20308_50648# vdd pmos_6p0 w=1.22u l=1u
X6921 a_29916_44279# a_29828_44376# vss vss nmos_6p0 w=0.82u l=1u
X6922 vdd a_32604_40008# a_32516_40052# vdd pmos_6p0 w=1.22u l=1u
X6923 a_17828_34264# cap_shunt_n a_17620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X6924 a_23072_6340# cap_series_gyn a_21748_6402# vss nmos_6p0 w=0.82u l=0.6u
X6925 a_21540_25564# cap_shunt_n a_21748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X6926 a_30428_19668# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X6927 a_13460_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X6928 vss tune_shunt[6] a_3828_45240# vss nmos_6p0 w=0.51u l=0.6u
X6929 a_6532_29076# cap_shunt_n a_6740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X6930 a_29492_23996# cap_shunt_p a_29700_23650# vdd pmos_6p0 w=1.2u l=0.5u
X6931 a_1924_4472# cap_shunt_p a_1716_3988# vdd pmos_6p0 w=1.2u l=0.5u
X6932 vss cap_shunt_p a_33936_37700# vss nmos_6p0 w=0.82u l=0.6u
X6933 a_29916_41143# a_29828_41240# vss vss nmos_6p0 w=0.82u l=1u
X6934 a_33732_35832# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X6935 vss tune_shunt[7] a_20740_34264# vss nmos_6p0 w=0.51u l=0.6u
X6936 a_9428_17378# cap_shunt_p a_9220_17724# vdd pmos_6p0 w=1.2u l=0.5u
X6937 a_34144_47108# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6938 a_17828_31128# cap_shunt_n a_17620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X6939 a_6508_55255# a_6420_55352# vss vss nmos_6p0 w=0.82u l=1u
X6940 a_21540_22428# cap_shunt_p a_21748_22082# vdd pmos_6p0 w=1.2u l=0.5u
X6941 a_3380_51512# cap_shunt_n a_3172_51028# vdd pmos_6p0 w=1.2u l=0.5u
X6942 a_6292_50306# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6943 vss tune_shunt[6] a_3828_42104# vss nmos_6p0 w=0.51u l=0.6u
X6944 a_36384_50648# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X6945 vdd tune_shunt[5] a_2500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X6946 a_15568_38968# cap_shunt_n a_13460_38968# vss nmos_6p0 w=0.82u l=0.6u
X6947 vdd a_19836_55255# a_19748_55352# vdd pmos_6p0 w=1.22u l=1u
X6948 a_36524_28599# a_36436_28696# vss vss nmos_6p0 w=0.82u l=1u
X6949 vss tune_shunt[7] a_20740_31128# vss nmos_6p0 w=0.51u l=0.6u
X6950 a_11592_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6951 vss cap_series_gyp a_21056_7608# vss nmos_6p0 w=0.82u l=0.6u
X6952 a_15700_6402# cap_series_gyp a_16632_6340# vss nmos_6p0 w=0.82u l=0.6u
X6953 a_3620_46324# cap_shunt_p a_3828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X6954 vss cap_shunt_n a_25984_42404# vss nmos_6p0 w=0.82u l=0.6u
X6955 a_32604_32168# a_32516_32212# vss vss nmos_6p0 w=0.82u l=1u
X6956 vdd a_32156_32168# a_32068_32212# vdd pmos_6p0 w=1.22u l=1u
X6957 vss cap_shunt_n a_14784_29560# vss nmos_6p0 w=0.82u l=0.6u
X6958 a_9316_22082# cap_shunt_p a_10248_22020# vss nmos_6p0 w=0.82u l=0.6u
X6959 vdd a_34844_8648# a_34756_8692# vdd pmos_6p0 w=1.22u l=1u
X6960 a_22436_11828# cap_series_gyn a_22644_12312# vdd pmos_6p0 w=1.2u l=0.5u
X6961 vdd a_19836_52119# a_19748_52216# vdd pmos_6p0 w=1.22u l=1u
X6962 a_24764_50984# a_24676_51028# vss vss nmos_6p0 w=0.82u l=1u
X6963 vdd a_2140_43144# a_2052_43188# vdd pmos_6p0 w=1.22u l=1u
X6964 vdd tune_shunt[7] a_24452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X6965 vdd a_6508_30167# a_6420_30264# vdd pmos_6p0 w=1.22u l=1u
X6966 a_36524_25463# a_36436_25560# vss vss nmos_6p0 w=0.82u l=1u
X6967 vdd tune_shunt[5] a_28484_32212# vdd pmos_6p0 w=1.2u l=0.5u
X6968 a_35740_3511# a_35652_3608# vss vss nmos_6p0 w=0.82u l=1u
X6969 a_3828_45240# cap_shunt_p a_4760_45240# vss nmos_6p0 w=0.82u l=0.6u
X6970 a_6532_38484# cap_shunt_n a_6740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X6971 vdd tune_shunt[6] a_24452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X6972 vss cap_shunt_n a_14784_26424# vss nmos_6p0 w=0.82u l=0.6u
X6973 vdd a_34844_5512# a_34756_5556# vdd pmos_6p0 w=1.22u l=1u
X6974 a_18404_3988# cap_series_gyp a_18612_4472# vdd pmos_6p0 w=1.2u l=0.5u
X6975 a_3828_24856# cap_shunt_p a_3620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X6976 vdd a_27228_28599# a_27140_28696# vdd pmos_6p0 w=1.22u l=1u
X6977 a_10808_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X6978 a_32156_27464# a_32068_27508# vss vss nmos_6p0 w=0.82u l=1u
X6979 a_3828_42104# cap_shunt_p a_4760_42104# vss nmos_6p0 w=0.82u l=0.6u
X6980 a_6740_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X6981 a_17620_43188# cap_shunt_p a_17828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X6982 a_6532_35348# cap_shunt_n a_6740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X6983 vdd tune_series_gy[3] a_28484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X6984 vss tune_shunt[3] a_25780_43672# vss nmos_6p0 w=0.51u l=0.6u
X6985 vdd tune_shunt[6] a_24452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X6986 vdd tune_series_gy[5] a_18404_9884# vdd pmos_6p0 w=1.2u l=0.5u
X6987 a_3828_21720# cap_shunt_p a_3620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X6988 vdd a_22412_53687# a_22324_53784# vdd pmos_6p0 w=1.22u l=1u
X6989 a_30812_22327# a_30724_22424# vss vss nmos_6p0 w=0.82u l=1u
X6990 vss cap_shunt_p a_14112_13880# vss nmos_6p0 w=0.82u l=0.6u
X6991 vdd tune_shunt[4] a_20532_16532# vdd pmos_6p0 w=1.2u l=0.5u
X6992 a_9428_20514# cap_shunt_p a_10360_20452# vss nmos_6p0 w=0.82u l=0.6u
X6993 a_9876_53080# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X6994 a_32156_24328# a_32068_24372# vss vss nmos_6p0 w=0.82u l=1u
X6995 a_6084_19292# cap_shunt_p a_6292_18946# vdd pmos_6p0 w=1.2u l=0.5u
X6996 a_6084_49084# cap_shunt_p a_6292_48738# vdd pmos_6p0 w=1.2u l=0.5u
X6997 vss tune_shunt[3] a_5844_11106# vss nmos_6p0 w=0.51u l=0.6u
X6998 a_6420_14588# cap_shunt_p a_6628_14242# vdd pmos_6p0 w=1.2u l=0.5u
X6999 vdd tune_shunt[0] a_28484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X7000 vss tune_shunt[6] a_14580_43672# vss nmos_6p0 w=0.51u l=0.6u
X7001 vss tune_shunt[5] a_25780_40536# vss nmos_6p0 w=0.51u l=0.6u
X7002 a_29700_39330# cap_shunt_p a_29492_39676# vdd pmos_6p0 w=1.2u l=0.5u
X7003 vss tune_series_gy[2] a_11780_6040# vss nmos_6p0 w=0.51u l=0.6u
X7004 vdd tune_series_gy[4] a_18404_6748# vdd pmos_6p0 w=1.2u l=0.5u
X7005 vdd a_11212_53687# a_11124_53784# vdd pmos_6p0 w=1.22u l=1u
X7006 vdd a_22412_50551# a_22324_50648# vdd pmos_6p0 w=1.22u l=1u
X7007 vss tune_series_gy[5] a_21748_14242# vss nmos_6p0 w=0.51u l=0.6u
X7008 vss tune_series_gygy[4] a_34516_15810# vss nmos_6p0 w=0.51u l=0.6u
X7009 vss cap_shunt_n a_19152_23288# vss nmos_6p0 w=0.82u l=0.6u
X7010 a_9464_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7011 a_32612_33058# cap_shunt_n a_34328_32996# vss nmos_6p0 w=0.82u l=0.6u
X7012 a_35692_3988# tune_series_gygy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7013 a_6084_16156# cap_shunt_p a_6292_15810# vdd pmos_6p0 w=1.2u l=0.5u
X7014 a_31260_42711# a_31172_42808# vss vss nmos_6p0 w=0.82u l=1u
X7015 a_21748_37762# cap_shunt_n a_21540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X7016 vdd a_31820_55688# a_31732_55732# vdd pmos_6p0 w=1.22u l=1u
X7017 vss tune_shunt[6] a_14580_40536# vss nmos_6p0 w=0.51u l=0.6u
X7018 a_13252_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7019 a_21540_19292# cap_shunt_p a_21748_18946# vdd pmos_6p0 w=1.2u l=0.5u
X7020 a_33732_32696# cap_shunt_n a_33524_32212# vdd pmos_6p0 w=1.2u l=0.5u
X7021 a_13796_17378# cap_shunt_p a_14728_17316# vss nmos_6p0 w=0.82u l=0.6u
X7022 vss tune_series_gy[5] a_21748_11106# vss nmos_6p0 w=0.51u l=0.6u
X7023 a_6628_12674# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7024 vdd a_34396_13352# a_34308_13396# vdd pmos_6p0 w=1.22u l=1u
X7025 a_18032_18884# cap_shunt_p a_16708_18946# vss nmos_6p0 w=0.82u l=0.6u
X7026 a_24452_8316# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7027 a_21748_22082# cap_shunt_p a_23464_22020# vss nmos_6p0 w=0.82u l=0.6u
X7028 a_33024_43972# cap_shunt_gyn a_33024_44376# vdd pmos_6p0 w=1.215u l=0.5u
X7029 a_33732_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7030 a_17828_24856# cap_shunt_n a_17620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7031 vdd a_32268_17623# a_32180_17720# vdd pmos_6p0 w=1.22u l=1u
X7032 a_13252_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7033 a_21540_16156# cap_series_gyn a_21748_15810# vdd pmos_6p0 w=1.2u l=0.5u
X7034 a_22644_7608# cap_series_gyp a_23576_7608# vss nmos_6p0 w=0.82u l=0.6u
X7035 a_31436_6748# cap_series_gygyn a_31624_6748# vdd pmos_6p0 w=1.2u l=0.5u
X7036 a_36384_44376# tune_shunt_gy[3] vdd vdd pmos_6p0 w=1.215u l=0.5u
X7037 a_29492_14588# cap_series_gyp a_29700_14242# vdd pmos_6p0 w=1.2u l=0.5u
X7038 vdd tune_shunt_gy[0] a_37444_33400# vdd pmos_6p0 w=1.215u l=0.5u
X7039 a_18032_15748# cap_shunt_p a_16708_15810# vss nmos_6p0 w=0.82u l=0.6u
X7040 a_25572_14964# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7041 a_13588_28700# cap_shunt_n a_13796_28354# vdd pmos_6p0 w=1.2u l=0.5u
X7042 a_3640_4772# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7043 vss cap_shunt_n a_22064_43672# vss nmos_6p0 w=0.82u l=0.6u
X7044 vdd tune_shunt[7] a_10452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X7045 a_21540_20860# cap_shunt_p a_21748_20514# vdd pmos_6p0 w=1.2u l=0.5u
X7046 a_17828_21720# cap_shunt_p a_17620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X7047 vss cap_shunt_p a_25984_36132# vss nmos_6p0 w=0.82u l=0.6u
X7048 a_20532_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7049 vdd a_30028_54120# a_29940_54164# vdd pmos_6p0 w=1.22u l=1u
X7050 a_34328_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7051 a_22680_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7052 a_4380_55688# a_4292_55732# vss vss nmos_6p0 w=0.82u l=1u
X7053 vdd a_21740_47848# a_21652_47892# vdd pmos_6p0 w=1.22u l=1u
X7054 a_25572_11828# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7055 a_24360_12312# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7056 a_13588_34972# cap_shunt_n a_13796_34626# vdd pmos_6p0 w=1.2u l=0.5u
X7057 vss tune_series_gy[4] a_18724_6040# vss nmos_6p0 w=0.51u l=0.6u
X7058 vdd a_14460_11351# a_14372_11448# vdd pmos_6p0 w=1.22u l=1u
X7059 a_36688_21720# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X7060 vss cap_shunt_p a_22064_40536# vss nmos_6p0 w=0.82u l=0.6u
X7061 a_8184_7908# cap_series_gyn a_7768_8316# vss nmos_6p0 w=0.82u l=0.6u
X7062 a_20532_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7063 a_32604_22760# a_32516_22804# vss vss nmos_6p0 w=0.82u l=1u
X7064 vdd a_30028_50984# a_29940_51028# vdd pmos_6p0 w=1.22u l=1u
X7065 a_27496_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X7066 vss cap_shunt_n a_4256_9176# vss nmos_6p0 w=0.82u l=0.6u
X7067 a_30428_19668# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7068 a_13588_31836# cap_shunt_n a_13796_31490# vdd pmos_6p0 w=1.2u l=0.5u
X7069 a_6740_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7070 vdd a_15356_19624# a_15268_19668# vdd pmos_6p0 w=1.22u l=1u
X7071 a_6532_29076# cap_shunt_n a_6740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X7072 a_24652_52119# a_24564_52216# vss vss nmos_6p0 w=0.82u l=1u
X7073 a_11884_50551# a_11796_50648# vss vss nmos_6p0 w=0.82u l=1u
X7074 vdd tune_shunt[7] a_24452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X7075 a_22436_7124# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7076 a_28692_10744# cap_series_gyp a_28484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X7077 vdd a_10540_44712# a_10452_44756# vdd pmos_6p0 w=1.22u l=1u
X7078 a_32156_18056# a_32068_18100# vss vss nmos_6p0 w=0.82u l=1u
X7079 vdd a_27228_19191# a_27140_19288# vdd pmos_6p0 w=1.22u l=1u
X7080 a_32432_20452# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X7081 a_35264_49080# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X7082 vdd tune_shunt[5] a_2500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X7083 a_6740_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7084 a_9668_13396# cap_shunt_p a_9876_13880# vdd pmos_6p0 w=1.2u l=0.5u
X7085 a_9876_48376# cap_shunt_p a_9668_47892# vdd pmos_6p0 w=1.2u l=0.5u
X7086 vss tune_shunt[6] a_25780_34264# vss nmos_6p0 w=0.51u l=0.6u
X7087 a_2708_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7088 a_11780_6040# cap_series_gyn a_11572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X7089 a_15120_12612# cap_shunt_p a_13796_12674# vss nmos_6p0 w=0.82u l=0.6u
X7090 a_15904_50244# cap_shunt_p a_13796_50306# vss nmos_6p0 w=0.82u l=0.6u
X7091 vdd a_32716_16055# a_32628_16152# vdd pmos_6p0 w=1.22u l=1u
X7092 a_7540_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7093 a_18388_3266# cap_series_gyn a_19320_3204# vss nmos_6p0 w=0.82u l=0.6u
X7094 a_32156_14920# a_32068_14964# vss vss nmos_6p0 w=0.82u l=1u
X7095 vdd a_1692_33736# a_1604_33780# vdd pmos_6p0 w=1.22u l=1u
X7096 vss tune_series_gygy[5] a_35880_25940# vss nmos_6p0 w=0.51u l=0.6u
X7097 vss cap_shunt_p a_27104_4472# vss nmos_6p0 w=0.82u l=0.6u
X7098 vdd tune_shunt_gy[1] a_37444_40053# vdd pmos_6p0 w=1.215u l=0.5u
X7099 vdd a_33164_39575# a_33076_39672# vdd pmos_6p0 w=1.22u l=1u
X7100 a_29720_9884# cap_series_gyn a_29532_9884# vdd pmos_6p0 w=1.2u l=0.5u
X7101 a_22436_11828# cap_series_gyn a_22644_12312# vdd pmos_6p0 w=1.2u l=0.5u
X7102 a_9876_18584# cap_shunt_p a_10808_18584# vss nmos_6p0 w=0.82u l=0.6u
X7103 vdd a_31820_49416# a_31732_49460# vdd pmos_6p0 w=1.22u l=1u
X7104 vss tune_shunt[7] a_25780_31128# vss nmos_6p0 w=0.51u l=0.6u
X7105 a_12768_39268# cap_shunt_n a_10660_39330# vss nmos_6p0 w=0.82u l=0.6u
X7106 vdd tune_shunt[5] a_28484_32212# vdd pmos_6p0 w=1.2u l=0.5u
X7107 vdd a_26892_55255# a_26804_55352# vdd pmos_6p0 w=1.22u l=1u
X7108 a_5544_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7109 vdd a_32716_12919# a_32628_13016# vdd pmos_6p0 w=1.22u l=1u
X7110 a_35692_36916# cap_series_gygyp a_35880_36916# vdd pmos_6p0 w=1.2u l=0.5u
X7111 vdd a_36748_32168# a_36660_32212# vdd pmos_6p0 w=1.22u l=1u
X7112 vdd a_1692_30600# a_1604_30644# vdd pmos_6p0 w=1.22u l=1u
X7113 a_15804_11784# a_15716_11828# vss vss nmos_6p0 w=0.82u l=1u
X7114 a_9876_15448# cap_shunt_p a_10808_15448# vss nmos_6p0 w=0.82u l=0.6u
X7115 vdd a_31820_46280# a_31732_46324# vdd pmos_6p0 w=1.22u l=1u
X7116 a_33948_41143# a_33860_41240# vss vss nmos_6p0 w=0.82u l=1u
X7117 a_29700_34626# cap_shunt_p a_29492_34972# vdd pmos_6p0 w=1.2u l=0.5u
X7118 a_21636_6040# cap_series_gyp a_21428_5556# vdd pmos_6p0 w=1.2u l=0.5u
X7119 a_31024_37700# cap_shunt_n a_29700_37762# vss nmos_6p0 w=0.82u l=0.6u
X7120 vdd a_26892_52119# a_26804_52216# vdd pmos_6p0 w=1.22u l=1u
X7121 a_28124_20759# a_28036_20856# vss vss nmos_6p0 w=0.82u l=1u
X7122 a_28484_10260# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7123 a_25572_10260# cap_series_gyn a_25780_10744# vdd pmos_6p0 w=1.2u l=0.5u
X7124 a_35880_14964# cap_series_gygyn a_35692_14964# vdd pmos_6p0 w=1.2u l=0.5u
X7125 a_28692_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7126 a_19388_52552# a_19300_52596# vss vss nmos_6p0 w=0.82u l=1u
X7127 vdd tune_shunt[4] a_20532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X7128 a_35040_44757# cap_shunt_gyp a_35040_45302# vdd pmos_6p0 w=1.215u l=0.5u
X7129 vdd tune_shunt[6] a_3620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X7130 a_29700_31490# cap_shunt_p a_29492_31836# vdd pmos_6p0 w=1.2u l=0.5u
X7131 a_36748_27464# a_36660_27508# vss vss nmos_6p0 w=0.82u l=1u
X7132 a_16708_44034# cap_shunt_p a_18424_43972# vss nmos_6p0 w=0.82u l=0.6u
X7133 a_6508_39575# a_6420_39672# vss vss nmos_6p0 w=0.82u l=1u
X7134 a_9540_12674# cap_shunt_p a_9332_13020# vdd pmos_6p0 w=1.2u l=0.5u
X7135 a_16500_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7136 a_6084_49084# cap_shunt_p a_6292_48738# vdd pmos_6p0 w=1.2u l=0.5u
X7137 a_26768_43972# cap_shunt_p a_24660_44034# vss nmos_6p0 w=0.82u l=0.6u
X7138 vss tune_series_gy[5] a_18612_12674# vss nmos_6p0 w=0.51u l=0.6u
X7139 a_22680_14180# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7140 a_16708_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7141 vss cap_shunt_p a_4816_32996# vss nmos_6p0 w=0.82u l=0.6u
X7142 a_25780_42104# cap_shunt_n a_25572_41620# vdd pmos_6p0 w=1.2u l=0.5u
X7143 a_28692_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7144 a_35880_11828# cap_series_gygyp a_35692_11828# vdd pmos_6p0 w=1.2u l=0.5u
X7145 vss cap_shunt_n a_22064_34264# vss nmos_6p0 w=0.82u l=0.6u
X7146 a_30016_9176# cap_series_gyn a_28692_9176# vss nmos_6p0 w=0.82u l=0.6u
X7147 a_5844_9176# cap_shunt_p a_6776_9176# vss nmos_6p0 w=0.82u l=0.6u
X7148 a_21540_11452# cap_series_gyn a_21748_11106# vdd pmos_6p0 w=1.2u l=0.5u
X7149 vdd a_29692_21192# a_29604_21236# vdd pmos_6p0 w=1.22u l=1u
X7150 a_16708_40898# cap_shunt_n a_18424_40836# vss nmos_6p0 w=0.82u l=0.6u
X7151 a_5844_9176# cap_shunt_p a_5636_8692# vdd pmos_6p0 w=1.2u l=0.5u
X7152 a_26768_40836# cap_shunt_n a_24660_40898# vss nmos_6p0 w=0.82u l=0.6u
X7153 a_20532_24372# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7154 a_22680_11044# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7155 vdd a_12668_52119# a_12580_52216# vdd pmos_6p0 w=1.22u l=1u
X7156 a_10340_25940# cap_shunt_n a_10548_26424# vdd pmos_6p0 w=1.2u l=0.5u
X7157 vdd a_15804_53687# a_15716_53784# vdd pmos_6p0 w=1.22u l=1u
X7158 a_14580_42104# cap_shunt_n a_14372_41620# vdd pmos_6p0 w=1.2u l=0.5u
X7159 a_13588_25564# cap_shunt_n a_13796_25218# vdd pmos_6p0 w=1.2u l=0.5u
X7160 a_36688_12312# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X7161 vss cap_shunt_n a_22064_31128# vss nmos_6p0 w=0.82u l=0.6u
X7162 a_7768_5180# cap_series_gyn a_7580_5180# vdd pmos_6p0 w=1.2u l=0.5u
X7163 a_4492_8215# a_4404_8312# vss vss nmos_6p0 w=0.82u l=1u
X7164 vss tune_shunt[7] a_10660_26786# vss nmos_6p0 w=0.51u l=0.6u
X7165 a_32404_38108# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7166 vdd tune_shunt[6] a_25572_36916# vdd pmos_6p0 w=1.2u l=0.5u
X7167 a_32948_45540# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7168 a_21748_42466# cap_shunt_n a_21540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X7169 a_20532_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7170 a_20740_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7171 vss tune_shunt[6] a_25780_37400# vss nmos_6p0 w=0.51u l=0.6u
X7172 a_1924_7970# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X7173 a_6740_46808# cap_shunt_p a_6532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X7174 a_10340_22804# cap_shunt_n a_10548_23288# vdd pmos_6p0 w=1.2u l=0.5u
X7175 a_13588_22428# cap_shunt_n a_13796_22082# vdd pmos_6p0 w=1.2u l=0.5u
X7176 a_14484_3988# cap_series_gyp a_14692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X7177 a_35292_19624# a_35204_19668# vss vss nmos_6p0 w=0.82u l=1u
X7178 a_15512_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7179 a_26712_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7180 a_8120_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7181 a_34308_5180# cap_series_gygyp a_34516_4834# vdd pmos_6p0 w=1.2u l=0.5u
X7182 a_25572_18100# cap_series_gyn a_25780_18584# vdd pmos_6p0 w=1.2u l=0.5u
X7183 a_34308_23996# cap_series_gygyp a_34516_23650# vdd pmos_6p0 w=1.2u l=0.5u
X7184 a_28692_4472# cap_series_gyp a_29624_4472# vss nmos_6p0 w=0.82u l=0.6u
X7185 vdd a_26556_45847# a_26468_45944# vdd pmos_6p0 w=1.22u l=1u
X7186 vss tune_shunt[6] a_2708_40898# vss nmos_6p0 w=0.51u l=0.6u
X7187 a_26376_9476# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7188 a_1924_4834# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X7189 a_36720_47893# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X7190 a_13588_28700# cap_shunt_n a_13796_28354# vdd pmos_6p0 w=1.2u l=0.5u
X7191 vss tune_shunt[7] a_16708_15810# vss nmos_6p0 w=0.51u l=0.6u
X7192 a_2588_52552# a_2500_52596# vss vss nmos_6p0 w=0.82u l=1u
X7193 a_23308_36872# a_23220_36916# vss vss nmos_6p0 w=0.82u l=1u
X7194 a_15512_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7195 a_6292_17016# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7196 a_22188_55688# a_22100_55732# vss vss nmos_6p0 w=0.82u l=1u
X7197 a_34396_7080# a_34308_7124# vss vss nmos_6p0 w=0.82u l=1u
X7198 a_14112_20152# cap_shunt_p a_12788_20152# vss nmos_6p0 w=0.82u l=0.6u
X7199 vss cap_shunt_n a_23072_32996# vss nmos_6p0 w=0.82u l=0.6u
X7200 a_18612_4472# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7201 a_25780_21720# cap_shunt_p a_26712_21720# vss nmos_6p0 w=0.82u l=0.6u
X7202 a_33524_35348# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7203 vdd a_26892_48983# a_26804_49080# vdd pmos_6p0 w=1.22u l=1u
X7204 a_5544_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7205 a_35692_24372# cap_series_gygyp a_35880_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7206 a_36972_3511# a_36884_3608# vss vss nmos_6p0 w=0.82u l=1u
X7207 a_2724_8692# cap_shunt_n a_2932_9176# vdd pmos_6p0 w=1.2u l=0.5u
X7208 vdd a_26444_54120# a_26356_54164# vdd pmos_6p0 w=1.22u l=1u
X7209 vss cap_shunt_p a_10640_50244# vss nmos_6p0 w=0.82u l=0.6u
X7210 vdd tune_series_gy[5] a_19524_11828# vdd pmos_6p0 w=1.2u l=0.5u
X7211 vdd a_1692_24328# a_1604_24372# vdd pmos_6p0 w=1.22u l=1u
X7212 vss cap_shunt_n a_35840_34264# vss nmos_6p0 w=0.82u l=0.6u
X7213 a_2724_10260# cap_shunt_n a_2932_10744# vdd pmos_6p0 w=1.2u l=0.5u
X7214 vdd tune_shunt[7] a_6420_13020# vdd pmos_6p0 w=1.2u l=0.5u
X7215 vss tune_series_gygy[5] a_35880_16532# vss nmos_6p0 w=0.51u l=0.6u
X7216 a_19152_37400# cap_shunt_n a_17828_37400# vss nmos_6p0 w=0.82u l=0.6u
X7217 a_20740_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7218 a_5544_26424# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7219 vss cap_series_gyp a_16016_7608# vss nmos_6p0 w=0.82u l=0.6u
X7220 vss cap_series_gyp a_25984_4772# vss nmos_6p0 w=0.82u l=0.6u
X7221 a_35692_21236# cap_series_gygyp a_35880_21236# vdd pmos_6p0 w=1.2u l=0.5u
X7222 vdd a_26444_50984# a_26356_51028# vdd pmos_6p0 w=1.22u l=1u
X7223 a_28124_14487# a_28036_14584# vss vss nmos_6p0 w=0.82u l=1u
X7224 vss cap_shunt_n a_15904_20452# vss nmos_6p0 w=0.82u l=0.6u
X7225 vdd a_1692_21192# a_1604_21236# vdd pmos_6p0 w=1.22u l=1u
X7226 vss cap_shunt_n a_35840_31128# vss nmos_6p0 w=0.82u l=0.6u
X7227 a_7336_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7228 vdd a_27676_34871# a_27588_34968# vdd pmos_6p0 w=1.22u l=1u
X7229 a_24660_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7230 a_29700_25218# cap_shunt_p a_29492_25564# vdd pmos_6p0 w=1.2u l=0.5u
X7231 a_14124_54120# a_14036_54164# vss vss nmos_6p0 w=0.82u l=1u
X7232 a_6084_16532# cap_shunt_p a_6292_17016# vdd pmos_6p0 w=1.2u l=0.5u
X7233 a_34396_55255# a_34308_55352# vss vss nmos_6p0 w=0.82u l=1u
X7234 a_5844_9538# cap_shunt_p a_5636_9884# vdd pmos_6p0 w=1.2u l=0.5u
X7235 a_18612_6402# cap_series_gyn a_20328_6340# vss nmos_6p0 w=0.82u l=0.6u
X7236 a_28124_11351# a_28036_11448# vss vss nmos_6p0 w=0.82u l=1u
X7237 a_10864_15748# cap_shunt_p a_9540_15810# vss nmos_6p0 w=0.82u l=0.6u
X7238 a_28692_18584# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7239 a_8568_53380# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7240 a_14896_49944# cap_shunt_n a_12788_49944# vss nmos_6p0 w=0.82u l=0.6u
X7241 a_6292_51512# cap_shunt_p a_8008_51512# vss nmos_6p0 w=0.82u l=0.6u
X7242 vdd a_29132_47848# a_29044_47892# vdd pmos_6p0 w=1.22u l=1u
X7243 a_16708_34626# cap_shunt_n a_18424_34564# vss nmos_6p0 w=0.82u l=0.6u
X7244 a_26768_34564# cap_shunt_p a_24660_34626# vss nmos_6p0 w=0.82u l=0.6u
X7245 vdd a_33500_3511# a_33412_3608# vdd pmos_6p0 w=1.22u l=1u
X7246 a_20496_3204# cap_series_gyn a_18388_3266# vss nmos_6p0 w=0.82u l=0.6u
X7247 a_21748_29922# cap_shunt_n a_21540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X7248 vss cap_shunt_p a_4816_23588# vss nmos_6p0 w=0.82u l=0.6u
X7249 a_22436_11828# cap_series_gyn a_22644_12312# vdd pmos_6p0 w=1.2u l=0.5u
X7250 a_15176_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7251 a_5636_3612# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7252 a_16800_10744# cap_series_gyn a_14692_10744# vss nmos_6p0 w=0.82u l=0.6u
X7253 a_28692_15448# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7254 vss cap_shunt_p a_8400_50244# vss nmos_6p0 w=0.82u l=0.6u
X7255 a_31932_43144# a_31844_43188# vss vss nmos_6p0 w=0.82u l=1u
X7256 a_25780_32696# cap_shunt_p a_25572_32212# vdd pmos_6p0 w=1.2u l=0.5u
X7257 a_1716_6748# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7258 a_13588_19292# cap_shunt_p a_13796_18946# vdd pmos_6p0 w=1.2u l=0.5u
X7259 vdd tune_shunt[6] a_9668_49460# vdd pmos_6p0 w=1.2u l=0.5u
X7260 a_35600_49461# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X7261 a_5844_9538# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X7262 a_14484_10260# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7263 vdd a_29132_44712# a_29044_44756# vdd pmos_6p0 w=1.22u l=1u
X7264 a_16708_31490# cap_shunt_n a_18424_31428# vss nmos_6p0 w=0.82u l=0.6u
X7265 a_34516_4834# tune_series_gygy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X7266 a_21748_36194# cap_shunt_n a_21540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X7267 a_26768_31428# cap_shunt_p a_24660_31490# vss nmos_6p0 w=0.82u l=0.6u
X7268 a_13796_42466# cap_shunt_n a_13588_42812# vdd pmos_6p0 w=1.2u l=0.5u
X7269 a_27496_27992# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7270 a_8848_20152# cap_shunt_p a_6740_20152# vss nmos_6p0 w=0.82u l=0.6u
X7271 a_29700_34626# cap_shunt_p a_29492_34972# vdd pmos_6p0 w=1.2u l=0.5u
X7272 a_10640_48676# cap_shunt_p a_9316_48738# vss nmos_6p0 w=0.82u l=0.6u
X7273 a_6740_15448# cap_shunt_p a_6532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X7274 a_13588_16156# cap_shunt_p a_13796_15810# vdd pmos_6p0 w=1.2u l=0.5u
X7275 a_35600_46325# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X7276 a_9668_52596# cap_shunt_n a_9876_53080# vdd pmos_6p0 w=1.2u l=0.5u
X7277 a_3620_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7278 a_37420_38007# a_37332_38104# vss vss nmos_6p0 w=0.82u l=1u
X7279 vdd tune_shunt[7] a_25572_27508# vdd pmos_6p0 w=1.2u l=0.5u
X7280 vdd tune_shunt[2] a_1716_7124# vdd pmos_6p0 w=1.2u l=0.5u
X7281 a_25572_10260# cap_series_gyn a_25780_10744# vdd pmos_6p0 w=1.2u l=0.5u
X7282 a_9668_52596# cap_shunt_n a_9876_53080# vdd pmos_6p0 w=1.2u l=0.5u
X7283 a_21748_33058# cap_shunt_n a_21540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X7284 a_6956_55255# a_6868_55352# vss vss nmos_6p0 w=0.82u l=1u
X7285 a_27496_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7286 a_29700_31490# cap_shunt_p a_29492_31836# vdd pmos_6p0 w=1.2u l=0.5u
X7287 a_24452_44380# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7288 a_21540_9884# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7289 a_21748_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7290 a_6740_12312# cap_shunt_p a_6532_11828# vdd pmos_6p0 w=1.2u l=0.5u
X7291 a_11800_8692# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7292 vss tune_series_gy[3] a_21524_3266# vss nmos_6p0 w=0.51u l=0.6u
X7293 a_2708_45602# cap_shunt_p a_2500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X7294 a_25780_42104# cap_shunt_n a_25572_41620# vdd pmos_6p0 w=1.2u l=0.5u
X7295 a_33524_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7296 vdd a_14012_5079# a_13924_5176# vdd pmos_6p0 w=1.22u l=1u
X7297 a_36512_41621# cap_shunt_gyn a_36532_42104# vss nmos_6p0 w=0.82u l=0.6u
X7298 a_24452_41244# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7299 a_21540_6748# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7300 a_6740_53080# cap_shunt_n a_8456_53080# vss nmos_6p0 w=0.82u l=0.6u
X7301 a_21748_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7302 vdd a_6956_30167# a_6868_30264# vdd pmos_6p0 w=1.22u l=1u
X7303 vss tune_shunt[7] a_16708_29922# vss nmos_6p0 w=0.51u l=0.6u
X7304 a_25780_12312# cap_series_gyp a_26712_12312# vss nmos_6p0 w=0.82u l=0.6u
X7305 a_11668_43672# cap_shunt_n a_13384_43672# vss nmos_6p0 w=0.82u l=0.6u
X7306 a_10340_25940# cap_shunt_n a_10548_26424# vdd pmos_6p0 w=1.2u l=0.5u
X7307 vss cap_shunt_p a_23072_23588# vss nmos_6p0 w=0.82u l=0.6u
X7308 a_14580_42104# cap_shunt_n a_14372_41620# vdd pmos_6p0 w=1.2u l=0.5u
X7309 a_9204_51874# cap_shunt_n a_10136_51812# vss nmos_6p0 w=0.82u l=0.6u
X7310 a_34516_12674# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7311 a_12376_45540# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7312 vss cap_series_gygyp a_37080_24856# vss nmos_6p0 w=0.82u l=0.6u
X7313 a_31624_22428# cap_series_gygyn a_31648_22020# vss nmos_6p0 w=0.82u l=0.6u
X7314 a_34536_8316# cap_series_gygyp a_35344_7908# vss nmos_6p0 w=0.82u l=0.6u
X7315 a_12788_20152# cap_shunt_p a_12580_19668# vdd pmos_6p0 w=1.2u l=0.5u
X7316 a_6084_50652# cap_shunt_p a_6292_50306# vdd pmos_6p0 w=1.2u l=0.5u
X7317 a_3828_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7318 vss cap_shunt_p a_15904_14180# vss nmos_6p0 w=0.82u l=0.6u
X7319 vdd a_27676_28599# a_27588_28696# vdd pmos_6p0 w=1.22u l=1u
X7320 a_6740_46808# cap_shunt_p a_6532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X7321 a_11668_40536# cap_shunt_n a_13384_40536# vss nmos_6p0 w=0.82u l=0.6u
X7322 a_10340_22804# cap_shunt_n a_10548_23288# vdd pmos_6p0 w=1.2u l=0.5u
X7323 vss tune_shunt[7] a_10548_32696# vss nmos_6p0 w=0.51u l=0.6u
X7324 a_12376_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7325 vdd tune_shunt[7] a_13252_33780# vdd pmos_6p0 w=1.2u l=0.5u
X7326 a_34308_23996# cap_series_gygyp a_34516_23650# vdd pmos_6p0 w=1.2u l=0.5u
X7327 vdd a_22860_53687# a_22772_53784# vdd pmos_6p0 w=1.22u l=1u
X7328 a_3828_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7329 vdd tune_shunt[7] a_3172_16532# vdd pmos_6p0 w=1.2u l=0.5u
X7330 a_17620_46324# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7331 vss cap_series_gyp a_22848_3204# vss nmos_6p0 w=0.82u l=0.6u
X7332 a_24660_17378# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7333 a_30800_4472# cap_series_gyp a_28692_4472# vss nmos_6p0 w=0.82u l=0.6u
X7334 a_36188_50984# a_36100_51028# vss vss nmos_6p0 w=0.82u l=1u
X7335 a_16708_28354# cap_shunt_n a_18424_28292# vss nmos_6p0 w=0.82u l=0.6u
X7336 vdd a_35292_25896# a_35204_25940# vdd pmos_6p0 w=1.22u l=1u
X7337 a_16252_16488# a_16164_16532# vss vss nmos_6p0 w=0.82u l=1u
X7338 vss cap_shunt_p a_19936_45240# vss nmos_6p0 w=0.82u l=0.6u
X7339 a_26768_28292# cap_shunt_n a_24660_28354# vss nmos_6p0 w=0.82u l=0.6u
X7340 vss tune_shunt[6] a_7748_40898# vss nmos_6p0 w=0.51u l=0.6u
X7341 vdd tune_shunt[7] a_13252_30644# vdd pmos_6p0 w=1.2u l=0.5u
X7342 a_22436_8692# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7343 vdd a_11660_53687# a_11572_53784# vdd pmos_6p0 w=1.22u l=1u
X7344 vdd a_22860_50551# a_22772_50648# vdd pmos_6p0 w=1.22u l=1u
X7345 a_15176_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7346 a_34516_4834# cap_series_gygyp a_34308_5180# vdd pmos_6p0 w=1.2u l=0.5u
X7347 a_14012_55255# a_13924_55352# vss vss nmos_6p0 w=0.82u l=1u
X7348 a_14372_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7349 a_22848_32696# cap_shunt_n a_20740_32696# vss nmos_6p0 w=0.82u l=0.6u
X7350 a_16708_25218# cap_shunt_n a_18424_25156# vss nmos_6p0 w=0.82u l=0.6u
X7351 vdd a_35292_22760# a_35204_22804# vdd pmos_6p0 w=1.22u l=1u
X7352 vss tune_series_gy[0] a_29384_3612# vss nmos_6p0 w=0.51u l=0.6u
X7353 a_10452_45948# cap_shunt_n a_10660_45602# vdd pmos_6p0 w=1.2u l=0.5u
X7354 vss cap_shunt_n a_19936_42104# vss nmos_6p0 w=0.82u l=0.6u
X7355 a_13796_36194# cap_shunt_n a_13588_36540# vdd pmos_6p0 w=1.2u l=0.5u
X7356 a_26768_25156# cap_shunt_p a_24660_25218# vss nmos_6p0 w=0.82u l=0.6u
X7357 a_2932_12312# cap_shunt_n a_2724_11828# vdd pmos_6p0 w=1.2u l=0.5u
X7358 a_6628_12674# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7359 vdd tune_shunt[7] a_6420_13020# vdd pmos_6p0 w=1.2u l=0.5u
X7360 a_8064_35832# cap_shunt_n a_6740_35832# vss nmos_6p0 w=0.82u l=0.6u
X7361 a_15176_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7362 a_31436_6748# tune_series_gygy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7363 a_6084_49460# cap_shunt_p a_6292_49944# vdd pmos_6p0 w=1.2u l=0.5u
X7364 vdd tune_shunt[5] a_29492_38108# vdd pmos_6p0 w=1.2u l=0.5u
X7365 a_22644_13880# cap_series_gyn a_22436_13396# vdd pmos_6p0 w=1.2u l=0.5u
X7366 vdd a_2588_55688# a_2500_55732# vdd pmos_6p0 w=1.22u l=1u
X7367 a_10548_32696# cap_shunt_n a_11480_32696# vss nmos_6p0 w=0.82u l=0.6u
X7368 vss cap_shunt_p a_8848_48376# vss nmos_6p0 w=0.82u l=0.6u
X7369 a_30688_45944# cap_shunt_gyn a_30500_45944# vdd pmos_6p0 w=1.215u l=0.5u
X7370 a_13796_33058# cap_shunt_n a_13588_33404# vdd pmos_6p0 w=1.2u l=0.5u
X7371 a_21748_26786# cap_shunt_n a_21540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X7372 a_16500_23996# cap_shunt_n a_16708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X7373 a_27496_18584# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7374 a_29700_25218# cap_shunt_p a_29492_25564# vdd pmos_6p0 w=1.2u l=0.5u
X7375 vdd a_19836_54120# a_19748_54164# vdd pmos_6p0 w=1.22u l=1u
X7376 vdd tune_shunt[7] a_21540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X7377 a_6084_16532# cap_shunt_p a_6292_17016# vdd pmos_6p0 w=1.2u l=0.5u
X7378 vss cap_series_gyn a_30920_9476# vss nmos_6p0 w=0.82u l=0.6u
X7379 vdd a_2140_9783# a_2052_9880# vdd pmos_6p0 w=1.22u l=1u
X7380 a_35180_14487# a_35092_14584# vss vss nmos_6p0 w=0.82u l=1u
X7381 a_27496_15448# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X7382 a_20620_44279# a_20532_44376# vss vss nmos_6p0 w=0.82u l=1u
X7383 a_2708_39330# cap_shunt_n a_2500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X7384 a_31624_6748# tune_series_gygy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X7385 a_23856_7908# cap_series_gyp a_21748_7970# vss nmos_6p0 w=0.82u l=0.6u
X7386 vdd a_30476_54120# a_30388_54164# vdd pmos_6p0 w=1.22u l=1u
X7387 a_36636_52552# a_36548_52596# vss vss nmos_6p0 w=0.82u l=1u
X7388 vdd tune_shunt[7] a_17620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X7389 vdd a_9420_53687# a_9332_53784# vdd pmos_6p0 w=1.22u l=1u
X7390 vdd a_19836_50984# a_19748_51028# vdd pmos_6p0 w=1.22u l=1u
X7391 a_36160_43734# cap_shunt_gyn a_36160_43189# vdd pmos_6p0 w=1.215u l=0.5u
X7392 a_21748_14242# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7393 a_21180_54120# a_21092_54164# vss vss nmos_6p0 w=0.82u l=1u
X7394 vdd a_2140_18056# a_2052_18100# vdd pmos_6p0 w=1.22u l=1u
X7395 vdd a_19388_49416# a_19300_49460# vdd pmos_6p0 w=1.22u l=1u
X7396 a_16028_21192# a_15940_21236# vss vss nmos_6p0 w=0.82u l=1u
X7397 a_20620_41143# a_20532_41240# vss vss nmos_6p0 w=0.82u l=1u
X7398 a_25780_32696# cap_shunt_p a_25572_32212# vdd pmos_6p0 w=1.2u l=0.5u
X7399 vss cap_series_gyp a_13888_4472# vss nmos_6p0 w=0.82u l=0.6u
X7400 a_35180_11351# a_35092_11448# vss vss nmos_6p0 w=0.82u l=1u
X7401 vdd a_30476_50984# a_30388_51028# vdd pmos_6p0 w=1.22u l=1u
X7402 a_2708_9538# cap_shunt_n a_3640_9476# vss nmos_6p0 w=0.82u l=0.6u
X7403 vss cap_series_gygyn a_37080_18584# vss nmos_6p0 w=0.82u l=0.6u
X7404 a_27788_55255# a_27700_55352# vss vss nmos_6p0 w=0.82u l=1u
X7405 vss tune_shunt[7] a_10548_35832# vss nmos_6p0 w=0.51u l=0.6u
X7406 vdd tune_shunt[7] a_17620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X7407 a_34144_44376# cap_shunt_gyp a_34144_43972# vdd pmos_6p0 w=1.215u l=0.5u
X7408 a_29492_30268# cap_shunt_p a_29700_29922# vdd pmos_6p0 w=1.2u l=0.5u
X7409 a_22436_7124# cap_series_gyp a_22644_7608# vdd pmos_6p0 w=1.2u l=0.5u
X7410 a_21748_11106# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7411 vdd a_10540_55255# a_10452_55352# vdd pmos_6p0 w=1.22u l=1u
X7412 a_13796_42466# cap_shunt_n a_13588_42812# vdd pmos_6p0 w=1.2u l=0.5u
X7413 a_35880_22804# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7414 a_25780_7608# cap_series_gyn a_25572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X7415 vss tune_series_gy[5] a_24660_12674# vss nmos_6p0 w=0.51u l=0.6u
X7416 a_15700_7970# cap_series_gyn a_17416_7908# vss nmos_6p0 w=0.82u l=0.6u
X7417 a_15700_7970# cap_series_gyn a_15492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X7418 vss cap_series_gyn a_24752_13880# vss nmos_6p0 w=0.82u l=0.6u
X7419 a_22644_9176# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7420 vss cap_series_gygyn a_37080_15448# vss nmos_6p0 w=0.82u l=0.6u
X7421 a_14236_52552# a_14148_52596# vss vss nmos_6p0 w=0.82u l=1u
X7422 a_12376_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7423 a_25572_10260# cap_series_gyn a_25780_10744# vdd pmos_6p0 w=1.2u l=0.5u
X7424 a_17620_18100# cap_shunt_p a_17828_18584# vdd pmos_6p0 w=1.2u l=0.5u
X7425 a_10988_44712# a_10900_44756# vss vss nmos_6p0 w=0.82u l=1u
X7426 a_30408_35832# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7427 vdd a_27676_19191# a_27588_19288# vdd pmos_6p0 w=1.22u l=1u
X7428 a_6644_53788# cap_shunt_n a_6852_53442# vdd pmos_6p0 w=1.2u l=0.5u
X7429 a_25572_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7430 a_13588_20860# cap_shunt_n a_13796_20514# vdd pmos_6p0 w=1.2u l=0.5u
X7431 vss tune_shunt[7] a_10548_23288# vss nmos_6p0 w=0.51u l=0.6u
X7432 vss cap_series_gyp a_24752_10744# vss nmos_6p0 w=0.82u l=0.6u
X7433 a_13720_13880# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7434 vdd tune_shunt[7] a_13252_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7435 a_32612_37762# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X7436 a_2708_45602# cap_shunt_p a_2500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X7437 a_10988_41576# a_10900_41620# vss vss nmos_6p0 w=0.82u l=1u
X7438 vdd a_1692_41143# a_1604_41240# vdd pmos_6p0 w=1.22u l=1u
X7439 a_25572_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7440 vdd a_35292_16488# a_35204_16532# vdd pmos_6p0 w=1.22u l=1u
X7441 a_10452_39676# cap_shunt_n a_10660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X7442 a_24660_33058# cap_shunt_p a_25592_32996# vss nmos_6p0 w=0.82u l=0.6u
X7443 a_13588_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7444 vdd tune_shunt[7] a_13252_21236# vdd pmos_6p0 w=1.2u l=0.5u
X7445 a_32612_34626# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7446 a_33936_32996# cap_shunt_n a_32612_33058# vss nmos_6p0 w=0.82u l=0.6u
X7447 a_8064_29560# cap_shunt_n a_6740_29560# vss nmos_6p0 w=0.82u l=0.6u
X7448 a_9668_51028# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7449 vdd a_5948_11784# a_5860_11828# vdd pmos_6p0 w=1.22u l=1u
X7450 vdd a_2588_49416# a_2500_49460# vdd pmos_6p0 w=1.22u l=1u
X7451 a_4816_37700# cap_shunt_n a_2708_37762# vss nmos_6p0 w=0.82u l=0.6u
X7452 a_22848_23288# cap_shunt_p a_20740_23288# vss nmos_6p0 w=0.82u l=0.6u
X7453 a_2500_23996# cap_shunt_p a_2708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X7454 a_1924_6040# cap_shunt_p a_2856_6040# vss nmos_6p0 w=0.82u l=0.6u
X7455 a_12788_20152# cap_shunt_p a_12580_19668# vdd pmos_6p0 w=1.2u l=0.5u
X7456 vdd a_8300_55255# a_8212_55352# vdd pmos_6p0 w=1.22u l=1u
X7457 a_6084_50652# cap_shunt_p a_6292_50306# vdd pmos_6p0 w=1.2u l=0.5u
X7458 a_29492_38108# cap_shunt_n a_29700_37762# vdd pmos_6p0 w=1.2u l=0.5u
X7459 vdd tune_series_gy[5] a_25572_13396# vdd pmos_6p0 w=1.2u l=0.5u
X7460 a_13796_26786# cap_shunt_n a_13588_27132# vdd pmos_6p0 w=1.2u l=0.5u
X7461 a_20060_55688# a_19972_55732# vss vss nmos_6p0 w=0.82u l=1u
X7462 vss tune_series_gy[5] a_15720_11452# vss nmos_6p0 w=0.51u l=0.6u
X7463 a_10660_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7464 a_8064_26424# cap_shunt_n a_6740_26424# vss nmos_6p0 w=0.82u l=0.6u
X7465 a_28572_20759# a_28484_20856# vss vss nmos_6p0 w=0.82u l=1u
X7466 vdd a_32604_42711# a_32516_42808# vdd pmos_6p0 w=1.22u l=1u
X7467 a_6760_3988# cap_series_gyp a_6572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X7468 a_8860_3511# a_8772_3608# vss vss nmos_6p0 w=0.82u l=1u
X7469 vdd a_2588_46280# a_2500_46324# vdd pmos_6p0 w=1.22u l=1u
X7470 a_35692_25940# cap_series_gygyp a_35880_25940# vdd pmos_6p0 w=1.2u l=0.5u
X7471 a_10548_23288# cap_shunt_n a_11480_23288# vss nmos_6p0 w=0.82u l=0.6u
X7472 a_8736_14180# cap_shunt_p a_6628_14242# vss nmos_6p0 w=0.82u l=0.6u
X7473 a_37632_33400# cap_shunt_gyp a_37652_32996# vss nmos_6p0 w=0.82u l=0.6u
X7474 a_32612_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7475 vss tune_series_gy[3] a_14692_6040# vss nmos_6p0 w=0.51u l=0.6u
X7476 a_16500_14588# cap_shunt_p a_16708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X7477 a_6956_39575# a_6868_39672# vss vss nmos_6p0 w=0.82u l=1u
X7478 vss cap_shunt_n a_9856_29860# vss nmos_6p0 w=0.82u l=0.6u
X7479 vss cap_shunt_p a_3248_4472# vss nmos_6p0 w=0.82u l=0.6u
X7480 a_28484_8692# cap_series_gyn a_28692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X7481 a_5844_11106# cap_shunt_n a_5636_11452# vdd pmos_6p0 w=1.2u l=0.5u
X7482 vdd a_18044_7080# a_17956_7124# vdd pmos_6p0 w=1.22u l=1u
X7483 a_10660_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7484 a_18404_9884# cap_series_gyp a_18612_9538# vdd pmos_6p0 w=1.2u l=0.5u
X7485 vdd tune_series_gy[5] a_21540_14588# vdd pmos_6p0 w=1.2u l=0.5u
X7486 a_33500_25896# a_33412_25940# vss vss nmos_6p0 w=0.82u l=1u
X7487 vdd a_19276_23895# a_19188_23992# vdd pmos_6p0 w=1.22u l=1u
X7488 a_35692_22804# cap_series_gygyp a_35880_22804# vdd pmos_6p0 w=1.2u l=0.5u
X7489 a_5488_49944# cap_shunt_p a_3380_49944# vss nmos_6p0 w=0.82u l=0.6u
X7490 a_20620_34871# a_20532_34968# vss vss nmos_6p0 w=0.82u l=1u
X7491 vss cap_shunt_n a_9856_26724# vss nmos_6p0 w=0.82u l=0.6u
X7492 a_28484_5556# cap_shunt_n a_28692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X7493 vdd a_24204_14920# a_24116_14964# vdd pmos_6p0 w=1.22u l=1u
X7494 a_11460_44756# cap_shunt_n a_11668_45240# vdd pmos_6p0 w=1.2u l=0.5u
X7495 a_27788_48983# a_27700_49080# vss vss nmos_6p0 w=0.82u l=1u
X7496 a_16708_45602# cap_shunt_p a_16500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X7497 vdd tune_shunt[7] a_17620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7498 a_18404_6748# cap_series_gyn a_18612_6402# vdd pmos_6p0 w=1.2u l=0.5u
X7499 vss cap_series_gyp a_19936_7908# vss nmos_6p0 w=0.82u l=0.6u
X7500 a_10452_45948# cap_shunt_n a_10660_45602# vdd pmos_6p0 w=1.2u l=0.5u
X7501 vss tune_shunt[7] a_10548_29560# vss nmos_6p0 w=0.51u l=0.6u
X7502 vdd a_19276_20759# a_19188_20856# vdd pmos_6p0 w=1.22u l=1u
X7503 a_20532_40052# cap_shunt_p a_20740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X7504 vss tune_shunt[5] a_28692_32696# vss nmos_6p0 w=0.51u l=0.6u
X7505 a_13796_36194# cap_shunt_n a_13588_36540# vdd pmos_6p0 w=1.2u l=0.5u
X7506 a_11480_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7507 a_20620_31735# a_20532_31832# vss vss nmos_6p0 w=0.82u l=1u
X7508 a_22456_3204# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X7509 a_28484_13396# cap_series_gyp a_28692_13880# vdd pmos_6p0 w=1.2u l=0.5u
X7510 vss cap_shunt_p a_10752_20452# vss nmos_6p0 w=0.82u l=0.6u
X7511 vdd a_13788_52552# a_13700_52596# vdd pmos_6p0 w=1.22u l=1u
X7512 a_6084_49460# cap_shunt_p a_6292_49944# vdd pmos_6p0 w=1.2u l=0.5u
X7513 a_2588_38440# a_2500_38484# vss vss nmos_6p0 w=0.82u l=1u
X7514 a_22644_13880# cap_series_gyn a_22436_13396# vdd pmos_6p0 w=1.2u l=0.5u
X7515 a_30016_27992# cap_shunt_p a_28692_27992# vss nmos_6p0 w=0.82u l=0.6u
X7516 vdd tune_shunt[7] a_17620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X7517 a_20172_30167# a_20084_30264# vss vss nmos_6p0 w=0.82u l=1u
X7518 a_30408_29560# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7519 vss tune_shunt[7] a_10548_26424# vss nmos_6p0 w=0.51u l=0.6u
X7520 a_8008_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7521 vss tune_shunt[6] a_7748_37762# vss nmos_6p0 w=0.51u l=0.6u
X7522 vdd a_28460_3511# a_28372_3608# vdd pmos_6p0 w=1.22u l=1u
X7523 a_34396_3511# a_34308_3608# vss vss nmos_6p0 w=0.82u l=1u
X7524 a_13796_33058# cap_shunt_n a_13588_33404# vdd pmos_6p0 w=1.2u l=0.5u
X7525 a_11480_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7526 a_10660_23650# cap_shunt_n a_10452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X7527 vss cap_series_gyp a_12768_4772# vss nmos_6p0 w=0.82u l=0.6u
X7528 a_24660_17378# cap_series_gyp a_24452_17724# vdd pmos_6p0 w=1.2u l=0.5u
X7529 a_30016_24856# cap_shunt_p a_28692_24856# vss nmos_6p0 w=0.82u l=0.6u
X7530 a_20172_27031# a_20084_27128# vss vss nmos_6p0 w=0.82u l=1u
X7531 a_30408_26424# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7532 a_10660_6402# cap_series_gyn a_10452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X7533 a_12580_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7534 a_23756_36872# a_23668_36916# vss vss nmos_6p0 w=0.82u l=1u
X7535 vss tune_shunt[7] a_7748_34626# vss nmos_6p0 w=0.51u l=0.6u
X7536 a_2708_39330# cap_shunt_n a_2500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X7537 a_25572_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7538 vdd tune_series_gy[3] a_24452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X7539 a_37280_51029# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X7540 vss cap_shunt_gyp a_35868_48376# vss nmos_6p0 w=0.82u l=0.6u
X7541 a_16184_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7542 a_31624_22428# cap_series_gygyn a_31436_22428# vdd pmos_6p0 w=1.2u l=0.5u
X7543 a_3620_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7544 a_13588_39676# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7545 vdd tune_series_gy[4] a_14484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X7546 vdd a_26892_54120# a_26804_54164# vdd pmos_6p0 w=1.22u l=1u
X7547 a_32612_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7548 a_10472_12612# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7549 vdd a_19052_50551# a_18964_50648# vdd pmos_6p0 w=1.22u l=1u
X7550 vdd tune_shunt[6] a_20532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X7551 a_22064_38968# cap_shunt_n a_20740_38968# vss nmos_6p0 w=0.82u l=0.6u
X7552 a_29492_30268# cap_shunt_p a_29700_29922# vdd pmos_6p0 w=1.2u l=0.5u
X7553 a_24660_23650# cap_shunt_p a_25592_23588# vss nmos_6p0 w=0.82u l=0.6u
X7554 vss cap_shunt_n a_15904_43672# vss nmos_6p0 w=0.82u l=0.6u
X7555 a_31708_3944# a_31620_3988# vss vss nmos_6p0 w=0.82u l=1u
X7556 a_2500_9884# cap_shunt_n a_2708_9538# vdd pmos_6p0 w=1.2u l=0.5u
X7557 vdd a_26892_50984# a_26804_51028# vdd pmos_6p0 w=1.22u l=1u
X7558 a_32612_25218# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7559 a_1924_3266# cap_shunt_n a_1716_3612# vdd pmos_6p0 w=1.2u l=0.5u
X7560 a_28572_14487# a_28484_14584# vss vss nmos_6p0 w=0.82u l=1u
X7561 a_33948_54120# a_33860_54164# vss vss nmos_6p0 w=0.82u l=1u
X7562 vdd tune_shunt[7] a_29492_28700# vdd pmos_6p0 w=1.2u l=0.5u
X7563 a_30528_9476# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7564 vdd a_23868_54120# a_23780_54164# vdd pmos_6p0 w=1.22u l=1u
X7565 a_5936_48376# cap_shunt_p a_3828_48376# vss nmos_6p0 w=0.82u l=0.6u
X7566 a_13796_45602# cap_shunt_p a_14728_45540# vss nmos_6p0 w=0.82u l=0.6u
X7567 a_18612_11106# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7568 a_2708_20514# cap_shunt_p a_4424_20452# vss nmos_6p0 w=0.82u l=0.6u
X7569 a_34480_47893# cap_shunt_gyp a_34480_48438# vdd pmos_6p0 w=1.215u l=0.5u
X7570 a_34720_36132# cap_shunt_n a_32612_36194# vss nmos_6p0 w=0.82u l=0.6u
X7571 a_1924_6402# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X7572 a_2500_14588# cap_shunt_n a_2708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X7573 vdd tune_shunt[6] a_7540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X7574 a_14572_54120# a_14484_54164# vss vss nmos_6p0 w=0.82u l=1u
X7575 vss cap_shunt_n a_15904_40536# vss nmos_6p0 w=0.82u l=0.6u
X7576 a_37080_21720# cap_series_gygyp a_35880_21236# vss nmos_6p0 w=0.82u l=0.6u
X7577 a_6644_53788# cap_shunt_n a_6852_53442# vdd pmos_6p0 w=1.2u l=0.5u
X7578 a_10660_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7579 a_28572_11351# a_28484_11448# vss vss nmos_6p0 w=0.82u l=1u
X7580 a_21540_44380# cap_shunt_n a_21748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X7581 vdd a_23868_50984# a_23780_51028# vdd pmos_6p0 w=1.22u l=1u
X7582 a_13796_42466# cap_shunt_n a_14728_42404# vss nmos_6p0 w=0.82u l=0.6u
X7583 a_35692_16532# cap_series_gygyn a_35880_16532# vdd pmos_6p0 w=1.2u l=0.5u
X7584 a_18032_43972# cap_shunt_p a_16708_44034# vss nmos_6p0 w=0.82u l=0.6u
X7585 a_24452_34972# cap_shunt_p a_24660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X7586 a_16708_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7587 vdd a_29580_47848# a_29492_47892# vdd pmos_6p0 w=1.22u l=1u
X7588 vdd tune_shunt[6] a_7540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X7589 a_20620_28599# a_20532_28696# vss vss nmos_6p0 w=0.82u l=1u
X7590 a_16708_39330# cap_shunt_n a_16500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X7591 a_10660_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7592 a_26712_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X7593 a_21540_41244# cap_shunt_p a_21748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X7594 a_10452_39676# cap_shunt_n a_10660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X7595 vdd a_19276_14487# a_19188_14584# vdd pmos_6p0 w=1.22u l=1u
X7596 a_2708_48738# cap_shunt_p a_3640_48676# vss nmos_6p0 w=0.82u l=0.6u
X7597 a_33500_16488# a_33412_16532# vss vss nmos_6p0 w=0.82u l=1u
X7598 a_18032_40836# cap_shunt_n a_16708_40898# vss nmos_6p0 w=0.82u l=0.6u
X7599 a_24452_31836# cap_shunt_p a_24660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X7600 vss tune_shunt[7] a_6740_21720# vss nmos_6p0 w=0.51u l=0.6u
X7601 vdd a_29580_44712# a_29492_44756# vdd pmos_6p0 w=1.22u l=1u
X7602 a_20620_25463# a_20532_25560# vss vss nmos_6p0 w=0.82u l=1u
X7603 vss tune_shunt[4] a_28692_23288# vss nmos_6p0 w=0.51u l=0.6u
X7604 a_13796_26786# cap_shunt_n a_13588_27132# vdd pmos_6p0 w=1.2u l=0.5u
X7605 a_6532_25940# cap_shunt_n a_6740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X7606 a_35880_21236# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7607 vss tune_series_gy[4] a_18612_4472# vss nmos_6p0 w=0.51u l=0.6u
X7608 vdd tune_shunt[7] a_13588_23996# vdd pmos_6p0 w=1.2u l=0.5u
X7609 vdd a_15356_47848# a_15268_47892# vdd pmos_6p0 w=1.22u l=1u
X7610 a_6740_38968# cap_shunt_n a_8456_38968# vss nmos_6p0 w=0.82u l=0.6u
X7611 a_35692_8692# cap_series_gygyn a_35880_8692# vdd pmos_6p0 w=1.2u l=0.5u
X7612 a_31624_19292# cap_series_gygyn a_31436_19292# vdd pmos_6p0 w=1.2u l=0.5u
X7613 a_10548_34264# cap_shunt_n a_10340_33780# vdd pmos_6p0 w=1.2u l=0.5u
X7614 a_30016_18584# cap_series_gyp a_28692_18584# vss nmos_6p0 w=0.82u l=0.6u
X7615 vss tune_shunt[7] a_2708_15810# vss nmos_6p0 w=0.51u l=0.6u
X7616 a_21540_17724# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7617 a_29468_52119# a_29380_52216# vss vss nmos_6p0 w=0.82u l=1u
X7618 vss tune_shunt[7] a_7748_28354# vss nmos_6p0 w=0.51u l=0.6u
X7619 a_6532_22804# cap_shunt_p a_6740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X7620 a_3172_18100# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7621 a_1692_47415# a_1604_47512# vss vss nmos_6p0 w=0.82u l=1u
X7622 a_35692_5556# cap_series_gygyn a_35880_5556# vdd pmos_6p0 w=1.2u l=0.5u
X7623 a_10548_31128# cap_shunt_n a_10340_30644# vdd pmos_6p0 w=1.2u l=0.5u
X7624 a_1716_3988# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7625 a_30016_15448# cap_series_gyn a_28692_15448# vss nmos_6p0 w=0.82u l=0.6u
X7626 a_13452_55688# a_13364_55732# vss vss nmos_6p0 w=0.82u l=1u
X7627 a_30408_17016# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7628 a_20172_17623# a_20084_17720# vss vss nmos_6p0 w=0.82u l=1u
X7629 vss tune_shunt[7] a_7748_25218# vss nmos_6p0 w=0.51u l=0.6u
X7630 a_11460_44756# cap_shunt_n a_11668_45240# vdd pmos_6p0 w=1.2u l=0.5u
X7631 vdd a_35740_41143# a_35652_41240# vdd pmos_6p0 w=1.22u l=1u
X7632 a_3828_40536# cap_shunt_n a_3620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X7633 a_13252_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7634 a_10452_45948# cap_shunt_n a_10660_45602# vdd pmos_6p0 w=1.2u l=0.5u
X7635 vdd a_27228_44279# a_27140_44376# vdd pmos_6p0 w=1.22u l=1u
X7636 a_3620_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7637 a_6292_51512# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7638 a_36076_36439# a_35988_36536# vss vss nmos_6p0 w=0.82u l=1u
X7639 a_34308_23996# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7640 vdd tune_series_gygy[4] a_34308_13020# vdd pmos_6p0 w=1.2u l=0.5u
X7641 vdd a_33500_8648# a_33412_8692# vdd pmos_6p0 w=1.22u l=1u
X7642 a_2708_14242# cap_shunt_n a_4424_14180# vss nmos_6p0 w=0.82u l=0.6u
X7643 a_29720_16156# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7644 a_10428_55688# a_10340_55732# vss vss nmos_6p0 w=0.82u l=1u
X7645 vdd tune_shunt[7] a_20532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X7646 a_32156_40008# a_32068_40052# vss vss nmos_6p0 w=0.82u l=1u
X7647 vss cap_shunt_n a_18032_22020# vss nmos_6p0 w=0.82u l=0.6u
X7648 vdd a_31260_14920# a_31172_14964# vdd pmos_6p0 w=1.22u l=1u
X7649 a_2140_12919# a_2052_13016# vss vss nmos_6p0 w=0.82u l=1u
X7650 vss cap_shunt_gyp a_37548_51512# vss nmos_6p0 w=0.82u l=0.6u
X7651 a_27340_49416# a_27252_49460# vss vss nmos_6p0 w=0.82u l=1u
X7652 a_10660_23650# cap_shunt_n a_10452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X7653 a_26376_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7654 vdd a_33500_5512# a_33412_5556# vdd pmos_6p0 w=1.22u l=1u
X7655 a_13796_36194# cap_shunt_n a_14728_36132# vss nmos_6p0 w=0.82u l=0.6u
X7656 a_2708_11106# cap_shunt_n a_4424_11044# vss nmos_6p0 w=0.82u l=0.6u
X7657 a_24660_17378# cap_series_gyp a_24452_17724# vdd pmos_6p0 w=1.2u l=0.5u
X7658 a_19544_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X7659 vdd a_31260_11784# a_31172_11828# vdd pmos_6p0 w=1.22u l=1u
X7660 a_29916_53687# a_29828_53784# vss vss nmos_6p0 w=0.82u l=1u
X7661 a_27340_46280# a_27252_46324# vss vss nmos_6p0 w=0.82u l=1u
X7662 a_37080_12312# cap_series_gygyp a_35880_11828# vss nmos_6p0 w=0.82u l=0.6u
X7663 a_24316_49416# a_24228_49460# vss vss nmos_6p0 w=0.82u l=1u
X7664 vss cap_series_gygyn a_31816_21720# vss nmos_6p0 w=0.82u l=0.6u
X7665 vdd tune_series_gy[3] a_10492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X7666 a_1716_5556# cap_shunt_p a_1924_6040# vdd pmos_6p0 w=1.2u l=0.5u
X7667 a_14460_55255# a_14372_55352# vss vss nmos_6p0 w=0.82u l=1u
X7668 a_18032_34564# cap_shunt_n a_16708_34626# vss nmos_6p0 w=0.82u l=0.6u
X7669 vss cap_shunt_n a_12768_43972# vss nmos_6p0 w=0.82u l=0.6u
X7670 a_24452_25564# cap_shunt_p a_24660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X7671 a_9540_15810# cap_shunt_p a_9332_16156# vdd pmos_6p0 w=1.2u l=0.5u
X7672 vdd tune_shunt[5] a_3172_51028# vdd pmos_6p0 w=1.2u l=0.5u
X7673 a_29916_50551# a_29828_50648# vss vss nmos_6p0 w=0.82u l=1u
X7674 a_25572_33780# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7675 a_12788_49944# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7676 a_17828_40536# cap_shunt_n a_17620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X7677 a_29384_3612# tune_series_gy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X7678 a_2708_39330# cap_shunt_n a_3640_39268# vss nmos_6p0 w=0.82u l=0.6u
X7679 a_29492_30268# cap_shunt_p a_29700_29922# vdd pmos_6p0 w=1.2u l=0.5u
X7680 a_18032_31428# cap_shunt_n a_16708_31490# vss nmos_6p0 w=0.82u l=0.6u
X7681 a_18760_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7682 a_11436_55255# a_11348_55352# vss vss nmos_6p0 w=0.82u l=1u
X7683 vss cap_shunt_n a_12768_40836# vss nmos_6p0 w=0.82u l=0.6u
X7684 a_24452_22428# cap_shunt_p a_24660_22082# vdd pmos_6p0 w=1.2u l=0.5u
X7685 a_25592_9476# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7686 vss tune_shunt[7] a_6740_12312# vss nmos_6p0 w=0.51u l=0.6u
X7687 a_36636_38440# a_36548_38484# vss vss nmos_6p0 w=0.82u l=1u
X7688 a_14692_10744# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7689 a_25572_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7690 a_18612_4472# cap_series_gyp a_18404_3988# vdd pmos_6p0 w=1.2u l=0.5u
X7691 vss tune_shunt[6] a_6740_35832# vss nmos_6p0 w=0.51u l=0.6u
X7692 a_24660_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7693 a_29468_45847# a_29380_45944# vss vss nmos_6p0 w=0.82u l=1u
X7694 a_18760_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7695 vss cap_series_gyp a_27888_6040# vss nmos_6p0 w=0.82u l=0.6u
X7696 a_35880_11828# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7697 vss cap_shunt_n a_15568_27992# vss nmos_6p0 w=0.82u l=0.6u
X7698 a_13588_50652# cap_shunt_p a_13796_50306# vdd pmos_6p0 w=1.2u l=0.5u
X7699 vdd tune_shunt[7] a_13588_14588# vdd pmos_6p0 w=1.2u l=0.5u
X7700 a_10548_24856# cap_shunt_n a_10340_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7701 a_12788_15448# cap_shunt_p a_12580_14964# vdd pmos_6p0 w=1.2u l=0.5u
X7702 a_24660_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7703 a_31036_41576# a_30948_41620# vss vss nmos_6p0 w=0.82u l=1u
X7704 a_24452_34972# cap_shunt_p a_24660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X7705 a_29468_42711# a_29380_42808# vss vss nmos_6p0 w=0.82u l=1u
X7706 a_7748_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7707 a_6308_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7708 a_10452_39676# cap_shunt_n a_10660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X7709 vss cap_shunt_n a_15568_24856# vss nmos_6p0 w=0.82u l=0.6u
X7710 a_16476_21192# a_16388_21236# vss vss nmos_6p0 w=0.82u l=1u
X7711 a_8008_49944# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7712 a_2500_47516# cap_shunt_p a_2708_47170# vdd pmos_6p0 w=1.2u l=0.5u
X7713 a_6740_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7714 a_12788_12312# cap_shunt_p a_12580_11828# vdd pmos_6p0 w=1.2u l=0.5u
X7715 a_24452_31836# cap_shunt_p a_24660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X7716 vss tune_series_gy[5] a_28692_13880# vss nmos_6p0 w=0.51u l=0.6u
X7717 a_32156_33736# a_32068_33780# vss vss nmos_6p0 w=0.82u l=1u
X7718 a_8960_53380# cap_shunt_n a_6852_53442# vss nmos_6p0 w=0.82u l=0.6u
X7719 vss cap_shunt_gyp a_37548_45240# vss nmos_6p0 w=0.82u l=0.6u
X7720 a_6740_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7721 vdd a_21292_55688# a_21204_55732# vdd pmos_6p0 w=1.22u l=1u
X7722 a_14684_52552# a_14596_52596# vss vss nmos_6p0 w=0.82u l=1u
X7723 a_25592_37700# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7724 a_17416_6340# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X7725 a_10452_5180# cap_series_gyp a_10660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X7726 a_2708_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7727 vss tune_series_gy[4] a_28692_10744# vss nmos_6p0 w=0.51u l=0.6u
X7728 a_17596_13352# a_17508_13396# vss vss nmos_6p0 w=0.82u l=1u
X7729 vss cap_shunt_p a_14112_20152# vss nmos_6p0 w=0.82u l=0.6u
X7730 a_1716_6748# cap_shunt_n a_1924_6402# vdd pmos_6p0 w=1.2u l=0.5u
X7731 a_22456_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7732 a_32156_30600# a_32068_30644# vss vss nmos_6p0 w=0.82u l=1u
X7733 a_25572_3988# cap_shunt_p a_25780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X7734 a_17620_36916# cap_shunt_n a_17828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X7735 vss tune_shunt[7] a_20740_27992# vss nmos_6p0 w=0.51u l=0.6u
X7736 a_3172_18100# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7737 vss tune_shunt[7] a_6404_22082# vss nmos_6p0 w=0.51u l=0.6u
X7738 a_21748_9538# cap_series_gyp a_21540_9884# vdd pmos_6p0 w=1.2u l=0.5u
X7739 a_17596_10216# a_17508_10260# vss vss nmos_6p0 w=0.82u l=1u
X7740 a_18032_28292# cap_shunt_n a_16708_28354# vss nmos_6p0 w=0.82u l=0.6u
X7741 a_2500_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7742 a_24452_19292# cap_series_gyn a_24660_18946# vdd pmos_6p0 w=1.2u l=0.5u
X7743 a_13252_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7744 vss cap_shunt_p a_34720_29860# vss nmos_6p0 w=0.82u l=0.6u
X7745 vss tune_shunt[5] a_20740_24856# vss nmos_6p0 w=0.51u l=0.6u
X7746 vdd a_5388_5512# a_5300_5556# vdd pmos_6p0 w=1.22u l=1u
X7747 a_21748_6402# cap_series_gyn a_21540_6748# vdd pmos_6p0 w=1.2u l=0.5u
X7748 a_18032_25156# cap_shunt_n a_16708_25218# vss nmos_6p0 w=0.82u l=0.6u
X7749 a_24452_16156# cap_series_gyn a_24660_15810# vdd pmos_6p0 w=1.2u l=0.5u
X7750 a_35532_48676# cap_shunt_gyn a_35264_48676# vss nmos_6p0 w=0.82u l=0.6u
X7751 a_2708_34626# cap_shunt_n a_2500_34972# vdd pmos_6p0 w=1.2u l=0.5u
X7752 vss cap_shunt_n a_12768_34564# vss nmos_6p0 w=0.82u l=0.6u
X7753 vdd a_31708_25896# a_31620_25940# vdd pmos_6p0 w=1.22u l=1u
X7754 a_32380_3511# a_32292_3608# vss vss nmos_6p0 w=0.82u l=1u
X7755 a_15512_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7756 a_25572_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7757 a_35692_8692# cap_series_gygyn a_35880_8692# vdd pmos_6p0 w=1.2u l=0.5u
X7758 vdd tune_shunt[3] a_5636_11452# vdd pmos_6p0 w=1.2u l=0.5u
X7759 vss tune_shunt[7] a_6740_29560# vss nmos_6p0 w=0.51u l=0.6u
X7760 vss cap_shunt_p a_34720_26724# vss nmos_6p0 w=0.82u l=0.6u
X7761 vdd a_25100_53687# a_25012_53784# vdd pmos_6p0 w=1.22u l=1u
X7762 a_34348_8316# cap_series_gygyp a_34536_8316# vdd pmos_6p0 w=1.2u l=0.5u
X7763 vss cap_series_gyp a_24752_7608# vss nmos_6p0 w=0.82u l=0.6u
X7764 a_18760_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7765 vss cap_shunt_n a_12768_31428# vss nmos_6p0 w=0.82u l=0.6u
X7766 a_35880_22804# cap_series_gygyp a_35904_23288# vss nmos_6p0 w=0.82u l=0.6u
X7767 vdd a_31708_22760# a_31620_22804# vdd pmos_6p0 w=1.22u l=1u
X7768 a_28692_40536# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7769 a_2708_31490# cap_shunt_p a_2500_31836# vdd pmos_6p0 w=1.2u l=0.5u
X7770 a_15512_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7771 a_35692_5556# cap_series_gygyn a_35880_5556# vdd pmos_6p0 w=1.2u l=0.5u
X7772 a_25572_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7773 a_35308_45240# cap_shunt_gyp a_35040_45302# vss nmos_6p0 w=0.82u l=0.6u
X7774 a_13588_44380# cap_shunt_n a_13796_44034# vdd pmos_6p0 w=1.2u l=0.5u
X7775 vss tune_shunt[7] a_6740_26424# vss nmos_6p0 w=0.51u l=0.6u
X7776 vdd a_2140_8648# a_2052_8692# vdd pmos_6p0 w=1.22u l=1u
X7777 a_24660_14242# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7778 a_9668_18100# cap_shunt_p a_9876_18584# vdd pmos_6p0 w=1.2u l=0.5u
X7779 vdd a_25100_50551# a_25012_50648# vdd pmos_6p0 w=1.22u l=1u
X7780 a_11984_32996# cap_shunt_n a_10660_33058# vss nmos_6p0 w=0.82u l=0.6u
X7781 a_9668_18100# cap_shunt_p a_9876_18584# vdd pmos_6p0 w=1.2u l=0.5u
X7782 a_20532_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7783 a_18760_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7784 a_31820_54120# a_31732_54164# vss vss nmos_6p0 w=0.82u l=1u
X7785 vss tune_shunt[3] a_32612_37762# vss nmos_6p0 w=0.51u l=0.6u
X7786 vss cap_shunt_p a_31024_39268# vss nmos_6p0 w=0.82u l=0.6u
X7787 vss cap_series_gygyn a_35840_18884# vss nmos_6p0 w=0.82u l=0.6u
X7788 a_13588_41244# cap_shunt_n a_13796_40898# vdd pmos_6p0 w=1.2u l=0.5u
X7789 a_6628_14242# cap_shunt_p a_6420_14588# vdd pmos_6p0 w=1.2u l=0.5u
X7790 vss cap_series_gyn a_26768_6340# vss nmos_6p0 w=0.82u l=0.6u
X7791 a_24660_11106# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7792 a_15532_11452# cap_series_gyp a_15720_11452# vdd pmos_6p0 w=1.2u l=0.5u
X7793 vdd a_24652_14920# a_24564_14964# vdd pmos_6p0 w=1.22u l=1u
X7794 vss tune_shunt[6] a_10660_42466# vss nmos_6p0 w=0.51u l=0.6u
X7795 a_24452_25564# cap_shunt_p a_24660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X7796 a_15532_11452# cap_series_gyp a_15720_11452# vdd pmos_6p0 w=1.2u l=0.5u
X7797 a_20740_37400# cap_shunt_n a_22456_37400# vss nmos_6p0 w=0.82u l=0.6u
X7798 vss tune_series_gy[2] a_14468_3266# vss nmos_6p0 w=0.51u l=0.6u
X7799 vss tune_shunt[5] a_32612_34626# vss nmos_6p0 w=0.51u l=0.6u
X7800 vdd a_10540_54120# a_10452_54164# vdd pmos_6p0 w=1.22u l=1u
X7801 a_24660_7970# cap_series_gyp a_24452_8316# vdd pmos_6p0 w=1.2u l=0.5u
X7802 vss cap_series_gygyn a_35840_15748# vss nmos_6p0 w=0.82u l=0.6u
X7803 a_2500_38108# cap_shunt_n a_2708_37762# vdd pmos_6p0 w=1.2u l=0.5u
X7804 vdd a_36524_14487# a_36436_14584# vdd pmos_6p0 w=1.22u l=1u
X7805 a_31372_49416# a_31284_49460# vss vss nmos_6p0 w=0.82u l=1u
X7806 vss cap_shunt_p a_26768_3204# vss nmos_6p0 w=0.82u l=0.6u
X7807 a_24452_22428# cap_shunt_p a_24660_22082# vdd pmos_6p0 w=1.2u l=0.5u
X7808 a_19732_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7809 a_33524_32212# cap_shunt_n a_33732_32696# vdd pmos_6p0 w=1.2u l=0.5u
X7810 a_2708_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7811 a_15120_22020# cap_shunt_n a_13796_22082# vss nmos_6p0 w=0.82u l=0.6u
X7812 vss tune_shunt[0] a_29700_4834# vss nmos_6p0 w=0.51u l=0.6u
X7813 a_12788_48376# cap_shunt_p a_12580_47892# vdd pmos_6p0 w=1.2u l=0.5u
X7814 vdd tune_series_gy[3] a_24452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X7815 a_2932_10744# cap_shunt_n a_4648_10744# vss nmos_6p0 w=0.82u l=0.6u
X7816 vdd a_36524_11351# a_36436_11448# vdd pmos_6p0 w=1.22u l=1u
X7817 a_6628_12674# cap_shunt_p a_7560_12612# vss nmos_6p0 w=0.82u l=0.6u
X7818 a_18816_20452# cap_shunt_p a_16708_20514# vss nmos_6p0 w=0.82u l=0.6u
X7819 a_33948_53687# a_33860_53784# vss vss nmos_6p0 w=0.82u l=1u
X7820 a_21516_47415# a_21428_47512# vss vss nmos_6p0 w=0.82u l=1u
X7821 a_31372_46280# a_31284_46324# vss vss nmos_6p0 w=0.82u l=1u
X7822 a_21672_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7823 a_9204_51874# cap_shunt_n a_8996_52220# vdd pmos_6p0 w=1.2u l=0.5u
X7824 a_19732_10744# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7825 a_17828_46808# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7826 a_5544_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7827 a_7768_8316# cap_series_gyn a_7580_8316# vdd pmos_6p0 w=1.2u l=0.5u
X7828 vdd a_29244_19624# a_29156_19668# vdd pmos_6p0 w=1.22u l=1u
X7829 a_24452_34972# cap_shunt_p a_24660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X7830 a_30408_9176# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X7831 vdd a_1692_40008# a_1604_40052# vdd pmos_6p0 w=1.22u l=1u
X7832 a_33948_50551# a_33860_50648# vss vss nmos_6p0 w=0.82u l=1u
X7833 vdd a_10092_46280# a_10004_46324# vdd pmos_6p0 w=1.22u l=1u
X7834 vss cap_shunt_n a_11872_32696# vss nmos_6p0 w=0.82u l=0.6u
X7835 a_9876_51512# cap_shunt_n a_9668_51028# vdd pmos_6p0 w=1.2u l=0.5u
X7836 a_17620_27508# cap_shunt_n a_17828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X7837 vss tune_shunt[7] a_20740_18584# vss nmos_6p0 w=0.51u l=0.6u
X7838 a_9532_3511# a_9444_3608# vss vss nmos_6p0 w=0.82u l=1u
X7839 a_5544_42104# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7840 a_24452_31836# cap_shunt_p a_24660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X7841 vss cap_shunt_n a_12768_28292# vss nmos_6p0 w=0.82u l=0.6u
X7842 a_2500_14588# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7843 a_27340_52119# a_27252_52216# vss vss nmos_6p0 w=0.82u l=1u
X7844 vss cap_shunt_p a_30800_27992# vss nmos_6p0 w=0.82u l=0.6u
X7845 a_35880_24372# cap_series_gygyp a_35692_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7846 a_24660_42466# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7847 a_6060_38007# a_5972_38104# vss vss nmos_6p0 w=0.82u l=1u
X7848 vss tune_shunt[5] a_3380_49944# vss nmos_6p0 w=0.51u l=0.6u
X7849 vss tune_series_gy[5] a_20740_15448# vss nmos_6p0 w=0.51u l=0.6u
X7850 a_11144_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7851 a_14484_3988# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7852 vss tune_shunt[6] a_20740_38968# vss nmos_6p0 w=0.51u l=0.6u
X7853 vss cap_shunt_n a_12768_25156# vss nmos_6p0 w=0.82u l=0.6u
X7854 vdd a_31708_16488# a_31620_16532# vdd pmos_6p0 w=1.22u l=1u
X7855 a_2708_25218# cap_shunt_p a_2500_25564# vdd pmos_6p0 w=1.2u l=0.5u
X7856 vss cap_shunt_p a_30800_24856# vss nmos_6p0 w=0.82u l=0.6u
X7857 vss cap_series_gyp a_30016_4472# vss nmos_6p0 w=0.82u l=0.6u
X7858 a_23072_7908# cap_series_gyp a_21748_7970# vss nmos_6p0 w=0.82u l=0.6u
X7859 a_35880_21236# cap_series_gygyp a_35692_21236# vdd pmos_6p0 w=1.2u l=0.5u
X7860 a_28692_34264# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7861 a_33164_23895# a_33076_23992# vss vss nmos_6p0 w=0.82u l=1u
X7862 a_16708_17378# cap_shunt_p a_16500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X7863 vss tune_shunt[6] a_3828_46808# vss nmos_6p0 w=0.51u l=0.6u
X7864 a_36748_33736# a_36660_33780# vss vss nmos_6p0 w=0.82u l=1u
X7865 a_20532_19668# cap_shunt_p a_20740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X7866 a_1692_32168# a_1604_32212# vss vss nmos_6p0 w=0.82u l=1u
X7867 a_21636_6040# cap_series_gyp a_23352_6040# vss nmos_6p0 w=0.82u l=0.6u
X7868 a_31820_47848# a_31732_47892# vss vss nmos_6p0 w=0.82u l=1u
X7869 a_2708_22082# cap_shunt_p a_2500_22428# vdd pmos_6p0 w=1.2u l=0.5u
X7870 a_5844_9538# cap_shunt_p a_7560_9476# vss nmos_6p0 w=0.82u l=0.6u
X7871 a_24660_37762# cap_shunt_p a_24452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X7872 a_6740_34264# cap_shunt_n a_6532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X7873 a_28692_31128# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7874 a_2932_10744# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X7875 a_15512_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7876 vdd a_32156_36872# a_32068_36916# vdd pmos_6p0 w=1.22u l=1u
X7877 a_36748_30600# a_36660_30644# vss vss nmos_6p0 w=0.82u l=1u
X7878 vss tune_shunt[7] a_10660_36194# vss nmos_6p0 w=0.51u l=0.6u
X7879 vss cap_shunt_n a_8064_35832# vss nmos_6p0 w=0.82u l=0.6u
X7880 a_11984_23588# cap_shunt_n a_10660_23650# vss nmos_6p0 w=0.82u l=0.6u
X7881 a_24452_19292# cap_series_gyn a_24660_18946# vdd pmos_6p0 w=1.2u l=0.5u
X7882 vdd a_29916_20759# a_29828_20856# vdd pmos_6p0 w=1.22u l=1u
X7883 a_27496_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7884 vdd a_6508_34871# a_6420_34968# vdd pmos_6p0 w=1.22u l=1u
X7885 vss cap_shunt_n a_18816_37700# vss nmos_6p0 w=0.82u l=0.6u
X7886 vdd tune_shunt[6] a_28484_36916# vdd pmos_6p0 w=1.2u l=0.5u
X7887 a_6532_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7888 a_3828_32696# cap_shunt_p a_5544_32696# vss nmos_6p0 w=0.82u l=0.6u
X7889 a_10340_32212# cap_shunt_n a_10548_32696# vdd pmos_6p0 w=1.2u l=0.5u
X7890 vss tune_shunt[7] a_32612_28354# vss nmos_6p0 w=0.51u l=0.6u
X7891 a_15700_7970# cap_series_gyn a_16632_7908# vss nmos_6p0 w=0.82u l=0.6u
X7892 a_6740_31128# cap_shunt_n a_6532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X7893 a_20740_26424# cap_shunt_n a_20532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X7894 a_18404_11452# cap_series_gyn a_18612_11106# vdd pmos_6p0 w=1.2u l=0.5u
X7895 a_30800_35832# cap_shunt_p a_28692_35832# vss nmos_6p0 w=0.82u l=0.6u
X7896 a_11668_46808# cap_shunt_n a_11460_46324# vdd pmos_6p0 w=1.2u l=0.5u
X7897 vss tune_shunt[7] a_10660_33058# vss nmos_6p0 w=0.51u l=0.6u
X7898 a_6196_22428# cap_shunt_p a_6404_22082# vdd pmos_6p0 w=1.2u l=0.5u
X7899 a_24452_16156# cap_series_gyn a_24660_15810# vdd pmos_6p0 w=1.2u l=0.5u
X7900 a_16296_43672# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7901 a_27496_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7902 a_6532_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7903 a_3828_46808# cap_shunt_p a_4760_46808# vss nmos_6p0 w=0.82u l=0.6u
X7904 vss tune_shunt[4] a_32612_25218# vss nmos_6p0 w=0.51u l=0.6u
X7905 a_19524_7124# cap_series_gyp a_19732_7608# vdd pmos_6p0 w=1.2u l=0.5u
X7906 vss tune_shunt[5] a_6292_18946# vss nmos_6p0 w=0.51u l=0.6u
X7907 a_21672_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7908 a_20740_23288# cap_shunt_p a_20532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X7909 a_18816_14180# cap_shunt_p a_16708_14242# vss nmos_6p0 w=0.82u l=0.6u
X7910 a_13588_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7911 a_29532_13020# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7912 vdd a_15356_55255# a_15268_55352# vdd pmos_6p0 w=1.22u l=1u
X7913 a_9540_11106# cap_shunt_p a_9332_11452# vdd pmos_6p0 w=1.2u l=0.5u
X7914 a_16296_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7915 a_16364_12919# a_16276_13016# vss vss nmos_6p0 w=0.82u l=1u
X7916 a_8008_51812# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7917 vdd a_16924_25896# a_16836_25940# vdd pmos_6p0 w=1.22u l=1u
X7918 a_21672_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7919 vss tune_shunt[6] a_16708_45602# vss nmos_6p0 w=0.51u l=0.6u
X7920 a_13588_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X7921 vss tune_shunt[7] a_21748_18946# vss nmos_6p0 w=0.51u l=0.6u
X7922 vdd a_15356_52119# a_15268_52216# vdd pmos_6p0 w=1.22u l=1u
X7923 a_20284_50984# a_20196_51028# vss vss nmos_6p0 w=0.82u l=1u
X7924 vss tune_series_gygy[5] a_31624_22428# vss nmos_6p0 w=0.51u l=0.6u
X7925 vdd a_32604_38440# a_32516_38484# vdd pmos_6p0 w=1.22u l=1u
X7926 a_21748_29922# cap_shunt_n a_23464_29860# vss nmos_6p0 w=0.82u l=0.6u
X7927 a_29700_37762# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7928 a_24452_25564# cap_shunt_p a_24660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X7929 vdd a_16924_22760# a_16836_22804# vdd pmos_6p0 w=1.22u l=1u
X7930 a_13796_12674# cap_shunt_p a_13588_13020# vdd pmos_6p0 w=1.2u l=0.5u
X7931 vdd a_27676_44279# a_27588_44376# vdd pmos_6p0 w=1.22u l=1u
X7932 vdd a_16028_52552# a_15940_52596# vdd pmos_6p0 w=1.22u l=1u
X7933 a_24660_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7934 a_28692_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7935 vss cap_shunt_n a_11872_23288# vss nmos_6p0 w=0.82u l=0.6u
X7936 a_6740_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X7937 a_10876_55688# a_10788_55732# vss vss nmos_6p0 w=0.82u l=1u
X7938 a_2140_35304# a_2052_35348# vss vss nmos_6p0 w=0.82u l=1u
X7939 vdd a_32604_35304# a_32516_35348# vdd pmos_6p0 w=1.22u l=1u
X7940 a_21748_26786# cap_shunt_n a_23464_26724# vss nmos_6p0 w=0.82u l=0.6u
X7941 vss tune_series_gy[2] a_7768_6748# vss nmos_6p0 w=0.51u l=0.6u
X7942 a_29720_16156# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X7943 a_29700_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7944 a_24452_22428# cap_shunt_p a_24660_22082# vdd pmos_6p0 w=1.2u l=0.5u
X7945 a_2708_18946# cap_shunt_p a_2500_19292# vdd pmos_6p0 w=1.2u l=0.5u
X7946 vss cap_series_gyp a_30800_18584# vss nmos_6p0 w=0.82u l=0.6u
X7947 a_6292_48738# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X7948 a_24316_45847# a_24228_45944# vss vss nmos_6p0 w=0.82u l=1u
X7949 a_24660_33058# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X7950 a_25780_4472# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X7951 vdd a_27900_55688# a_27812_55732# vdd pmos_6p0 w=1.22u l=1u
X7952 a_10452_34972# cap_shunt_n a_10660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X7953 vdd tune_series_gy[3] a_21316_3988# vdd pmos_6p0 w=1.2u l=0.5u
X7954 a_12788_48376# cap_shunt_p a_12580_47892# vdd pmos_6p0 w=1.2u l=0.5u
X7955 a_4032_20452# cap_shunt_p a_2708_20514# vss nmos_6p0 w=0.82u l=0.6u
X7956 a_5276_52552# a_5188_52596# vss vss nmos_6p0 w=0.82u l=1u
X7957 a_11592_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7958 a_2708_15810# cap_shunt_p a_2500_16156# vdd pmos_6p0 w=1.2u l=0.5u
X7959 a_7748_34626# cap_shunt_n a_7540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X7960 vss cap_series_gyn a_30800_15448# vss nmos_6p0 w=0.82u l=0.6u
X7961 a_35904_37400# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X7962 a_10452_31836# cap_shunt_n a_10660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X7963 vss cap_shunt_n a_8064_29560# vss nmos_6p0 w=0.82u l=0.6u
X7964 vdd a_29132_54120# a_29044_54164# vdd pmos_6p0 w=1.22u l=1u
X7965 a_1692_22760# a_1604_22804# vss vss nmos_6p0 w=0.82u l=1u
X7966 a_34844_13352# a_34756_13396# vss vss nmos_6p0 w=0.82u l=1u
X7967 a_4760_13880# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X7968 a_24764_49416# a_24676_49460# vss vss nmos_6p0 w=0.82u l=1u
X7969 vss tune_shunt[5] a_6292_17378# vss nmos_6p0 w=0.51u l=0.6u
X7970 vdd a_6508_28599# a_6420_28696# vdd pmos_6p0 w=1.22u l=1u
X7971 vss tune_series_gy[4] a_21748_6402# vss nmos_6p0 w=0.51u l=0.6u
X7972 a_11592_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7973 a_7748_31490# cap_shunt_n a_7540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X7974 a_20732_52552# a_20644_52596# vss vss nmos_6p0 w=0.82u l=1u
X7975 a_30800_29560# cap_shunt_p a_28692_29560# vss nmos_6p0 w=0.82u l=0.6u
X7976 vdd a_32156_27464# a_32068_27508# vdd pmos_6p0 w=1.22u l=1u
X7977 a_6740_24856# cap_shunt_p a_6532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X7978 vss cap_shunt_n a_8064_26424# vss nmos_6p0 w=0.82u l=0.6u
X7979 vdd a_29132_50984# a_29044_51028# vdd pmos_6p0 w=1.22u l=1u
X7980 a_34844_10216# a_34756_10260# vss vss nmos_6p0 w=0.82u l=1u
X7981 a_27496_34264# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7982 vdd tune_shunt[7] a_28484_27508# vdd pmos_6p0 w=1.2u l=0.5u
X7983 vss cap_shunt_p a_26768_20452# vss nmos_6p0 w=0.82u l=0.6u
X7984 vdd tune_shunt[6] a_13588_47516# vdd pmos_6p0 w=1.2u l=0.5u
X7985 a_3828_23288# cap_shunt_p a_5544_23288# vss nmos_6p0 w=0.82u l=0.6u
X7986 a_11884_55255# a_11796_55352# vss vss nmos_6p0 w=0.82u l=1u
X7987 a_33500_50984# a_33412_51028# vss vss nmos_6p0 w=0.82u l=1u
X7988 a_2500_28700# cap_shunt_n a_2708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X7989 a_30800_26424# cap_shunt_p a_28692_26424# vss nmos_6p0 w=0.82u l=0.6u
X7990 a_20740_17016# cap_shunt_p a_20532_16532# vdd pmos_6p0 w=1.2u l=0.5u
X7991 a_6740_21720# cap_shunt_p a_6532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X7992 a_13460_21720# cap_shunt_n a_15176_21720# vss nmos_6p0 w=0.82u l=0.6u
X7993 a_3828_20152# cap_shunt_p a_3620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X7994 a_28692_15448# cap_series_gyn a_28484_14964# vdd pmos_6p0 w=1.2u l=0.5u
X7995 a_10660_37762# cap_shunt_n a_10452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X7996 vdd a_14460_5079# a_14372_5176# vdd pmos_6p0 w=1.22u l=1u
X7997 a_27496_31128# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X7998 a_9428_18946# cap_shunt_p a_10360_18884# vss nmos_6p0 w=0.82u l=0.6u
X7999 a_15400_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8000 a_25780_13880# cap_series_gyn a_27496_13880# vss nmos_6p0 w=0.82u l=0.6u
X8001 a_9668_10260# cap_shunt_p a_9876_10744# vdd pmos_6p0 w=1.2u l=0.5u
X8002 vdd tune_shunt[6] a_14372_41620# vdd pmos_6p0 w=1.2u l=0.5u
X8003 vss tune_shunt[6] a_25780_38968# vss nmos_6p0 w=0.51u l=0.6u
X8004 a_7540_38108# cap_shunt_n a_7748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X8005 a_13588_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8006 vss tune_shunt[6] a_16708_39330# vss nmos_6p0 w=0.51u l=0.6u
X8007 vss tune_shunt[7] a_24660_31490# vss nmos_6p0 w=0.51u l=0.6u
X8008 a_12444_10216# a_12356_10260# vss vss nmos_6p0 w=0.82u l=1u
X8009 a_28692_12312# cap_series_gyn a_28484_11828# vdd pmos_6p0 w=1.2u l=0.5u
X8010 a_31484_41576# a_31396_41620# vss vss nmos_6p0 w=0.82u l=1u
X8011 a_24660_37762# cap_shunt_p a_24452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X8012 a_9876_48376# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8013 a_34516_22082# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8014 a_25780_10744# cap_series_gyn a_27496_10744# vss nmos_6p0 w=0.82u l=0.6u
X8015 vdd a_35740_40008# a_35652_40052# vdd pmos_6p0 w=1.22u l=1u
X8016 a_13252_25940# cap_shunt_n a_13460_26424# vdd pmos_6p0 w=1.2u l=0.5u
X8017 a_24452_19292# cap_series_gyn a_24660_18946# vdd pmos_6p0 w=1.2u l=0.5u
X8018 a_3620_25940# cap_shunt_p a_3828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X8019 a_13588_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8020 a_21672_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8021 vdd tune_shunt[6] a_28484_36916# vdd pmos_6p0 w=1.2u l=0.5u
X8022 a_6292_17378# cap_shunt_p a_8008_17316# vss nmos_6p0 w=0.82u l=0.6u
X8023 a_10340_32212# cap_shunt_n a_10548_32696# vdd pmos_6p0 w=1.2u l=0.5u
X8024 a_24660_42466# cap_shunt_n a_24452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X8025 vss tune_shunt[7] a_10660_23650# vss nmos_6p0 w=0.51u l=0.6u
X8026 a_18404_11452# cap_series_gyn a_18612_11106# vdd pmos_6p0 w=1.2u l=0.5u
X8027 vdd tune_shunt[5] a_6532_52596# vdd pmos_6p0 w=1.2u l=0.5u
X8028 a_11668_46808# cap_shunt_n a_11460_46324# vdd pmos_6p0 w=1.2u l=0.5u
X8029 a_2140_29032# a_2052_29076# vss vss nmos_6p0 w=0.82u l=1u
X8030 vdd a_32604_29032# a_32516_29076# vdd pmos_6p0 w=1.22u l=1u
X8031 a_13252_22804# cap_shunt_n a_13460_23288# vdd pmos_6p0 w=1.2u l=0.5u
X8032 a_24452_16156# cap_series_gyn a_24660_15810# vdd pmos_6p0 w=1.2u l=0.5u
X8033 a_35600_48438# cap_shunt_gyp a_35600_47893# vdd pmos_6p0 w=1.215u l=0.5u
X8034 a_29700_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8035 a_33732_27992# cap_shunt_p a_33524_27508# vdd pmos_6p0 w=1.2u l=0.5u
X8036 a_3620_22804# cap_shunt_p a_3828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X8037 vss cap_shunt_p a_15120_12612# vss nmos_6p0 w=0.82u l=0.6u
X8038 a_9644_55255# a_9556_55352# vss vss nmos_6p0 w=0.82u l=1u
X8039 a_35692_3988# cap_series_gygyp a_35880_3988# vdd pmos_6p0 w=1.2u l=0.5u
X8040 a_6740_12312# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8041 a_4032_14180# cap_shunt_n a_2708_14242# vss nmos_6p0 w=0.82u l=0.6u
X8042 a_28484_14964# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8043 a_25572_14964# cap_series_gyp a_25780_15448# vdd pmos_6p0 w=1.2u l=0.5u
X8044 vss tune_shunt[6] a_11668_43672# vss nmos_6p0 w=0.51u l=0.6u
X8045 a_2140_25896# a_2052_25940# vss vss nmos_6p0 w=0.82u l=1u
X8046 a_29700_4834# cap_shunt_p a_29492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X8047 a_29700_4834# cap_shunt_p a_31416_4772# vss nmos_6p0 w=0.82u l=0.6u
X8048 a_29532_13020# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8049 a_21748_17378# cap_shunt_p a_23464_17316# vss nmos_6p0 w=0.82u l=0.6u
X8050 a_29700_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8051 a_17640_22020# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8052 a_19732_7608# cap_series_gyp a_21448_7608# vss nmos_6p0 w=0.82u l=0.6u
X8053 a_9540_11106# cap_shunt_p a_9332_11452# vdd pmos_6p0 w=1.2u l=0.5u
X8054 a_17828_20152# cap_shunt_p a_17620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X8055 vdd tune_shunt[7] a_21540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X8056 vdd a_16700_49416# a_16612_49460# vdd pmos_6p0 w=1.22u l=1u
X8057 a_10452_25564# cap_shunt_n a_10660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X8058 vdd tune_series_gygy[5] a_34308_22428# vdd pmos_6p0 w=1.2u l=0.5u
X8059 vss tune_series_gy[0] a_29384_3612# vss nmos_6p0 w=0.51u l=0.6u
X8060 a_22680_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8061 a_4032_11044# cap_shunt_n a_2708_11106# vss nmos_6p0 w=0.82u l=0.6u
X8062 a_28484_11828# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8063 a_25572_11828# cap_series_gyp a_25780_12312# vdd pmos_6p0 w=1.2u l=0.5u
X8064 vss tune_shunt[6] a_11668_40536# vss nmos_6p0 w=0.51u l=0.6u
X8065 a_22644_12312# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8066 vss tune_shunt[7] a_6404_22082# vss nmos_6p0 w=0.51u l=0.6u
X8067 a_19388_54120# a_19300_54164# vss vss nmos_6p0 w=0.82u l=1u
X8068 a_8064_45240# cap_shunt_p a_6740_45240# vss nmos_6p0 w=0.82u l=0.6u
X8069 vss cap_shunt_n a_22064_38968# vss nmos_6p0 w=0.82u l=0.6u
X8070 a_7748_25218# cap_shunt_n a_7540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X8071 a_3932_52119# a_3844_52216# vss vss nmos_6p0 w=0.82u l=1u
X8072 a_35880_3988# tune_series_gygy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X8073 a_22680_15748# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8074 a_13796_12674# cap_shunt_p a_13588_13020# vdd pmos_6p0 w=1.2u l=0.5u
X8075 a_3380_18584# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8076 vss cap_series_gyn a_26768_14180# vss nmos_6p0 w=0.82u l=0.6u
X8077 a_8064_42104# cap_shunt_n a_6740_42104# vss nmos_6p0 w=0.82u l=0.6u
X8078 a_11884_48983# a_11796_49080# vss vss nmos_6p0 w=0.82u l=1u
X8079 a_13460_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8080 vdd a_15804_18056# a_15716_18100# vdd pmos_6p0 w=1.22u l=1u
X8081 a_2708_48738# cap_shunt_p a_2500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X8082 vss cap_shunt_p a_9856_45540# vss nmos_6p0 w=0.82u l=0.6u
X8083 a_16500_30268# cap_shunt_n a_16708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X8084 a_7748_28354# cap_shunt_n a_7540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X8085 a_31624_6748# tune_series_gygy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X8086 a_1716_3988# cap_shunt_p a_1924_4472# vdd pmos_6p0 w=1.2u l=0.5u
X8087 a_32432_18884# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X8088 vdd a_24204_33736# a_24116_33780# vdd pmos_6p0 w=1.22u l=1u
X8089 a_35292_24328# a_35204_24372# vss vss nmos_6p0 w=0.82u l=1u
X8090 a_12580_13396# cap_shunt_p a_12788_13880# vdd pmos_6p0 w=1.2u l=0.5u
X8091 vdd tune_shunt[7] a_13588_38108# vdd pmos_6p0 w=1.2u l=0.5u
X8092 a_7768_6748# cap_series_gyp a_7580_6748# vdd pmos_6p0 w=1.2u l=0.5u
X8093 vss cap_series_gyp a_26768_11044# vss nmos_6p0 w=0.82u l=0.6u
X8094 a_34480_48438# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8095 a_16708_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8096 vdd tune_shunt[7] a_21540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X8097 a_33500_41576# a_33412_41620# vss vss nmos_6p0 w=0.82u l=1u
X8098 a_34516_12674# cap_series_gygyp a_35448_12612# vss nmos_6p0 w=0.82u l=0.6u
X8099 a_30800_17016# cap_series_gyn a_28692_17016# vss nmos_6p0 w=0.82u l=0.6u
X8100 a_13588_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8101 a_15904_48676# cap_shunt_n a_13796_48738# vss nmos_6p0 w=0.82u l=0.6u
X8102 vss cap_shunt_n a_9856_42404# vss nmos_6p0 w=0.82u l=0.6u
X8103 vdd a_24204_30600# a_24116_30644# vdd pmos_6p0 w=1.22u l=1u
X8104 a_15512_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8105 vdd tune_shunt_gy[1] a_37444_38485# vdd pmos_6p0 w=1.215u l=0.5u
X8106 vdd tune_shunt[6] a_17620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X8107 a_20740_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8108 a_13588_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8109 a_9072_43972# cap_shunt_p a_7748_44034# vss nmos_6p0 w=0.82u l=0.6u
X8110 a_34480_46870# cap_shunt_gyn a_34480_46325# vdd pmos_6p0 w=1.215u l=0.5u
X8111 a_3828_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8112 vss tune_shunt[7] a_24660_22082# vss nmos_6p0 w=0.51u l=0.6u
X8113 vss tune_shunt[7] a_9540_12674# vss nmos_6p0 w=0.51u l=0.6u
X8114 vdd a_28124_38007# a_28036_38104# vdd pmos_6p0 w=1.22u l=1u
X8115 a_24660_36194# cap_shunt_p a_24452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X8116 a_2588_54120# a_2500_54164# vss vss nmos_6p0 w=0.82u l=1u
X8117 a_32612_34626# cap_shunt_n a_32404_34972# vdd pmos_6p0 w=1.2u l=0.5u
X8118 a_6404_22082# cap_shunt_p a_8120_22020# vss nmos_6p0 w=0.82u l=0.6u
X8119 vss cap_shunt_p a_11200_13880# vss nmos_6p0 w=0.82u l=0.6u
X8120 a_20740_24856# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8121 vss cap_shunt_n a_4816_9476# vss nmos_6p0 w=0.82u l=0.6u
X8122 a_20172_45847# a_20084_45944# vss vss nmos_6p0 w=0.82u l=1u
X8123 a_21540_42812# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8124 a_18268_55688# a_18180_55732# vss vss nmos_6p0 w=0.82u l=1u
X8125 a_9072_40836# cap_shunt_n a_7748_40898# vss nmos_6p0 w=0.82u l=0.6u
X8126 vss tune_series_gy[2] a_10660_4834# vss nmos_6p0 w=0.51u l=0.6u
X8127 a_28348_19624# a_28260_19668# vss vss nmos_6p0 w=0.82u l=1u
X8128 vdd tune_shunt[7] a_28484_27508# vdd pmos_6p0 w=1.2u l=0.5u
X8129 a_24660_33058# cap_shunt_p a_24452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X8130 vdd a_36748_27464# a_36660_27508# vdd pmos_6p0 w=1.22u l=1u
X8131 a_28124_19191# a_28036_19288# vss vss nmos_6p0 w=0.82u l=1u
X8132 vdd tune_series_gygy[5] a_34308_19292# vdd pmos_6p0 w=1.2u l=0.5u
X8133 a_6404_47170# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8134 a_2500_28700# cap_shunt_n a_2708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X8135 a_3828_43672# cap_shunt_p a_3620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X8136 a_11872_37400# cap_shunt_n a_10548_37400# vss nmos_6p0 w=0.82u l=0.6u
X8137 a_32612_31490# cap_shunt_n a_32404_31836# vdd pmos_6p0 w=1.2u l=0.5u
X8138 a_2724_11828# cap_shunt_n a_2932_12312# vdd pmos_6p0 w=1.2u l=0.5u
X8139 vdd tune_shunt[6] a_6532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X8140 a_30016_40536# cap_shunt_p a_28692_40536# vss nmos_6p0 w=0.82u l=0.6u
X8141 vss cap_shunt_p a_11200_10744# vss nmos_6p0 w=0.82u l=0.6u
X8142 a_20172_42711# a_20084_42808# vss vss nmos_6p0 w=0.82u l=1u
X8143 a_10660_37762# cap_shunt_n a_10452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X8144 vdd tune_series_gy[2] a_7580_8316# vdd pmos_6p0 w=1.2u l=0.5u
X8145 a_28484_8692# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8146 a_9220_17724# cap_shunt_p a_9428_17378# vdd pmos_6p0 w=1.2u l=0.5u
X8147 a_21964_47415# a_21876_47512# vss vss nmos_6p0 w=0.82u l=1u
X8148 a_31060_44757# cap_shunt_gyn a_31248_44757# vdd pmos_6p0 w=1.215u l=0.5u
X8149 a_36296_23288# cap_series_gygyp a_35880_22804# vss nmos_6p0 w=0.82u l=0.6u
X8150 vdd a_32156_8648# a_32068_8692# vdd pmos_6p0 w=1.22u l=1u
X8151 vdd tune_series_gygy[4] a_34308_16156# vdd pmos_6p0 w=1.2u l=0.5u
X8152 a_28124_16055# a_28036_16152# vss vss nmos_6p0 w=0.82u l=1u
X8153 a_19936_21720# cap_shunt_p a_17828_21720# vss nmos_6p0 w=0.82u l=0.6u
X8154 a_10360_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8155 a_13720_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8156 a_7540_38108# cap_shunt_n a_7748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X8157 a_2140_16488# a_2052_16532# vss vss nmos_6p0 w=0.82u l=1u
X8158 vss cap_series_gyn a_20048_6040# vss nmos_6p0 w=0.82u l=0.6u
X8159 vss tune_shunt[7] a_13796_12674# vss nmos_6p0 w=0.51u l=0.6u
X8160 a_33052_3511# a_32964_3608# vss vss nmos_6p0 w=0.82u l=1u
X8161 vdd a_29692_19624# a_29604_19668# vdd pmos_6p0 w=1.22u l=1u
X8162 vdd a_32604_55255# a_32516_55352# vdd pmos_6p0 w=1.22u l=1u
X8163 a_28484_5556# tune_shunt[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8164 a_7768_5180# cap_series_gyn a_7580_5180# vdd pmos_6p0 w=1.2u l=0.5u
X8165 a_33612_12919# a_33524_13016# vss vss nmos_6p0 w=0.82u l=1u
X8166 a_8848_27992# cap_shunt_n a_6740_27992# vss nmos_6p0 w=0.82u l=0.6u
X8167 a_13252_25940# cap_shunt_n a_13460_26424# vdd pmos_6p0 w=1.2u l=0.5u
X8168 vdd a_32156_5512# a_32068_5556# vdd pmos_6p0 w=1.22u l=1u
X8169 a_18612_7970# cap_series_gyp a_20328_7908# vss nmos_6p0 w=0.82u l=0.6u
X8170 vss tune_shunt[5] a_29700_31490# vss nmos_6p0 w=0.51u l=0.6u
X8171 a_2932_9176# cap_shunt_n a_4648_9176# vss nmos_6p0 w=0.82u l=0.6u
X8172 a_25780_37400# cap_shunt_p a_25572_36916# vdd pmos_6p0 w=1.2u l=0.5u
X8173 a_32404_38108# cap_shunt_p a_32612_37762# vdd pmos_6p0 w=1.2u l=0.5u
X8174 a_14484_3988# cap_series_gyp a_14692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X8175 a_11200_21720# cap_shunt_p a_9876_21720# vss nmos_6p0 w=0.82u l=0.6u
X8176 vdd a_32604_52119# a_32516_52216# vdd pmos_6p0 w=1.22u l=1u
X8177 a_24660_42466# cap_shunt_n a_24452_42812# vdd pmos_6p0 w=1.2u l=0.5u
X8178 a_20532_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8179 a_2500_30268# cap_shunt_n a_2708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X8180 a_8848_24856# cap_shunt_p a_6740_24856# vss nmos_6p0 w=0.82u l=0.6u
X8181 a_13252_22804# cap_shunt_n a_13460_23288# vdd pmos_6p0 w=1.2u l=0.5u
X8182 vss tune_series_gygy[3] a_35880_8692# vss nmos_6p0 w=0.51u l=0.6u
X8183 a_2932_9176# cap_shunt_n a_2724_8692# vdd pmos_6p0 w=1.2u l=0.5u
X8184 vdd a_18492_7080# a_18404_7124# vdd pmos_6p0 w=1.22u l=1u
X8185 a_35292_18056# a_35204_18100# vss vss nmos_6p0 w=0.82u l=1u
X8186 a_10660_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8187 a_34664_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8188 a_28484_25940# cap_shunt_p a_28692_26424# vdd pmos_6p0 w=1.2u l=0.5u
X8189 a_25572_14964# cap_series_gyp a_25780_15448# vdd pmos_6p0 w=1.2u l=0.5u
X8190 a_16500_28700# cap_shunt_n a_16708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X8191 a_13460_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8192 a_21448_12312# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8193 vss cap_shunt_p a_14896_17016# vss nmos_6p0 w=0.82u l=0.6u
X8194 a_24452_20860# cap_shunt_p a_24660_20514# vdd pmos_6p0 w=1.2u l=0.5u
X8195 vdd a_5724_54120# a_5636_54164# vdd pmos_6p0 w=1.22u l=1u
X8196 vdd a_32156_47415# a_32068_47512# vdd pmos_6p0 w=1.22u l=1u
X8197 vss cap_shunt_n a_9856_36132# vss nmos_6p0 w=0.82u l=0.6u
X8198 vdd a_24204_24328# a_24116_24372# vdd pmos_6p0 w=1.22u l=1u
X8199 a_35292_14920# a_35204_14964# vss vss nmos_6p0 w=0.82u l=1u
X8200 a_28484_22804# cap_shunt_p a_28692_23288# vdd pmos_6p0 w=1.2u l=0.5u
X8201 a_33524_35348# cap_shunt_n a_33732_35832# vdd pmos_6p0 w=1.2u l=0.5u
X8202 vdd a_19276_30167# a_19188_30264# vdd pmos_6p0 w=1.22u l=1u
X8203 a_16708_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8204 a_25572_11828# cap_series_gyp a_25780_12312# vdd pmos_6p0 w=1.2u l=0.5u
X8205 a_14112_18584# cap_shunt_p a_12788_18584# vss nmos_6p0 w=0.82u l=0.6u
X8206 a_13564_52119# a_13476_52216# vss vss nmos_6p0 w=0.82u l=1u
X8207 a_3828_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8208 a_1716_3612# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8209 a_15904_39268# cap_shunt_n a_13796_39330# vss nmos_6p0 w=0.82u l=0.6u
X8210 a_35880_10260# cap_series_gygyp a_35692_10260# vdd pmos_6p0 w=1.2u l=0.5u
X8211 vss cap_shunt_p a_10640_48676# vss nmos_6p0 w=0.82u l=0.6u
X8212 a_5636_9884# cap_shunt_p a_5844_9538# vdd pmos_6p0 w=1.2u l=0.5u
X8213 vdd a_37420_17623# a_37332_17720# vdd pmos_6p0 w=1.22u l=1u
X8214 vdd a_24204_21192# a_24116_21236# vdd pmos_6p0 w=1.22u l=1u
X8215 a_2588_47848# a_2500_47892# vss vss nmos_6p0 w=0.82u l=1u
X8216 a_30632_39268# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8217 vdd a_6956_34871# a_6868_34968# vdd pmos_6p0 w=1.22u l=1u
X8218 a_12264_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8219 a_21748_6402# cap_series_gyn a_23464_6340# vss nmos_6p0 w=0.82u l=0.6u
X8220 a_18940_11784# a_18852_11828# vss vss nmos_6p0 w=0.82u l=1u
X8221 a_20740_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8222 a_21540_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8223 a_14112_15448# cap_shunt_p a_12788_15448# vss nmos_6p0 w=0.82u l=0.6u
X8224 a_9072_34564# cap_shunt_n a_7748_34626# vss nmos_6p0 w=0.82u l=0.6u
X8225 vdd a_12108_9783# a_12020_9880# vdd pmos_6p0 w=1.22u l=1u
X8226 a_6532_41620# cap_shunt_n a_6740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X8227 a_3828_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8228 a_18044_8648# a_17956_8692# vss vss nmos_6p0 w=0.82u l=1u
X8229 vss tune_series_gygy[2] a_34536_6748# vss nmos_6p0 w=0.51u l=0.6u
X8230 a_35692_19668# cap_series_gygyp a_35880_19668# vdd pmos_6p0 w=1.2u l=0.5u
X8231 a_24660_26786# cap_shunt_p a_24452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X8232 a_32612_25218# cap_shunt_p a_32404_25564# vdd pmos_6p0 w=1.2u l=0.5u
X8233 vss cap_shunt_p a_15904_18884# vss nmos_6p0 w=0.82u l=0.6u
X8234 vdd a_1692_19624# a_1604_19668# vdd pmos_6p0 w=1.22u l=1u
X8235 a_30016_34264# cap_shunt_p a_28692_34264# vss nmos_6p0 w=0.82u l=0.6u
X8236 a_23632_3204# cap_series_gyp a_21524_3266# vss nmos_6p0 w=0.82u l=0.6u
X8237 a_20740_15448# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8238 vdd a_30140_41576# a_30052_41620# vdd pmos_6p0 w=1.22u l=1u
X8239 a_20172_36439# a_20084_36536# vss vss nmos_6p0 w=0.82u l=1u
X8240 a_21540_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8241 vss tune_shunt[6] a_7748_44034# vss nmos_6p0 w=0.51u l=0.6u
X8242 vss tune_shunt_gy[1] a_37632_38485# vss nmos_6p0 w=0.51u l=0.6u
X8243 a_9072_31428# cap_shunt_n a_7748_31490# vss nmos_6p0 w=0.82u l=0.6u
X8244 vdd a_20732_49416# a_20644_49460# vdd pmos_6p0 w=1.22u l=1u
X8245 a_2708_48738# cap_shunt_p a_2500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X8246 a_10660_29922# cap_shunt_n a_10452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X8247 vdd tune_series_gygy[3] a_35692_8692# vdd pmos_6p0 w=1.2u l=0.5u
X8248 a_3036_13352# a_2948_13396# vss vss nmos_6p0 w=0.82u l=1u
X8249 a_3828_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8250 vss tune_shunt[7] a_17828_32696# vss nmos_6p0 w=0.51u l=0.6u
X8251 vss cap_shunt_p a_15904_15748# vss nmos_6p0 w=0.82u l=0.6u
X8252 a_13588_49084# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8253 a_30016_31128# cap_shunt_n a_28692_31128# vss nmos_6p0 w=0.82u l=0.6u
X8254 a_37280_43734# tune_shunt_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X8255 a_6292_49944# cap_shunt_p a_8008_49944# vss nmos_6p0 w=0.82u l=0.6u
X8256 a_12580_49460# cap_shunt_n a_12788_49944# vdd pmos_6p0 w=1.2u l=0.5u
X8257 vdd a_32604_48983# a_32516_49080# vdd pmos_6p0 w=1.22u l=1u
X8258 a_10660_37762# cap_shunt_n a_11592_37700# vss nmos_6p0 w=0.82u l=0.6u
X8259 a_11572_5556# cap_series_gyn a_11780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X8260 vdd tune_series_gygy[2] a_35692_5556# vdd pmos_6p0 w=1.2u l=0.5u
X8261 vss tune_shunt[3] a_2932_10744# vss nmos_6p0 w=0.51u l=0.6u
X8262 vdd a_31260_33736# a_31172_33780# vdd pmos_6p0 w=1.22u l=1u
X8263 a_3828_15448# cap_shunt_p a_3620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X8264 vss cap_shunt_p a_8400_48676# vss nmos_6p0 w=0.82u l=0.6u
X8265 a_35692_36916# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8266 a_14484_10260# cap_series_gyn a_14692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X8267 vdd a_18940_53687# a_18852_53784# vdd pmos_6p0 w=1.22u l=1u
X8268 a_24660_36194# cap_shunt_p a_24452_36540# vdd pmos_6p0 w=1.2u l=0.5u
X8269 vss cap_shunt_n a_19936_46808# vss nmos_6p0 w=0.82u l=0.6u
X8270 a_28692_12312# cap_series_gyn a_30408_12312# vss nmos_6p0 w=0.82u l=0.6u
X8271 vdd a_16476_52552# a_16388_52596# vdd pmos_6p0 w=1.22u l=1u
X8272 a_32612_34626# cap_shunt_n a_32404_34972# vdd pmos_6p0 w=1.2u l=0.5u
X8273 a_19276_48983# a_19188_49080# vss vss nmos_6p0 w=0.82u l=1u
X8274 a_6760_7124# cap_series_gyp a_6572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X8275 vdd a_31260_30600# a_31172_30644# vdd pmos_6p0 w=1.22u l=1u
X8276 a_25780_27992# cap_shunt_p a_25572_27508# vdd pmos_6p0 w=1.2u l=0.5u
X8277 a_11200_12312# cap_shunt_p a_9876_12312# vss nmos_6p0 w=0.82u l=0.6u
X8278 a_24660_33058# cap_shunt_p a_24452_33404# vdd pmos_6p0 w=1.2u l=0.5u
X8279 vdd a_35180_38007# a_35092_38104# vdd pmos_6p0 w=1.22u l=1u
X8280 a_31416_34564# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8281 a_17828_32696# cap_shunt_n a_18760_32696# vss nmos_6p0 w=0.82u l=0.6u
X8282 a_32612_31490# cap_shunt_n a_32404_31836# vdd pmos_6p0 w=1.2u l=0.5u
X8283 a_24764_45847# a_24676_45944# vss vss nmos_6p0 w=0.82u l=1u
X8284 a_24452_44380# cap_shunt_p a_24660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X8285 a_8848_15448# cap_shunt_p a_6740_15448# vss nmos_6p0 w=0.82u l=0.6u
X8286 a_16500_20860# cap_shunt_p a_16708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X8287 vss tune_shunt[1] a_25780_4472# vss nmos_6p0 w=0.51u l=0.6u
X8288 a_16708_48738# cap_shunt_p a_16500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X8289 vdd a_37868_9783# a_37780_9880# vdd pmos_6p0 w=1.22u l=1u
X8290 a_28484_16532# cap_series_gyn a_28692_17016# vdd pmos_6p0 w=1.2u l=0.5u
X8291 a_33524_29076# cap_shunt_p a_33732_29560# vdd pmos_6p0 w=1.2u l=0.5u
X8292 a_11668_42104# cap_shunt_n a_11460_41620# vdd pmos_6p0 w=1.2u l=0.5u
X8293 a_31416_31428# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8294 a_24452_5180# cap_series_gyp a_24660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X8295 a_24452_11452# cap_series_gyp a_24660_11106# vdd pmos_6p0 w=1.2u l=0.5u
X8296 a_24452_41244# cap_shunt_n a_24660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X8297 vdd a_29580_54120# a_29492_54164# vdd pmos_6p0 w=1.22u l=1u
X8298 a_4424_9476# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8299 a_24452_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8300 vdd a_6956_28599# a_6868_28696# vdd pmos_6p0 w=1.22u l=1u
X8301 a_23576_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X8302 vdd a_37868_6647# a_37780_6744# vdd pmos_6p0 w=1.22u l=1u
X8303 a_21748_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8304 a_7540_42812# cap_shunt_n a_7748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X8305 a_9072_28292# cap_shunt_n a_7748_28354# vss nmos_6p0 w=0.82u l=0.6u
X8306 a_36160_45302# tune_shunt_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X8307 a_18760_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8308 a_25780_37400# cap_shunt_p a_25572_36916# vdd pmos_6p0 w=1.2u l=0.5u
X8309 vdd a_29580_50984# a_29492_51028# vdd pmos_6p0 w=1.22u l=1u
X8310 a_32404_38108# cap_shunt_p a_32612_37762# vdd pmos_6p0 w=1.2u l=0.5u
X8311 vdd tune_shunt[7] a_10340_33780# vdd pmos_6p0 w=1.2u l=0.5u
X8312 a_36624_23588# cap_series_gygyp a_34516_23650# vss nmos_6p0 w=0.82u l=0.6u
X8313 a_36636_54120# a_36548_54164# vss vss nmos_6p0 w=0.82u l=1u
X8314 a_6740_48376# cap_shunt_p a_8456_48376# vss nmos_6p0 w=0.82u l=0.6u
X8315 a_12264_23288# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8316 vdd a_37868_3511# a_37780_3608# vdd pmos_6p0 w=1.22u l=1u
X8317 vdd a_20620_23895# a_20532_23992# vdd pmos_6p0 w=1.22u l=1u
X8318 a_21540_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8319 a_6532_32212# cap_shunt_n a_6740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X8320 a_9072_25156# cap_shunt_n a_7748_25218# vss nmos_6p0 w=0.82u l=0.6u
X8321 a_18760_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8322 vss cap_shunt_n a_11984_32996# vss nmos_6p0 w=0.82u l=0.6u
X8323 a_3380_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8324 vdd tune_shunt[7] a_10340_30644# vdd pmos_6p0 w=1.2u l=0.5u
X8325 a_28484_25940# cap_shunt_p a_28692_26424# vdd pmos_6p0 w=1.2u l=0.5u
X8326 a_10492_8316# cap_series_gyp a_10680_8316# vdd pmos_6p0 w=1.2u l=0.5u
X8327 vss tune_shunt[7] a_12788_13880# vss nmos_6p0 w=0.51u l=0.6u
X8328 vdd tune_shunt[7] a_13588_30268# vdd pmos_6p0 w=1.2u l=0.5u
X8329 a_25572_14964# cap_series_gyp a_25780_15448# vdd pmos_6p0 w=1.2u l=0.5u
X8330 a_34516_4834# cap_series_gygyp a_34308_5180# vdd pmos_6p0 w=1.2u l=0.5u
X8331 vdd a_20620_20759# a_20532_20856# vdd pmos_6p0 w=1.22u l=1u
X8332 vss cap_series_gyn a_19712_3204# vss nmos_6p0 w=0.82u l=0.6u
X8333 a_4256_9176# cap_shunt_n a_2932_9176# vss nmos_6p0 w=0.82u l=0.6u
X8334 a_30924_50984# a_30836_51028# vss vss nmos_6p0 w=0.82u l=1u
X8335 a_28484_22804# cap_shunt_p a_28692_23288# vdd pmos_6p0 w=1.2u l=0.5u
X8336 a_12892_10216# a_12804_10260# vss vss nmos_6p0 w=0.82u l=1u
X8337 a_33524_35348# cap_shunt_n a_33732_35832# vdd pmos_6p0 w=1.2u l=0.5u
X8338 vss tune_shunt[7] a_17828_23288# vss nmos_6p0 w=0.51u l=0.6u
X8339 a_25572_11828# cap_series_gyp a_25780_12312# vdd pmos_6p0 w=1.2u l=0.5u
X8340 a_18404_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8341 a_10988_46280# a_10900_46324# vss vss nmos_6p0 w=0.82u l=1u
X8342 vdd a_1692_45847# a_1604_45944# vdd pmos_6p0 w=1.22u l=1u
X8343 a_35880_10260# cap_series_gygyp a_35692_10260# vdd pmos_6p0 w=1.2u l=0.5u
X8344 a_18404_3988# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8345 a_6628_12674# cap_shunt_p a_6420_13020# vdd pmos_6p0 w=1.2u l=0.5u
X8346 vss cap_shunt_p a_27888_32696# vss nmos_6p0 w=0.82u l=0.6u
X8347 vdd tune_shunt[7] a_10452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X8348 vdd a_31260_24328# a_31172_24372# vdd pmos_6p0 w=1.22u l=1u
X8349 vss tune_series_gy[3] a_21524_4472# vss nmos_6p0 w=0.51u l=0.6u
X8350 a_2140_22327# a_2052_22424# vss vss nmos_6p0 w=0.82u l=1u
X8351 a_19388_53687# a_19300_53784# vss vss nmos_6p0 w=0.82u l=1u
X8352 a_9876_53080# cap_shunt_n a_10808_53080# vss nmos_6p0 w=0.82u l=0.6u
X8353 vdd a_25548_47415# a_25460_47512# vdd pmos_6p0 w=1.22u l=1u
X8354 a_7540_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8355 vdd a_1692_42711# a_1604_42808# vdd pmos_6p0 w=1.22u l=1u
X8356 a_24660_26786# cap_shunt_p a_24452_27132# vdd pmos_6p0 w=1.2u l=0.5u
X8357 a_12788_13880# cap_shunt_p a_13720_13880# vss nmos_6p0 w=0.82u l=0.6u
X8358 a_31416_28292# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8359 a_32612_25218# cap_shunt_p a_32404_25564# vdd pmos_6p0 w=1.2u l=0.5u
X8360 a_21748_23650# cap_shunt_p a_21540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X8361 a_19276_39575# a_19188_39672# vss vss nmos_6p0 w=0.82u l=1u
X8362 a_10660_29922# cap_shunt_n a_10452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X8363 a_5844_9538# cap_shunt_p a_6776_9476# vss nmos_6p0 w=0.82u l=0.6u
X8364 vss tune_shunt[5] a_20740_43672# vss nmos_6p0 w=0.51u l=0.6u
X8365 vdd a_36076_31735# a_35988_31832# vdd pmos_6p0 w=1.22u l=1u
X8366 a_1924_7608# cap_shunt_n a_2856_7608# vss nmos_6p0 w=0.82u l=0.6u
X8367 vss cap_shunt_p a_23856_39268# vss nmos_6p0 w=0.82u l=0.6u
X8368 a_31416_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8369 a_17828_23288# cap_shunt_n a_18760_23288# vss nmos_6p0 w=0.82u l=0.6u
X8370 vdd a_37868_36439# a_37780_36536# vdd pmos_6p0 w=1.22u l=1u
X8371 a_16140_55688# a_16052_55732# vss vss nmos_6p0 w=0.82u l=1u
X8372 a_22644_12312# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8373 vss tune_shunt[6] a_20740_40536# vss nmos_6p0 w=0.51u l=0.6u
X8374 a_7540_36540# cap_shunt_n a_7748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X8375 vss tune_series_gy[4] a_14692_7608# vss nmos_6p0 w=0.51u l=0.6u
X8376 a_14484_10260# cap_series_gyn a_14692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X8377 a_2708_50306# cap_shunt_n a_2500_50652# vdd pmos_6p0 w=1.2u l=0.5u
X8378 a_4424_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8379 a_15512_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8380 a_16708_42466# cap_shunt_n a_16500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X8381 a_25572_40052# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8382 vss tune_shunt[6] a_6740_45240# vss nmos_6p0 w=0.51u l=0.6u
X8383 a_20532_44756# cap_shunt_n a_20740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X8384 a_11480_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8385 vss tune_shunt[5] a_6292_51874# vss nmos_6p0 w=0.51u l=0.6u
X8386 a_7540_33404# cap_shunt_n a_7748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X8387 a_18760_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8388 a_25780_27992# cap_shunt_p a_25572_27508# vdd pmos_6p0 w=1.2u l=0.5u
X8389 vdd tune_shunt[7] a_10340_24372# vdd pmos_6p0 w=1.2u l=0.5u
X8390 a_6760_3988# cap_series_gyp a_7568_4472# vss nmos_6p0 w=0.82u l=0.6u
X8391 a_6776_9176# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8392 a_2588_53687# a_2500_53784# vss vss nmos_6p0 w=0.82u l=1u
X8393 vdd a_11996_20759# a_11908_20856# vdd pmos_6p0 w=1.22u l=1u
X8394 a_15512_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8395 a_14372_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8396 vss tune_shunt[6] a_6740_42104# vss nmos_6p0 w=0.51u l=0.6u
X8397 vdd a_24652_33736# a_24564_33780# vdd pmos_6p0 w=1.22u l=1u
X8398 vdd a_20620_14487# a_20532_14584# vdd pmos_6p0 w=1.22u l=1u
X8399 a_24452_44380# cap_shunt_p a_24660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X8400 a_33732_35832# cap_shunt_n a_35448_35832# vss nmos_6p0 w=0.82u l=0.6u
X8401 a_16500_20860# cap_shunt_p a_16708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X8402 a_18760_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8403 a_35628_30167# a_35540_30264# vss vss nmos_6p0 w=0.82u l=1u
X8404 a_1716_7124# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8405 a_28484_3988# tune_series_gy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8406 vss tune_shunt[7] a_13796_29922# vss nmos_6p0 w=0.51u l=0.6u
X8407 vss cap_shunt_n a_11984_23588# vss nmos_6p0 w=0.82u l=0.6u
X8408 vss cap_shunt_n a_15568_34264# vss nmos_6p0 w=0.82u l=0.6u
X8409 a_23968_12312# cap_series_gyn a_22644_12312# vss nmos_6p0 w=0.82u l=0.6u
X8410 a_28484_16532# cap_series_gyn a_28692_17016# vdd pmos_6p0 w=1.2u l=0.5u
X8411 a_33524_29076# cap_shunt_p a_33732_29560# vdd pmos_6p0 w=1.2u l=0.5u
X8412 a_20532_14964# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8413 vss cap_shunt_p a_5488_17016# vss nmos_6p0 w=0.82u l=0.6u
X8414 a_9220_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8415 vdd a_24652_30600# a_24564_30644# vdd pmos_6p0 w=1.22u l=1u
X8416 vss tune_series_gy[3] a_24660_6402# vss nmos_6p0 w=0.51u l=0.6u
X8417 a_24452_41244# cap_shunt_n a_24660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X8418 vdd tune_series_gy[4] a_24452_9884# vdd pmos_6p0 w=1.2u l=0.5u
X8419 vdd a_1692_39575# a_1604_39672# vdd pmos_6p0 w=1.22u l=1u
X8420 a_2708_9538# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X8421 a_35628_27031# a_35540_27128# vss vss nmos_6p0 w=0.82u l=1u
X8422 a_4704_18584# cap_shunt_p a_3380_18584# vss nmos_6p0 w=0.82u l=0.6u
X8423 vdd a_17596_3944# a_17508_3988# vdd pmos_6p0 w=1.22u l=1u
X8424 vss cap_shunt_n a_15568_31128# vss nmos_6p0 w=0.82u l=0.6u
X8425 vdd a_13900_3511# a_13812_3608# vdd pmos_6p0 w=1.22u l=1u
X8426 vdd a_28572_38007# a_28484_38104# vdd pmos_6p0 w=1.22u l=1u
X8427 vdd a_36524_30167# a_36436_30264# vdd pmos_6p0 w=1.22u l=1u
X8428 a_21524_4472# cap_series_gyn a_21316_3988# vdd pmos_6p0 w=1.2u l=0.5u
X8429 vdd tune_series_gy[3] a_24452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X8430 a_30812_52119# a_30724_52216# vss vss nmos_6p0 w=0.82u l=1u
X8431 vdd a_1692_36439# a_1604_36536# vdd pmos_6p0 w=1.22u l=1u
X8432 vdd tune_shunt[7] a_10340_33780# vdd pmos_6p0 w=1.2u l=0.5u
X8433 a_14784_32696# cap_shunt_n a_13460_32696# vss nmos_6p0 w=0.82u l=0.6u
X8434 a_29624_27992# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8435 vss cap_shunt_p a_27888_23288# vss nmos_6p0 w=0.82u l=0.6u
X8436 vss cap_shunt_n a_30800_6040# vss nmos_6p0 w=0.82u l=0.6u
X8437 a_28796_19624# a_28708_19668# vss vss nmos_6p0 w=0.82u l=1u
X8438 a_13564_6647# a_13476_6744# vss vss nmos_6p0 w=0.82u l=1u
X8439 a_28572_19191# a_28484_19288# vss vss nmos_6p0 w=0.82u l=1u
X8440 a_18612_6402# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X8441 vdd a_29916_8215# a_29828_8312# vdd pmos_6p0 w=1.22u l=1u
X8442 a_6292_51874# cap_shunt_p a_8008_51812# vss nmos_6p0 w=0.82u l=0.6u
X8443 a_17620_46324# cap_shunt_n a_17828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X8444 vdd tune_shunt[7] a_10340_30644# vdd pmos_6p0 w=1.2u l=0.5u
X8445 a_28484_25940# cap_shunt_p a_28692_26424# vdd pmos_6p0 w=1.2u l=0.5u
X8446 vdd a_36076_25463# a_35988_25560# vdd pmos_6p0 w=1.22u l=1u
X8447 a_29624_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8448 a_14728_12612# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8449 a_21748_14242# cap_series_gyn a_21540_14588# vdd pmos_6p0 w=1.2u l=0.5u
X8450 a_11612_8692# cap_series_gyp a_11800_8692# vdd pmos_6p0 w=1.2u l=0.5u
X8451 a_28572_16055# a_28484_16152# vss vss nmos_6p0 w=0.82u l=1u
X8452 a_8456_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8453 vss tune_shunt[7] a_20740_34264# vss nmos_6p0 w=0.51u l=0.6u
X8454 a_28484_22804# cap_shunt_p a_28692_23288# vdd pmos_6p0 w=1.2u l=0.5u
X8455 vdd tune_shunt[6] a_9668_49460# vdd pmos_6p0 w=1.2u l=0.5u
X8456 a_33732_35832# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X8457 vdd tune_shunt[6] a_7540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X8458 a_19732_13880# cap_series_gyn a_19524_13396# vdd pmos_6p0 w=1.2u l=0.5u
X8459 a_2500_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8460 a_2708_44034# cap_shunt_p a_2500_44380# vdd pmos_6p0 w=1.2u l=0.5u
X8461 vdd a_37868_27031# a_37780_27128# vdd pmos_6p0 w=1.22u l=1u
X8462 a_21540_45948# cap_shunt_p a_21748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X8463 a_16708_36194# cap_shunt_n a_16500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X8464 a_20532_38484# cap_shunt_n a_20740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X8465 a_2932_9176# cap_shunt_n a_2724_8692# vdd pmos_6p0 w=1.2u l=0.5u
X8466 a_34536_9884# cap_series_gygyn a_34348_9884# vdd pmos_6p0 w=1.2u l=0.5u
X8467 vss cap_shunt_n a_34720_36132# vss nmos_6p0 w=0.82u l=0.6u
X8468 vss tune_shunt[7] a_20740_31128# vss nmos_6p0 w=0.51u l=0.6u
X8469 a_7540_27132# cap_shunt_n a_7748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X8470 vss cap_shunt_p a_10752_18884# vss nmos_6p0 w=0.82u l=0.6u
X8471 vdd a_31708_32168# a_31620_32212# vdd pmos_6p0 w=1.22u l=1u
X8472 a_16500_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8473 a_2708_40898# cap_shunt_p a_2500_41244# vdd pmos_6p0 w=1.2u l=0.5u
X8474 a_19320_3204# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8475 a_28484_3988# cap_series_gyp a_28692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X8476 vdd tune_shunt[7] a_17620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X8477 vss cap_shunt_p a_30800_40536# vss nmos_6p0 w=0.82u l=0.6u
X8478 a_15512_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8479 a_16708_33058# cap_shunt_n a_16500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X8480 a_20532_35348# cap_shunt_n a_20740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X8481 a_34536_6748# cap_series_gygyp a_34348_6748# vdd pmos_6p0 w=1.2u l=0.5u
X8482 a_25548_52552# a_25460_52596# vss vss nmos_6p0 w=0.82u l=1u
X8483 a_33732_29560# cap_shunt_p a_35448_29560# vss nmos_6p0 w=0.82u l=0.6u
X8484 a_21748_23650# cap_shunt_p a_21540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X8485 a_25780_26424# cap_shunt_p a_25572_25940# vdd pmos_6p0 w=1.2u l=0.5u
X8486 a_10092_54120# a_10004_54164# vss vss nmos_6p0 w=0.82u l=1u
X8487 a_3828_48376# cap_shunt_p a_3620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X8488 a_31708_27464# a_31620_27508# vss vss nmos_6p0 w=0.82u l=1u
X8489 vdd a_24652_24328# a_24564_24372# vdd pmos_6p0 w=1.22u l=1u
X8490 vdd a_22524_52552# a_22436_52596# vdd pmos_6p0 w=1.22u l=1u
X8491 vdd a_31708_7080# a_31620_7124# vdd pmos_6p0 w=1.22u l=1u
X8492 vss cap_series_gygyn a_32824_20452# vss nmos_6p0 w=0.82u l=0.6u
X8493 a_6532_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8494 a_25780_23288# cap_shunt_p a_25572_22804# vdd pmos_6p0 w=1.2u l=0.5u
X8495 vdd tune_series_gy[5] a_21540_8316# vdd pmos_6p0 w=1.2u l=0.5u
X8496 a_13796_12674# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8497 a_20740_42104# cap_shunt_p a_20532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X8498 a_9428_18946# cap_shunt_p a_9220_19292# vdd pmos_6p0 w=1.2u l=0.5u
X8499 a_3828_45240# cap_shunt_p a_3620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X8500 a_31708_24328# a_31620_24372# vss vss nmos_6p0 w=0.82u l=1u
X8501 a_14484_10260# cap_series_gyn a_14692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X8502 a_13796_12674# cap_shunt_p a_15512_12612# vss nmos_6p0 w=0.82u l=0.6u
X8503 vdd a_24652_21192# a_24564_21236# vdd pmos_6p0 w=1.22u l=1u
X8504 a_13252_36916# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8505 vss tune_shunt[3] a_5844_11106# vss nmos_6p0 w=0.51u l=0.6u
X8506 a_23856_12612# cap_series_gyn a_21748_12674# vss nmos_6p0 w=0.82u l=0.6u
X8507 vss cap_shunt_n a_18032_29860# vss nmos_6p0 w=0.82u l=0.6u
X8508 a_3620_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8509 a_26376_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8510 vdd tune_series_gygy[5] a_34308_17724# vdd pmos_6p0 w=1.2u l=0.5u
X8511 a_7728_22020# cap_shunt_p a_6404_22082# vss nmos_6p0 w=0.82u l=0.6u
X8512 a_31372_55688# a_31284_55732# vss vss nmos_6p0 w=0.82u l=1u
X8513 a_36188_52119# a_36100_52216# vss vss nmos_6p0 w=0.82u l=1u
X8514 a_13588_50652# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8515 a_21672_45240# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8516 a_32404_36540# cap_shunt_n a_32612_36194# vdd pmos_6p0 w=1.2u l=0.5u
X8517 vss cap_shunt_n a_5936_35832# vss nmos_6p0 w=0.82u l=0.6u
X8518 a_29700_4834# cap_shunt_p a_30632_4772# vss nmos_6p0 w=0.82u l=0.6u
X8519 a_2708_18946# cap_shunt_p a_4424_18884# vss nmos_6p0 w=0.82u l=0.6u
X8520 a_30812_42711# a_30724_42808# vss vss nmos_6p0 w=0.82u l=1u
X8521 vss tune_shunt[6] a_21748_37762# vss nmos_6p0 w=0.51u l=0.6u
X8522 vdd tune_shunt[6] a_20532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X8523 vdd a_1692_27031# a_1604_27128# vdd pmos_6p0 w=1.22u l=1u
X8524 vdd tune_shunt[7] a_10340_24372# vdd pmos_6p0 w=1.2u l=0.5u
X8525 a_25572_7124# cap_series_gyn a_25780_7608# vdd pmos_6p0 w=1.2u l=0.5u
X8526 a_14784_23288# cap_shunt_n a_13460_23288# vss nmos_6p0 w=0.82u l=0.6u
X8527 vdd tune_series_gygy[3] a_34348_8316# vdd pmos_6p0 w=1.2u l=0.5u
X8528 vss cap_shunt_n a_18032_26724# vss nmos_6p0 w=0.82u l=0.6u
X8529 a_15492_8316# cap_series_gyn a_15700_7970# vdd pmos_6p0 w=1.2u l=0.5u
X8530 a_29624_18584# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X8531 a_24452_44380# cap_shunt_p a_24660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X8532 a_26376_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8533 vdd tune_series_gy[3] a_21316_3612# vdd pmos_6p0 w=1.2u l=0.5u
X8534 a_19724_38007# a_19636_38104# vss vss nmos_6p0 w=0.82u l=1u
X8535 vdd a_33948_13352# a_33860_13396# vdd pmos_6p0 w=1.22u l=1u
X8536 a_21672_42104# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8537 a_32404_33404# cap_shunt_n a_32612_33058# vdd pmos_6p0 w=1.2u l=0.5u
X8538 a_2708_15810# cap_shunt_p a_4424_15748# vss nmos_6p0 w=0.82u l=0.6u
X8539 vss tune_shunt[6] a_21748_34626# vss nmos_6p0 w=0.51u l=0.6u
X8540 a_21748_33058# cap_shunt_n a_22680_32996# vss nmos_6p0 w=0.82u l=0.6u
X8541 a_33732_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8542 a_9980_3511# a_9892_3608# vss vss nmos_6p0 w=0.82u l=1u
X8543 a_28484_16532# cap_series_gyn a_28692_17016# vdd pmos_6p0 w=1.2u l=0.5u
X8544 a_29624_15448# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8545 a_9220_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8546 vdd tune_shunt[6] a_7540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X8547 a_21748_45602# cap_shunt_p a_23464_45540# vss nmos_6p0 w=0.82u l=0.6u
X8548 a_24452_41244# cap_shunt_n a_24660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X8549 a_17828_48376# cap_shunt_p a_17620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X8550 a_8456_12312# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8551 a_21540_39676# cap_shunt_p a_21748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X8552 a_13460_35832# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8553 vss tune_shunt[3] a_2932_10744# vss nmos_6p0 w=0.51u l=0.6u
X8554 vdd a_31260_41143# a_31172_41240# vdd pmos_6p0 w=1.22u l=1u
X8555 vdd a_12444_17623# a_12356_17720# vdd pmos_6p0 w=1.22u l=1u
X8556 a_20740_21720# cap_shunt_p a_21672_21720# vss nmos_6p0 w=0.82u l=0.6u
X8557 vdd tune_shunt[7] a_16500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X8558 a_29916_55255# a_29828_55352# vss vss nmos_6p0 w=0.82u l=1u
X8559 a_2140_50984# a_2052_51028# vss vss nmos_6p0 w=0.82u l=1u
X8560 a_21292_47848# a_21204_47892# vss vss nmos_6p0 w=0.82u l=1u
X8561 a_21748_42466# cap_shunt_n a_23464_42404# vss nmos_6p0 w=0.82u l=0.6u
X8562 a_17828_45240# cap_shunt_p a_17620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X8563 vss cap_shunt_p a_30800_34264# vss nmos_6p0 w=0.82u l=0.6u
X8564 a_16708_26786# cap_shunt_n a_16500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X8565 vss tune_series_gy[5] a_19732_9176# vss nmos_6p0 w=0.51u l=0.6u
X8566 a_3932_55688# a_3844_55732# vss vss nmos_6p0 w=0.82u l=1u
X8567 a_20532_29076# cap_shunt_n a_20740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X8568 a_22680_43972# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8569 a_35692_25940# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8570 a_24204_47415# a_24116_47512# vss vss nmos_6p0 w=0.82u l=1u
X8571 a_36636_53687# a_36548_53784# vss vss nmos_6p0 w=0.82u l=1u
X8572 vss cap_shunt_n a_30800_31128# vss nmos_6p0 w=0.82u l=0.6u
X8573 a_36232_20452# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X8574 a_6572_3988# cap_series_gyp a_6760_3988# vdd pmos_6p0 w=1.2u l=0.5u
X8575 vss cap_shunt_p a_8064_45240# vss nmos_6p0 w=0.82u l=0.6u
X8576 a_22680_40836# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8577 a_21748_14242# cap_series_gyn a_21540_14588# vdd pmos_6p0 w=1.2u l=0.5u
X8578 a_17828_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8579 vdd a_6508_44279# a_6420_44376# vdd pmos_6p0 w=1.22u l=1u
X8580 a_35692_22804# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8581 a_25780_17016# cap_series_gyp a_25572_16532# vdd pmos_6p0 w=1.2u l=0.5u
X8582 vss cap_shunt_p a_8512_22020# vss nmos_6p0 w=0.82u l=0.6u
X8583 a_9876_13880# cap_shunt_p a_11592_13880# vss nmos_6p0 w=0.82u l=0.6u
X8584 a_6740_40536# cap_shunt_n a_6532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X8585 vss cap_shunt_p a_10864_9476# vss nmos_6p0 w=0.82u l=0.6u
X8586 vss cap_shunt_n a_8064_42104# vss nmos_6p0 w=0.82u l=0.6u
X8587 a_3828_38968# cap_shunt_n a_3620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X8588 a_28692_34264# cap_shunt_p a_28484_33780# vdd pmos_6p0 w=1.2u l=0.5u
X8589 vss cap_series_gyn a_27888_7608# vss nmos_6p0 w=0.82u l=0.6u
X8590 a_31708_18056# a_31620_18100# vss vss nmos_6p0 w=0.82u l=1u
X8591 vss cap_shunt_gyn a_34188_43672# vss nmos_6p0 w=0.82u l=0.6u
X8592 a_17260_50551# a_17172_50648# vss vss nmos_6p0 w=0.82u l=1u
X8593 a_6532_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8594 a_11800_8692# cap_series_gyp a_11612_8692# vdd pmos_6p0 w=1.2u l=0.5u
X8595 a_34516_12674# cap_series_gygyp a_34308_13020# vdd pmos_6p0 w=1.2u l=0.5u
X8596 a_6292_49944# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8597 a_7580_5180# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8598 a_9876_10744# cap_shunt_p a_11592_10744# vss nmos_6p0 w=0.82u l=0.6u
X8599 a_20740_32696# cap_shunt_n a_20532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X8600 a_13588_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8601 a_3828_35832# cap_shunt_n a_3620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X8602 vss cap_shunt_p a_31808_32996# vss nmos_6p0 w=0.82u l=0.6u
X8603 a_28692_31128# cap_shunt_n a_28484_30644# vdd pmos_6p0 w=1.2u l=0.5u
X8604 vss cap_shunt_n a_5936_29560# vss nmos_6p0 w=0.82u l=0.6u
X8605 a_31708_14920# a_31620_14964# vss vss nmos_6p0 w=0.82u l=1u
X8606 a_13252_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8607 vdd a_32716_39575# a_32628_39672# vdd pmos_6p0 w=1.22u l=1u
X8608 a_22456_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8609 a_32156_38440# a_32068_38484# vss vss nmos_6p0 w=0.82u l=1u
X8610 a_17828_37400# cap_shunt_n a_19544_37400# vss nmos_6p0 w=0.82u l=0.6u
X8611 a_6740_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8612 a_3620_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8613 vdd a_29468_22327# a_29380_22424# vdd pmos_6p0 w=1.22u l=1u
X8614 a_34396_21192# a_34308_21236# vss vss nmos_6p0 w=0.82u l=1u
X8615 a_27888_37400# cap_shunt_p a_25780_37400# vss nmos_6p0 w=0.82u l=0.6u
X8616 vss tune_shunt[7] a_3828_32696# vss nmos_6p0 w=0.51u l=0.6u
X8617 a_13588_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8618 vss tune_shunt[7] a_21748_28354# vss nmos_6p0 w=0.51u l=0.6u
X8619 a_32404_27132# cap_shunt_p a_32612_26786# vdd pmos_6p0 w=1.2u l=0.5u
X8620 vss cap_shunt_p a_5936_26424# vss nmos_6p0 w=0.82u l=0.6u
X8621 a_25780_26424# cap_shunt_p a_25572_25940# vdd pmos_6p0 w=1.2u l=0.5u
X8622 a_13888_4472# cap_series_gyp a_11780_4472# vss nmos_6p0 w=0.82u l=0.6u
X8623 a_12580_18100# cap_shunt_p a_12788_18584# vdd pmos_6p0 w=1.2u l=0.5u
X8624 a_36720_46870# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8625 vdd tune_shunt[7] a_20532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X8626 vss cap_shunt_p a_9072_43972# vss nmos_6p0 w=0.82u l=0.6u
X8627 a_22456_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8628 a_3620_13396# cap_shunt_n a_3828_13880# vdd pmos_6p0 w=1.2u l=0.5u
X8629 vss cap_shunt_p a_7728_47108# vss nmos_6p0 w=0.82u l=0.6u
X8630 a_12580_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8631 vss cap_shunt_p a_18032_17316# vss nmos_6p0 w=0.82u l=0.6u
X8632 vdd a_16924_32168# a_16836_32212# vdd pmos_6p0 w=1.22u l=1u
X8633 a_26376_17316# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X8634 a_13460_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8635 a_10452_6748# cap_series_gyn a_10660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X8636 a_2932_9176# cap_shunt_n a_2724_8692# vdd pmos_6p0 w=1.2u l=0.5u
X8637 vdd a_17372_55688# a_17284_55732# vdd pmos_6p0 w=1.22u l=1u
X8638 a_3620_41620# cap_shunt_p a_3828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X8639 vss tune_shunt[5] a_21748_25218# vss nmos_6p0 w=0.51u l=0.6u
X8640 a_21748_23650# cap_shunt_p a_22680_23588# vss nmos_6p0 w=0.82u l=0.6u
X8641 a_25780_23288# cap_shunt_p a_25572_22804# vdd pmos_6p0 w=1.2u l=0.5u
X8642 a_17416_7908# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8643 a_1924_6402# cap_shunt_n a_2856_6340# vss nmos_6p0 w=0.82u l=0.6u
X8644 vdd a_18940_52552# a_18852_52596# vdd pmos_6p0 w=1.22u l=1u
X8645 a_28124_44279# a_28036_44376# vss vss nmos_6p0 w=0.82u l=1u
X8646 vss cap_shunt_n a_9072_40836# vss nmos_6p0 w=0.82u l=0.6u
X8647 a_25572_33780# cap_shunt_p a_25780_34264# vdd pmos_6p0 w=1.2u l=0.5u
X8648 a_6776_11044# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8649 a_28484_33780# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8650 a_12580_11828# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8651 vss tune_shunt[7] a_9876_21720# vss nmos_6p0 w=0.51u l=0.6u
X8652 a_2140_44712# a_2052_44756# vss vss nmos_6p0 w=0.82u l=1u
X8653 a_21748_36194# cap_shunt_n a_23464_36132# vss nmos_6p0 w=0.82u l=0.6u
X8654 a_21540_13020# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8655 a_29916_48983# a_29828_49080# vss vss nmos_6p0 w=0.82u l=1u
X8656 a_17828_38968# cap_shunt_n a_17620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X8657 a_13252_36916# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8658 a_13460_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8659 a_29492_11452# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8660 vss tune_series_gy[5] a_18612_12674# vss nmos_6p0 w=0.51u l=0.6u
X8661 vdd a_37868_47848# a_37780_47892# vdd pmos_6p0 w=1.22u l=1u
X8662 a_10452_44380# cap_shunt_n a_10660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X8663 a_16924_27464# a_16836_27508# vss vss nmos_6p0 w=0.82u l=1u
X8664 a_1924_3266# cap_shunt_n a_2856_3204# vss nmos_6p0 w=0.82u l=0.6u
X8665 a_21840_12312# cap_series_gyn a_19732_12312# vss nmos_6p0 w=0.82u l=0.6u
X8666 vdd a_14348_55688# a_14260_55732# vdd pmos_6p0 w=1.22u l=1u
X8667 vdd a_25996_47415# a_25908_47512# vdd pmos_6p0 w=1.22u l=1u
X8668 vdd tune_shunt_gy[5] a_37444_47512# vdd pmos_6p0 w=1.215u l=0.5u
X8669 a_28124_41143# a_28036_41240# vss vss nmos_6p0 w=0.82u l=1u
X8670 a_25572_30644# cap_shunt_p a_25780_31128# vdd pmos_6p0 w=1.2u l=0.5u
X8671 a_28484_30644# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8672 vss cap_shunt_p a_3248_4772# vss nmos_6p0 w=0.82u l=0.6u
X8673 a_8344_12612# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8674 a_2140_41576# a_2052_41620# vss vss nmos_6p0 w=0.82u l=1u
X8675 a_32404_36540# cap_shunt_n a_32612_36194# vdd pmos_6p0 w=1.2u l=0.5u
X8676 a_17828_35832# cap_shunt_n a_17620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X8677 vss cap_shunt_p a_10864_14180# vss nmos_6p0 w=0.82u l=0.6u
X8678 vdd a_18044_55255# a_17956_55352# vdd pmos_6p0 w=1.22u l=1u
X8679 a_7748_44034# cap_shunt_p a_7540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X8680 a_11460_40052# cap_shunt_n a_11668_40536# vdd pmos_6p0 w=1.2u l=0.5u
X8681 a_21540_34972# cap_shunt_p a_21748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X8682 a_1716_3612# cap_shunt_n a_1924_3266# vdd pmos_6p0 w=1.2u l=0.5u
X8683 a_10452_41244# cap_shunt_n a_10660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X8684 a_22680_34564# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8685 a_16924_24328# a_16836_24372# vss vss nmos_6p0 w=0.82u l=1u
X8686 a_27228_12919# a_27140_13016# vss vss nmos_6p0 w=0.82u l=1u
X8687 a_35692_16532# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8688 vdd tune_shunt[7] a_3620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X8689 a_32404_33404# cap_shunt_n a_32612_33058# vdd pmos_6p0 w=1.2u l=0.5u
X8690 vss cap_shunt_p a_10864_11044# vss nmos_6p0 w=0.82u l=0.6u
X8691 a_7748_40898# cap_shunt_n a_7540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X8692 a_21540_31836# cap_shunt_n a_21748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X8693 a_24660_18946# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X8694 vdd a_18044_52119# a_17956_52216# vdd pmos_6p0 w=1.22u l=1u
X8695 a_2856_6040# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8696 a_17620_14964# cap_shunt_p a_17828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X8697 a_20532_44756# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8698 a_22680_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8699 a_17828_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8700 vdd tune_shunt[1] a_5636_3612# vdd pmos_6p0 w=1.2u l=0.5u
X8701 a_34844_19624# a_34756_19668# vss vss nmos_6p0 w=0.82u l=1u
X8702 a_4760_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8703 a_9332_9884# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8704 a_13588_45948# cap_shunt_p a_13796_45602# vdd pmos_6p0 w=1.2u l=0.5u
X8705 vss tune_shunt[6] a_2708_40898# vss nmos_6p0 w=0.51u l=0.6u
X8706 a_3828_29560# cap_shunt_n a_3620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X8707 vdd tune_shunt[7] a_16500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X8708 a_15120_29860# cap_shunt_n a_13796_29922# vss nmos_6p0 w=0.82u l=0.6u
X8709 a_28692_24856# cap_shunt_p a_28484_24372# vdd pmos_6p0 w=1.2u l=0.5u
X8710 vdd a_4492_6647# a_4404_6744# vdd pmos_6p0 w=1.22u l=1u
X8711 a_27004_45847# a_26916_45944# vss vss nmos_6p0 w=0.82u l=1u
X8712 a_35292_40008# a_35204_40052# vss vss nmos_6p0 w=0.82u l=1u
X8713 vss cap_series_gyp a_26768_7908# vss nmos_6p0 w=0.82u l=0.6u
X8714 a_9204_51874# cap_shunt_n a_8996_52220# vdd pmos_6p0 w=1.2u l=0.5u
X8715 vdd tune_shunt[6] a_24452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X8716 vss cap_shunt_p a_31808_23588# vss nmos_6p0 w=0.82u l=0.6u
X8717 a_15120_26724# cap_shunt_n a_13796_26786# vss nmos_6p0 w=0.82u l=0.6u
X8718 vss cap_shunt_p a_14112_18584# vss nmos_6p0 w=0.82u l=0.6u
X8719 vdd a_4492_3511# a_4404_3608# vdd pmos_6p0 w=1.22u l=1u
X8720 vdd tune_series_gy[4] a_24452_9884# vdd pmos_6p0 w=1.2u l=0.5u
X8721 a_22456_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8722 vdd a_1692_47848# a_1604_47892# vdd pmos_6p0 w=1.22u l=1u
X8723 a_34396_11784# a_34308_11828# vss vss nmos_6p0 w=0.82u l=1u
X8724 a_25780_20152# cap_series_gyp a_27496_20152# vss nmos_6p0 w=0.82u l=0.6u
X8725 a_20740_43672# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8726 vss tune_shunt[7] a_3828_23288# vss nmos_6p0 w=0.51u l=0.6u
X8727 a_3172_18100# cap_shunt_p a_3380_18584# vdd pmos_6p0 w=1.2u l=0.5u
X8728 a_25780_17016# cap_series_gyp a_25572_16532# vdd pmos_6p0 w=1.2u l=0.5u
X8729 vss tune_shunt[7] a_9428_17378# vss nmos_6p0 w=0.51u l=0.6u
X8730 a_3380_51512# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8731 vss cap_series_gygyp a_35840_4772# vss nmos_6p0 w=0.82u l=0.6u
X8732 a_25236_3612# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8733 vdd tune_shunt[7] a_17620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X8734 vss cap_shunt_p a_14112_15448# vss nmos_6p0 w=0.82u l=0.6u
X8735 vss tune_shunt[7] a_13460_21720# vss nmos_6p0 w=0.51u l=0.6u
X8736 vdd a_25548_49416# a_25460_49460# vdd pmos_6p0 w=1.22u l=1u
X8737 vss cap_shunt_n a_9072_34564# vss nmos_6p0 w=0.82u l=0.6u
X8738 vdd tune_series_gy[3] a_24452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X8739 a_22456_15448# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8740 a_23420_52552# a_23332_52596# vss vss nmos_6p0 w=0.82u l=1u
X8741 a_31260_47415# a_31172_47512# vss vss nmos_6p0 w=0.82u l=1u
X8742 vdd a_1692_44712# a_1604_44756# vdd pmos_6p0 w=1.22u l=1u
X8743 vss cap_shunt_n a_15904_43972# vss nmos_6p0 w=0.82u l=0.6u
X8744 vss tune_series_gy[5] a_22644_12312# vss nmos_6p0 w=0.51u l=0.6u
X8745 a_33948_55255# a_33860_55352# vss vss nmos_6p0 w=0.82u l=1u
X8746 a_20740_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8747 a_13252_32212# cap_shunt_n a_13460_32696# vdd pmos_6p0 w=1.2u l=0.5u
X8748 a_12768_4772# cap_series_gyp a_10660_4834# vss nmos_6p0 w=0.82u l=0.6u
X8749 vss tune_series_gy[5] a_25780_13880# vss nmos_6p0 w=0.51u l=0.6u
X8750 a_16252_49416# a_16164_49460# vss vss nmos_6p0 w=0.82u l=1u
X8751 a_3620_32212# cap_shunt_p a_3828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X8752 vss cap_shunt_n a_15120_22020# vss nmos_6p0 w=0.82u l=0.6u
X8753 a_34516_12674# cap_series_gygyp a_34308_13020# vdd pmos_6p0 w=1.2u l=0.5u
X8754 a_5544_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8755 a_28124_34871# a_28036_34968# vss vss nmos_6p0 w=0.82u l=1u
X8756 vdd tune_series_gy[2] a_14260_3612# vdd pmos_6p0 w=1.2u l=0.5u
X8757 a_30920_9476# cap_series_gyn a_29720_9884# vss nmos_6p0 w=0.82u l=0.6u
X8758 vdd a_25548_46280# a_25460_46324# vdd pmos_6p0 w=1.22u l=1u
X8759 vss cap_shunt_n a_9072_31428# vss nmos_6p0 w=0.82u l=0.6u
X8760 a_25572_24372# cap_shunt_p a_25780_24856# vdd pmos_6p0 w=1.2u l=0.5u
X8761 a_28484_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8762 vss cap_shunt_n a_15904_40836# vss nmos_6p0 w=0.82u l=0.6u
X8763 vss tune_shunt[7] a_9876_12312# vss nmos_6p0 w=0.51u l=0.6u
X8764 vss tune_shunt[7] a_13796_31490# vss nmos_6p0 w=0.51u l=0.6u
X8765 a_17828_29560# cap_shunt_n a_17620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X8766 vss tune_series_gy[4] a_25780_10744# vss nmos_6p0 w=0.51u l=0.6u
X8767 a_16500_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8768 a_13252_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8769 vss cap_shunt_n a_4256_10744# vss nmos_6p0 w=0.82u l=0.6u
X8770 a_28124_31735# a_28036_31832# vss vss nmos_6p0 w=0.82u l=1u
X8771 a_22680_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8772 a_18424_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8773 a_25572_21236# cap_shunt_p a_25780_21720# vdd pmos_6p0 w=1.2u l=0.5u
X8774 vdd a_34396_53687# a_34308_53784# vdd pmos_6p0 w=1.22u l=1u
X8775 a_28692_38968# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8776 a_32404_27132# cap_shunt_p a_32612_26786# vdd pmos_6p0 w=1.2u l=0.5u
X8777 a_18516_5556# cap_series_gyn a_18724_6040# vdd pmos_6p0 w=1.2u l=0.5u
X8778 a_3640_9476# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8779 a_12580_18100# cap_shunt_p a_12788_18584# vdd pmos_6p0 w=1.2u l=0.5u
X8780 a_25572_19668# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8781 a_21540_25564# cap_shunt_n a_21748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X8782 vss tune_series_gy[4] a_32632_14588# vss nmos_6p0 w=0.51u l=0.6u
X8783 a_16500_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8784 a_12992_45240# cap_shunt_n a_11668_45240# vss nmos_6p0 w=0.82u l=0.6u
X8785 a_31268_45240# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X8786 a_20532_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8787 a_22680_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8788 a_8848_43672# cap_shunt_p a_6740_43672# vss nmos_6p0 w=0.82u l=0.6u
X8789 a_20740_43672# cap_shunt_n a_20532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X8790 vdd a_34396_50551# a_34308_50648# vdd pmos_6p0 w=1.22u l=1u
X8791 a_13588_39676# cap_shunt_n a_13796_39330# vdd pmos_6p0 w=1.2u l=0.5u
X8792 a_36688_26424# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X8793 a_15532_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8794 a_21540_22428# cap_shunt_p a_21748_22082# vdd pmos_6p0 w=1.2u l=0.5u
X8795 vss tune_series_gy[3] a_32632_11452# vss nmos_6p0 w=0.51u l=0.6u
X8796 a_25572_33780# cap_shunt_p a_25780_34264# vdd pmos_6p0 w=1.2u l=0.5u
X8797 a_3380_51512# cap_shunt_n a_3172_51028# vdd pmos_6p0 w=1.2u l=0.5u
X8798 a_12992_42104# cap_shunt_n a_11668_42104# vss nmos_6p0 w=0.82u l=0.6u
X8799 a_20532_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8800 a_8848_40536# cap_shunt_n a_6740_40536# vss nmos_6p0 w=0.82u l=0.6u
X8801 a_21748_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8802 a_10340_36916# cap_shunt_n a_10548_37400# vdd pmos_6p0 w=1.2u l=0.5u
X8803 vss tune_series_gy[1] a_6760_3988# vss nmos_6p0 w=0.51u l=0.6u
X8804 vdd tune_shunt[7] a_7540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X8805 a_25572_30644# cap_shunt_p a_25780_31128# vdd pmos_6p0 w=1.2u l=0.5u
X8806 a_34516_22082# cap_series_gygyp a_35448_22020# vss nmos_6p0 w=0.82u l=0.6u
X8807 a_25996_52552# a_25908_52596# vss vss nmos_6p0 w=0.82u l=1u
X8808 a_21748_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8809 vss tune_shunt[7] a_16708_29922# vss nmos_6p0 w=0.51u l=0.6u
X8810 a_16700_47848# a_16612_47892# vss vss nmos_6p0 w=0.82u l=1u
X8811 vdd a_24204_40008# a_24116_40052# vdd pmos_6p0 w=1.22u l=1u
X8812 a_18816_18884# cap_shunt_p a_16708_18946# vss nmos_6p0 w=0.82u l=0.6u
X8813 a_18724_6040# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X8814 a_25780_35832# cap_shunt_p a_26712_35832# vss nmos_6p0 w=0.82u l=0.6u
X8815 vdd tune_shunt[7] a_7540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X8816 a_33524_27508# cap_shunt_p a_33732_27992# vdd pmos_6p0 w=1.2u l=0.5u
X8817 a_35056_35832# cap_shunt_n a_33732_35832# vss nmos_6p0 w=0.82u l=0.6u
X8818 a_3828_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8819 vdd tune_shunt[4] a_29492_23996# vdd pmos_6p0 w=1.2u l=0.5u
X8820 a_9316_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8821 a_15120_17316# cap_shunt_p a_13796_17378# vss nmos_6p0 w=0.82u l=0.6u
X8822 vdd a_22972_52552# a_22884_52596# vdd pmos_6p0 w=1.22u l=1u
X8823 a_32156_44279# a_32068_44376# vss vss nmos_6p0 w=0.82u l=1u
X8824 vss cap_shunt_n a_9072_28292# vss nmos_6p0 w=0.82u l=0.6u
X8825 vdd a_1692_38440# a_1604_38484# vdd pmos_6p0 w=1.22u l=1u
X8826 vss cap_series_gyp a_27104_9176# vss nmos_6p0 w=0.82u l=0.6u
X8827 a_18816_15748# cap_shunt_p a_16708_15810# vss nmos_6p0 w=0.82u l=0.6u
X8828 a_20740_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8829 a_28692_18584# cap_series_gyp a_28484_18100# vdd pmos_6p0 w=1.2u l=0.5u
X8830 vss cap_shunt_p a_5152_32696# vss nmos_6p0 w=0.82u l=0.6u
X8831 vss tune_series_gy[4] a_18612_6402# vss nmos_6p0 w=0.51u l=0.6u
X8832 a_3828_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8833 vss cap_shunt_n a_4032_12612# vss nmos_6p0 w=0.82u l=0.6u
X8834 a_32156_41143# a_32068_41240# vss vss nmos_6p0 w=0.82u l=1u
X8835 a_28124_28599# a_28036_28696# vss vss nmos_6p0 w=0.82u l=1u
X8836 vss cap_shunt_n a_9072_25156# vss nmos_6p0 w=0.82u l=0.6u
X8837 vss cap_shunt_n a_5488_51512# vss nmos_6p0 w=0.82u l=0.6u
X8838 vdd a_1692_35304# a_1604_35348# vdd pmos_6p0 w=1.22u l=1u
X8839 vss cap_shunt_n a_15904_34564# vss nmos_6p0 w=0.82u l=0.6u
X8840 vdd a_34844_25896# a_34756_25940# vdd pmos_6p0 w=1.22u l=1u
X8841 a_15804_16488# a_15716_16532# vss vss nmos_6p0 w=0.82u l=1u
X8842 a_13796_17378# cap_shunt_p a_13588_17724# vdd pmos_6p0 w=1.2u l=0.5u
X8843 vss cap_shunt_p a_11200_20152# vss nmos_6p0 w=0.82u l=0.6u
X8844 a_29700_39330# cap_shunt_p a_29492_39676# vdd pmos_6p0 w=1.2u l=0.5u
X8845 a_20740_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8846 vss cap_shunt_gyp a_35532_45540# vss nmos_6p0 w=0.82u l=0.6u
X8847 a_6740_13880# cap_shunt_p a_6532_13396# vdd pmos_6p0 w=1.2u l=0.5u
X8848 a_11144_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8849 a_12656_35832# cap_shunt_n a_10548_35832# vss nmos_6p0 w=0.82u l=0.6u
X8850 a_24204_32168# a_24116_32212# vss vss nmos_6p0 w=0.82u l=1u
X8851 a_9668_10260# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8852 a_28124_25463# a_28036_25560# vss vss nmos_6p0 w=0.82u l=1u
X8853 a_18424_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8854 vss cap_shunt_n a_15904_31428# vss nmos_6p0 w=0.82u l=0.6u
X8855 vdd a_34844_22760# a_34756_22804# vdd pmos_6p0 w=1.22u l=1u
X8856 a_3828_34264# cap_shunt_n a_3620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X8857 vss tune_shunt[7] a_13796_22082# vss nmos_6p0 w=0.51u l=0.6u
X8858 a_35880_19668# cap_series_gygyp a_35692_19668# vdd pmos_6p0 w=1.2u l=0.5u
X8859 a_17828_26424# cap_shunt_n a_17620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X8860 vss cap_shunt_gyn a_35532_42404# vss nmos_6p0 w=0.82u l=0.6u
X8861 a_21540_19292# cap_shunt_p a_21748_18946# vdd pmos_6p0 w=1.2u l=0.5u
X8862 a_16708_48738# cap_shunt_p a_18424_48676# vss nmos_6p0 w=0.82u l=0.6u
X8863 a_16500_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8864 a_30616_21236# cap_series_gygyn a_30428_21236# vdd pmos_6p0 w=1.2u l=0.5u
X8865 a_10340_3612# cap_series_gyn a_10548_3266# vdd pmos_6p0 w=1.2u l=0.5u
X8866 a_3172_18100# cap_shunt_p a_3380_18584# vdd pmos_6p0 w=1.2u l=0.5u
X8867 a_3828_31128# cap_shunt_n a_3620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X8868 a_17828_23288# cap_shunt_n a_17620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X8869 a_19732_7608# cap_series_gyp a_19524_7124# vdd pmos_6p0 w=1.2u l=0.5u
X8870 a_2708_12674# cap_shunt_n a_2500_13020# vdd pmos_6p0 w=1.2u l=0.5u
X8871 a_21540_16156# cap_series_gyn a_21748_15810# vdd pmos_6p0 w=1.2u l=0.5u
X8872 a_16500_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8873 a_20532_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8874 a_5276_54120# a_5188_54164# vss vss nmos_6p0 w=0.82u l=1u
X8875 vdd a_14012_53687# a_13924_53784# vdd pmos_6p0 w=1.22u l=1u
X8876 a_8848_34264# cap_shunt_n a_6740_34264# vss nmos_6p0 w=0.82u l=0.6u
X8877 a_13252_32212# cap_shunt_n a_13460_32696# vdd pmos_6p0 w=1.2u l=0.5u
X8878 vdd a_12892_17623# a_12804_17720# vdd pmos_6p0 w=1.22u l=1u
X8879 a_14580_46808# cap_shunt_p a_14372_46324# vdd pmos_6p0 w=1.2u l=0.5u
X8880 a_6760_3988# cap_series_gyp a_6784_4472# vss nmos_6p0 w=0.82u l=0.6u
X8881 a_36688_17016# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X8882 a_1716_7124# cap_shunt_n a_1924_7608# vdd pmos_6p0 w=1.2u l=0.5u
X8883 a_25572_24372# cap_shunt_p a_25780_24856# vdd pmos_6p0 w=1.2u l=0.5u
X8884 a_10092_5512# a_10004_5556# vss vss nmos_6p0 w=0.82u l=1u
X8885 vdd a_28348_41576# a_28260_41620# vdd pmos_6p0 w=1.22u l=1u
X8886 a_27496_38968# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X8887 a_13460_37400# cap_shunt_n a_14392_37400# vss nmos_6p0 w=0.82u l=0.6u
X8888 a_8848_31128# cap_shunt_n a_6740_31128# vss nmos_6p0 w=0.82u l=0.6u
X8889 a_21748_14242# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8890 a_10340_27508# cap_shunt_n a_10548_27992# vdd pmos_6p0 w=1.2u l=0.5u
X8891 a_20732_54120# a_20644_54164# vss vss nmos_6p0 w=0.82u l=1u
X8892 a_21748_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8893 a_35448_4772# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X8894 a_28484_32212# cap_shunt_p a_28692_32696# vdd pmos_6p0 w=1.2u l=0.5u
X8895 a_24652_47415# a_24564_47512# vss vss nmos_6p0 w=0.82u l=1u
X8896 a_25780_29560# cap_shunt_p a_26712_29560# vss nmos_6p0 w=0.82u l=0.6u
X8897 vdd tune_shunt[7] a_24452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X8898 vdd tune_shunt[7] a_7540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X8899 a_28692_9176# cap_series_gyn a_29624_9176# vss nmos_6p0 w=0.82u l=0.6u
X8900 a_25572_21236# cap_shunt_p a_25780_21720# vdd pmos_6p0 w=1.2u l=0.5u
X8901 a_35180_34871# a_35092_34968# vss vss nmos_6p0 w=0.82u l=1u
X8902 a_35056_29560# cap_shunt_p a_33732_29560# vss nmos_6p0 w=0.82u l=0.6u
X8903 a_21748_11106# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X8904 a_31808_37700# cap_shunt_n a_29700_37762# vss nmos_6p0 w=0.82u l=0.6u
X8905 a_3620_43188# cap_shunt_p a_3828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X8906 a_21748_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X8907 a_29492_23996# cap_shunt_p a_29700_23650# vdd pmos_6p0 w=1.2u l=0.5u
X8908 a_9668_14964# cap_shunt_p a_9876_15448# vdd pmos_6p0 w=1.2u l=0.5u
X8909 vdd a_12220_55688# a_12132_55732# vdd pmos_6p0 w=1.22u l=1u
X8910 vdd a_6956_44279# a_6868_44376# vdd pmos_6p0 w=1.22u l=1u
X8911 a_25780_26424# cap_shunt_p a_26712_26424# vss nmos_6p0 w=0.82u l=0.6u
X8912 vdd a_12556_9783# a_12468_9880# vdd pmos_6p0 w=1.22u l=1u
X8913 a_20284_49416# a_20196_49460# vss vss nmos_6p0 w=0.82u l=1u
X8914 a_7580_5180# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8915 a_18492_8648# a_18404_8692# vss vss nmos_6p0 w=0.82u l=1u
X8916 a_35180_31735# a_35092_31832# vss vss nmos_6p0 w=0.82u l=1u
X8917 a_15532_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8918 a_35264_45944# cap_shunt_gyp a_35264_45540# vdd pmos_6p0 w=1.215u l=0.5u
X8919 a_24540_3944# a_24452_3988# vss vss nmos_6p0 w=0.82u l=1u
X8920 vdd tune_series_gy[5] a_29492_14588# vdd pmos_6p0 w=1.2u l=0.5u
X8921 a_9856_32996# cap_shunt_n a_7748_33058# vss nmos_6p0 w=0.82u l=0.6u
X8922 a_25572_33780# cap_shunt_p a_25780_34264# vdd pmos_6p0 w=1.2u l=0.5u
X8923 vdd a_1692_29032# a_1604_29076# vdd pmos_6p0 w=1.22u l=1u
X8924 vss cap_shunt_n a_15904_28292# vss nmos_6p0 w=0.82u l=0.6u
X8925 a_9668_11828# cap_shunt_p a_9876_12312# vdd pmos_6p0 w=1.2u l=0.5u
X8926 vdd a_32716_47848# a_32628_47892# vdd pmos_6p0 w=1.22u l=1u
X8927 a_27888_6040# cap_series_gyp a_25780_6040# vss nmos_6p0 w=0.82u l=0.6u
X8928 vdd a_27788_53687# a_27700_53784# vdd pmos_6p0 w=1.22u l=1u
X8929 a_10340_36916# cap_shunt_n a_10548_37400# vdd pmos_6p0 w=1.2u l=0.5u
X8930 a_12656_29560# cap_shunt_n a_10548_29560# vss nmos_6p0 w=0.82u l=0.6u
X8931 vss cap_shunt_p a_5152_23288# vss nmos_6p0 w=0.82u l=0.6u
X8932 vss cap_series_gyn a_25984_9476# vss nmos_6p0 w=0.82u l=0.6u
X8933 a_35264_42808# cap_shunt_gyn a_35264_42404# vdd pmos_6p0 w=1.215u l=0.5u
X8934 vdd tune_shunt[7] a_9668_13396# vdd pmos_6p0 w=1.2u l=0.5u
X8935 a_22644_10744# cap_series_gyp a_22436_10260# vdd pmos_6p0 w=1.2u l=0.5u
X8936 a_3620_13396# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8937 a_25572_30644# cap_shunt_p a_25780_31128# vdd pmos_6p0 w=1.2u l=0.5u
X8938 a_17640_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8939 vss cap_shunt_n a_15904_25156# vss nmos_6p0 w=0.82u l=0.6u
X8940 a_24452_8316# cap_series_gyp a_24660_7970# vdd pmos_6p0 w=1.2u l=0.5u
X8941 vdd a_34844_16488# a_34756_16532# vdd pmos_6p0 w=1.22u l=1u
X8942 vss cap_series_gyn a_23968_12312# vss nmos_6p0 w=0.82u l=0.6u
X8943 vdd a_8412_54120# a_8324_54164# vdd pmos_6p0 w=1.22u l=1u
X8944 vdd a_27788_50551# a_27700_50648# vdd pmos_6p0 w=1.22u l=1u
X8945 a_12656_26424# cap_shunt_n a_10548_26424# vss nmos_6p0 w=0.82u l=0.6u
X8946 a_24204_22760# a_24116_22804# vss vss nmos_6p0 w=0.82u l=1u
X8947 a_16500_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8948 a_4032_18884# cap_shunt_p a_2708_18946# vss nmos_6p0 w=0.82u l=0.6u
X8949 vss cap_series_gyp a_23744_6040# vss nmos_6p0 w=0.82u l=0.6u
X8950 a_3036_19624# a_2948_19668# vss vss nmos_6p0 w=0.82u l=1u
X8951 a_17640_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X8952 a_3828_24856# cap_shunt_p a_3620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X8953 a_24452_5180# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8954 a_17828_17016# cap_shunt_p a_17620_16532# vdd pmos_6p0 w=1.2u l=0.5u
X8955 a_16252_52119# a_16164_52216# vss vss nmos_6p0 w=0.82u l=1u
X8956 vdd a_35292_36872# a_35204_36916# vdd pmos_6p0 w=1.22u l=1u
X8957 vss cap_series_gyp a_33048_14180# vss nmos_6p0 w=0.82u l=0.6u
X8958 a_16708_39330# cap_shunt_n a_18424_39268# vss nmos_6p0 w=0.82u l=0.6u
X8959 a_16500_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8960 a_4032_15748# cap_shunt_p a_2708_15810# vss nmos_6p0 w=0.82u l=0.6u
X8961 vdd a_20172_31735# a_20084_31832# vdd pmos_6p0 w=1.22u l=1u
X8962 a_30140_43144# a_30052_43188# vss vss nmos_6p0 w=0.82u l=1u
X8963 a_17620_43188# cap_shunt_p a_17828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X8964 a_26768_39268# cap_shunt_p a_24660_39330# vss nmos_6p0 w=0.82u l=0.6u
X8965 a_28572_44279# a_28484_44376# vss vss nmos_6p0 w=0.82u l=1u
X8966 vdd a_31260_40008# a_31172_40052# vdd pmos_6p0 w=1.22u l=1u
X8967 a_3828_21720# cap_shunt_p a_3620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X8968 a_32404_36540# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8969 vss cap_series_gyp a_33048_11044# vss nmos_6p0 w=0.82u l=0.6u
X8970 a_13796_17378# cap_shunt_p a_13588_17724# vdd pmos_6p0 w=1.2u l=0.5u
X8971 a_13796_47170# cap_shunt_p a_13588_47516# vdd pmos_6p0 w=1.2u l=0.5u
X8972 a_29700_39330# cap_shunt_p a_29492_39676# vdd pmos_6p0 w=1.2u l=0.5u
X8973 a_16708_22082# cap_shunt_n a_17640_22020# vss nmos_6p0 w=0.82u l=0.6u
X8974 vss cap_series_gyn a_26768_18884# vss nmos_6p0 w=0.82u l=0.6u
X8975 vdd a_14796_55688# a_14708_55732# vdd pmos_6p0 w=1.22u l=1u
X8976 vdd a_37868_55255# a_37780_55352# vdd pmos_6p0 w=1.22u l=1u
X8977 a_8064_46808# cap_shunt_p a_6740_46808# vss nmos_6p0 w=0.82u l=0.6u
X8978 a_28572_41143# a_28484_41240# vss vss nmos_6p0 w=0.82u l=1u
X8979 a_36188_3511# a_36100_3608# vss vss nmos_6p0 w=0.82u l=1u
X8980 a_6740_13880# cap_shunt_p a_6532_13396# vdd pmos_6p0 w=1.2u l=0.5u
X8981 a_33500_49416# a_33412_49460# vss vss nmos_6p0 w=0.82u l=1u
X8982 a_6740_20152# cap_shunt_p a_6532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X8983 a_32404_33404# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X8984 vdd a_23420_49416# a_23332_49460# vdd pmos_6p0 w=1.22u l=1u
X8985 vdd a_18492_55255# a_18404_55352# vdd pmos_6p0 w=1.22u l=1u
X8986 a_21748_37762# cap_shunt_n a_21540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X8987 a_35180_28599# a_35092_28696# vss vss nmos_6p0 w=0.82u l=1u
X8988 vss tune_series_gy[3] a_18388_3266# vss nmos_6p0 w=0.51u l=0.6u
X8989 vss cap_series_gyn a_26768_15748# vss nmos_6p0 w=0.82u l=0.6u
X8990 vdd a_37868_52119# a_37780_52216# vdd pmos_6p0 w=1.22u l=1u
X8991 vdd tune_shunt[4] a_17620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X8992 a_18388_3266# cap_series_gyn a_20104_3204# vss nmos_6p0 w=0.82u l=0.6u
X8993 a_5844_10744# cap_shunt_p a_6776_10744# vss nmos_6p0 w=0.82u l=0.6u
X8994 a_27676_12919# a_27588_13016# vss vss nmos_6p0 w=0.82u l=1u
X8995 a_33500_46280# a_33412_46324# vss vss nmos_6p0 w=0.82u l=1u
X8996 a_21748_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X8997 a_5844_3266# cap_shunt_n a_5636_3612# vdd pmos_6p0 w=1.2u l=0.5u
X8998 vdd a_33500_10216# a_33412_10260# vdd pmos_6p0 w=1.22u l=1u
X8999 a_30616_21236# cap_series_gygyn a_30428_21236# vdd pmos_6p0 w=1.2u l=0.5u
X9000 a_31260_32168# a_31172_32212# vss vss nmos_6p0 w=0.82u l=1u
X9001 vdd a_18492_52119# a_18404_52216# vdd pmos_6p0 w=1.22u l=1u
X9002 a_16028_35304# a_15940_35348# vss vss nmos_6p0 w=0.82u l=1u
X9003 a_35180_25463# a_35092_25560# vss vss nmos_6p0 w=0.82u l=1u
X9004 vss tune_series_gygy[1] a_34516_4834# vss nmos_6p0 w=0.51u l=0.6u
X9005 a_16700_53687# a_16612_53784# vss vss nmos_6p0 w=0.82u l=1u
X9006 vdd tune_shunt[6] a_17620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X9007 vdd a_35740_38440# a_35652_38484# vdd pmos_6p0 w=1.22u l=1u
X9008 a_29492_14588# cap_series_gyp a_29700_14242# vdd pmos_6p0 w=1.2u l=0.5u
X9009 a_21748_25218# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9010 vss cap_series_gygyn a_31032_20152# vss nmos_6p0 w=0.82u l=0.6u
X9011 a_24752_7608# cap_series_gyp a_22644_7608# vss nmos_6p0 w=0.82u l=0.6u
X9012 a_15700_4834# cap_series_gyn a_15492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X9013 a_25780_17016# cap_series_gyp a_26712_17016# vss nmos_6p0 w=0.82u l=0.6u
X9014 vss tune_shunt[7] a_24660_26786# vss nmos_6p0 w=0.51u l=0.6u
X9015 a_18180_3612# cap_series_gyn a_18388_3266# vdd pmos_6p0 w=1.2u l=0.5u
X9016 a_6740_53080# cap_shunt_n a_6532_52596# vdd pmos_6p0 w=1.2u l=0.5u
X9017 a_21524_3266# cap_series_gyp a_21316_3612# vdd pmos_6p0 w=1.2u l=0.5u
X9018 a_14580_46808# cap_shunt_p a_14372_46324# vdd pmos_6p0 w=1.2u l=0.5u
X9019 a_6572_7124# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9020 a_34516_17378# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9021 a_20532_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9022 a_25572_24372# cap_shunt_p a_25780_24856# vdd pmos_6p0 w=1.2u l=0.5u
X9023 a_9856_23588# cap_shunt_p a_7748_23650# vss nmos_6p0 w=0.82u l=0.6u
X9024 vdd a_20620_30167# a_20532_30264# vdd pmos_6p0 w=1.22u l=1u
X9025 a_27452_45847# a_27364_45944# vss vss nmos_6p0 w=0.82u l=1u
X9026 a_10340_27508# cap_shunt_n a_10548_27992# vdd pmos_6p0 w=1.2u l=0.5u
X9027 vss tune_series_gy[4] a_11800_8692# vss nmos_6p0 w=0.51u l=0.6u
X9028 a_13588_34972# cap_shunt_n a_13796_34626# vdd pmos_6p0 w=1.2u l=0.5u
X9029 a_7540_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9030 a_21524_3266# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X9031 vss tune_shunt[6] a_13796_45602# vss nmos_6p0 w=0.51u l=0.6u
X9032 vdd tune_shunt[7] a_13252_38484# vdd pmos_6p0 w=1.2u l=0.5u
X9033 a_28484_32212# cap_shunt_p a_28692_32696# vdd pmos_6p0 w=1.2u l=0.5u
X9034 a_26768_6340# cap_series_gyn a_24660_6402# vss nmos_6p0 w=0.82u l=0.6u
X9035 a_11256_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9036 vss tune_shunt[5] a_12788_20152# vss nmos_6p0 w=0.51u l=0.6u
X9037 a_25780_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9038 a_20532_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9039 a_25572_21236# cap_shunt_p a_25780_21720# vdd pmos_6p0 w=1.2u l=0.5u
X9040 vdd a_18604_50551# a_18516_50648# vdd pmos_6p0 w=1.22u l=1u
X9041 a_10660_29922# cap_shunt_n a_12376_29860# vss nmos_6p0 w=0.82u l=0.6u
X9042 a_30800_9176# cap_series_gyn a_28692_9176# vss nmos_6p0 w=0.82u l=0.6u
X9043 a_36188_55688# a_36100_55732# vss vss nmos_6p0 w=0.82u l=1u
X9044 vdd a_1692_55255# a_1604_55352# vdd pmos_6p0 w=1.22u l=1u
X9045 a_13588_31836# cap_shunt_n a_13796_31490# vdd pmos_6p0 w=1.2u l=0.5u
X9046 a_36720_49461# cap_shunt_gyp a_36720_50006# vdd pmos_6p0 w=1.215u l=0.5u
X9047 vdd a_20172_25463# a_20084_25560# vdd pmos_6p0 w=1.22u l=1u
X9048 vss tune_shunt[7] a_9428_17378# vss nmos_6p0 w=0.51u l=0.6u
X9049 a_26768_3204# cap_shunt_p a_25444_3266# vss nmos_6p0 w=0.82u l=0.6u
X9050 a_11256_11044# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9051 a_25780_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9052 vdd tune_shunt[7] a_13252_35348# vdd pmos_6p0 w=1.2u l=0.5u
X9053 a_17640_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9054 vdd a_25996_49416# a_25908_49460# vdd pmos_6p0 w=1.22u l=1u
X9055 a_10660_26786# cap_shunt_n a_12376_26724# vss nmos_6p0 w=0.82u l=0.6u
X9056 a_2708_44034# cap_shunt_p a_4424_43972# vss nmos_6p0 w=0.82u l=0.6u
X9057 a_2500_20860# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9058 vdd a_1692_52119# a_1604_52216# vdd pmos_6p0 w=1.22u l=1u
X9059 a_36720_46325# cap_shunt_gyp a_36720_46870# vdd pmos_6p0 w=1.215u l=0.5u
X9060 a_2708_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9061 vdd a_20172_22327# a_20084_22424# vdd pmos_6p0 w=1.22u l=1u
X9062 vdd tune_shunt[7] a_10452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X9063 a_6740_32696# cap_shunt_n a_7672_32696# vss nmos_6p0 w=0.82u l=0.6u
X9064 vdd a_25996_46280# a_25908_46324# vdd pmos_6p0 w=1.22u l=1u
X9065 a_28572_34871# a_28484_34968# vss vss nmos_6p0 w=0.82u l=1u
X9066 a_2708_40898# cap_shunt_p a_4424_40836# vss nmos_6p0 w=0.82u l=0.6u
X9067 a_32404_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9068 a_7768_6748# cap_series_gyp a_7580_6748# vdd pmos_6p0 w=1.2u l=0.5u
X9069 a_7540_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9070 a_9332_14588# cap_shunt_p a_9540_14242# vdd pmos_6p0 w=1.2u l=0.5u
X9071 a_1692_33303# a_1604_33400# vss vss nmos_6p0 w=0.82u l=1u
X9072 a_12788_20152# cap_shunt_p a_13720_20152# vss nmos_6p0 w=0.82u l=0.6u
X9073 a_29624_40536# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9074 vdd a_18044_54120# a_17956_54164# vdd pmos_6p0 w=1.22u l=1u
X9075 a_13796_37762# cap_shunt_n a_13588_38108# vdd pmos_6p0 w=1.2u l=0.5u
X9076 a_21748_29922# cap_shunt_n a_21540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X9077 a_28572_31735# a_28484_31832# vss vss nmos_6p0 w=0.82u l=1u
X9078 a_22644_9176# cap_series_gyp a_22436_8692# vdd pmos_6p0 w=1.2u l=0.5u
X9079 a_35692_36916# cap_series_gygyp a_35880_36916# vdd pmos_6p0 w=1.2u l=0.5u
X9080 a_8748_55688# a_8660_55732# vss vss nmos_6p0 w=0.82u l=1u
X9081 a_16028_29032# a_15940_29076# vss vss nmos_6p0 w=0.82u l=1u
X9082 a_21316_3988# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9083 vdd tune_series_gy[4] a_11612_8692# vdd pmos_6p0 w=1.2u l=0.5u
X9084 vdd a_18044_50984# a_17956_51028# vdd pmos_6p0 w=1.22u l=1u
X9085 a_20620_48983# a_20532_49080# vss vss nmos_6p0 w=0.82u l=1u
X9086 vdd tune_shunt[6] a_16500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X9087 a_29700_14242# cap_series_gyp a_31416_14180# vss nmos_6p0 w=0.82u l=0.6u
X9088 vdd tune_shunt[6] a_17620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X9089 vdd a_19276_34871# a_19188_34968# vdd pmos_6p0 w=1.22u l=1u
X9090 a_16708_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9091 vdd a_3036_25896# a_2948_25940# vdd pmos_6p0 w=1.22u l=1u
X9092 vdd tune_series_gygy[5] a_35692_18100# vdd pmos_6p0 w=1.2u l=0.5u
X9093 a_31260_22760# a_31172_22804# vss vss nmos_6p0 w=0.82u l=1u
X9094 a_28484_10260# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9095 a_16028_25896# a_15940_25940# vss vss nmos_6p0 w=0.82u l=1u
X9096 a_35880_14964# cap_series_gygyn a_35692_14964# vdd pmos_6p0 w=1.2u l=0.5u
X9097 vss tune_shunt[7] a_2708_15810# vss nmos_6p0 w=0.51u l=0.6u
X9098 vdd a_28236_47415# a_28148_47512# vdd pmos_6p0 w=1.22u l=1u
X9099 a_37868_23895# a_37780_23992# vss vss nmos_6p0 w=0.82u l=1u
X9100 a_29700_11106# cap_series_gyp a_31416_11044# vss nmos_6p0 w=0.82u l=0.6u
X9101 vdd tune_shunt[7] a_17620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X9102 a_6084_49084# cap_shunt_p a_6292_48738# vdd pmos_6p0 w=1.2u l=0.5u
X9103 a_34748_46808# cap_shunt_gyn a_34480_46870# vss nmos_6p0 w=0.82u l=0.6u
X9104 vdd a_3036_22760# a_2948_22804# vdd pmos_6p0 w=1.22u l=1u
X9105 vdd a_4492_5512# a_4404_5556# vdd pmos_6p0 w=1.22u l=1u
X9106 a_13796_47170# cap_shunt_p a_13588_47516# vdd pmos_6p0 w=1.2u l=0.5u
X9107 a_19544_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9108 a_23352_6040# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X9109 vss tune_series_gy[5] a_24660_17378# vss nmos_6p0 w=0.51u l=0.6u
X9110 a_35880_11828# cap_series_gygyp a_35692_11828# vdd pmos_6p0 w=1.2u l=0.5u
X9111 a_6740_43672# cap_shunt_p a_6532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X9112 a_25780_42104# cap_shunt_n a_25572_41620# vdd pmos_6p0 w=1.2u l=0.5u
X9113 a_13796_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9114 a_14692_7608# cap_series_gyp a_14484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X9115 a_13104_4472# cap_series_gyp a_11780_4472# vss nmos_6p0 w=0.82u l=0.6u
X9116 vss tune_shunt[7] a_13796_39330# vss nmos_6p0 w=0.51u l=0.6u
X9117 a_35292_5512# a_35204_5556# vss vss nmos_6p0 w=0.82u l=1u
X9118 vdd a_2588_13352# a_2500_13396# vdd pmos_6p0 w=1.22u l=1u
X9119 a_30016_38968# cap_shunt_n a_28692_38968# vss nmos_6p0 w=0.82u l=0.6u
X9120 a_5152_37400# cap_shunt_n a_3828_37400# vss nmos_6p0 w=0.82u l=0.6u
X9121 vss cap_shunt_p a_30016_32696# vss nmos_6p0 w=0.82u l=0.6u
X9122 a_21748_7970# cap_series_gyp a_23464_7908# vss nmos_6p0 w=0.82u l=0.6u
X9123 a_20532_24372# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9124 a_7952_9176# cap_shunt_p a_5844_9176# vss nmos_6p0 w=0.82u l=0.6u
X9125 a_14692_10744# cap_series_gyn a_16408_10744# vss nmos_6p0 w=0.82u l=0.6u
X9126 vdd a_24652_40008# a_24564_40052# vdd pmos_6p0 w=1.22u l=1u
X9127 a_20284_52119# a_20196_52216# vss vss nmos_6p0 w=0.82u l=1u
X9128 a_10340_25940# cap_shunt_n a_10548_26424# vdd pmos_6p0 w=1.2u l=0.5u
X9129 vdd a_1692_48983# a_1604_49080# vdd pmos_6p0 w=1.22u l=1u
X9130 a_13588_25564# cap_shunt_n a_13796_25218# vdd pmos_6p0 w=1.2u l=0.5u
X9131 a_14580_42104# cap_shunt_n a_14372_41620# vdd pmos_6p0 w=1.2u l=0.5u
X9132 a_35628_36439# a_35540_36536# vss vss nmos_6p0 w=0.82u l=1u
X9133 a_13720_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9134 a_27004_55688# a_26916_55732# vss vss nmos_6p0 w=0.82u l=1u
X9135 vdd tune_shunt[7] a_13252_29076# vdd pmos_6p0 w=1.2u l=0.5u
X9136 a_25780_12312# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9137 a_20532_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9138 a_31708_40008# a_31620_40052# vss vss nmos_6p0 w=0.82u l=1u
X9139 a_10340_22804# cap_shunt_n a_10548_23288# vdd pmos_6p0 w=1.2u l=0.5u
X9140 vss tune_shunt[4] a_33732_35832# vss nmos_6p0 w=0.51u l=0.6u
X9141 a_13588_22428# cap_shunt_n a_13796_22082# vdd pmos_6p0 w=1.2u l=0.5u
X9142 vss cap_shunt_p a_22848_20152# vss nmos_6p0 w=0.82u l=0.6u
X9143 vdd a_20172_16055# a_20084_16152# vdd pmos_6p0 w=1.22u l=1u
X9144 vss cap_shunt_p a_18032_45540# vss nmos_6p0 w=0.82u l=0.6u
X9145 a_13720_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9146 vss tune_shunt[5] a_6292_50306# vss nmos_6p0 w=0.51u l=0.6u
X9147 a_28572_28599# a_28484_28696# vss vss nmos_6p0 w=0.82u l=1u
X9148 vdd a_17708_12919# a_17620_13016# vdd pmos_6p0 w=1.22u l=1u
X9149 a_9204_51874# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9150 a_2708_34626# cap_shunt_n a_4424_34564# vss nmos_6p0 w=0.82u l=0.6u
X9151 a_5636_3612# cap_shunt_n a_5844_3266# vdd pmos_6p0 w=1.2u l=0.5u
X9152 a_2500_11452# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9153 a_29624_34264# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9154 a_14728_22020# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9155 vss cap_shunt_n a_18032_42404# vss nmos_6p0 w=0.82u l=0.6u
X9156 a_24652_32168# a_24564_32212# vss vss nmos_6p0 w=0.82u l=1u
X9157 vss tune_shunt[7] a_29700_26786# vss nmos_6p0 w=0.51u l=0.6u
X9158 a_6740_23288# cap_shunt_p a_7672_23288# vss nmos_6p0 w=0.82u l=0.6u
X9159 a_26376_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9160 a_28572_25463# a_28484_25560# vss vss nmos_6p0 w=0.82u l=1u
X9161 a_2708_31490# cap_shunt_p a_4424_31428# vss nmos_6p0 w=0.82u l=0.6u
X9162 a_28484_32212# cap_shunt_p a_28692_32696# vdd pmos_6p0 w=1.2u l=0.5u
X9163 a_1692_23895# a_1604_23992# vss vss nmos_6p0 w=0.82u l=1u
X9164 a_19732_7608# cap_series_gyp a_19524_7124# vdd pmos_6p0 w=1.2u l=0.5u
X9165 a_35880_3988# cap_series_gygyp a_35692_3988# vdd pmos_6p0 w=1.2u l=0.5u
X9166 vdd a_34396_52552# a_34308_52596# vdd pmos_6p0 w=1.22u l=1u
X9167 a_29624_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9168 a_16708_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9169 a_21748_28354# cap_shunt_n a_21540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X9170 a_2724_10260# cap_shunt_n a_2932_10744# vdd pmos_6p0 w=1.2u l=0.5u
X9171 vdd tune_shunt[7] a_16500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X9172 a_28692_4472# cap_series_gyp a_28484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X9173 vdd a_8412_9783# a_8324_9880# vdd pmos_6p0 w=1.22u l=1u
X9174 a_29492_5180# cap_shunt_p a_29700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X9175 a_20732_53687# a_20644_53784# vss vss nmos_6p0 w=0.82u l=1u
X9176 a_13788_50984# a_13700_51028# vss vss nmos_6p0 w=0.82u l=1u
X9177 a_29700_29922# cap_shunt_p a_30632_29860# vss nmos_6p0 w=0.82u l=0.6u
X9178 vdd a_19276_28599# a_19188_28696# vdd pmos_6p0 w=1.22u l=1u
X9179 a_6292_18584# cap_shunt_p a_7224_18584# vss nmos_6p0 w=0.82u l=0.6u
X9180 a_9108_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9181 a_24452_9884# cap_series_gyn a_24660_9538# vdd pmos_6p0 w=1.2u l=0.5u
X9182 vss tune_shunt[6] a_6740_35832# vss nmos_6p0 w=0.51u l=0.6u
X9183 a_20620_39575# a_20532_39672# vss vss nmos_6p0 w=0.82u l=1u
X9184 vdd tune_shunt[7] a_16500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X9185 a_20740_18584# cap_shunt_p a_20532_18100# vdd pmos_6p0 w=1.2u l=0.5u
X9186 a_11592_53080# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9187 a_10548_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9188 vdd tune_shunt[7] a_12580_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9189 a_9876_17016# cap_shunt_p a_9668_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9190 vdd a_24204_19624# a_24116_19668# vdd pmos_6p0 w=1.22u l=1u
X9191 vdd a_14460_53687# a_14372_53784# vdd pmos_6p0 w=1.22u l=1u
X9192 vdd tune_shunt[7] a_17620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X9193 a_33500_52119# a_33412_52216# vss vss nmos_6p0 w=0.82u l=1u
X9194 a_29700_26786# cap_shunt_p a_30632_26724# vss nmos_6p0 w=0.82u l=0.6u
X9195 a_14504_13880# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9196 a_16708_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9197 a_24452_6748# cap_series_gyn a_24660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X9198 vdd a_8412_3511# a_8324_3608# vdd pmos_6p0 w=1.22u l=1u
X9199 a_14692_6040# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X9200 a_33732_34264# cap_shunt_n a_33524_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9201 a_9332_14588# cap_shunt_p a_9540_14242# vdd pmos_6p0 w=1.2u l=0.5u
X9202 vdd a_28796_41576# a_28708_41620# vdd pmos_6p0 w=1.22u l=1u
X9203 a_7748_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9204 vss tune_shunt[7] a_2708_29922# vss nmos_6p0 w=0.51u l=0.6u
X9205 a_34516_15810# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9206 a_19544_23288# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9207 a_13796_37762# cap_shunt_n a_13588_38108# vdd pmos_6p0 w=1.2u l=0.5u
X9208 a_6532_36916# cap_shunt_n a_6740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X9209 a_21748_29922# cap_shunt_n a_21540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X9210 a_37444_50648# cap_shunt_gyn a_37632_50648# vdd pmos_6p0 w=1.215u l=0.5u
X9211 a_25780_32696# cap_shunt_p a_25572_32212# vdd pmos_6p0 w=1.2u l=0.5u
X9212 a_13588_19292# cap_shunt_p a_13796_18946# vdd pmos_6p0 w=1.2u l=0.5u
X9213 a_13796_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9214 a_33732_31128# cap_shunt_n a_33524_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9215 vss cap_shunt_p a_30016_23288# vss nmos_6p0 w=0.82u l=0.6u
X9216 a_11460_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9217 a_36300_35304# a_36212_35348# vss vss nmos_6p0 w=0.82u l=1u
X9218 a_11984_4772# cap_series_gyp a_10660_4834# vss nmos_6p0 w=0.82u l=0.6u
X9219 vdd tune_shunt[6] a_16500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X9220 a_31708_33736# a_31620_33780# vss vss nmos_6p0 w=0.82u l=1u
X9221 a_13796_22082# cap_shunt_n a_15512_22020# vss nmos_6p0 w=0.82u l=0.6u
X9222 vdd a_35740_55255# a_35652_55352# vdd pmos_6p0 w=1.22u l=1u
X9223 a_10452_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9224 a_23856_22020# cap_shunt_p a_21748_22082# vss nmos_6p0 w=0.82u l=0.6u
X9225 vss tune_shunt[7] a_33732_29560# vss nmos_6p0 w=0.51u l=0.6u
X9226 a_13588_16156# cap_shunt_p a_13796_15810# vdd pmos_6p0 w=1.2u l=0.5u
X9227 a_36512_41621# cap_shunt_gyn a_36324_41621# vdd pmos_6p0 w=1.215u l=0.5u
X9228 vdd tune_series_gygy[5] a_35692_18100# vdd pmos_6p0 w=1.2u l=0.5u
X9229 a_3620_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9230 vdd a_29468_41143# a_29380_41240# vdd pmos_6p0 w=1.22u l=1u
X9231 a_2140_30167# a_2052_30264# vss vss nmos_6p0 w=0.82u l=1u
X9232 a_9668_52596# cap_shunt_n a_9876_53080# vdd pmos_6p0 w=1.2u l=0.5u
X9233 a_22436_8692# cap_series_gyp a_22644_9176# vdd pmos_6p0 w=1.2u l=0.5u
X9234 a_35880_14964# cap_series_gygyn a_35692_14964# vdd pmos_6p0 w=1.2u l=0.5u
X9235 vss cap_shunt_p a_5936_45240# vss nmos_6p0 w=0.82u l=0.6u
X9236 a_31708_30600# a_31620_30644# vss vss nmos_6p0 w=0.82u l=1u
X9237 a_2708_28354# cap_shunt_n a_4424_28292# vss nmos_6p0 w=0.82u l=0.6u
X9238 vdd a_35740_52119# a_35652_52216# vdd pmos_6p0 w=1.22u l=1u
X9239 vdd tune_shunt[4] a_20532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X9240 a_31624_8316# cap_series_gygyn a_31436_8316# vdd pmos_6p0 w=1.2u l=0.5u
X9241 a_18180_3612# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9242 a_13588_20860# cap_shunt_n a_13796_20514# vdd pmos_6p0 w=1.2u l=0.5u
X9243 a_6084_49084# cap_shunt_p a_6292_48738# vdd pmos_6p0 w=1.2u l=0.5u
X9244 a_22456_43672# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9245 vss cap_shunt_n a_18032_36132# vss nmos_6p0 w=0.82u l=0.6u
X9246 a_19524_13396# cap_series_gyn a_19732_13880# vdd pmos_6p0 w=1.2u l=0.5u
X9247 vdd a_22076_54120# a_21988_54164# vdd pmos_6p0 w=1.22u l=1u
X9248 a_2140_27031# a_2052_27128# vss vss nmos_6p0 w=0.82u l=1u
X9249 a_3640_12612# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9250 a_28236_52552# a_28148_52596# vss vss nmos_6p0 w=0.82u l=1u
X9251 a_26376_36132# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9252 a_1924_7970# cap_shunt_n a_1716_8316# vdd pmos_6p0 w=1.2u l=0.5u
X9253 a_31708_8648# a_31620_8692# vss vss nmos_6p0 w=0.82u l=1u
X9254 a_35880_11828# cap_series_gygyp a_35692_11828# vdd pmos_6p0 w=1.2u l=0.5u
X9255 vss cap_shunt_p a_5936_42104# vss nmos_6p0 w=0.82u l=0.6u
X9256 a_25780_42104# cap_shunt_n a_25572_41620# vdd pmos_6p0 w=1.2u l=0.5u
X9257 a_2708_25218# cap_shunt_p a_4424_25156# vss nmos_6p0 w=0.82u l=0.6u
X9258 a_29700_4834# tune_shunt[0] vss vss nmos_6p0 w=0.51u l=0.6u
X9259 vss tune_shunt[5] a_21748_44034# vss nmos_6p0 w=0.51u l=0.6u
X9260 a_37632_33781# cap_shunt_gyn a_37444_33781# vdd pmos_6p0 w=1.215u l=0.5u
X9261 vdd a_21516_55255# a_21428_55352# vdd pmos_6p0 w=1.22u l=1u
X9262 a_22456_40536# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9263 a_24452_5180# cap_series_gyp a_24660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X9264 vdd a_8860_54120# a_8772_54164# vdd pmos_6p0 w=1.22u l=1u
X9265 vdd a_22076_50984# a_21988_51028# vdd pmos_6p0 w=1.22u l=1u
X9266 a_24652_22760# a_24564_22804# vss vss nmos_6p0 w=0.82u l=1u
X9267 vss tune_series_gy[4] a_29700_17378# vss nmos_6p0 w=0.51u l=0.6u
X9268 a_19388_55255# a_19300_55352# vss vss nmos_6p0 w=0.82u l=1u
X9269 a_17620_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9270 a_37080_26424# cap_series_gygyp a_35880_25940# vss nmos_6p0 w=0.82u l=0.6u
X9271 vss cap_shunt_p a_11536_20452# vss nmos_6p0 w=0.82u l=0.6u
X9272 a_13796_47170# cap_shunt_p a_14728_47108# vss nmos_6p0 w=0.82u l=0.6u
X9273 a_14580_42104# cap_shunt_n a_14372_41620# vdd pmos_6p0 w=1.2u l=0.5u
X9274 vdd a_21516_52119# a_21428_52216# vdd pmos_6p0 w=1.22u l=1u
X9275 a_18032_48676# cap_shunt_p a_16708_48738# vss nmos_6p0 w=0.82u l=0.6u
X9276 a_24452_39676# cap_shunt_p a_24660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X9277 a_2500_23996# cap_shunt_p a_2708_23650# vdd pmos_6p0 w=1.2u l=0.5u
X9278 vss tune_shunt[7] a_6740_29560# vss nmos_6p0 w=0.51u l=0.6u
X9279 vdd tune_shunt[7] a_16500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X9280 vdd a_8860_50984# a_8772_51028# vdd pmos_6p0 w=1.22u l=1u
X9281 a_24660_12674# cap_series_gyn a_26376_12612# vss nmos_6p0 w=0.82u l=0.6u
X9282 vdd a_19276_19191# a_19188_19288# vdd pmos_6p0 w=1.22u l=1u
X9283 a_28484_7124# cap_series_gyp a_28692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X9284 vss tune_shunt[7] a_6740_26424# vss nmos_6p0 w=0.51u l=0.6u
X9285 a_31416_4772# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9286 a_18404_8316# cap_series_gyp a_18612_7970# vdd pmos_6p0 w=1.2u l=0.5u
X9287 vdd tune_shunt[6] a_3620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9288 vdd a_7404_55688# a_7316_55732# vdd pmos_6p0 w=1.22u l=1u
X9289 a_10548_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9290 a_33500_42711# a_33412_42808# vss vss nmos_6p0 w=0.82u l=1u
X9291 a_24660_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9292 a_29700_17378# cap_series_gyp a_30632_17316# vss nmos_6p0 w=0.82u l=0.6u
X9293 vss tune_shunt[3] a_32612_37762# vss nmos_6p0 w=0.51u l=0.6u
X9294 a_17620_33780# cap_shunt_n a_17828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X9295 a_18760_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9296 vss tune_shunt_gy[3] a_37632_44376# vss nmos_6p0 w=0.51u l=0.6u
X9297 a_35880_25940# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9298 a_37444_44376# cap_shunt_gyp a_37632_44376# vdd pmos_6p0 w=1.215u l=0.5u
X9299 vdd tune_shunt[7] a_3620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9300 vss cap_shunt_n a_12992_45240# vss nmos_6p0 w=0.82u l=0.6u
X9301 a_14372_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9302 a_9868_53687# a_9780_53784# vss vss nmos_6p0 w=0.82u l=1u
X9303 vss tune_shunt[6] a_6740_46808# vss nmos_6p0 w=0.51u l=0.6u
X9304 a_10548_38968# cap_shunt_n a_10340_38484# vdd pmos_6p0 w=1.2u l=0.5u
X9305 a_24660_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9306 a_36300_29032# a_36212_29076# vss vss nmos_6p0 w=0.82u l=1u
X9307 vdd tune_shunt[7] a_16500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X9308 vss tune_shunt[5] a_32612_34626# vss nmos_6p0 w=0.51u l=0.6u
X9309 a_17620_30644# cap_shunt_n a_17828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X9310 a_10452_36540# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9311 a_6532_27508# cap_shunt_n a_6740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X9312 a_30924_49416# a_30836_49460# vss vss nmos_6p0 w=0.82u l=1u
X9313 vss tune_shunt_gy[2] a_37632_41240# vss nmos_6p0 w=0.51u l=0.6u
X9314 a_2588_55255# a_2500_55352# vss vss nmos_6p0 w=0.82u l=1u
X9315 vss cap_shunt_n a_15568_38968# vss nmos_6p0 w=0.82u l=0.6u
X9316 a_32632_11452# cap_series_gyp a_32444_11452# vdd pmos_6p0 w=1.2u l=0.5u
X9317 vss cap_shunt_n a_12992_42104# vss nmos_6p0 w=0.82u l=0.6u
X9318 a_23072_37700# cap_shunt_n a_21748_37762# vss nmos_6p0 w=0.82u l=0.6u
X9319 a_16476_35304# a_16388_35348# vss vss nmos_6p0 w=0.82u l=1u
X9320 a_29492_28700# cap_shunt_p a_29700_28354# vdd pmos_6p0 w=1.2u l=0.5u
X9321 a_18180_3612# cap_series_gyn a_18388_3266# vdd pmos_6p0 w=1.2u l=0.5u
X9322 a_5844_10744# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X9323 a_10548_35832# cap_shunt_n a_10340_35348# vdd pmos_6p0 w=1.2u l=0.5u
X9324 a_9876_20152# cap_shunt_p a_11592_20152# vss nmos_6p0 w=0.82u l=0.6u
X9325 a_9220_20860# cap_shunt_p a_9428_20514# vdd pmos_6p0 w=1.2u l=0.5u
X9326 a_37420_6647# a_37332_6744# vss vss nmos_6p0 w=0.82u l=1u
X9327 a_15720_11452# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9328 vdd tune_shunt[7] a_16500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X9329 vdd tune_series_gy[2] a_11572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X9330 a_28692_40536# cap_shunt_p a_28484_40052# vdd pmos_6p0 w=1.2u l=0.5u
X9331 a_10452_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9332 a_13452_3511# a_13364_3608# vss vss nmos_6p0 w=0.82u l=1u
X9333 a_9876_17016# cap_shunt_p a_9668_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9334 a_30924_46280# a_30836_46324# vss vss nmos_6p0 w=0.82u l=1u
X9335 a_15120_45540# cap_shunt_p a_13796_45602# vss nmos_6p0 w=0.82u l=0.6u
X9336 vss tune_shunt[7] a_28692_27992# vss nmos_6p0 w=0.51u l=0.6u
X9337 vdd a_27788_52552# a_27700_52596# vdd pmos_6p0 w=1.22u l=1u
X9338 a_18816_43972# cap_shunt_p a_16708_44034# vss nmos_6p0 w=0.82u l=0.6u
X9339 vdd a_36524_34871# a_36436_34968# vdd pmos_6p0 w=1.22u l=1u
X9340 a_37420_3511# a_37332_3608# vss vss nmos_6p0 w=0.82u l=1u
X9341 a_24660_23650# cap_shunt_p a_24452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X9342 a_15120_42404# cap_shunt_n a_13796_42466# vss nmos_6p0 w=0.82u l=0.6u
X9343 vdd tune_shunt[7] a_17620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9344 a_33732_34264# cap_shunt_n a_33524_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9345 vss tune_shunt[7] a_28692_24856# vss nmos_6p0 w=0.51u l=0.6u
X9346 a_18612_12674# cap_series_gyn a_18404_13020# vdd pmos_6p0 w=1.2u l=0.5u
X9347 vdd a_21516_48983# a_21428_49080# vdd pmos_6p0 w=1.22u l=1u
X9348 a_22456_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9349 vss cap_shunt_n a_35056_35832# vss nmos_6p0 w=0.82u l=0.6u
X9350 a_2140_17623# a_2052_17720# vss vss nmos_6p0 w=0.82u l=1u
X9351 a_9876_48376# cap_shunt_p a_10808_48376# vss nmos_6p0 w=0.82u l=0.6u
X9352 a_18816_40836# cap_shunt_n a_16708_40898# vss nmos_6p0 w=0.82u l=0.6u
X9353 a_7672_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9354 a_25780_32696# cap_shunt_p a_25572_32212# vdd pmos_6p0 w=1.2u l=0.5u
X9355 vss cap_series_gyp a_30800_7608# vss nmos_6p0 w=0.82u l=0.6u
X9356 vdd tune_shunt[7] a_17620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9357 a_33732_31128# cap_shunt_n a_33524_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9358 vss tune_shunt[7] a_7748_29922# vss nmos_6p0 w=0.51u l=0.6u
X9359 a_7168_10744# cap_shunt_p a_5844_10744# vss nmos_6p0 w=0.82u l=0.6u
X9360 a_5612_38007# a_5524_38104# vss vss nmos_6p0 w=0.82u l=1u
X9361 a_22456_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9362 a_13564_8215# a_13476_8312# vss vss nmos_6p0 w=0.82u l=1u
X9363 a_11648_9476# cap_shunt_p a_9540_9538# vss nmos_6p0 w=0.82u l=0.6u
X9364 a_4816_9476# cap_shunt_n a_2708_9538# vss nmos_6p0 w=0.82u l=0.6u
X9365 a_13796_42466# cap_shunt_n a_13588_42812# vdd pmos_6p0 w=1.2u l=0.5u
X9366 a_32404_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9367 a_37080_17016# cap_series_gygyn a_35880_16532# vss nmos_6p0 w=0.82u l=0.6u
X9368 vss tune_shunt[7] a_17828_37400# vss nmos_6p0 w=0.51u l=0.6u
X9369 vss tune_shunt[6] a_20740_38968# vss nmos_6p0 w=0.51u l=0.6u
X9370 a_36720_50006# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9371 a_25572_10260# cap_series_gyn a_25780_10744# vdd pmos_6p0 w=1.2u l=0.5u
X9372 a_32656_14180# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X9373 a_2500_14588# cap_shunt_n a_2708_14242# vdd pmos_6p0 w=1.2u l=0.5u
X9374 a_17620_18100# cap_shunt_p a_17828_18584# vdd pmos_6p0 w=1.2u l=0.5u
X9375 a_25572_40052# cap_shunt_n a_25780_40536# vdd pmos_6p0 w=1.2u l=0.5u
X9376 a_18032_39268# cap_shunt_n a_16708_39330# vss nmos_6p0 w=0.82u l=0.6u
X9377 a_32716_23895# a_32628_23992# vss vss nmos_6p0 w=0.82u l=1u
X9378 a_28484_40052# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9379 a_19732_10744# cap_series_gyn a_19524_10260# vdd pmos_6p0 w=1.2u l=0.5u
X9380 a_25572_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9381 a_7748_37762# cap_shunt_n a_9464_37700# vss nmos_6p0 w=0.82u l=0.6u
X9382 a_21540_44380# cap_shunt_n a_21748_44034# vdd pmos_6p0 w=1.2u l=0.5u
X9383 a_13588_20860# cap_shunt_n a_13796_20514# vdd pmos_6p0 w=1.2u l=0.5u
X9384 vdd a_35404_39575# a_35316_39672# vdd pmos_6p0 w=1.22u l=1u
X9385 a_16924_33736# a_16836_33780# vss vss nmos_6p0 w=0.82u l=1u
X9386 a_32656_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X9387 a_14372_40052# cap_shunt_n a_14580_40536# vdd pmos_6p0 w=1.2u l=0.5u
X9388 vdd a_31708_36872# a_31620_36916# vdd pmos_6p0 w=1.22u l=1u
X9389 a_27228_22327# a_27140_22424# vss vss nmos_6p0 w=0.82u l=1u
X9390 vss tune_shunt[5] a_6292_17016# vss nmos_6p0 w=0.51u l=0.6u
X9391 a_2708_45602# cap_shunt_p a_2500_45948# vdd pmos_6p0 w=1.2u l=0.5u
X9392 a_25572_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9393 vdd tune_shunt[7] a_3620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X9394 a_27104_21720# cap_shunt_p a_25780_21720# vss nmos_6p0 w=0.82u l=0.6u
X9395 vdd a_18492_54120# a_18404_54164# vdd pmos_6p0 w=1.22u l=1u
X9396 a_23464_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9397 a_2708_12674# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9398 a_21540_41244# cap_shunt_p a_21748_40898# vdd pmos_6p0 w=1.2u l=0.5u
X9399 a_24660_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9400 a_21316_3988# cap_series_gyn a_21524_4472# vdd pmos_6p0 w=1.2u l=0.5u
X9401 vss tune_shunt[7] a_32612_28354# vss nmos_6p0 w=0.51u l=0.6u
X9402 a_17620_24372# cap_shunt_n a_17828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X9403 vdd a_6060_33303# a_5972_33400# vdd pmos_6p0 w=1.22u l=1u
X9404 a_16924_30600# a_16836_30644# vss vss nmos_6p0 w=0.82u l=1u
X9405 vdd tune_series_gy[3] a_18180_3612# vdd pmos_6p0 w=1.2u l=0.5u
X9406 a_35880_16532# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9407 a_20532_14964# cap_series_gyn a_20740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X9408 a_6084_17724# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9409 a_16476_29032# a_16388_29076# vss vss nmos_6p0 w=0.82u l=1u
X9410 vdd tune_shunt[5] a_3620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X9411 a_35292_52552# a_35204_52596# vss vss nmos_6p0 w=0.82u l=1u
X9412 vdd a_18492_50984# a_18404_51028# vdd pmos_6p0 w=1.22u l=1u
X9413 a_32268_16055# a_32180_16152# vss vss nmos_6p0 w=0.82u l=1u
X9414 a_25548_54120# a_25460_54164# vss vss nmos_6p0 w=0.82u l=1u
X9415 a_10548_29560# cap_shunt_n a_10340_29076# vdd pmos_6p0 w=1.2u l=0.5u
X9416 a_24660_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9417 a_12788_20152# cap_shunt_p a_12580_19668# vdd pmos_6p0 w=1.2u l=0.5u
X9418 vdd a_15468_54120# a_15380_54164# vdd pmos_6p0 w=1.22u l=1u
X9419 a_24452_39676# cap_shunt_p a_24660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X9420 vss tune_shunt[4] a_32612_25218# vss nmos_6p0 w=0.51u l=0.6u
X9421 a_17620_21236# cap_shunt_p a_17828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X9422 a_29468_47415# a_29380_47512# vss vss nmos_6p0 w=0.82u l=1u
X9423 a_37280_44757# cap_shunt_gyp a_37280_45302# vdd pmos_6p0 w=1.215u l=0.5u
X9424 vdd tune_shunt[7] a_16500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X9425 a_4032_6040# cap_shunt_p a_1924_6040# vss nmos_6p0 w=0.82u l=0.6u
X9426 a_27104_6040# cap_series_gyp a_25780_6040# vss nmos_6p0 w=0.82u l=0.6u
X9427 a_10452_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9428 a_24660_4834# cap_series_gyp a_24452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X9429 vdd a_14908_55255# a_14820_55352# vdd pmos_6p0 w=1.22u l=1u
X9430 a_10548_34264# cap_shunt_n a_10340_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9431 vdd a_36524_28599# a_36436_28696# vdd pmos_6p0 w=1.22u l=1u
X9432 a_16476_25896# a_16388_25940# vss vss nmos_6p0 w=0.82u l=1u
X9433 a_32268_52552# a_32180_52596# vss vss nmos_6p0 w=0.82u l=1u
X9434 a_14692_7608# cap_series_gyp a_14484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X9435 a_35880_21236# cap_series_gygyp a_36688_21720# vss nmos_6p0 w=0.82u l=0.6u
X9436 vdd a_28684_47415# a_28596_47512# vdd pmos_6p0 w=1.22u l=1u
X9437 a_30640_20152# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X9438 a_15120_36132# cap_shunt_n a_13796_36194# vss nmos_6p0 w=0.82u l=0.6u
X9439 vss tune_series_gy[4] a_28692_18584# vss nmos_6p0 w=0.51u l=0.6u
X9440 vss tune_shunt[6] a_16708_45602# vss nmos_6p0 w=0.51u l=0.6u
X9441 vss cap_shunt_p a_35056_29560# vss nmos_6p0 w=0.82u l=0.6u
X9442 vdd a_14908_52119# a_14820_52216# vdd pmos_6p0 w=1.22u l=1u
X9443 a_18816_34564# cap_shunt_n a_16708_34626# vss nmos_6p0 w=0.82u l=0.6u
X9444 a_10548_31128# cap_shunt_n a_10340_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9445 vdd a_35740_3511# a_35652_3608# vdd pmos_6p0 w=1.22u l=1u
X9446 a_33544_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9447 a_24660_14242# cap_series_gyn a_24452_14588# vdd pmos_6p0 w=1.2u l=0.5u
X9448 vdd tune_shunt[7] a_17620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X9449 a_19936_12612# cap_series_gyn a_18612_12674# vss nmos_6p0 w=0.82u l=0.6u
X9450 a_23464_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X9451 vss tune_series_gy[4] a_28692_15448# vss nmos_6p0 w=0.51u l=0.6u
X9452 a_35168_44376# cap_shunt_gyn a_35188_43972# vss nmos_6p0 w=0.82u l=0.6u
X9453 vdd a_1692_54120# a_1604_54164# vdd pmos_6p0 w=1.22u l=1u
X9454 a_13796_36194# cap_shunt_n a_13588_36540# vdd pmos_6p0 w=1.2u l=0.5u
X9455 a_18816_31428# cap_shunt_n a_16708_31490# vss nmos_6p0 w=0.82u l=0.6u
X9456 a_1716_5556# cap_shunt_p a_1924_6040# vdd pmos_6p0 w=1.2u l=0.5u
X9457 a_21672_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9458 a_27452_55688# a_27364_55732# vss vss nmos_6p0 w=0.82u l=1u
X9459 a_6084_49460# cap_shunt_p a_6292_49944# vdd pmos_6p0 w=1.2u l=0.5u
X9460 a_32464_46870# cap_shunt_gyn a_32464_46325# vdd pmos_6p0 w=1.215u l=0.5u
X9461 a_33544_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9462 a_34536_9884# cap_series_gygyn a_34348_9884# vdd pmos_6p0 w=1.2u l=0.5u
X9463 a_32632_11452# cap_series_gyp a_32444_11452# vdd pmos_6p0 w=1.2u l=0.5u
X9464 a_22644_13880# cap_series_gyn a_22436_13396# vdd pmos_6p0 w=1.2u l=0.5u
X9465 a_29492_28700# cap_shunt_p a_29700_28354# vdd pmos_6p0 w=1.2u l=0.5u
X9466 vdd tune_shunt[7] a_17620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X9467 a_9220_20860# cap_shunt_p a_9428_20514# vdd pmos_6p0 w=1.2u l=0.5u
X9468 vdd a_30812_22327# a_30724_22424# vdd pmos_6p0 w=1.22u l=1u
X9469 a_18724_6040# cap_series_gyn a_18516_5556# vdd pmos_6p0 w=1.2u l=0.5u
X9470 vdd a_30812_8215# a_30724_8312# vdd pmos_6p0 w=1.22u l=1u
X9471 vdd a_1692_50984# a_1604_51028# vdd pmos_6p0 w=1.22u l=1u
X9472 vss cap_shunt_p a_15904_50244# vss nmos_6p0 w=0.82u l=0.6u
X9473 vdd a_34844_41576# a_34756_41620# vdd pmos_6p0 w=1.22u l=1u
X9474 a_13796_33058# cap_shunt_n a_13588_33404# vdd pmos_6p0 w=1.2u l=0.5u
X9475 a_10660_23650# cap_shunt_n a_10452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X9476 a_9876_17016# cap_shunt_p a_9668_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9477 a_4828_52552# a_4740_52596# vss vss nmos_6p0 w=0.82u l=1u
X9478 vss tune_series_gy[4] a_25780_20152# vss nmos_6p0 w=0.51u l=0.6u
X9479 a_4032_43972# cap_shunt_p a_2708_44034# vss nmos_6p0 w=0.82u l=0.6u
X9480 a_16500_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9481 a_34536_6748# cap_series_gygyp a_34348_6748# vdd pmos_6p0 w=1.2u l=0.5u
X9482 a_2708_15810# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9483 a_24428_55688# a_24340_55732# vss vss nmos_6p0 w=0.82u l=1u
X9484 vss cap_series_gyp a_17024_6340# vss nmos_6p0 w=0.82u l=0.6u
X9485 vdd a_19724_17623# a_19636_17720# vdd pmos_6p0 w=1.22u l=1u
X9486 a_7540_23996# cap_shunt_p a_7748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X9487 vss cap_shunt_n a_12768_39268# vss nmos_6p0 w=0.82u l=0.6u
X9488 a_2708_39330# cap_shunt_n a_2500_39676# vdd pmos_6p0 w=1.2u l=0.5u
X9489 vss cap_shunt_n a_30800_38968# vss nmos_6p0 w=0.82u l=0.6u
X9490 a_2724_10260# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9491 a_17828_42104# cap_shunt_n a_17620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X9492 a_25572_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9493 a_24660_23650# cap_shunt_p a_24452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X9494 a_6060_6647# a_5972_6744# vss vss nmos_6p0 w=0.82u l=1u
X9495 vdd a_31260_42711# a_31172_42808# vdd pmos_6p0 w=1.22u l=1u
X9496 a_16500_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9497 a_28692_26424# cap_shunt_p a_28484_25940# vdd pmos_6p0 w=1.2u l=0.5u
X9498 a_23308_19624# a_23220_19668# vss vss nmos_6p0 w=0.82u l=1u
X9499 a_8512_47108# cap_shunt_p a_6404_47170# vss nmos_6p0 w=0.82u l=0.6u
X9500 a_4032_40836# cap_shunt_p a_2708_40898# vss nmos_6p0 w=0.82u l=0.6u
X9501 a_8848_53080# cap_shunt_n a_6740_53080# vss nmos_6p0 w=0.82u l=0.6u
X9502 a_8680_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9503 vdd a_31708_27464# a_31620_27508# vdd pmos_6p0 w=1.22u l=1u
X9504 a_27104_12312# cap_series_gyp a_25780_12312# vss nmos_6p0 w=0.82u l=0.6u
X9505 a_13588_49084# cap_shunt_n a_13796_48738# vdd pmos_6p0 w=1.2u l=0.5u
X9506 a_6740_48376# cap_shunt_p a_6532_47892# vdd pmos_6p0 w=1.2u l=0.5u
X9507 a_13776_43672# cap_shunt_n a_11668_43672# vss nmos_6p0 w=0.82u l=0.6u
X9508 a_23464_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9509 a_25548_47848# a_25460_47892# vss vss nmos_6p0 w=0.82u l=1u
X9510 a_28692_23288# cap_shunt_p a_28484_22804# vdd pmos_6p0 w=1.2u l=0.5u
X9511 a_35692_13396# cap_series_gygyn a_35880_13396# vdd pmos_6p0 w=1.2u l=0.5u
X9512 vdd a_28236_49416# a_28148_49460# vdd pmos_6p0 w=1.22u l=1u
X9513 a_13796_42466# cap_shunt_n a_13588_42812# vdd pmos_6p0 w=1.2u l=0.5u
X9514 vdd a_31260_8648# a_31172_8692# vdd pmos_6p0 w=1.22u l=1u
X9515 vss cap_series_gygyn a_32824_18884# vss nmos_6p0 w=0.82u l=0.6u
X9516 a_25444_3266# cap_shunt_p a_25236_3612# vdd pmos_6p0 w=1.2u l=0.5u
X9517 a_19152_20152# cap_shunt_p a_17828_20152# vss nmos_6p0 w=0.82u l=0.6u
X9518 vss cap_shunt_p a_26768_43972# vss nmos_6p0 w=0.82u l=0.6u
X9519 a_8680_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9520 a_36636_55255# a_36548_55352# vss vss nmos_6p0 w=0.82u l=1u
X9521 vss tune_series_gygy[5] a_35880_22804# vss nmos_6p0 w=0.51u l=0.6u
X9522 a_28692_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9523 a_6740_45240# cap_shunt_p a_6532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X9524 a_13776_40536# cap_shunt_n a_11668_40536# vss nmos_6p0 w=0.82u l=0.6u
X9525 a_31024_14180# cap_series_gyp a_29700_14242# vss nmos_6p0 w=0.82u l=0.6u
X9526 a_10808_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9527 vdd a_24652_19624# a_24564_19668# vdd pmos_6p0 w=1.22u l=1u
X9528 vss cap_shunt_p a_8064_46808# vss nmos_6p0 w=0.82u l=0.6u
X9529 vdd tune_shunt[6] a_7540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X9530 a_25572_40052# cap_shunt_n a_25780_40536# vdd pmos_6p0 w=1.2u l=0.5u
X9531 a_10548_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9532 vdd a_28236_46280# a_28148_46324# vdd pmos_6p0 w=1.22u l=1u
X9533 vdd a_31260_5512# a_31172_5556# vdd pmos_6p0 w=1.22u l=1u
X9534 a_6644_53788# cap_shunt_n a_6852_53442# vdd pmos_6p0 w=1.2u l=0.5u
X9535 a_14260_3612# cap_series_gyn a_14468_3266# vdd pmos_6p0 w=1.2u l=0.5u
X9536 a_6532_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9537 a_34516_17378# cap_series_gygyn a_34308_17724# vdd pmos_6p0 w=1.2u l=0.5u
X9538 vss cap_shunt_n a_26768_40836# vss nmos_6p0 w=0.82u l=0.6u
X9539 vss tune_shunt[6] a_16708_39330# vss nmos_6p0 w=0.51u l=0.6u
X9540 a_28692_10744# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9541 a_20740_37400# cap_shunt_n a_20532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X9542 a_18816_28292# cap_shunt_n a_16708_28354# vss nmos_6p0 w=0.82u l=0.6u
X9543 a_25984_6340# cap_series_gyn a_24660_6402# vss nmos_6p0 w=0.82u l=0.6u
X9544 a_31024_11044# cap_series_gyp a_29700_11106# vss nmos_6p0 w=0.82u l=0.6u
X9545 a_10548_24856# cap_shunt_n a_10340_24372# vdd pmos_6p0 w=1.2u l=0.5u
X9546 vdd tune_shunt[6] a_7540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X9547 a_14372_40052# cap_shunt_n a_14580_40536# vdd pmos_6p0 w=1.2u l=0.5u
X9548 a_35880_11828# cap_series_gygyp a_36688_12312# vss nmos_6p0 w=0.82u l=0.6u
X9549 a_33544_28292# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9550 a_32156_53687# a_32068_53784# vss vss nmos_6p0 w=0.82u l=1u
X9551 a_7580_6748# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9552 a_35904_13880# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X9553 vdd tune_shunt[7] a_6532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X9554 a_13588_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9555 a_32732_45240# cap_shunt_gyp a_32464_45302# vss nmos_6p0 w=0.82u l=0.6u
X9556 a_18816_25156# cap_shunt_n a_16708_25218# vss nmos_6p0 w=0.82u l=0.6u
X9557 a_35880_18100# cap_series_gygyn a_35692_18100# vdd pmos_6p0 w=1.2u l=0.5u
X9558 a_14580_45240# cap_shunt_p a_15512_45240# vss nmos_6p0 w=0.82u l=0.6u
X9559 a_25780_42104# cap_shunt_n a_26712_42104# vss nmos_6p0 w=0.82u l=0.6u
X9560 a_6760_5556# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X9561 a_20532_14964# cap_series_gyn a_20740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X9562 a_6084_17724# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9563 vdd a_11884_50551# a_11796_50648# vdd pmos_6p0 w=1.22u l=1u
X9564 a_33544_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9565 vdd tune_shunt[7] a_29492_30268# vdd pmos_6p0 w=1.2u l=0.5u
X9566 vss cap_shunt_p a_4032_22020# vss nmos_6p0 w=0.82u l=0.6u
X9567 a_32156_50551# a_32068_50648# vss vss nmos_6p0 w=0.82u l=1u
X9568 a_31624_8316# cap_series_gygyn a_31436_8316# vdd pmos_6p0 w=1.2u l=0.5u
X9569 a_35904_10744# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X9570 vdd tune_shunt[7] a_6532_11828# vdd pmos_6p0 w=1.2u l=0.5u
X9571 vdd tune_shunt[5] a_3172_49460# vdd pmos_6p0 w=1.2u l=0.5u
X9572 a_24452_39676# cap_shunt_p a_24660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X9573 vdd a_16924_36872# a_16836_36916# vdd pmos_6p0 w=1.22u l=1u
X9574 a_13796_26786# cap_shunt_n a_13588_27132# vdd pmos_6p0 w=1.2u l=0.5u
X9575 vss cap_series_gyp a_23968_7608# vss nmos_6p0 w=0.82u l=0.6u
X9576 a_18612_6402# cap_series_gyn a_19544_6340# vss nmos_6p0 w=0.82u l=0.6u
X9577 vdd tune_series_gy[5] a_25572_13396# vdd pmos_6p0 w=1.2u l=0.5u
X9578 a_14580_42104# cap_shunt_n a_15512_42104# vss nmos_6p0 w=0.82u l=0.6u
X9579 a_6740_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9580 vdd tune_shunt[7] a_13588_23996# vdd pmos_6p0 w=1.2u l=0.5u
X9581 a_7768_6748# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X9582 a_2140_49416# a_2052_49460# vss vss nmos_6p0 w=0.82u l=1u
X9583 a_10548_34264# cap_shunt_n a_10340_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9584 a_21540_17724# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9585 a_17640_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9586 a_19712_3204# cap_series_gyn a_18388_3266# vss nmos_6p0 w=0.82u l=0.6u
X9587 a_37420_20759# a_37332_20856# vss vss nmos_6p0 w=0.82u l=1u
X9588 a_21636_6040# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9589 a_21316_3988# cap_series_gyn a_21524_4472# vdd pmos_6p0 w=1.2u l=0.5u
X9590 vdd a_35292_55688# a_35204_55732# vdd pmos_6p0 w=1.22u l=1u
X9591 a_28684_52552# a_28596_52596# vss vss nmos_6p0 w=0.82u l=1u
X9592 vss cap_shunt_n a_19152_37400# vss nmos_6p0 w=0.82u l=0.6u
X9593 a_1924_7970# cap_shunt_n a_2856_7908# vss nmos_6p0 w=0.82u l=0.6u
X9594 a_4032_34564# cap_shunt_n a_2708_34626# vss nmos_6p0 w=0.82u l=0.6u
X9595 vdd tune_shunt[4] a_2500_13020# vdd pmos_6p0 w=1.2u l=0.5u
X9596 a_2140_46280# a_2052_46324# vss vss nmos_6p0 w=0.82u l=1u
X9597 a_10548_31128# cap_shunt_n a_10340_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9598 vss tune_series_gygy[4] a_34516_15810# vss nmos_6p0 w=0.51u l=0.6u
X9599 a_17640_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9600 vss cap_series_gyn a_30016_9176# vss nmos_6p0 w=0.82u l=0.6u
X9601 vdd a_2140_10216# a_2052_10260# vdd pmos_6p0 w=1.22u l=1u
X9602 vdd a_21964_55255# a_21876_55352# vdd pmos_6p0 w=1.22u l=1u
X9603 a_11460_44756# cap_shunt_n a_11668_45240# vdd pmos_6p0 w=1.2u l=0.5u
X9604 a_3828_40536# cap_shunt_n a_3620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X9605 vdd a_28124_23895# a_28036_23992# vdd pmos_6p0 w=1.22u l=1u
X9606 a_17828_32696# cap_shunt_n a_17620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X9607 a_21428_5556# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9608 vdd a_8412_8648# a_8324_8692# vdd pmos_6p0 w=1.22u l=1u
X9609 a_24660_14242# cap_series_gyn a_24452_14588# vdd pmos_6p0 w=1.2u l=0.5u
X9610 a_36232_18884# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X9611 a_36384_50648# cap_shunt_gyp a_36384_50244# vdd pmos_6p0 w=1.215u l=0.5u
X9612 a_10452_45948# cap_shunt_n a_10660_45602# vdd pmos_6p0 w=1.2u l=0.5u
X9613 vdd a_10540_8648# a_10452_8692# vdd pmos_6p0 w=1.22u l=1u
X9614 vdd a_32268_55688# a_32180_55732# vdd pmos_6p0 w=1.22u l=1u
X9615 a_4032_31428# cap_shunt_p a_2708_31490# vss nmos_6p0 w=0.82u l=0.6u
X9616 a_4760_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9617 a_21748_6402# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9618 a_28692_17016# cap_series_gyn a_28484_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9619 a_13796_36194# cap_shunt_n a_13588_36540# vdd pmos_6p0 w=1.2u l=0.5u
X9620 a_19732_9176# cap_series_gyp a_19524_8692# vdd pmos_6p0 w=1.2u l=0.5u
X9621 a_37444_41621# cap_shunt_gyp a_37632_41621# vdd pmos_6p0 w=1.215u l=0.5u
X9622 vss cap_shunt_p a_10864_15748# vss nmos_6p0 w=0.82u l=0.6u
X9623 vdd a_21964_52119# a_21876_52216# vdd pmos_6p0 w=1.22u l=1u
X9624 a_7748_45602# cap_shunt_p a_7540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X9625 vdd a_28124_20759# a_28036_20856# vdd pmos_6p0 w=1.22u l=1u
X9626 a_6084_49460# cap_shunt_p a_6292_49944# vdd pmos_6p0 w=1.2u l=0.5u
X9627 a_6740_38968# cap_shunt_n a_6532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X9628 a_29492_28700# cap_shunt_p a_29700_28354# vdd pmos_6p0 w=1.2u l=0.5u
X9629 vss tune_series_gy[3] a_14692_6040# vss nmos_6p0 w=0.51u l=0.6u
X9630 vss cap_series_gyn a_21840_12312# vss nmos_6p0 w=0.82u l=0.6u
X9631 a_36232_15748# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X9632 a_6852_53442# cap_shunt_n a_8568_53380# vss nmos_6p0 w=0.82u l=0.6u
X9633 vdd a_10540_5512# a_10452_5556# vdd pmos_6p0 w=1.22u l=1u
X9634 vss cap_shunt_n a_14896_49944# vss nmos_6p0 w=0.82u l=0.6u
X9635 a_4760_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9636 a_34844_24328# a_34756_24372# vss vss nmos_6p0 w=0.82u l=1u
X9637 a_13796_33058# cap_shunt_n a_13588_33404# vdd pmos_6p0 w=1.2u l=0.5u
X9638 a_10660_23650# cap_shunt_n a_10452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X9639 a_6776_9476# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9640 vss cap_shunt_p a_26768_34564# vss nmos_6p0 w=0.82u l=0.6u
X9641 a_13460_35832# cap_shunt_n a_15176_35832# vss nmos_6p0 w=0.82u l=0.6u
X9642 a_6740_35832# cap_shunt_n a_6532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X9643 a_2856_7608# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9644 vdd tune_series_gy[4] a_25572_8692# vdd pmos_6p0 w=1.2u l=0.5u
X9645 a_10808_12312# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9646 a_7540_23996# cap_shunt_p a_7748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X9647 a_10548_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9648 a_2724_8692# cap_shunt_n a_2932_9176# vdd pmos_6p0 w=1.2u l=0.5u
X9649 vdd a_7852_55688# a_7764_55732# vdd pmos_6p0 w=1.22u l=1u
X9650 vdd a_27228_8215# a_27140_8312# vdd pmos_6p0 w=1.22u l=1u
X9651 a_34348_9884# cap_series_gygyn a_34536_9884# vdd pmos_6p0 w=1.2u l=0.5u
X9652 a_2724_10260# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9653 a_6532_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9654 vss cap_shunt_p a_26768_31428# vss nmos_6p0 w=0.82u l=0.6u
X9655 a_25780_27992# cap_shunt_p a_27496_27992# vss nmos_6p0 w=0.82u l=0.6u
X9656 a_28692_26424# cap_shunt_p a_28484_25940# vdd pmos_6p0 w=1.2u l=0.5u
X9657 vdd a_22188_47848# a_22100_47892# vdd pmos_6p0 w=1.22u l=1u
X9658 a_21748_44034# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9659 a_32604_36872# a_32516_36916# vss vss nmos_6p0 w=0.82u l=1u
X9660 a_20740_27992# cap_shunt_n a_20532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X9661 vdd tune_series_gy[3] a_25572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X9662 a_13588_39676# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9663 a_36624_4772# cap_series_gygyp a_34516_4834# vss nmos_6p0 w=0.82u l=0.6u
X9664 a_25984_32996# cap_shunt_p a_24660_33058# vss nmos_6p0 w=0.82u l=0.6u
X9665 a_34348_6748# cap_series_gygyp a_34536_6748# vdd pmos_6p0 w=1.2u l=0.5u
X9666 a_9540_15810# cap_shunt_p a_9332_16156# vdd pmos_6p0 w=1.2u l=0.5u
X9667 vdd a_4828_55688# a_4740_55732# vdd pmos_6p0 w=1.22u l=1u
X9668 a_16028_50984# a_15940_51028# vss vss nmos_6p0 w=0.82u l=1u
X9669 a_34144_47108# cap_shunt_gyp a_34144_47512# vdd pmos_6p0 w=1.215u l=0.5u
X9670 vdd a_23308_25896# a_23220_25940# vdd pmos_6p0 w=1.22u l=1u
X9671 a_25780_24856# cap_shunt_p a_27496_24856# vss nmos_6p0 w=0.82u l=0.6u
X9672 vdd a_35740_54120# a_35652_54164# vdd pmos_6p0 w=1.22u l=1u
X9673 a_32928_45944# cap_shunt_gyn a_32740_45944# vdd pmos_6p0 w=1.215u l=0.5u
X9674 a_28692_23288# cap_shunt_p a_28484_22804# vdd pmos_6p0 w=1.2u l=0.5u
X9675 a_29492_30268# cap_shunt_p a_29700_29922# vdd pmos_6p0 w=1.2u l=0.5u
X9676 a_11780_4472# cap_series_gyp a_11572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X9677 a_9668_21236# cap_shunt_p a_9876_21720# vdd pmos_6p0 w=1.2u l=0.5u
X9678 a_28348_43144# a_28260_43188# vss vss nmos_6p0 w=0.82u l=1u
X9679 vss cap_shunt_n a_15120_29860# vss nmos_6p0 w=0.82u l=0.6u
X9680 a_6292_51512# cap_shunt_p a_6084_51028# vdd pmos_6p0 w=1.2u l=0.5u
X9681 vss tune_shunt[4] a_24660_42466# vss nmos_6p0 w=0.51u l=0.6u
X9682 a_6740_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9683 a_7568_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X9684 a_15720_11452# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9685 vss tune_shunt[6] a_10660_37762# vss nmos_6p0 w=0.51u l=0.6u
X9686 a_24452_13020# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9687 vdd tune_shunt[4] a_33524_33780# vdd pmos_6p0 w=1.2u l=0.5u
X9688 vdd a_23308_22760# a_23220_22804# vdd pmos_6p0 w=1.22u l=1u
X9689 vdd a_35740_50984# a_35652_51028# vdd pmos_6p0 w=1.22u l=1u
X9690 a_13252_36916# cap_shunt_n a_13460_37400# vdd pmos_6p0 w=1.2u l=0.5u
X9691 vdd a_16924_27464# a_16836_27508# vdd pmos_6p0 w=1.22u l=1u
X9692 a_37420_14487# a_37332_14584# vss vss nmos_6p0 w=0.82u l=1u
X9693 a_25572_40052# cap_shunt_n a_25780_40536# vdd pmos_6p0 w=1.2u l=0.5u
X9694 vdd a_32716_54120# a_32628_54164# vdd pmos_6p0 w=1.22u l=1u
X9695 a_3620_36916# cap_shunt_n a_3828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X9696 vss cap_shunt_n a_15120_26724# vss nmos_6p0 w=0.82u l=0.6u
X9697 a_6740_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9698 a_34516_17378# cap_series_gygyn a_34308_17724# vdd pmos_6p0 w=1.2u l=0.5u
X9699 a_13588_50652# cap_shunt_p a_13796_50306# vdd pmos_6p0 w=1.2u l=0.5u
X9700 a_4032_28292# cap_shunt_n a_2708_28354# vss nmos_6p0 w=0.82u l=0.6u
X9701 vdd tune_shunt[7] a_13588_14588# vdd pmos_6p0 w=1.2u l=0.5u
X9702 vss tune_shunt[7] a_10660_34626# vss nmos_6p0 w=0.51u l=0.6u
X9703 vss tune_series_gy[4] a_29720_13020# vss nmos_6p0 w=0.51u l=0.6u
X9704 a_23420_54120# a_23332_54164# vss vss nmos_6p0 w=0.82u l=1u
X9705 vdd tune_shunt[4] a_33524_30644# vdd pmos_6p0 w=1.2u l=0.5u
X9706 a_10548_24856# cap_shunt_n a_10340_24372# vdd pmos_6p0 w=1.2u l=0.5u
X9707 vss cap_shunt_p a_7168_9176# vss nmos_6p0 w=0.82u l=0.6u
X9708 vdd a_36972_3511# a_36884_3608# vdd pmos_6p0 w=1.22u l=1u
X9709 a_37420_11351# a_37332_11448# vss vss nmos_6p0 w=0.82u l=1u
X9710 vdd a_21964_48983# a_21876_49080# vdd pmos_6p0 w=1.22u l=1u
X9711 a_27340_47415# a_27252_47512# vss vss nmos_6p0 w=0.82u l=1u
X9712 a_17640_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9713 vdd a_32716_50984# a_32628_51028# vdd pmos_6p0 w=1.22u l=1u
X9714 a_10660_45602# cap_shunt_n a_12376_45540# vss nmos_6p0 w=0.82u l=0.6u
X9715 a_25780_9176# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9716 vdd a_16252_14920# a_16164_14964# vdd pmos_6p0 w=1.22u l=1u
X9717 a_36384_44376# cap_shunt_gyp a_36384_43972# vdd pmos_6p0 w=1.215u l=0.5u
X9718 a_10452_39676# cap_shunt_n a_10660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X9719 a_4032_25156# cap_shunt_p a_2708_25218# vss nmos_6p0 w=0.82u l=0.6u
X9720 a_25444_3266# cap_shunt_p a_25236_3612# vdd pmos_6p0 w=1.2u l=0.5u
X9721 a_14692_9176# cap_series_gyn a_14484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X9722 vdd a_32268_49416# a_32180_49460# vdd pmos_6p0 w=1.22u l=1u
X9723 vdd a_20172_41143# a_20084_41240# vdd pmos_6p0 w=1.22u l=1u
X9724 a_32612_37762# cap_shunt_p a_34328_37700# vss nmos_6p0 w=0.82u l=0.6u
X9725 vdd tune_series_gy[4] a_32444_14588# vdd pmos_6p0 w=1.2u l=0.5u
X9726 a_17620_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9727 vdd a_13340_50984# a_13252_51028# vdd pmos_6p0 w=1.22u l=1u
X9728 a_7748_39330# cap_shunt_n a_7540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X9729 a_21316_3612# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9730 vdd a_28124_14487# a_28036_14584# vdd pmos_6p0 w=1.22u l=1u
X9731 a_20532_14964# cap_series_gyn a_20740_15448# vdd pmos_6p0 w=1.2u l=0.5u
X9732 a_10660_42466# cap_shunt_n a_12376_42404# vss nmos_6p0 w=0.82u l=0.6u
X9733 vdd a_16252_11784# a_16164_11828# vdd pmos_6p0 w=1.22u l=1u
X9734 a_14692_6040# cap_series_gyn a_14484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X9735 vdd a_34396_18056# a_34308_18100# vdd pmos_6p0 w=1.22u l=1u
X9736 a_34844_18056# a_34756_18100# vss vss nmos_6p0 w=0.82u l=1u
X9737 vdd a_29916_19191# a_29828_19288# vdd pmos_6p0 w=1.22u l=1u
X9738 vdd tune_shunt[3] a_25572_43188# vdd pmos_6p0 w=1.2u l=0.5u
X9739 a_13796_26786# cap_shunt_n a_13588_27132# vdd pmos_6p0 w=1.2u l=0.5u
X9740 vdd tune_shunt[3] a_2500_9884# vdd pmos_6p0 w=1.2u l=0.5u
X9741 a_11592_43972# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9742 vss tune_series_gy[4] a_15700_7970# vss nmos_6p0 w=0.51u l=0.6u
X9743 vss cap_shunt_n a_26768_28292# vss nmos_6p0 w=0.82u l=0.6u
X9744 vdd a_28124_11351# a_28036_11448# vdd pmos_6p0 w=1.22u l=1u
X9745 a_16708_17378# cap_shunt_p a_16500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X9746 a_6740_29560# cap_shunt_n a_6532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X9747 a_25548_53687# a_25460_53784# vss vss nmos_6p0 w=0.82u l=1u
X9748 vdd a_31708_47415# a_31620_47512# vdd pmos_6p0 w=1.22u l=1u
X9749 a_13460_29560# cap_shunt_n a_15176_29560# vss nmos_6p0 w=0.82u l=0.6u
X9750 a_9108_50652# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9751 a_12992_46808# cap_shunt_n a_11668_46808# vss nmos_6p0 w=0.82u l=0.6u
X9752 a_34844_14920# a_34756_14964# vss vss nmos_6p0 w=0.82u l=1u
X9753 vdd tune_shunt[6] a_14372_43188# vdd pmos_6p0 w=1.2u l=0.5u
X9754 a_4760_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9755 a_10092_55255# a_10004_55352# vss vss nmos_6p0 w=0.82u l=1u
X9756 a_11592_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9757 vss tune_series_gy[3] a_15700_4834# vss nmos_6p0 w=0.51u l=0.6u
X9758 a_35292_38440# a_35204_38484# vss vss nmos_6p0 w=0.82u l=1u
X9759 vss cap_shunt_p a_26768_25156# vss nmos_6p0 w=0.82u l=0.6u
X9760 vdd a_12332_47415# a_12244_47512# vdd pmos_6p0 w=1.22u l=1u
X9761 vdd a_33164_9783# a_33076_9880# vdd pmos_6p0 w=1.22u l=1u
X9762 a_33500_55688# a_33412_55732# vss vss nmos_6p0 w=0.82u l=1u
X9763 a_27676_22327# a_27588_22424# vss vss nmos_6p0 w=0.82u l=1u
X9764 a_25548_50551# a_25460_50648# vss vss nmos_6p0 w=0.82u l=1u
X9765 a_13460_26424# cap_shunt_n a_15176_26424# vss nmos_6p0 w=0.82u l=0.6u
X9766 a_18388_3266# cap_series_gyn a_18180_3612# vdd pmos_6p0 w=1.2u l=0.5u
X9767 vdd tune_shunt[4] a_2500_13020# vdd pmos_6p0 w=1.2u l=0.5u
X9768 a_35264_49080# cap_shunt_gyn a_35264_48676# vdd pmos_6p0 w=1.215u l=0.5u
X9769 vdd a_24204_44712# a_24116_44756# vdd pmos_6p0 w=1.22u l=1u
X9770 vdd tune_shunt_gy[1] a_36100_39672# vdd pmos_6p0 w=1.215u l=0.5u
X9771 a_14392_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9772 a_25780_18584# cap_series_gyn a_27496_18584# vss nmos_6p0 w=0.82u l=0.6u
X9773 a_16708_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9774 a_28692_17016# cap_series_gyn a_28484_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9775 vdd tune_shunt[6] a_14372_46324# vdd pmos_6p0 w=1.2u l=0.5u
X9776 vdd a_3036_41576# a_2948_41620# vdd pmos_6p0 w=1.22u l=1u
X9777 a_17828_15448# cap_shunt_p a_17620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X9778 a_7748_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9779 a_34308_23996# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9780 a_25996_54120# a_25908_54164# vss vss nmos_6p0 w=0.82u l=1u
X9781 a_3380_49944# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X9782 vss tune_shunt[6] a_24660_36194# vss nmos_6p0 w=0.51u l=0.6u
X9783 a_25984_23588# cap_shunt_p a_24660_23650# vss nmos_6p0 w=0.82u l=0.6u
X9784 vdd tune_shunt[3] a_5636_11452# vdd pmos_6p0 w=1.2u l=0.5u
X9785 a_33948_3944# a_33860_3988# vss vss nmos_6p0 w=0.82u l=1u
X9786 a_14392_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9787 vdd a_16700_13352# a_16612_13396# vdd pmos_6p0 w=1.22u l=1u
X9788 vdd a_23308_16488# a_23220_16532# vdd pmos_6p0 w=1.22u l=1u
X9789 a_25780_15448# cap_series_gyp a_27496_15448# vss nmos_6p0 w=0.82u l=0.6u
X9790 a_4816_20452# cap_shunt_p a_2708_20514# vss nmos_6p0 w=0.82u l=0.6u
X9791 a_20740_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9792 vss tune_series_gy[4] a_11800_8692# vss nmos_6p0 w=0.51u l=0.6u
X9793 a_3828_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9794 vss tune_shunt[6] a_24660_33058# vss nmos_6p0 w=0.51u l=0.6u
X9795 a_13588_44380# cap_shunt_n a_13796_44034# vdd pmos_6p0 w=1.2u l=0.5u
X9796 vss tune_shunt[7] a_10660_28354# vss nmos_6p0 w=0.51u l=0.6u
X9797 a_21524_3266# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X9798 a_13252_27508# cap_shunt_n a_13460_27992# vdd pmos_6p0 w=1.2u l=0.5u
X9799 a_9668_18100# cap_shunt_p a_9876_18584# vdd pmos_6p0 w=1.2u l=0.5u
X9800 a_20532_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9801 a_9332_11452# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9802 a_3620_27508# cap_shunt_n a_3828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X9803 a_9668_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9804 vss cap_shunt_p a_15120_17316# vss nmos_6p0 w=0.82u l=0.6u
X9805 a_18424_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9806 a_13588_41244# cap_shunt_n a_13796_40898# vdd pmos_6p0 w=1.2u l=0.5u
X9807 a_19936_35832# cap_shunt_n a_17828_35832# vss nmos_6p0 w=0.82u l=0.6u
X9808 vss tune_shunt[7] a_10660_25218# vss nmos_6p0 w=0.51u l=0.6u
X9809 a_6628_14242# cap_shunt_p a_6420_14588# vdd pmos_6p0 w=1.2u l=0.5u
X9810 a_25572_19668# cap_series_gyp a_25780_20152# vdd pmos_6p0 w=1.2u l=0.5u
X9811 vss tune_shunt[7] a_13796_26786# vss nmos_6p0 w=0.51u l=0.6u
X9812 a_9540_15810# cap_shunt_p a_9332_16156# vdd pmos_6p0 w=1.2u l=0.5u
X9813 a_10660_36194# cap_shunt_n a_12376_36132# vss nmos_6p0 w=0.82u l=0.6u
X9814 a_28692_35832# cap_shunt_p a_30408_35832# vss nmos_6p0 w=0.82u l=0.6u
X9815 a_18612_4834# cap_series_gyp a_18404_5180# vdd pmos_6p0 w=1.2u l=0.5u
X9816 a_9668_11828# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9817 a_18424_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9818 a_2140_52119# a_2052_52216# vss vss nmos_6p0 w=0.82u l=1u
X9819 a_2708_17378# cap_shunt_p a_2500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X9820 a_33524_32212# cap_shunt_n a_33732_32696# vdd pmos_6p0 w=1.2u l=0.5u
X9821 vss tune_shunt[7] a_9540_12674# vss nmos_6p0 w=0.51u l=0.6u
X9822 a_6292_51512# cap_shunt_p a_6084_51028# vdd pmos_6p0 w=1.2u l=0.5u
X9823 a_2708_50306# cap_shunt_n a_4424_50244# vss nmos_6p0 w=0.82u l=0.6u
X9824 a_35880_8692# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X9825 a_21540_13020# cap_series_gyn a_21748_12674# vdd pmos_6p0 w=1.2u l=0.5u
X9826 vdd tune_shunt[5] a_6084_19292# vdd pmos_6p0 w=1.2u l=0.5u
X9827 a_8848_38968# cap_shunt_n a_6740_38968# vss nmos_6p0 w=0.82u l=0.6u
X9828 a_13252_36916# cap_shunt_n a_13460_37400# vdd pmos_6p0 w=1.2u l=0.5u
X9829 a_11592_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9830 a_9204_51874# cap_shunt_n a_8996_52220# vdd pmos_6p0 w=1.2u l=0.5u
X9831 a_7748_34626# cap_shunt_n a_7540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X9832 vdd tune_shunt[5] a_6084_16156# vdd pmos_6p0 w=1.2u l=0.5u
X9833 a_16708_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9834 a_24452_34972# cap_shunt_p a_24660_34626# vdd pmos_6p0 w=1.2u l=0.5u
X9835 a_21748_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9836 vss cap_shunt_n a_4816_37700# vss nmos_6p0 w=0.82u l=0.6u
X9837 a_29384_3612# tune_series_gy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X9838 vdd a_24204_38440# a_24116_38484# vdd pmos_6p0 w=1.22u l=1u
X9839 a_11592_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9840 a_23756_19624# a_23668_19668# vss vss nmos_6p0 w=0.82u l=1u
X9841 a_7748_31490# cap_shunt_n a_7540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X9842 vdd a_9644_8648# a_9556_8692# vdd pmos_6p0 w=1.22u l=1u
X9843 a_28484_36916# cap_shunt_p a_28692_37400# vdd pmos_6p0 w=1.2u l=0.5u
X9844 a_31624_6748# cap_series_gygyn a_31436_6748# vdd pmos_6p0 w=1.2u l=0.5u
X9845 vdd a_4380_55255# a_4292_55352# vdd pmos_6p0 w=1.22u l=1u
X9846 vdd a_19276_44279# a_19188_44376# vdd pmos_6p0 w=1.22u l=1u
X9847 a_16708_36194# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9848 a_10092_7080# a_10004_7124# vss vss nmos_6p0 w=0.82u l=1u
X9849 a_34516_17378# cap_series_gygyn a_35448_17316# vss nmos_6p0 w=0.82u l=0.6u
X9850 a_24452_31836# cap_shunt_p a_24660_31490# vdd pmos_6p0 w=1.2u l=0.5u
X9851 vss tune_shunt[5] a_6292_51512# vss nmos_6p0 w=0.51u l=0.6u
X9852 a_25996_47848# a_25908_47892# vss vss nmos_6p0 w=0.82u l=1u
X9853 a_35880_24372# cap_series_gygyp a_35692_24372# vdd pmos_6p0 w=1.2u l=0.5u
X9854 vdd a_28684_49416# a_28596_49460# vdd pmos_6p0 w=1.22u l=1u
X9855 vdd a_24204_35304# a_24116_35348# vdd pmos_6p0 w=1.22u l=1u
X9856 vdd a_9644_5512# a_9556_5556# vdd pmos_6p0 w=1.22u l=1u
X9857 a_4816_14180# cap_shunt_n a_2708_14242# vss nmos_6p0 w=0.82u l=0.6u
X9858 a_16812_54120# a_16724_54164# vss vss nmos_6p0 w=0.82u l=1u
X9859 vdd a_4380_52119# a_4292_52216# vdd pmos_6p0 w=1.22u l=1u
X9860 a_16708_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X9861 vdd a_3036_32168# a_2948_32212# vdd pmos_6p0 w=1.22u l=1u
X9862 a_8968_4772# cap_series_gyn a_7768_5180# vss nmos_6p0 w=0.82u l=0.6u
X9863 a_35880_21236# cap_series_gygyp a_35692_21236# vdd pmos_6p0 w=1.2u l=0.5u
X9864 vdd a_28684_46280# a_28596_46324# vdd pmos_6p0 w=1.22u l=1u
X9865 a_21524_3266# cap_series_gyp a_23240_3204# vss nmos_6p0 w=0.82u l=0.6u
X9866 vdd tune_series_gy[4] a_29492_11452# vdd pmos_6p0 w=1.2u l=0.5u
X9867 a_16708_17378# cap_shunt_p a_16500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X9868 vss cap_shunt_p a_5488_49944# vss nmos_6p0 w=0.82u l=0.6u
X9869 a_4816_11044# cap_shunt_n a_2708_11106# vss nmos_6p0 w=0.82u l=0.6u
X9870 vdd a_35180_14487# a_35092_14584# vdd pmos_6p0 w=1.22u l=1u
X9871 vss cap_shunt_p a_11200_18584# vss nmos_6p0 w=0.82u l=0.6u
X9872 vss tune_shunt[6] a_2708_45602# vss nmos_6p0 w=0.51u l=0.6u
X9873 a_7580_6748# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9874 a_19936_29560# cap_shunt_n a_17828_29560# vss nmos_6p0 w=0.82u l=0.6u
X9875 a_7560_10744# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9876 a_24660_37762# cap_shunt_p a_24452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X9877 a_3036_27464# a_2948_27508# vss vss nmos_6p0 w=0.82u l=1u
X9878 a_35868_48376# cap_shunt_gyp a_35600_48438# vss nmos_6p0 w=0.82u l=0.6u
X9879 a_27888_7608# cap_series_gyn a_25780_7608# vss nmos_6p0 w=0.82u l=0.6u
X9880 a_10864_9476# cap_shunt_p a_9540_9538# vss nmos_6p0 w=0.82u l=0.6u
X9881 vdd a_35180_11351# a_35092_11448# vdd pmos_6p0 w=1.22u l=1u
X9882 vss cap_shunt_p a_11200_15448# vss nmos_6p0 w=0.82u l=0.6u
X9883 a_20172_47415# a_20084_47512# vss vss nmos_6p0 w=0.82u l=1u
X9884 vss cap_shunt_n a_23072_37700# vss nmos_6p0 w=0.82u l=0.6u
X9885 a_6532_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9886 vdd tune_series_gy[4] a_22436_7124# vdd pmos_6p0 w=1.2u l=0.5u
X9887 a_29744_9476# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X9888 a_10340_32212# cap_shunt_n a_10548_32696# vdd pmos_6p0 w=1.2u l=0.5u
X9889 a_28692_29560# cap_shunt_p a_30408_29560# vss nmos_6p0 w=0.82u l=0.6u
X9890 a_30616_19668# cap_series_gygyn a_30428_19668# vdd pmos_6p0 w=1.2u l=0.5u
X9891 a_19936_26424# cap_shunt_n a_17828_26424# vss nmos_6p0 w=0.82u l=0.6u
X9892 a_20740_26424# cap_shunt_n a_20532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X9893 a_3036_24328# a_2948_24372# vss vss nmos_6p0 w=0.82u l=1u
X9894 a_2140_45847# a_2052_45944# vss vss nmos_6p0 w=0.82u l=1u
X9895 a_24452_9884# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9896 a_22644_12312# cap_series_gyn a_22436_11828# vdd pmos_6p0 w=1.2u l=0.5u
X9897 vss tune_shunt[7] a_13796_17378# vss nmos_6p0 w=0.51u l=0.6u
X9898 a_6532_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9899 a_28692_26424# cap_shunt_p a_30408_26424# vss nmos_6p0 w=0.82u l=0.6u
X9900 vss tune_series_gy[4] a_14692_10744# vss nmos_6p0 w=0.51u l=0.6u
X9901 a_10660_4834# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X9902 a_33612_17623# a_33524_17720# vss vss nmos_6p0 w=0.82u l=1u
X9903 a_16708_29922# cap_shunt_n a_17640_29860# vss nmos_6p0 w=0.82u l=0.6u
X9904 vss tune_shunt[7] a_24660_23650# vss nmos_6p0 w=0.51u l=0.6u
X9905 a_20740_23288# cap_shunt_p a_20532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X9906 vss cap_shunt_p a_8848_21720# vss nmos_6p0 w=0.82u l=0.6u
X9907 a_2140_42711# a_2052_42808# vss vss nmos_6p0 w=0.82u l=1u
X9908 vss tune_shunt[5] a_29700_36194# vss nmos_6p0 w=0.51u l=0.6u
X9909 a_11592_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9910 a_24452_6748# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9911 vdd a_35628_31735# a_35540_31832# vdd pmos_6p0 w=1.22u l=1u
X9912 a_9540_12674# cap_shunt_p a_10472_12612# vss nmos_6p0 w=0.82u l=0.6u
X9913 a_13252_27508# cap_shunt_n a_13460_27992# vdd pmos_6p0 w=1.2u l=0.5u
X9914 a_16708_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X9915 a_16500_34972# cap_shunt_n a_16708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X9916 a_16708_26786# cap_shunt_n a_17640_26724# vss nmos_6p0 w=0.82u l=0.6u
X9917 vdd a_8860_9783# a_8772_9880# vdd pmos_6p0 w=1.22u l=1u
X9918 vss tune_shunt[5] a_29700_33058# vss nmos_6p0 w=0.51u l=0.6u
X9919 a_11592_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9920 vss tune_shunt[7] a_24660_20514# vss nmos_6p0 w=0.51u l=0.6u
X9921 a_7748_25218# cap_shunt_n a_7540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X9922 a_2856_6340# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9923 a_25572_19668# cap_series_gyp a_25780_20152# vdd pmos_6p0 w=1.2u l=0.5u
X9924 vdd a_28572_23895# a_28484_23992# vdd pmos_6p0 w=1.22u l=1u
X9925 a_18388_3266# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X9926 a_24452_25564# cap_shunt_p a_24660_25218# vdd pmos_6p0 w=1.2u l=0.5u
X9927 vss tune_shunt[6] a_6740_45240# vss nmos_6p0 w=0.51u l=0.6u
X9928 a_16500_31836# cap_shunt_n a_16708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X9929 vdd a_24204_29032# a_24116_29076# vdd pmos_6p0 w=1.22u l=1u
X9930 vdd a_33500_14920# a_33412_14964# vdd pmos_6p0 w=1.22u l=1u
X9931 a_29700_36194# cap_shunt_n a_30632_36132# vss nmos_6p0 w=0.82u l=0.6u
X9932 a_28484_27508# cap_shunt_p a_28692_27992# vdd pmos_6p0 w=1.2u l=0.5u
X9933 a_2856_3204# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X9934 vdd a_28572_20759# a_28484_20856# vdd pmos_6p0 w=1.22u l=1u
X9935 vdd a_38092_32168# a_38004_32212# vdd pmos_6p0 w=1.22u l=1u
X9936 a_24452_22428# cap_shunt_p a_24660_22082# vdd pmos_6p0 w=1.2u l=0.5u
X9937 a_1716_8316# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9938 vss tune_shunt[6] a_6740_42104# vss nmos_6p0 w=0.51u l=0.6u
X9939 vdd a_8860_3511# a_8772_3608# vdd pmos_6p0 w=1.22u l=1u
X9940 a_6292_51512# cap_shunt_p a_6084_51028# vdd pmos_6p0 w=1.2u l=0.5u
X9941 a_12580_13396# cap_shunt_p a_12788_13880# vdd pmos_6p0 w=1.2u l=0.5u
X9942 a_35292_41143# a_35204_41240# vss vss nmos_6p0 w=0.82u l=1u
X9943 a_25780_9176# cap_series_gyp a_25572_8692# vdd pmos_6p0 w=1.2u l=0.5u
X9944 a_21540_13020# cap_series_gyn a_21748_12674# vdd pmos_6p0 w=1.2u l=0.5u
X9945 a_5636_8692# cap_shunt_p a_5844_9176# vdd pmos_6p0 w=1.2u l=0.5u
X9946 a_34348_9884# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9947 vdd a_33500_11784# a_33412_11828# vdd pmos_6p0 w=1.22u l=1u
X9948 vdd tune_shunt[5] a_6084_19292# vdd pmos_6p0 w=1.2u l=0.5u
X9949 a_12788_48376# cap_shunt_p a_12580_47892# vdd pmos_6p0 w=1.2u l=0.5u
X9950 vss tune_shunt[6] a_2708_39330# vss nmos_6p0 w=0.51u l=0.6u
X9951 a_37632_33400# cap_shunt_gyp a_37444_33400# vdd pmos_6p0 w=1.215u l=0.5u
X9952 a_15700_9538# cap_series_gyn a_15492_9884# vdd pmos_6p0 w=1.2u l=0.5u
X9953 a_14504_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9954 vss cap_shunt_p a_27104_21720# vss nmos_6p0 w=0.82u l=0.6u
X9955 a_9204_51874# cap_shunt_n a_8996_52220# vdd pmos_6p0 w=1.2u l=0.5u
X9956 a_6532_46324# cap_shunt_p a_6740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X9957 a_9072_39268# cap_shunt_n a_7748_39330# vss nmos_6p0 w=0.82u l=0.6u
X9958 a_12444_20759# a_12356_20856# vss vss nmos_6p0 w=0.82u l=1u
X9959 a_9316_47170# cap_shunt_p a_9108_47516# vdd pmos_6p0 w=1.2u l=0.5u
X9960 a_7748_34626# cap_shunt_n a_7540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X9961 a_16700_55255# a_16612_55352# vss vss nmos_6p0 w=0.82u l=1u
X9962 a_22680_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X9963 a_25780_6040# cap_series_gyp a_25572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X9964 a_38092_27464# a_38004_27508# vss vss nmos_6p0 w=0.82u l=1u
X9965 a_34348_6748# tune_series_gygy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9966 vdd tune_shunt[5] a_6084_16156# vdd pmos_6p0 w=1.2u l=0.5u
X9967 vdd a_20620_34871# a_20532_34968# vdd pmos_6p0 w=1.22u l=1u
X9968 a_15700_6402# cap_series_gyp a_15492_6748# vdd pmos_6p0 w=1.2u l=0.5u
X9969 vss tune_series_gy[2] a_14468_3266# vss nmos_6p0 w=0.51u l=0.6u
X9970 vdd a_37084_52552# a_36996_52596# vdd pmos_6p0 w=1.22u l=1u
X9971 a_21540_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X9972 a_7748_31490# cap_shunt_n a_7540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X9973 a_28484_36916# cap_shunt_p a_28692_37400# vdd pmos_6p0 w=1.2u l=0.5u
X9974 a_16476_50984# a_16388_51028# vss vss nmos_6p0 w=0.82u l=1u
X9975 a_35880_36916# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X9976 vdd a_23756_25896# a_23668_25940# vdd pmos_6p0 w=1.22u l=1u
X9977 a_35880_24372# cap_series_gygyp a_35692_24372# vdd pmos_6p0 w=1.2u l=0.5u
X9978 a_6572_5556# cap_series_gyp a_6760_5556# vdd pmos_6p0 w=1.2u l=0.5u
X9979 a_21540_8316# cap_series_gyp a_21748_7970# vdd pmos_6p0 w=1.2u l=0.5u
X9980 a_28796_43144# a_28708_43188# vss vss nmos_6p0 w=0.82u l=1u
X9981 a_34536_6748# tune_series_gygy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X9982 vdd a_34396_3511# a_34308_3608# vdd pmos_6p0 w=1.22u l=1u
X9983 a_26768_7908# cap_series_gyp a_24660_7970# vss nmos_6p0 w=0.82u l=0.6u
X9984 a_11256_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9985 a_19936_17016# cap_shunt_p a_17828_17016# vss nmos_6p0 w=0.82u l=0.6u
X9986 vdd a_31260_38440# a_31172_38484# vdd pmos_6p0 w=1.22u l=1u
X9987 a_9108_22428# cap_shunt_p a_9316_22082# vdd pmos_6p0 w=1.2u l=0.5u
X9988 vss tune_series_gy[5] a_19732_7608# vss nmos_6p0 w=0.51u l=0.6u
X9989 a_3036_14920# a_2948_14964# vss vss nmos_6p0 w=0.82u l=1u
X9990 a_20740_17016# cap_shunt_p a_20532_16532# vdd pmos_6p0 w=1.2u l=0.5u
X9991 a_2140_36439# a_2052_36536# vss vss nmos_6p0 w=0.82u l=1u
X9992 vdd a_35628_25463# a_35540_25560# vdd pmos_6p0 w=1.22u l=1u
X9993 a_3640_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X9994 a_3828_20152# cap_shunt_p a_3620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X9995 vdd a_23756_22760# a_23668_22804# vdd pmos_6p0 w=1.22u l=1u
X9996 a_37548_51512# cap_shunt_gyp a_37280_51574# vss nmos_6p0 w=0.82u l=0.6u
X9997 a_35880_21236# cap_series_gygyp a_35692_21236# vdd pmos_6p0 w=1.2u l=0.5u
X9998 a_28692_17016# cap_series_gyn a_30408_17016# vss nmos_6p0 w=0.82u l=0.6u
X9999 vss tune_shunt[7] a_10548_37400# vss nmos_6p0 w=0.51u l=0.6u
X10000 vss tune_shunt[4] a_28692_40536# vss nmos_6p0 w=0.51u l=0.6u
X10001 vss cap_series_gyp a_16800_4472# vss nmos_6p0 w=0.82u l=0.6u
X10002 a_9668_10260# cap_shunt_p a_9876_10744# vdd pmos_6p0 w=1.2u l=0.5u
X10003 vss cap_shunt_p a_8848_12312# vss nmos_6p0 w=0.82u l=0.6u
X10004 a_11668_43672# cap_shunt_n a_11460_43188# vdd pmos_6p0 w=1.2u l=0.5u
X10005 vdd a_31260_35304# a_31172_35348# vdd pmos_6p0 w=1.22u l=1u
X10006 a_34536_9884# cap_series_gygyn a_34560_9476# vss nmos_6p0 w=0.82u l=0.6u
X10007 a_9668_10260# cap_shunt_p a_9876_10744# vdd pmos_6p0 w=1.2u l=0.5u
X10008 vss tune_series_gy[5] a_24660_14242# vss nmos_6p0 w=0.51u l=0.6u
X10009 vdd tune_shunt[7] a_9220_17724# vdd pmos_6p0 w=1.2u l=0.5u
X10010 a_28692_7608# cap_series_gyp a_28484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X10011 a_5836_3944# a_5748_3988# vss vss nmos_6p0 w=0.82u l=1u
X10012 a_11200_17016# cap_shunt_p a_9876_17016# vss nmos_6p0 w=0.82u l=0.6u
X10013 a_24660_37762# cap_shunt_p a_24452_38108# vdd pmos_6p0 w=1.2u l=0.5u
X10014 a_37632_40053# cap_shunt_gyn a_37444_40053# vdd pmos_6p0 w=1.215u l=0.5u
X10015 a_31416_39268# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10016 a_18612_7970# cap_series_gyp a_18404_8316# vdd pmos_6p0 w=1.2u l=0.5u
X10017 vss tune_shunt[6] a_7748_45602# vss nmos_6p0 w=0.51u l=0.6u
X10018 a_7748_44034# cap_shunt_p a_8680_43972# vss nmos_6p0 w=0.82u l=0.6u
X10019 a_16500_25564# cap_shunt_n a_16708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X10020 a_21316_3612# cap_series_gyp a_21524_3266# vdd pmos_6p0 w=1.2u l=0.5u
X10021 a_16708_17378# cap_shunt_p a_17640_17316# vss nmos_6p0 w=0.82u l=0.6u
X10022 a_24452_19292# cap_series_gyn a_24660_18946# vdd pmos_6p0 w=1.2u l=0.5u
X10023 vss tune_series_gy[4] a_25780_9176# vss nmos_6p0 w=0.51u l=0.6u
X10024 vss tune_series_gy[5] a_24660_11106# vss nmos_6p0 w=0.51u l=0.6u
X10025 a_2932_9176# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X10026 a_30616_19668# cap_series_gygyn a_30428_19668# vdd pmos_6p0 w=1.2u l=0.5u
X10027 a_22848_37400# cap_shunt_n a_20740_37400# vss nmos_6p0 w=0.82u l=0.6u
X10028 a_11800_7124# cap_series_gyp a_11612_7124# vdd pmos_6p0 w=1.2u l=0.5u
X10029 a_20740_26424# cap_shunt_n a_20532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X10030 a_24660_22082# cap_shunt_p a_26376_22020# vss nmos_6p0 w=0.82u l=0.6u
X10031 vdd a_23532_55688# a_23444_55732# vdd pmos_6p0 w=1.22u l=1u
X10032 a_11668_46808# cap_shunt_n a_11460_46324# vdd pmos_6p0 w=1.2u l=0.5u
X10033 vdd a_28572_14487# a_28484_14584# vdd pmos_6p0 w=1.22u l=1u
X10034 a_16924_52552# a_16836_52596# vss vss nmos_6p0 w=0.82u l=1u
X10035 a_7748_40898# cap_shunt_n a_8680_40836# vss nmos_6p0 w=0.82u l=0.6u
X10036 a_2500_30268# cap_shunt_n a_2708_29922# vdd pmos_6p0 w=1.2u l=0.5u
X10037 a_16500_22428# cap_shunt_n a_16708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X10038 a_24452_16156# cap_series_gyn a_24660_15810# vdd pmos_6p0 w=1.2u l=0.5u
X10039 a_10548_3266# cap_series_gyn a_10340_3612# vdd pmos_6p0 w=1.2u l=0.5u
X10040 vss tune_series_gy[5] a_19732_13880# vss nmos_6p0 w=0.51u l=0.6u
X10041 vss cap_series_gygyp a_36624_20452# vss nmos_6p0 w=0.82u l=0.6u
X10042 a_2708_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10043 a_10548_37400# cap_shunt_n a_11480_37400# vss nmos_6p0 w=0.82u l=0.6u
X10044 a_20740_23288# cap_shunt_p a_20532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X10045 a_28484_14964# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10046 a_16500_28700# cap_shunt_n a_16708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X10047 a_31436_8316# tune_series_gygy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10048 vdd a_28572_11351# a_28484_11448# vdd pmos_6p0 w=1.22u l=1u
X10049 a_25996_53687# a_25908_53784# vss vss nmos_6p0 w=0.82u l=1u
X10050 a_18760_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10051 vdd a_20508_55688# a_20420_55732# vdd pmos_6p0 w=1.22u l=1u
X10052 vdd tune_shunt[6] a_10340_38484# vdd pmos_6p0 w=1.2u l=0.5u
X10053 a_20532_33780# cap_shunt_n a_20740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X10054 vdd tune_shunt[6] a_3620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X10055 vdd tune_shunt[7] a_21540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X10056 vss tune_series_gy[5] a_19732_10744# vss nmos_6p0 w=0.51u l=0.6u
X10057 a_25592_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10058 a_25780_4472# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X10059 a_24660_44034# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X10060 vdd a_20620_28599# a_20532_28696# vdd pmos_6p0 w=1.22u l=1u
X10061 vdd a_24204_55255# a_24116_55352# vdd pmos_6p0 w=1.22u l=1u
X10062 a_16500_34972# cap_shunt_n a_16708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X10063 a_28484_11828# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10064 vss cap_series_gyp a_27104_12312# vss nmos_6p0 w=0.82u l=0.6u
X10065 vdd a_12780_47415# a_12692_47512# vdd pmos_6p0 w=1.22u l=1u
X10066 a_17620_40052# cap_shunt_n a_17828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X10067 a_25996_50551# a_25908_50648# vss vss nmos_6p0 w=0.82u l=1u
X10068 vss tune_shunt_gy[6] a_37632_50648# vss nmos_6p0 w=0.51u l=0.6u
X10069 vdd tune_shunt[7] a_10340_35348# vdd pmos_6p0 w=1.2u l=0.5u
X10070 a_20532_30644# cap_shunt_n a_20740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X10071 a_7748_25218# cap_shunt_n a_7540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X10072 vss cap_series_gygyn a_32040_22020# vss nmos_6p0 w=0.82u l=0.6u
X10073 vss tune_shunt[7] a_12788_18584# vss nmos_6p0 w=0.51u l=0.6u
X10074 a_25572_19668# cap_series_gyp a_25780_20152# vdd pmos_6p0 w=1.2u l=0.5u
X10075 vdd a_24652_44712# a_24564_44756# vdd pmos_6p0 w=1.22u l=1u
X10076 vdd a_24204_52119# a_24116_52216# vdd pmos_6p0 w=1.22u l=1u
X10077 a_16500_31836# cap_shunt_n a_16708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X10078 vss cap_shunt_n a_22848_27992# vss nmos_6p0 w=0.82u l=0.6u
X10079 a_30924_55688# a_30836_55732# vss vss nmos_6p0 w=0.82u l=1u
X10080 a_35292_7080# a_35204_7124# vss vss nmos_6p0 w=0.82u l=1u
X10081 a_28484_27508# cap_shunt_p a_28692_27992# vdd pmos_6p0 w=1.2u l=0.5u
X10082 vss tune_shunt[7] a_12788_15448# vss nmos_6p0 w=0.51u l=0.6u
X10083 a_29720_16156# cap_series_gyn a_29532_16156# vdd pmos_6p0 w=1.2u l=0.5u
X10084 a_37548_45240# cap_shunt_gyp a_37280_45302# vss nmos_6p0 w=0.82u l=0.6u
X10085 vss tune_shunt[2] a_1924_4472# vss nmos_6p0 w=0.51u l=0.6u
X10086 vdd a_23756_16488# a_23668_16532# vdd pmos_6p0 w=1.22u l=1u
X10087 a_14728_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10088 vss cap_shunt_n a_22848_24856# vss nmos_6p0 w=0.82u l=0.6u
X10089 a_5936_21720# cap_shunt_p a_3828_21720# vss nmos_6p0 w=0.82u l=0.6u
X10090 vss tune_shunt[6] a_28692_34264# vss nmos_6p0 w=0.51u l=0.6u
X10091 vdd a_31260_29032# a_31172_29076# vdd pmos_6p0 w=1.22u l=1u
X10092 a_9540_9538# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10093 a_30136_15748# cap_series_gyn a_29720_16156# vss nmos_6p0 w=0.82u l=0.6u
X10094 a_34308_20860# cap_series_gygyp a_34516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X10095 a_29624_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10096 a_24660_29922# cap_shunt_n a_24452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X10097 a_14728_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10098 a_12788_18584# cap_shunt_p a_13720_18584# vss nmos_6p0 w=0.82u l=0.6u
X10099 vdd tune_shunt[6] a_17620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X10100 vss tune_shunt[6] a_7748_39330# vss nmos_6p0 w=0.51u l=0.6u
X10101 vss tune_shunt[5] a_28692_31128# vss nmos_6p0 w=0.51u l=0.6u
X10102 a_18612_4834# cap_series_gyp a_18404_5180# vdd pmos_6p0 w=1.2u l=0.5u
X10103 a_16500_19292# cap_shunt_p a_16708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X10104 vdd a_30812_41143# a_30724_41240# vdd pmos_6p0 w=1.22u l=1u
X10105 a_8456_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10106 a_33524_32212# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10107 a_20844_47848# a_20756_47892# vss vss nmos_6p0 w=0.82u l=1u
X10108 vdd a_9644_43144# a_9556_43188# vdd pmos_6p0 w=1.22u l=1u
X10109 a_28484_36916# cap_shunt_p a_28692_37400# vdd pmos_6p0 w=1.2u l=0.5u
X10110 vss cap_shunt_p a_8736_12612# vss nmos_6p0 w=0.82u l=0.6u
X10111 vdd a_36076_36439# a_35988_36536# vdd pmos_6p0 w=1.22u l=1u
X10112 a_32612_34626# cap_shunt_n a_32404_34972# vdd pmos_6p0 w=1.2u l=0.5u
X10113 a_12788_15448# cap_shunt_p a_13720_15448# vss nmos_6p0 w=0.82u l=0.6u
X10114 a_24660_37762# cap_shunt_p a_25592_37700# vss nmos_6p0 w=0.82u l=0.6u
X10115 a_7748_34626# cap_shunt_n a_8680_34564# vss nmos_6p0 w=0.82u l=0.6u
X10116 a_21540_42812# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10117 a_16500_16156# cap_shunt_p a_16708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X10118 a_33936_37700# cap_shunt_p a_32612_37762# vss nmos_6p0 w=0.82u l=0.6u
X10119 a_20740_20152# cap_shunt_p a_22456_20152# vss nmos_6p0 w=0.82u l=0.6u
X10120 a_2500_28700# cap_shunt_n a_2708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X10121 a_35488_42166# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X10122 vdd a_19724_33303# a_19636_33400# vdd pmos_6p0 w=1.22u l=1u
X10123 a_32612_31490# cap_shunt_n a_32404_31836# vdd pmos_6p0 w=1.2u l=0.5u
X10124 a_9108_22428# cap_shunt_p a_9316_22082# vdd pmos_6p0 w=1.2u l=0.5u
X10125 a_29196_3612# cap_series_gyn a_29384_3612# vdd pmos_6p0 w=1.2u l=0.5u
X10126 a_2724_11828# cap_shunt_n a_2932_12312# vdd pmos_6p0 w=1.2u l=0.5u
X10127 a_20740_17016# cap_shunt_p a_20532_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10128 vdd tune_series_gy[4] a_25572_18100# vdd pmos_6p0 w=1.2u l=0.5u
X10129 a_7748_31490# cap_shunt_n a_8680_31428# vss nmos_6p0 w=0.82u l=0.6u
X10130 a_25592_14180# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X10131 a_20732_55255# a_20644_55352# vss vss nmos_6p0 w=0.82u l=1u
X10132 a_16708_47170# cap_shunt_n a_16500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X10133 a_17828_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10134 a_2708_22082# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10135 vdd a_29916_53687# a_29828_53784# vdd pmos_6p0 w=1.22u l=1u
X10136 vdd a_24204_48983# a_24116_49080# vdd pmos_6p0 w=1.22u l=1u
X10137 a_7540_38108# cap_shunt_n a_7748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X10138 a_10248_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10139 vdd tune_shunt[2] a_1716_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10140 a_10492_8316# cap_series_gyp a_10680_8316# vdd pmos_6p0 w=1.2u l=0.5u
X10141 a_6760_5556# cap_series_gyp a_6572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10142 a_35840_4772# cap_series_gygyp a_34516_4834# vss nmos_6p0 w=0.82u l=0.6u
X10143 a_8680_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10144 vdd tune_shunt[7] a_10340_29076# vdd pmos_6p0 w=1.2u l=0.5u
X10145 vdd tune_shunt[7] a_9220_17724# vdd pmos_6p0 w=1.2u l=0.5u
X10146 a_20532_24372# cap_shunt_n a_20740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X10147 a_25592_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X10148 a_15512_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10149 a_35880_3988# cap_series_gygyp a_36688_4472# vss nmos_6p0 w=0.82u l=0.6u
X10150 a_13252_25940# cap_shunt_n a_13460_26424# vdd pmos_6p0 w=1.2u l=0.5u
X10151 vdd a_20620_19191# a_20532_19288# vdd pmos_6p0 w=1.22u l=1u
X10152 a_16812_50551# a_16724_50648# vss vss nmos_6p0 w=0.82u l=1u
X10153 vdd a_24652_38440# a_24564_38484# vdd pmos_6p0 w=1.22u l=1u
X10154 a_13796_29922# cap_shunt_n a_15512_29860# vss nmos_6p0 w=0.82u l=0.6u
X10155 vdd a_29916_50551# a_29828_50648# vdd pmos_6p0 w=1.22u l=1u
X10156 a_7540_42812# cap_shunt_n a_7748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X10157 a_23856_29860# cap_shunt_n a_21748_29922# vss nmos_6p0 w=0.82u l=0.6u
X10158 a_16500_25564# cap_shunt_n a_16708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X10159 a_25780_37400# cap_shunt_p a_25572_36916# vdd pmos_6p0 w=1.2u l=0.5u
X10160 a_3620_25940# cap_shunt_p a_3828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X10161 a_8680_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10162 a_13796_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10163 a_14692_7608# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X10164 a_6784_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X10165 a_20532_21236# cap_shunt_p a_20740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X10166 a_20532_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10167 vss tune_shunt[6] a_28692_37400# vss nmos_6p0 w=0.51u l=0.6u
X10168 a_13252_22804# cap_shunt_n a_13460_23288# vdd pmos_6p0 w=1.2u l=0.5u
X10169 a_31708_38440# a_31620_38484# vss vss nmos_6p0 w=0.82u l=1u
X10170 vdd a_24652_35304# a_24564_35348# vdd pmos_6p0 w=1.22u l=1u
X10171 a_13796_26786# cap_shunt_n a_15512_26724# vss nmos_6p0 w=0.82u l=0.6u
X10172 a_23856_26724# cap_shunt_n a_21748_26786# vss nmos_6p0 w=0.82u l=0.6u
X10173 a_16500_22428# cap_shunt_n a_16708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X10174 vss cap_shunt_p a_22848_18584# vss nmos_6p0 w=0.82u l=0.6u
X10175 a_33948_21192# a_33860_21236# vss vss nmos_6p0 w=0.82u l=1u
X10176 a_37280_51029# cap_shunt_gyp a_37280_51574# vdd pmos_6p0 w=1.215u l=0.5u
X10177 a_3620_22804# cap_shunt_p a_3828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X10178 a_28484_18100# cap_series_gyp a_28692_18584# vdd pmos_6p0 w=1.2u l=0.5u
X10179 vss tune_shunt[7] a_3828_32696# vss nmos_6p0 w=0.51u l=0.6u
X10180 vdd tune_shunt[5] a_6084_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10181 vdd a_29468_45847# a_29380_45944# vdd pmos_6p0 w=1.22u l=1u
X10182 vss tune_shunt[5] a_6292_48738# vss nmos_6p0 w=0.51u l=0.6u
X10183 vdd tune_shunt[7] a_6532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X10184 vdd tune_shunt[7] a_9668_13396# vdd pmos_6p0 w=1.2u l=0.5u
X10185 a_10660_28354# cap_shunt_n a_10452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X10186 vdd tune_shunt[6] a_10340_38484# vdd pmos_6p0 w=1.2u l=0.5u
X10187 a_20532_33780# cap_shunt_n a_20740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X10188 vss cap_series_gyn a_22848_15448# vss nmos_6p0 w=0.82u l=0.6u
X10189 a_21316_3612# cap_series_gyp a_21524_3266# vdd pmos_6p0 w=1.2u l=0.5u
X10190 vdd a_29468_42711# a_29380_42808# vdd pmos_6p0 w=1.22u l=1u
X10191 vss cap_shunt_p a_25984_32996# vss nmos_6p0 w=0.82u l=0.6u
X10192 a_34328_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10193 vdd tune_shunt[7] a_6532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X10194 a_8456_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10195 vss cap_shunt_p a_5936_46808# vss nmos_6p0 w=0.82u l=0.6u
X10196 vdd tune_shunt[7] a_10340_35348# vdd pmos_6p0 w=1.2u l=0.5u
X10197 a_20532_30644# cap_shunt_n a_20740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X10198 a_24660_6402# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X10199 vdd tune_shunt[7] a_9332_13020# vdd pmos_6p0 w=1.2u l=0.5u
X10200 a_14728_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10201 a_7748_28354# cap_shunt_n a_8680_28292# vss nmos_6p0 w=0.82u l=0.6u
X10202 a_24452_9884# cap_series_gyn a_24660_9538# vdd pmos_6p0 w=1.2u l=0.5u
X10203 a_21540_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10204 a_29196_3612# tune_series_gy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10205 a_28236_54120# a_28148_54164# vss vss nmos_6p0 w=0.82u l=1u
X10206 a_29492_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10207 a_8456_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10208 a_9316_22082# cap_shunt_p a_11032_22020# vss nmos_6p0 w=0.82u l=0.6u
X10209 vdd a_31260_55255# a_31172_55352# vdd pmos_6p0 w=1.22u l=1u
X10210 a_20740_35832# cap_shunt_n a_21672_35832# vss nmos_6p0 w=0.82u l=0.6u
X10211 a_3828_32696# cap_shunt_p a_4760_32696# vss nmos_6p0 w=0.82u l=0.6u
X10212 vss cap_shunt_p a_18816_20452# vss nmos_6p0 w=0.82u l=0.6u
X10213 a_28484_27508# cap_shunt_p a_28692_27992# vdd pmos_6p0 w=1.2u l=0.5u
X10214 vdd a_36076_27031# a_35988_27128# vdd pmos_6p0 w=1.22u l=1u
X10215 a_7748_25218# cap_shunt_n a_8680_25156# vss nmos_6p0 w=0.82u l=0.6u
X10216 a_32612_25218# cap_shunt_p a_32404_25564# vdd pmos_6p0 w=1.2u l=0.5u
X10217 a_24452_6748# cap_series_gyn a_24660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X10218 a_2708_12674# cap_shunt_n a_3640_12612# vss nmos_6p0 w=0.82u l=0.6u
X10219 a_2500_20860# cap_shunt_p a_2708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X10220 a_21540_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10221 vdd tune_shunt[7] a_24452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X10222 a_29720_16156# cap_series_gyn a_29532_16156# vdd pmos_6p0 w=1.2u l=0.5u
X10223 a_15568_21720# cap_shunt_n a_13460_21720# vss nmos_6p0 w=0.82u l=0.6u
X10224 a_2708_48738# cap_shunt_p a_2500_49084# vdd pmos_6p0 w=1.2u l=0.5u
X10225 a_29492_31836# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10226 a_10660_29922# cap_shunt_n a_10452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X10227 a_12788_13880# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10228 vdd a_13788_10216# a_13700_10260# vdd pmos_6p0 w=1.22u l=1u
X10229 vdd a_31260_52119# a_31172_52216# vdd pmos_6p0 w=1.22u l=1u
X10230 a_4032_50244# cap_shunt_n a_2708_50306# vss nmos_6p0 w=0.82u l=0.6u
X10231 a_27888_13880# cap_series_gyn a_25780_13880# vss nmos_6p0 w=0.82u l=0.6u
X10232 a_34308_20860# cap_series_gygyp a_34516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X10233 a_22524_50984# a_22436_51028# vss vss nmos_6p0 w=0.82u l=1u
X10234 a_11592_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10235 a_7540_30268# cap_shunt_n a_7748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X10236 vss tune_shunt[7] a_16708_31490# vss nmos_6p0 w=0.51u l=0.6u
X10237 vss tune_shunt[7] a_6628_14242# vss nmos_6p0 w=0.51u l=0.6u
X10238 vdd a_11996_19191# a_11908_19288# vdd pmos_6p0 w=1.22u l=1u
X10239 a_16708_37762# cap_shunt_n a_16500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X10240 a_24660_29922# cap_shunt_n a_24452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X10241 a_17828_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10242 vdd a_29916_44279# a_29828_44376# vdd pmos_6p0 w=1.22u l=1u
X10243 a_7540_36540# cap_shunt_n a_7748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X10244 a_28692_32696# cap_shunt_p a_28484_32212# vdd pmos_6p0 w=1.2u l=0.5u
X10245 a_16500_19292# cap_shunt_p a_16708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X10246 a_4760_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10247 a_27888_10744# cap_series_gyn a_25780_10744# vss nmos_6p0 w=0.82u l=0.6u
X10248 vdd a_4380_54120# a_4292_54164# vdd pmos_6p0 w=1.22u l=1u
X10249 a_33024_43972# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10250 a_35692_36916# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10251 a_8680_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10252 a_21636_6040# cap_series_gyp a_21428_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10253 a_16708_42466# cap_shunt_n a_16500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X10254 a_9316_47170# cap_shunt_p a_10248_47108# vss nmos_6p0 w=0.82u l=0.6u
X10255 vdd a_32380_3511# a_32292_3608# vdd pmos_6p0 w=1.22u l=1u
X10256 a_18612_11106# cap_series_gyn a_20328_11044# vss nmos_6p0 w=0.82u l=0.6u
X10257 a_9220_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10258 vdd a_24652_29032# a_24564_29076# vdd pmos_6p0 w=1.22u l=1u
X10259 a_10660_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10260 vdd tune_shunt[5] a_6084_50652# vdd pmos_6p0 w=1.2u l=0.5u
X10261 a_34844_40008# a_34756_40052# vss vss nmos_6p0 w=0.82u l=1u
X10262 a_7540_33404# cap_shunt_n a_7748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X10263 a_16500_16156# cap_shunt_p a_16708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X10264 a_4760_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10265 a_25780_27992# cap_shunt_p a_25572_27508# vdd pmos_6p0 w=1.2u l=0.5u
X10266 a_6060_14487# a_5972_14584# vss vss nmos_6p0 w=0.82u l=1u
X10267 a_13796_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10268 vss cap_shunt_n a_12992_46808# vss nmos_6p0 w=0.82u l=0.6u
X10269 a_6532_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10270 a_20740_46808# cap_shunt_p a_20532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X10271 a_13796_17378# cap_shunt_p a_15512_17316# vss nmos_6p0 w=0.82u l=0.6u
X10272 a_33948_11784# a_33860_11828# vss vss nmos_6p0 w=0.82u l=1u
X10273 a_3864_12312# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10274 a_23856_17316# cap_shunt_p a_21748_17378# vss nmos_6p0 w=0.82u l=0.6u
X10275 vdd tune_shunt[7] a_13588_28700# vdd pmos_6p0 w=1.2u l=0.5u
X10276 vdd tune_shunt[7] a_21540_20860# vdd pmos_6p0 w=1.2u l=0.5u
X10277 vss tune_shunt[7] a_3828_23288# vss nmos_6p0 w=0.51u l=0.6u
X10278 a_12892_20759# a_12804_20856# vss vss nmos_6p0 w=0.82u l=1u
X10279 a_25780_43672# cap_shunt_p a_27496_43672# vss nmos_6p0 w=0.82u l=0.6u
X10280 vdd tune_shunt[7] a_6532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X10281 a_37420_8215# a_37332_8312# vss vss nmos_6p0 w=0.82u l=1u
X10282 a_30812_47415# a_30724_47512# vss vss nmos_6p0 w=0.82u l=1u
X10283 vdd tune_shunt[7] a_10340_29076# vdd pmos_6p0 w=1.2u l=0.5u
X10284 a_20532_24372# cap_shunt_n a_20740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X10285 a_27228_5079# a_27140_5176# vss vss nmos_6p0 w=0.82u l=1u
X10286 vss tune_series_gy[5] a_22644_12312# vss nmos_6p0 w=0.51u l=0.6u
X10287 a_22456_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10288 a_15804_49416# a_15716_49460# vss vss nmos_6p0 w=0.82u l=1u
X10289 vdd a_23308_41576# a_23220_41620# vdd pmos_6p0 w=1.22u l=1u
X10290 a_13252_25940# cap_shunt_n a_13460_26424# vdd pmos_6p0 w=1.2u l=0.5u
X10291 vss cap_shunt_p a_25984_23588# vss nmos_6p0 w=0.82u l=0.6u
X10292 a_28692_12312# cap_series_gyn a_29624_12312# vss nmos_6p0 w=0.82u l=0.6u
X10293 vdd a_32156_13352# a_32068_13396# vdd pmos_6p0 w=1.22u l=1u
X10294 a_28236_47848# a_28148_47892# vss vss nmos_6p0 w=0.82u l=1u
X10295 a_14580_43672# cap_shunt_n a_16296_43672# vss nmos_6p0 w=0.82u l=0.6u
X10296 a_25780_40536# cap_shunt_n a_27496_40536# vss nmos_6p0 w=0.82u l=0.6u
X10297 vss tune_series_gy[2] a_10660_4834# vss nmos_6p0 w=0.51u l=0.6u
X10298 a_21540_8316# cap_series_gyp a_21748_7970# vdd pmos_6p0 w=1.2u l=0.5u
X10299 a_35904_20152# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X10300 vdd tune_shunt[7] a_6532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X10301 vss cap_shunt_p a_11536_18884# vss nmos_6p0 w=0.82u l=0.6u
X10302 vss tune_shunt[5] a_3380_18584# vss nmos_6p0 w=0.51u l=0.6u
X10303 vss cap_shunt_p a_15120_45540# vss nmos_6p0 w=0.82u l=0.6u
X10304 a_6740_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10305 a_32404_38108# cap_shunt_p a_32612_37762# vdd pmos_6p0 w=1.2u l=0.5u
X10306 a_25780_37400# cap_shunt_p a_25572_36916# vdd pmos_6p0 w=1.2u l=0.5u
X10307 vdd tune_series_gy[5] a_28484_13396# vdd pmos_6p0 w=1.2u l=0.5u
X10308 vss cap_shunt_p a_18816_14180# vss nmos_6p0 w=0.82u l=0.6u
X10309 vdd a_31260_48983# a_31172_49080# vdd pmos_6p0 w=1.22u l=1u
X10310 a_34412_43972# cap_shunt_gyp a_34144_43972# vss nmos_6p0 w=0.82u l=0.6u
X10311 a_20740_29560# cap_shunt_n a_21672_29560# vss nmos_6p0 w=0.82u l=0.6u
X10312 a_20532_21236# cap_shunt_p a_20740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X10313 a_34144_44376# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X10314 a_13252_22804# cap_shunt_n a_13460_23288# vdd pmos_6p0 w=1.2u l=0.5u
X10315 a_14580_40536# cap_shunt_n a_16296_40536# vss nmos_6p0 w=0.82u l=0.6u
X10316 a_21540_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10317 vss tune_shunt[7] a_13460_32696# vss nmos_6p0 w=0.51u l=0.6u
X10318 a_29492_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10319 vss cap_shunt_n a_15120_42404# vss nmos_6p0 w=0.82u l=0.6u
X10320 a_21636_6040# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X10321 a_6740_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10322 vdd tune_shunt[7] a_13588_30268# vdd pmos_6p0 w=1.2u l=0.5u
X10323 a_20740_26424# cap_shunt_n a_21672_26424# vss nmos_6p0 w=0.82u l=0.6u
X10324 a_3828_23288# cap_shunt_p a_4760_23288# vss nmos_6p0 w=0.82u l=0.6u
X10325 a_25572_14964# cap_series_gyp a_25780_15448# vdd pmos_6p0 w=1.2u l=0.5u
X10326 vdd tune_shunt[5] a_6084_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10327 vdd a_33948_53687# a_33860_53784# vdd pmos_6p0 w=1.22u l=1u
X10328 a_18424_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10329 a_27228_30167# a_27140_30264# vss vss nmos_6p0 w=0.82u l=1u
X10330 a_2500_11452# cap_shunt_n a_2708_11106# vdd pmos_6p0 w=1.2u l=0.5u
X10331 vdd tune_series_gy[5] a_24452_14588# vdd pmos_6p0 w=1.2u l=0.5u
X10332 a_2140_55688# a_2052_55732# vss vss nmos_6p0 w=0.82u l=1u
X10333 a_10660_28354# cap_shunt_n a_10452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X10334 a_20532_33780# cap_shunt_n a_20740_34264# vdd pmos_6p0 w=1.2u l=0.5u
X10335 vdd a_8860_8648# a_8772_8692# vdd pmos_6p0 w=1.22u l=1u
X10336 vdd a_5612_17623# a_5524_17720# vdd pmos_6p0 w=1.22u l=1u
X10337 a_20844_50551# a_20756_50648# vss vss nmos_6p0 w=0.82u l=1u
X10338 a_16924_38440# a_16836_38484# vss vss nmos_6p0 w=0.82u l=1u
X10339 a_25572_11828# cap_series_gyp a_25780_12312# vdd pmos_6p0 w=1.2u l=0.5u
X10340 vdd a_33948_50551# a_33860_50648# vdd pmos_6p0 w=1.22u l=1u
X10341 a_14372_44756# cap_shunt_p a_14580_45240# vdd pmos_6p0 w=1.2u l=0.5u
X10342 a_18424_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10343 a_27228_27031# a_27140_27128# vss vss nmos_6p0 w=0.82u l=1u
X10344 a_9540_9538# cap_shunt_p a_9332_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10345 a_19732_12312# cap_series_gyn a_19524_11828# vdd pmos_6p0 w=1.2u l=0.5u
X10346 vss tune_shunt[7] a_16708_22082# vss nmos_6p0 w=0.51u l=0.6u
X10347 a_2708_42466# cap_shunt_p a_2500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X10348 a_20532_30644# cap_shunt_n a_20740_31128# vdd pmos_6p0 w=1.2u l=0.5u
X10349 vdd a_9532_3511# a_9444_3608# vdd pmos_6p0 w=1.22u l=1u
X10350 a_21540_45948# cap_shunt_p a_21748_45602# vdd pmos_6p0 w=1.2u l=0.5u
X10351 a_16708_36194# cap_shunt_n a_16500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X10352 vdd a_28124_30167# a_28036_30264# vdd pmos_6p0 w=1.22u l=1u
X10353 a_9540_12674# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10354 a_22412_52119# a_22324_52216# vss vss nmos_6p0 w=0.82u l=1u
X10355 a_4760_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10356 a_7540_27132# cap_shunt_n a_7748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X10357 vdd tune_shunt[7] a_6308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X10358 a_25444_3266# cap_shunt_p a_27160_3204# vss nmos_6p0 w=0.82u l=0.6u
X10359 vdd a_23980_55688# a_23892_55732# vdd pmos_6p0 w=1.22u l=1u
X10360 a_16708_33058# cap_shunt_n a_16500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X10361 a_9876_18584# cap_shunt_p a_11592_18584# vss nmos_6p0 w=0.82u l=0.6u
X10362 a_29532_9884# cap_series_gyn a_29720_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10363 a_12788_17016# cap_shunt_p a_12580_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10364 a_2500_20860# cap_shunt_p a_2708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X10365 vdd a_9196_55255# a_9108_55352# vdd pmos_6p0 w=1.22u l=1u
X10366 vdd a_27676_8215# a_27588_8312# vdd pmos_6p0 w=1.22u l=1u
X10367 a_19732_9176# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10368 a_29720_16156# cap_series_gyn a_29532_16156# vdd pmos_6p0 w=1.2u l=0.5u
X10369 a_28692_38968# cap_shunt_n a_28484_38484# vdd pmos_6p0 w=1.2u l=0.5u
X10370 a_4760_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10371 a_24660_9538# cap_series_gyn a_24452_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10372 a_35880_36916# cap_series_gygyp a_35904_37400# vss nmos_6p0 w=0.82u l=0.6u
X10373 a_10660_29922# cap_shunt_n a_10452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X10374 a_35292_54120# a_35204_54164# vss vss nmos_6p0 w=0.82u l=1u
X10375 vss tune_shunt_gy[3] a_35168_44376# vss nmos_6p0 w=0.51u l=0.6u
X10376 a_7952_9476# cap_shunt_p a_5844_9538# vss nmos_6p0 w=0.82u l=0.6u
X10377 a_9876_15448# cap_shunt_p a_11592_15448# vss nmos_6p0 w=0.82u l=0.6u
X10378 a_17828_34264# cap_shunt_n a_17620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X10379 vdd a_34396_8648# a_34308_8692# vdd pmos_6p0 w=1.22u l=1u
X10380 a_13588_49084# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10381 a_31708_44279# a_31620_44376# vss vss nmos_6p0 w=0.82u l=1u
X10382 a_7540_30268# cap_shunt_n a_7748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X10383 a_4032_7608# cap_shunt_n a_1924_7608# vss nmos_6p0 w=0.82u l=0.6u
X10384 a_27104_7608# cap_series_gyn a_25780_7608# vss nmos_6p0 w=0.82u l=0.6u
X10385 a_28692_35832# cap_shunt_p a_28484_35348# vdd pmos_6p0 w=1.2u l=0.5u
X10386 a_24660_6402# cap_series_gyn a_24452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X10387 vdd a_24652_55255# a_24564_55352# vdd pmos_6p0 w=1.22u l=1u
X10388 a_35292_3511# a_35204_3608# vss vss nmos_6p0 w=0.82u l=1u
X10389 vdd tune_series_gy[5] a_21540_11452# vdd pmos_6p0 w=1.2u l=0.5u
X10390 a_18940_50984# a_18852_51028# vss vss nmos_6p0 w=0.82u l=1u
X10391 a_25780_34264# cap_shunt_p a_27496_34264# vss nmos_6p0 w=0.82u l=0.6u
X10392 a_34396_25896# a_34308_25940# vss vss nmos_6p0 w=0.82u l=1u
X10393 a_32268_54120# a_32180_54164# vss vss nmos_6p0 w=0.82u l=1u
X10394 a_28692_32696# cap_shunt_p a_28484_32212# vdd pmos_6p0 w=1.2u l=0.5u
X10395 vdd a_34396_5512# a_34308_5556# vdd pmos_6p0 w=1.22u l=1u
X10396 a_7748_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10397 a_32464_44757# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X10398 a_31708_41143# a_31620_41240# vss vss nmos_6p0 w=0.82u l=1u
X10399 a_17828_31128# cap_shunt_n a_17620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X10400 vss tune_shunt[7] a_13460_35832# vss nmos_6p0 w=0.51u l=0.6u
X10401 a_32404_30268# cap_shunt_p a_32612_29922# vdd pmos_6p0 w=1.2u l=0.5u
X10402 vdd a_24652_52119# a_24564_52216# vdd pmos_6p0 w=1.22u l=1u
X10403 a_16708_42466# cap_shunt_n a_16500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X10404 a_9220_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10405 vdd a_23308_32168# a_23220_32212# vdd pmos_6p0 w=1.22u l=1u
X10406 a_25780_31128# cap_shunt_p a_27496_31128# vss nmos_6p0 w=0.82u l=0.6u
X10407 a_12580_19668# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10408 vdd tune_shunt[5] a_6084_50652# vdd pmos_6p0 w=1.2u l=0.5u
X10409 a_32612_31490# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X10410 a_11824_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X10411 a_30616_19668# cap_series_gygyn a_30640_20152# vss nmos_6p0 w=0.82u l=0.6u
X10412 vss tune_shunt[7] a_25780_27992# vss nmos_6p0 w=0.51u l=0.6u
X10413 a_11612_8692# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10414 a_3620_46324# cap_shunt_p a_3828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X10415 vss cap_shunt_n a_15120_36132# vss nmos_6p0 w=0.82u l=0.6u
X10416 a_25780_27992# cap_shunt_p a_25572_27508# vdd pmos_6p0 w=1.2u l=0.5u
X10417 a_36720_48438# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10418 a_26712_32696# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10419 a_29720_9884# cap_series_gyn a_30528_9476# vss nmos_6p0 w=0.82u l=0.6u
X10420 a_23464_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X10421 vss tune_shunt[6] a_10660_44034# vss nmos_6p0 w=0.51u l=0.6u
X10422 a_25572_38484# cap_shunt_p a_25780_38968# vdd pmos_6p0 w=1.2u l=0.5u
X10423 a_28484_38484# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10424 vdd tune_shunt[2] a_1716_3988# vdd pmos_6p0 w=1.2u l=0.5u
X10425 a_16500_20860# cap_shunt_p a_16708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X10426 vss tune_shunt[7] a_25780_24856# vss nmos_6p0 w=0.51u l=0.6u
X10427 vss tune_shunt[7] a_13460_23288# vss nmos_6p0 w=0.51u l=0.6u
X10428 a_23308_27464# a_23220_27508# vss vss nmos_6p0 w=0.82u l=1u
X10429 a_32604_3944# a_32516_3988# vss vss nmos_6p0 w=0.82u l=1u
X10430 a_20740_17016# cap_shunt_p a_21672_17016# vss nmos_6p0 w=0.82u l=0.6u
X10431 a_18424_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10432 a_11780_4472# cap_series_gyp a_13496_4472# vss nmos_6p0 w=0.82u l=0.6u
X10433 a_25572_35348# cap_shunt_p a_25780_35832# vdd pmos_6p0 w=1.2u l=0.5u
X10434 a_28484_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10435 vdd tune_shunt[5] a_32404_34972# vdd pmos_6p0 w=1.2u l=0.5u
X10436 vss tune_shunt[6] a_13796_42466# vss nmos_6p0 w=0.51u l=0.6u
X10437 a_2708_36194# cap_shunt_n a_2500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X10438 a_4828_54120# a_4740_54164# vss vss nmos_6p0 w=0.82u l=1u
X10439 a_21540_39676# cap_shunt_p a_21748_39330# vdd pmos_6p0 w=1.2u l=0.5u
X10440 a_20532_24372# cap_shunt_n a_20740_24856# vdd pmos_6p0 w=1.2u l=0.5u
X10441 a_1716_8316# cap_shunt_n a_1924_7970# vdd pmos_6p0 w=1.2u l=0.5u
X10442 a_16500_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10443 a_23308_24328# a_23220_24372# vss vss nmos_6p0 w=0.82u l=1u
X10444 a_6292_18946# cap_shunt_p a_7224_18884# vss nmos_6p0 w=0.82u l=0.6u
X10445 vss cap_series_gyn a_17024_7908# vss nmos_6p0 w=0.82u l=0.6u
X10446 a_22680_39268# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10447 a_18424_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10448 a_2500_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10449 a_19152_27992# cap_shunt_n a_17828_27992# vss nmos_6p0 w=0.82u l=0.6u
X10450 vdd tune_shunt[4] a_32404_31836# vdd pmos_6p0 w=1.2u l=0.5u
X10451 a_27228_17623# a_27140_17720# vss vss nmos_6p0 w=0.82u l=1u
X10452 a_2724_11828# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10453 vdd tune_shunt[5] a_3620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X10454 a_32404_38108# cap_shunt_p a_32612_37762# vdd pmos_6p0 w=1.2u l=0.5u
X10455 a_2708_33058# cap_shunt_p a_2500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X10456 a_6060_8215# a_5972_8312# vss vss nmos_6p0 w=0.82u l=1u
X10457 vdd tune_series_gy[5] a_28484_13396# vdd pmos_6p0 w=1.2u l=0.5u
X10458 a_20740_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10459 a_11200_51512# cap_shunt_n a_9876_51512# vss nmos_6p0 w=0.82u l=0.6u
X10460 a_16708_26786# cap_shunt_n a_16500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X10461 a_20532_21236# cap_shunt_p a_20740_21720# vdd pmos_6p0 w=1.2u l=0.5u
X10462 a_6292_15810# cap_shunt_p a_7224_15748# vss nmos_6p0 w=0.82u l=0.6u
X10463 vss tune_shunt[1] a_25780_4472# vss nmos_6p0 w=0.51u l=0.6u
X10464 a_17620_19668# cap_shunt_p a_17828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X10465 a_19152_24856# cap_shunt_n a_17828_24856# vss nmos_6p0 w=0.82u l=0.6u
X10466 vdd a_24316_45847# a_24228_45944# vdd pmos_6p0 w=1.22u l=1u
X10467 a_21748_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10468 vss cap_shunt_p a_11424_50244# vss nmos_6p0 w=0.82u l=0.6u
X10469 a_13460_34264# cap_shunt_n a_13252_33780# vdd pmos_6p0 w=1.2u l=0.5u
X10470 a_3380_17016# cap_shunt_p a_3172_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10471 a_1924_6040# cap_shunt_p a_1716_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10472 vdd tune_series_gy[1] a_6572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10473 a_2500_11452# cap_shunt_n a_2708_11106# vdd pmos_6p0 w=1.2u l=0.5u
X10474 a_28692_29560# cap_shunt_p a_28484_29076# vdd pmos_6p0 w=1.2u l=0.5u
X10475 a_21748_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10476 vdd a_24652_48983# a_24564_49080# vdd pmos_6p0 w=1.22u l=1u
X10477 a_13460_31128# cap_shunt_n a_13252_30644# vdd pmos_6p0 w=1.2u l=0.5u
X10478 vdd tune_series_gy[4] a_21540_5180# vdd pmos_6p0 w=1.2u l=0.5u
X10479 a_8120_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10480 a_14112_48376# cap_shunt_p a_12788_48376# vss nmos_6p0 w=0.82u l=0.6u
X10481 a_32268_47848# a_32180_47892# vss vss nmos_6p0 w=0.82u l=1u
X10482 vdd tune_shunt[6] a_7540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X10483 a_14372_44756# cap_shunt_p a_14580_45240# vdd pmos_6p0 w=1.2u l=0.5u
X10484 a_11984_37700# cap_shunt_n a_10660_37762# vss nmos_6p0 w=0.82u l=0.6u
X10485 a_7748_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10486 a_17828_24856# cap_shunt_n a_17620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X10487 vss tune_shunt[7] a_13460_29560# vss nmos_6p0 w=0.51u l=0.6u
X10488 vss cap_shunt_n a_4032_29860# vss nmos_6p0 w=0.82u l=0.6u
X10489 a_16708_36194# cap_shunt_n a_16500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X10490 a_14392_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10491 a_10136_51812# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10492 a_25984_7908# cap_series_gyp a_24660_7970# vss nmos_6p0 w=0.82u l=0.6u
X10493 a_34396_16488# a_34308_16532# vss vss nmos_6p0 w=0.82u l=1u
X10494 a_4312_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10495 a_31648_22020# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X10496 a_17828_21720# cap_shunt_p a_17620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X10497 vss tune_shunt[7] a_13460_26424# vss nmos_6p0 w=0.51u l=0.6u
X10498 vss cap_shunt_p a_11648_14180# vss nmos_6p0 w=0.82u l=0.6u
X10499 vss cap_shunt_p a_4032_26724# vss nmos_6p0 w=0.82u l=0.6u
X10500 vdd tune_shunt[7] a_17620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X10501 a_32156_55255# a_32068_55352# vss vss nmos_6p0 w=0.82u l=1u
X10502 vss cap_shunt_n a_9072_39268# vss nmos_6p0 w=0.82u l=0.6u
X10503 a_16708_33058# cap_shunt_n a_16500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X10504 vss cap_shunt_n a_15904_48676# vss nmos_6p0 w=0.82u l=0.6u
X10505 a_14392_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10506 a_28236_53687# a_28148_53784# vss vss nmos_6p0 w=0.82u l=1u
X10507 a_32732_46808# cap_shunt_gyn a_32464_46870# vss nmos_6p0 w=0.82u l=0.6u
X10508 vdd a_35180_30167# a_35092_30264# vdd pmos_6p0 w=1.22u l=1u
X10509 a_21748_23650# cap_shunt_p a_21540_23996# vdd pmos_6p0 w=1.2u l=0.5u
X10510 a_14580_46808# cap_shunt_p a_15512_46808# vss nmos_6p0 w=0.82u l=0.6u
X10511 a_18404_5180# cap_series_gyp a_18612_4834# vdd pmos_6p0 w=1.2u l=0.5u
X10512 vss tune_series_gy[4] a_25780_18584# vss nmos_6p0 w=0.51u l=0.6u
X10513 vdd tune_shunt[5] a_6644_53788# vdd pmos_6p0 w=1.2u l=0.5u
X10514 a_6760_7124# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X10515 vss cap_shunt_p a_11648_11044# vss nmos_6p0 w=0.82u l=0.6u
X10516 a_18424_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10517 a_26712_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10518 a_9108_50652# cap_shunt_p a_9316_50306# vdd pmos_6p0 w=1.2u l=0.5u
X10519 a_19936_45240# cap_shunt_p a_17828_45240# vss nmos_6p0 w=0.82u l=0.6u
X10520 a_28124_39575# a_28036_39672# vss vss nmos_6p0 w=0.82u l=1u
X10521 a_25572_29076# cap_shunt_p a_25780_29560# vdd pmos_6p0 w=1.2u l=0.5u
X10522 a_9540_9538# cap_shunt_p a_9332_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10523 a_15804_52119# a_15716_52216# vss vss nmos_6p0 w=0.82u l=1u
X10524 a_3036_43144# a_2948_43188# vss vss nmos_6p0 w=0.82u l=1u
X10525 vdd a_34844_36872# a_34756_36916# vdd pmos_6p0 w=1.22u l=1u
X10526 a_28484_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10527 a_18612_7970# cap_series_gyp a_19544_7908# vss nmos_6p0 w=0.82u l=0.6u
X10528 vss tune_shunt[7] a_9876_17016# vss nmos_6p0 w=0.51u l=0.6u
X10529 a_28236_50551# a_28148_50648# vss vss nmos_6p0 w=0.82u l=1u
X10530 a_3828_48376# cap_shunt_p a_3620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X10531 vss tune_shunt[7] a_13796_36194# vss nmos_6p0 w=0.51u l=0.6u
X10532 vss tune_series_gy[5] a_25780_15448# vss nmos_6p0 w=0.51u l=0.6u
X10533 a_6532_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10534 a_16500_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10535 a_29720_9884# cap_series_gyn a_29532_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10536 a_23308_18056# a_23220_18100# vss vss nmos_6p0 w=0.82u l=1u
X10537 a_9668_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10538 a_18424_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10539 vdd tune_shunt[7] a_2500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X10540 a_19936_42104# cap_shunt_n a_17828_42104# vss nmos_6p0 w=0.82u l=0.6u
X10541 a_20740_42104# cap_shunt_p a_20532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X10542 a_3036_40008# a_2948_40052# vss vss nmos_6p0 w=0.82u l=1u
X10543 vdd tune_shunt[4] a_32404_25564# vdd pmos_6p0 w=1.2u l=0.5u
X10544 a_14484_10260# cap_series_gyn a_14692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X10545 vdd a_2140_14920# a_2052_14964# vdd pmos_6p0 w=1.22u l=1u
X10546 a_3828_45240# cap_shunt_p a_3620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X10547 a_17828_37400# cap_shunt_n a_17620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X10548 vss tune_shunt[7] a_13796_33058# vss nmos_6p0 w=0.51u l=0.6u
X10549 a_2708_26786# cap_shunt_p a_2500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X10550 vss cap_shunt_n a_11872_37400# vss nmos_6p0 w=0.82u l=0.6u
X10551 a_10660_4834# cap_series_gyp a_10452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X10552 a_28684_54120# a_28596_54164# vss vss nmos_6p0 w=0.82u l=1u
X10553 a_32404_30268# cap_shunt_p a_32612_29922# vdd pmos_6p0 w=1.2u l=0.5u
X10554 a_10660_4834# cap_series_gyp a_12376_4772# vss nmos_6p0 w=0.82u l=0.6u
X10555 a_23308_14920# a_23220_14964# vss vss nmos_6p0 w=0.82u l=1u
X10556 a_8848_48376# cap_shunt_p a_6740_48376# vss nmos_6p0 w=0.82u l=0.6u
X10557 a_16708_45602# cap_shunt_p a_17640_45540# vss nmos_6p0 w=0.82u l=0.6u
X10558 a_25780_4472# cap_shunt_p a_25572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X10559 a_19152_18584# cap_shunt_p a_17828_18584# vss nmos_6p0 w=0.82u l=0.6u
X10560 vss cap_series_gygyp a_36296_23288# vss nmos_6p0 w=0.82u l=0.6u
X10561 vdd a_2140_11784# a_2052_11828# vdd pmos_6p0 w=1.22u l=1u
X10562 a_7748_44034# cap_shunt_p a_7540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X10563 a_11460_40052# cap_shunt_n a_11668_40536# vdd pmos_6p0 w=1.2u l=0.5u
X10564 a_25572_38484# cap_shunt_p a_25780_38968# vdd pmos_6p0 w=1.2u l=0.5u
X10565 a_12376_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10566 a_17620_14964# cap_shunt_p a_17828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X10567 a_3828_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10568 vdd a_28348_55688# a_28260_55732# vdd pmos_6p0 w=1.22u l=1u
X10569 a_24452_44380# cap_shunt_p a_24660_44034# vdd pmos_6p0 w=1.2u l=0.5u
X10570 a_16708_42466# cap_shunt_n a_17640_42404# vss nmos_6p0 w=0.82u l=0.6u
X10571 a_21748_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10572 a_19152_15448# cap_shunt_p a_17828_15448# vss nmos_6p0 w=0.82u l=0.6u
X10573 a_13460_24856# cap_shunt_n a_13252_24372# vdd pmos_6p0 w=1.2u l=0.5u
X10574 a_31624_22428# cap_series_gygyn a_32432_22020# vss nmos_6p0 w=0.82u l=0.6u
X10575 a_7748_40898# cap_shunt_n a_7540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X10576 vss tune_series_gy[4] a_14692_7608# vss nmos_6p0 w=0.51u l=0.6u
X10577 a_22972_50984# a_22884_51028# vss vss nmos_6p0 w=0.82u l=1u
X10578 vdd tune_shunt[6] a_7540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X10579 a_1692_36872# a_1604_36916# vss vss nmos_6p0 w=0.82u l=1u
X10580 a_25572_35348# cap_shunt_p a_25780_35832# vdd pmos_6p0 w=1.2u l=0.5u
X10581 a_17820_3511# a_17732_3608# vss vss nmos_6p0 w=0.82u l=1u
X10582 a_24452_41244# cap_shunt_n a_24660_40898# vdd pmos_6p0 w=1.2u l=0.5u
X10583 a_21748_25218# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10584 vss cap_shunt_n a_19936_32696# vss nmos_6p0 w=0.82u l=0.6u
X10585 a_13460_21720# cap_shunt_n a_13252_21236# vdd pmos_6p0 w=1.2u l=0.5u
X10586 a_30136_9476# cap_series_gyn a_29720_9884# vss nmos_6p0 w=0.82u l=0.6u
X10587 a_6084_17724# cap_shunt_p a_6292_17378# vdd pmos_6p0 w=1.2u l=0.5u
X10588 a_9876_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10589 vss tune_shunt[7] a_6516_20514# vss nmos_6p0 w=0.51u l=0.6u
X10590 a_33732_32696# cap_shunt_n a_34664_32696# vss nmos_6p0 w=0.82u l=0.6u
X10591 vdd a_21180_52552# a_21092_52596# vdd pmos_6p0 w=1.22u l=1u
X10592 a_2724_11828# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10593 a_25780_13880# cap_series_gyn a_25572_13396# vdd pmos_6p0 w=1.2u l=0.5u
X10594 a_32156_48983# a_32068_49080# vss vss nmos_6p0 w=0.82u l=1u
X10595 a_3828_37400# cap_shunt_n a_5544_37400# vss nmos_6p0 w=0.82u l=0.6u
X10596 a_16708_26786# cap_shunt_n a_16500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X10597 vdd a_37420_38007# a_37332_38104# vdd pmos_6p0 w=1.22u l=1u
X10598 vss cap_shunt_n a_5040_10744# vss nmos_6p0 w=0.82u l=0.6u
X10599 a_13796_23650# cap_shunt_n a_13588_23996# vdd pmos_6p0 w=1.2u l=0.5u
X10600 a_20664_13880# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X10601 a_13460_34264# cap_shunt_n a_13252_33780# vdd pmos_6p0 w=1.2u l=0.5u
X10602 a_6292_15810# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10603 a_3380_17016# cap_shunt_p a_3172_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10604 a_24452_17724# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10605 vss tune_series_gy[3] a_24660_6402# vss nmos_6p0 w=0.51u l=0.6u
X10606 vss cap_shunt_p a_4032_17316# vss nmos_6p0 w=0.82u l=0.6u
X10607 a_37420_19191# a_37332_19288# vss vss nmos_6p0 w=0.82u l=1u
X10608 vss cap_shunt_n a_15904_39268# vss nmos_6p0 w=0.82u l=0.6u
X10609 a_19524_8692# cap_series_gyp a_19732_9176# vdd pmos_6p0 w=1.2u l=0.5u
X10610 a_21748_14242# cap_series_gyn a_21540_14588# vdd pmos_6p0 w=1.2u l=0.5u
X10611 a_6084_18100# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10612 a_10548_32696# cap_shunt_n a_12264_32696# vss nmos_6p0 w=0.82u l=0.6u
X10613 vdd a_18044_3944# a_17956_3988# vdd pmos_6p0 w=1.22u l=1u
X10614 a_20664_10744# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X10615 a_13460_31128# cap_shunt_n a_13252_30644# vdd pmos_6p0 w=1.2u l=0.5u
X10616 a_3036_33736# a_2948_33780# vss vss nmos_6p0 w=0.82u l=1u
X10617 a_37420_16055# a_37332_16152# vss vss nmos_6p0 w=0.82u l=1u
X10618 a_3828_38968# cap_shunt_n a_3620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X10619 vdd a_10988_40008# a_10900_40052# vdd pmos_6p0 w=1.22u l=1u
X10620 vdd a_23756_41576# a_23668_41620# vdd pmos_6p0 w=1.22u l=1u
X10621 a_28684_47848# a_28596_47892# vss vss nmos_6p0 w=0.82u l=1u
X10622 vss cap_shunt_gyn a_35532_47108# vss nmos_6p0 w=0.82u l=0.6u
X10623 vdd a_36188_40008# a_36100_40052# vdd pmos_6p0 w=1.22u l=1u
X10624 a_6532_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10625 a_14012_6647# a_13924_6744# vss vss nmos_6p0 w=0.82u l=1u
X10626 vdd a_20172_45847# a_20084_45944# vdd pmos_6p0 w=1.22u l=1u
X10627 a_20740_32696# cap_shunt_n a_20532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X10628 a_3036_30600# a_2948_30644# vss vss nmos_6p0 w=0.82u l=1u
X10629 vdd tune_series_gy[3] a_32444_11452# vdd pmos_6p0 w=1.2u l=0.5u
X10630 a_3828_35832# cap_shunt_n a_3620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X10631 a_17828_27992# cap_shunt_n a_17620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X10632 a_1924_6040# cap_shunt_p a_1716_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10633 vdd a_20172_42711# a_20084_42808# vdd pmos_6p0 w=1.22u l=1u
X10634 a_10640_22020# cap_shunt_p a_9316_22082# vss nmos_6p0 w=0.82u l=0.6u
X10635 a_7580_8316# cap_series_gyn a_7768_8316# vdd pmos_6p0 w=1.2u l=0.5u
X10636 a_16500_44380# cap_shunt_p a_16708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X10637 a_16708_36194# cap_shunt_n a_17640_36132# vss nmos_6p0 w=0.82u l=0.6u
X10638 a_27676_30167# a_27588_30264# vss vss nmos_6p0 w=0.82u l=1u
X10639 a_2724_10260# cap_shunt_n a_2932_10744# vdd pmos_6p0 w=1.2u l=0.5u
X10640 a_25572_29076# cap_shunt_p a_25780_29560# vdd pmos_6p0 w=1.2u l=0.5u
X10641 a_12376_23588# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10642 a_35880_3988# cap_series_gygyp a_35904_4472# vss nmos_6p0 w=0.82u l=0.6u
X10643 a_9108_50652# cap_shunt_p a_9316_50306# vdd pmos_6p0 w=1.2u l=0.5u
X10644 a_3828_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10645 vdd a_33052_3511# a_32964_3608# vdd pmos_6p0 w=1.22u l=1u
X10646 a_12580_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10647 a_9428_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10648 a_16500_41244# cap_shunt_n a_16708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X10649 a_35292_53687# a_35204_53784# vss vss nmos_6p0 w=0.82u l=1u
X10650 a_27676_27031# a_27588_27128# vss vss nmos_6p0 w=0.82u l=1u
X10651 a_25548_55255# a_25460_55352# vss vss nmos_6p0 w=0.82u l=1u
X10652 vss tune_shunt[6] a_11668_45240# vss nmos_6p0 w=0.51u l=0.6u
X10653 vdd a_33500_24328# a_33412_24372# vdd pmos_6p0 w=1.22u l=1u
X10654 vdd tune_shunt[7] a_2500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X10655 a_28484_33780# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10656 a_22436_7124# cap_series_gyp a_22644_7608# vdd pmos_6p0 w=1.2u l=0.5u
X10657 a_34516_4834# tune_series_gygy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X10658 vdd tune_series_gy[3] a_14484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X10659 a_20740_42104# cap_shunt_p a_20532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X10660 vdd a_28572_30167# a_28484_30264# vdd pmos_6p0 w=1.22u l=1u
X10661 a_4032_6340# cap_shunt_n a_1924_6402# vss nmos_6p0 w=0.82u l=0.6u
X10662 a_12580_11828# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10663 a_25780_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10664 vdd a_32380_43144# a_32292_43188# vdd pmos_6p0 w=1.22u l=1u
X10665 a_15624_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X10666 a_22860_52119# a_22772_52216# vss vss nmos_6p0 w=0.82u l=1u
X10667 a_29700_34626# cap_shunt_p a_31416_34564# vss nmos_6p0 w=0.82u l=0.6u
X10668 a_35692_13396# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10669 a_35292_50551# a_35204_50648# vss vss nmos_6p0 w=0.82u l=1u
X10670 vss cap_shunt_n a_19936_23288# vss nmos_6p0 w=0.82u l=0.6u
X10671 a_9876_12312# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10672 vss tune_shunt[6] a_11668_42104# vss nmos_6p0 w=0.51u l=0.6u
X10673 a_9668_19668# cap_shunt_p a_9876_20152# vdd pmos_6p0 w=1.2u l=0.5u
X10674 vdd a_33500_21192# a_33412_21236# vdd pmos_6p0 w=1.22u l=1u
X10675 a_28484_30644# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10676 a_4032_3204# cap_shunt_n a_1924_3266# vss nmos_6p0 w=0.82u l=0.6u
X10677 a_25780_10744# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X10678 a_7748_44034# cap_shunt_p a_7540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X10679 a_29700_31490# cap_shunt_p a_31416_31428# vss nmos_6p0 w=0.82u l=0.6u
X10680 a_25236_3612# cap_shunt_p a_25444_3266# vdd pmos_6p0 w=1.2u l=0.5u
X10681 a_6084_52220# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10682 a_25572_38484# cap_shunt_p a_25780_38968# vdd pmos_6p0 w=1.2u l=0.5u
X10683 a_34720_32996# cap_shunt_n a_32612_33058# vss nmos_6p0 w=0.82u l=0.6u
X10684 a_18404_8316# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10685 vdd a_20620_44279# a_20532_44376# vdd pmos_6p0 w=1.22u l=1u
X10686 a_13796_14242# cap_shunt_p a_13588_14588# vdd pmos_6p0 w=1.2u l=0.5u
X10687 vdd tune_shunt[7] a_3620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X10688 a_13460_24856# cap_shunt_n a_13252_24372# vdd pmos_6p0 w=1.2u l=0.5u
X10689 a_7748_40898# cap_shunt_n a_7540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X10690 a_11668_45240# cap_shunt_n a_12600_45240# vss nmos_6p0 w=0.82u l=0.6u
X10691 a_25780_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10692 a_14468_3266# cap_series_gyn a_14260_3612# vdd pmos_6p0 w=1.2u l=0.5u
X10693 a_20532_44756# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10694 a_25572_35348# cap_shunt_p a_25780_35832# vdd pmos_6p0 w=1.2u l=0.5u
X10695 vdd tune_shunt[3] a_5636_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10696 vss tune_shunt[4] a_33732_35832# vss nmos_6p0 w=0.51u l=0.6u
X10697 a_9332_11452# cap_shunt_p a_9540_11106# vdd pmos_6p0 w=1.2u l=0.5u
X10698 vss cap_shunt_n a_22848_43672# vss nmos_6p0 w=0.82u l=0.6u
X10699 a_10548_23288# cap_shunt_n a_12264_23288# vss nmos_6p0 w=0.82u l=0.6u
X10700 vss cap_shunt_n a_5040_9176# vss nmos_6p0 w=0.82u l=0.6u
X10701 a_13588_45948# cap_shunt_p a_13796_45602# vdd pmos_6p0 w=1.2u l=0.5u
X10702 a_13460_21720# cap_shunt_n a_13252_21236# vdd pmos_6p0 w=1.2u l=0.5u
X10703 vdd a_20172_39575# a_20084_39672# vdd pmos_6p0 w=1.22u l=1u
X10704 a_11668_42104# cap_shunt_n a_12600_42104# vss nmos_6p0 w=0.82u l=0.6u
X10705 a_34536_6748# tune_series_gygy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X10706 a_6084_17724# cap_shunt_p a_6292_17378# vdd pmos_6p0 w=1.2u l=0.5u
X10707 a_28692_9176# cap_series_gyn a_28484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X10708 a_38092_30600# a_38004_30644# vss vss nmos_6p0 w=0.82u l=1u
X10709 a_3828_29560# cap_shunt_n a_3620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X10710 a_4828_53687# a_4740_53784# vss vss nmos_6p0 w=0.82u l=1u
X10711 a_2500_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10712 vdd a_23756_32168# a_23668_32212# vdd pmos_6p0 w=1.22u l=1u
X10713 a_18612_9538# cap_series_gyp a_18404_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10714 a_25780_13880# cap_series_gyn a_25572_13396# vdd pmos_6p0 w=1.2u l=0.5u
X10715 a_16500_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10716 a_25780_6040# cap_series_gyp a_27496_6040# vss nmos_6p0 w=0.82u l=0.6u
X10717 a_14728_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10718 vdd tune_shunt[6] a_11460_43188# vdd pmos_6p0 w=1.2u l=0.5u
X10719 vss cap_shunt_p a_22848_40536# vss nmos_6p0 w=0.82u l=0.6u
X10720 a_4424_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10721 a_17596_52552# a_17508_52596# vss vss nmos_6p0 w=0.82u l=1u
X10722 vdd a_20172_36439# a_20084_36536# vdd pmos_6p0 w=1.22u l=1u
X10723 vss tune_shunt[7] a_29700_29922# vss nmos_6p0 w=0.51u l=0.6u
X10724 a_13796_23650# cap_shunt_n a_13588_23996# vdd pmos_6p0 w=1.2u l=0.5u
X10725 a_28692_6040# cap_shunt_n a_28484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10726 vdd a_33948_52552# a_33860_52596# vdd pmos_6p0 w=1.22u l=1u
X10727 a_2500_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10728 a_18612_6402# cap_series_gyn a_18404_6748# vdd pmos_6p0 w=1.2u l=0.5u
X10729 a_21540_17724# cap_shunt_p a_21748_17378# vdd pmos_6p0 w=1.2u l=0.5u
X10730 a_36296_37400# cap_series_gygyp a_35880_36916# vss nmos_6p0 w=0.82u l=0.6u
X10731 vdd tune_series_gy[4] a_15492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X10732 a_14728_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10733 a_5152_13880# cap_shunt_n a_3828_13880# vss nmos_6p0 w=0.82u l=0.6u
X10734 a_23756_27464# a_23668_27508# vss vss nmos_6p0 w=0.82u l=1u
X10735 vdd tune_series_gy[2] a_11572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10736 a_6084_18100# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10737 vdd a_33948_7080# a_33860_7124# vdd pmos_6p0 w=1.22u l=1u
X10738 a_2708_12674# cap_shunt_n a_2500_13020# vdd pmos_6p0 w=1.2u l=0.5u
X10739 a_25548_48983# a_25460_49080# vss vss nmos_6p0 w=0.82u l=1u
X10740 a_32404_38108# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10741 vdd a_2140_31735# a_2052_31832# vdd pmos_6p0 w=1.22u l=1u
X10742 vss tune_shunt[7] a_13796_12674# vss nmos_6p0 w=0.51u l=0.6u
X10743 a_23756_24328# a_23668_24372# vss vss nmos_6p0 w=0.82u l=1u
X10744 a_29700_28354# cap_shunt_p a_31416_28292# vss nmos_6p0 w=0.82u l=0.6u
X10745 vss tune_series_gy[4] a_22644_7608# vss nmos_6p0 w=0.51u l=0.6u
X10746 a_32716_5079# a_32628_5176# vss vss nmos_6p0 w=0.82u l=1u
X10747 a_15904_12612# cap_shunt_p a_13796_12674# vss nmos_6p0 w=0.82u l=0.6u
X10748 a_34516_12674# cap_series_gygyp a_34308_13020# vdd pmos_6p0 w=1.2u l=0.5u
X10749 a_27676_17623# a_27588_17720# vss vss nmos_6p0 w=0.82u l=1u
X10750 a_2588_21192# a_2500_21236# vss vss nmos_6p0 w=0.82u l=1u
X10751 a_5844_11106# cap_shunt_n a_5636_11452# vdd pmos_6p0 w=1.2u l=0.5u
X10752 a_36076_33303# a_35988_33400# vss vss nmos_6p0 w=0.82u l=1u
X10753 a_20740_32696# cap_shunt_n a_20532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X10754 a_28484_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10755 vss tune_shunt[7] a_2708_29922# vss nmos_6p0 w=0.51u l=0.6u
X10756 a_29700_25218# cap_shunt_p a_31416_25156# vss nmos_6p0 w=0.82u l=0.6u
X10757 a_4816_18884# cap_shunt_p a_2708_18946# vss nmos_6p0 w=0.82u l=0.6u
X10758 vdd a_24764_45847# a_24676_45944# vdd pmos_6p0 w=1.22u l=1u
X10759 a_19524_8692# cap_series_gyp a_19732_9176# vdd pmos_6p0 w=1.2u l=0.5u
X10760 a_15720_11452# cap_series_gyp a_15744_11044# vss nmos_6p0 w=0.82u l=0.6u
X10761 vdd a_3036_36872# a_2948_36916# vdd pmos_6p0 w=1.22u l=1u
X10762 a_13460_37400# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10763 a_16500_44380# cap_shunt_p a_16708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X10764 a_21748_4834# cap_series_gyp a_21540_5180# vdd pmos_6p0 w=1.2u l=0.5u
X10765 a_13796_33058# cap_shunt_n a_14728_32996# vss nmos_6p0 w=0.82u l=0.6u
X10766 a_12580_18100# cap_shunt_p a_12788_18584# vdd pmos_6p0 w=1.2u l=0.5u
X10767 a_20532_40052# cap_shunt_p a_20740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X10768 a_4816_15748# cap_shunt_p a_2708_15810# vss nmos_6p0 w=0.82u l=0.6u
X10769 a_25780_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10770 a_20532_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10771 vss tune_shunt[7] a_33732_29560# vss nmos_6p0 w=0.51u l=0.6u
X10772 a_25572_29076# cap_shunt_p a_25780_29560# vdd pmos_6p0 w=1.2u l=0.5u
X10773 a_35692_7124# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10774 a_13796_45602# cap_shunt_p a_15512_45540# vss nmos_6p0 w=0.82u l=0.6u
X10775 vdd a_37420_55688# a_37332_55732# vdd pmos_6p0 w=1.22u l=1u
X10776 a_16500_41244# cap_shunt_n a_16708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X10777 a_23856_45540# cap_shunt_p a_21748_45602# vss nmos_6p0 w=0.82u l=0.6u
X10778 a_13588_39676# cap_shunt_n a_13796_39330# vdd pmos_6p0 w=1.2u l=0.5u
X10779 a_9428_17378# cap_shunt_p a_9220_17724# vdd pmos_6p0 w=1.2u l=0.5u
X10780 a_13796_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X10781 a_3620_41620# cap_shunt_p a_3828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X10782 a_3380_51512# cap_shunt_n a_3172_51028# vdd pmos_6p0 w=1.2u l=0.5u
X10783 a_25780_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10784 a_20532_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10785 a_22064_21720# cap_shunt_p a_20740_21720# vss nmos_6p0 w=0.82u l=0.6u
X10786 a_13796_42466# cap_shunt_n a_15512_42404# vss nmos_6p0 w=0.82u l=0.6u
X10787 vss tune_shunt[2] a_1924_4472# vss nmos_6p0 w=0.51u l=0.6u
X10788 a_10340_36916# cap_shunt_n a_10548_37400# vdd pmos_6p0 w=1.2u l=0.5u
X10789 vdd a_21628_54120# a_21540_54164# vdd pmos_6p0 w=1.22u l=1u
X10790 a_36160_43189# tune_shunt_gy[3] vdd vdd pmos_6p0 w=1.215u l=0.5u
X10791 a_23856_42404# cap_shunt_n a_21748_42466# vss nmos_6p0 w=0.82u l=0.6u
X10792 vss cap_shunt_n a_22848_34264# vss nmos_6p0 w=0.82u l=0.6u
X10793 a_4424_14180# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10794 a_3828_26424# cap_shunt_p a_3620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X10795 a_12332_54120# a_12244_54164# vss vss nmos_6p0 w=0.82u l=1u
X10796 a_2708_48738# cap_shunt_p a_4424_48676# vss nmos_6p0 w=0.82u l=0.6u
X10797 a_2500_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10798 a_28684_53687# a_28596_53784# vss vss nmos_6p0 w=0.82u l=1u
X10799 a_6084_52220# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10800 vdd a_21628_50984# a_21540_51028# vdd pmos_6p0 w=1.22u l=1u
X10801 a_14728_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10802 vss cap_shunt_n a_22848_31128# vss nmos_6p0 w=0.82u l=0.6u
X10803 a_4424_11044# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10804 vdd a_20172_27031# a_20084_27128# vdd pmos_6p0 w=1.22u l=1u
X10805 vdd a_27340_47848# a_27252_47892# vdd pmos_6p0 w=1.22u l=1u
X10806 a_33524_27508# cap_shunt_p a_33732_27992# vdd pmos_6p0 w=1.2u l=0.5u
X10807 a_3828_23288# cap_shunt_p a_3620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X10808 vdd tune_series_gy[3] a_29532_9884# vdd pmos_6p0 w=1.2u l=0.5u
X10809 a_13796_14242# cap_shunt_p a_13588_14588# vdd pmos_6p0 w=1.2u l=0.5u
X10810 vss cap_shunt_p a_4704_18584# vss nmos_6p0 w=0.82u l=0.6u
X10811 a_8456_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10812 a_28572_39575# a_28484_39672# vss vss nmos_6p0 w=0.82u l=1u
X10813 a_24660_6402# cap_series_gyn a_26376_6340# vss nmos_6p0 w=0.82u l=0.6u
X10814 a_2500_22428# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10815 a_28684_50551# a_28596_50648# vss vss nmos_6p0 w=0.82u l=1u
X10816 vdd a_2140_25463# a_2052_25560# vdd pmos_6p0 w=1.22u l=1u
X10817 a_12108_14487# a_12020_14584# vss vss nmos_6p0 w=0.82u l=1u
X10818 vss cap_shunt_n a_14784_32696# vss nmos_6p0 w=0.82u l=0.6u
X10819 a_11984_13880# cap_shunt_p a_9876_13880# vss nmos_6p0 w=0.82u l=0.6u
X10820 a_23756_18056# a_23668_18100# vss vss nmos_6p0 w=0.82u l=1u
X10821 vdd a_27340_44712# a_27252_44756# vdd pmos_6p0 w=1.22u l=1u
X10822 a_8456_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10823 a_25444_3266# cap_shunt_p a_26376_3204# vss nmos_6p0 w=0.82u l=0.6u
X10824 vdd a_2140_22327# a_2052_22424# vdd pmos_6p0 w=1.22u l=1u
X10825 vdd a_19388_53687# a_19300_53784# vdd pmos_6p0 w=1.22u l=1u
X10826 a_12108_11351# a_12020_11448# vss vss nmos_6p0 w=0.82u l=1u
X10827 vss tune_shunt[5] a_6292_49944# vss nmos_6p0 w=0.51u l=0.6u
X10828 a_17024_4772# cap_series_gyn a_15700_4834# vss nmos_6p0 w=0.82u l=0.6u
X10829 a_14484_8692# cap_series_gyn a_14692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X10830 vdd tune_shunt[5] a_16500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X10831 vdd tune_shunt[7] a_6196_22428# vdd pmos_6p0 w=1.2u l=0.5u
X10832 a_11984_10744# cap_shunt_p a_9876_10744# vss nmos_6p0 w=0.82u l=0.6u
X10833 a_23756_14920# a_23668_14964# vss vss nmos_6p0 w=0.82u l=1u
X10834 vdd tune_shunt[6] a_11460_43188# vdd pmos_6p0 w=1.2u l=0.5u
X10835 a_2856_7908# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10836 a_6740_21720# cap_shunt_p a_8456_21720# vss nmos_6p0 w=0.82u l=0.6u
X10837 vss tune_shunt[6] a_6740_46808# vss nmos_6p0 w=0.51u l=0.6u
X10838 a_14484_5556# cap_series_gyn a_14692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X10839 a_17828_26424# cap_shunt_n a_17620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X10840 vss tune_shunt[3] a_5844_9176# vss nmos_6p0 w=0.51u l=0.6u
X10841 a_35880_19668# cap_series_gygyp a_35692_19668# vdd pmos_6p0 w=1.2u l=0.5u
X10842 a_21540_17724# cap_shunt_p a_21748_17378# vdd pmos_6p0 w=1.2u l=0.5u
X10843 a_11032_50244# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10844 a_9464_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10845 vdd a_3036_27464# a_2948_27508# vdd pmos_6p0 w=1.22u l=1u
X10846 vdd a_37420_49416# a_37332_49460# vdd pmos_6p0 w=1.22u l=1u
X10847 a_5844_10744# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X10848 a_3172_18100# cap_shunt_p a_3380_18584# vdd pmos_6p0 w=1.2u l=0.5u
X10849 vdd a_33500_41143# a_33412_41240# vdd pmos_6p0 w=1.22u l=1u
X10850 a_17828_23288# cap_shunt_n a_17620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X10851 a_2708_12674# cap_shunt_n a_2500_13020# vdd pmos_6p0 w=1.2u l=0.5u
X10852 a_19724_20759# a_19636_20856# vss vss nmos_6p0 w=0.82u l=1u
X10853 a_13796_36194# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10854 a_13796_23650# cap_shunt_n a_14728_23588# vss nmos_6p0 w=0.82u l=0.6u
X10855 a_23532_47848# a_23444_47892# vss vss nmos_6p0 w=0.82u l=1u
X10856 a_20532_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10857 a_6532_25940# cap_shunt_n a_6740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X10858 a_13252_32212# cap_shunt_n a_13460_32696# vdd pmos_6p0 w=1.2u l=0.5u
X10859 vdd a_37420_46280# a_37332_46324# vdd pmos_6p0 w=1.22u l=1u
X10860 a_9464_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10861 a_13796_36194# cap_shunt_n a_15512_36132# vss nmos_6p0 w=0.82u l=0.6u
X10862 a_13588_13020# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10863 a_30364_20759# a_30276_20856# vss vss nmos_6p0 w=0.82u l=1u
X10864 a_23856_36132# cap_shunt_n a_21748_36194# vss nmos_6p0 w=0.82u l=0.6u
X10865 a_35692_25940# cap_series_gygyp a_35880_25940# vdd pmos_6p0 w=1.2u l=0.5u
X10866 vdd a_32268_23895# a_32180_23992# vdd pmos_6p0 w=1.22u l=1u
X10867 a_14580_46808# cap_shunt_p a_14372_46324# vdd pmos_6p0 w=1.2u l=0.5u
X10868 a_3620_32212# cap_shunt_p a_3828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X10869 a_34516_12674# cap_series_gygyp a_34308_13020# vdd pmos_6p0 w=1.2u l=0.5u
X10870 a_13796_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10871 vss tune_series_gy[0] a_28692_4472# vss nmos_6p0 w=0.51u l=0.6u
X10872 a_22680_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X10873 vdd a_29468_55255# a_29380_55352# vdd pmos_6p0 w=1.22u l=1u
X10874 a_12264_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10875 a_3640_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10876 a_7960_4472# cap_series_gyp a_6760_3988# vss nmos_6p0 w=0.82u l=0.6u
X10877 a_5844_11106# cap_shunt_n a_5636_11452# vdd pmos_6p0 w=1.2u l=0.5u
X10878 a_25780_17016# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10879 a_33920_45302# cap_shunt_gyn a_33920_44757# vdd pmos_6p0 w=1.215u l=0.5u
X10880 a_6532_22804# cap_shunt_p a_6740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X10881 vss cap_shunt_n a_33936_34564# vss nmos_6p0 w=0.82u l=0.6u
X10882 vdd a_2588_53687# a_2500_53784# vdd pmos_6p0 w=1.22u l=1u
X10883 a_2500_19292# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10884 a_13588_34972# cap_shunt_n a_13796_34626# vdd pmos_6p0 w=1.2u l=0.5u
X10885 a_33732_32696# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X10886 a_10340_27508# cap_shunt_n a_10548_27992# vdd pmos_6p0 w=1.2u l=0.5u
X10887 a_35692_22804# cap_series_gygyp a_35880_22804# vdd pmos_6p0 w=1.2u l=0.5u
X10888 vdd tune_shunt[7] a_10452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X10889 a_11780_4472# cap_series_gyp a_12712_4472# vss nmos_6p0 w=0.82u l=0.6u
X10890 vss cap_shunt_p a_7168_9476# vss nmos_6p0 w=0.82u l=0.6u
X10891 vdd a_29468_52119# a_29380_52216# vdd pmos_6p0 w=1.22u l=1u
X10892 a_4312_51512# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10893 a_34396_50984# a_34308_51028# vss vss nmos_6p0 w=0.82u l=1u
X10894 a_12580_47892# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10895 a_3640_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10896 vdd tune_shunt[6] a_6532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X10897 vss cap_shunt_n a_33936_31428# vss nmos_6p0 w=0.82u l=0.6u
X10898 a_2708_39330# cap_shunt_n a_4424_39268# vss nmos_6p0 w=0.82u l=0.6u
X10899 a_2500_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10900 a_20532_40052# cap_shunt_p a_20740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X10901 a_13588_31836# cap_shunt_n a_13796_31490# vdd pmos_6p0 w=1.2u l=0.5u
X10902 a_3620_43188# cap_shunt_p a_3828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X10903 vss tune_shunt[3] a_2708_9538# vss nmos_6p0 w=0.51u l=0.6u
X10904 a_9668_14964# cap_shunt_p a_9876_15448# vdd pmos_6p0 w=1.2u l=0.5u
X10905 vss cap_shunt_n a_18032_47108# vss nmos_6p0 w=0.82u l=0.6u
X10906 vss tune_shunt[7] a_17828_37400# vss nmos_6p0 w=0.51u l=0.6u
X10907 vdd tune_shunt[7] a_10452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X10908 vss cap_series_gyn a_23856_12612# vss nmos_6p0 w=0.82u l=0.6u
X10909 a_9668_14964# cap_shunt_p a_9876_15448# vdd pmos_6p0 w=1.2u l=0.5u
X10910 vss tune_series_gy[4] a_24660_18946# vss nmos_6p0 w=0.51u l=0.6u
X10911 a_19500_50551# a_19412_50648# vss vss nmos_6p0 w=0.82u l=1u
X10912 a_18404_3988# cap_series_gyp a_18612_4472# vdd pmos_6p0 w=1.2u l=0.5u
X10913 a_9428_17378# cap_shunt_p a_9220_17724# vdd pmos_6p0 w=1.2u l=0.5u
X10914 a_24660_29922# cap_shunt_n a_26376_29860# vss nmos_6p0 w=0.82u l=0.6u
X10915 vdd a_13564_9783# a_13476_9880# vdd pmos_6p0 w=1.22u l=1u
X10916 a_20740_45240# cap_shunt_n a_21672_45240# vss nmos_6p0 w=0.82u l=0.6u
X10917 vdd a_2140_16055# a_2052_16152# vdd pmos_6p0 w=1.22u l=1u
X10918 a_25572_33780# cap_shunt_p a_25780_34264# vdd pmos_6p0 w=1.2u l=0.5u
X10919 a_2708_22082# cap_shunt_p a_3640_22020# vss nmos_6p0 w=0.82u l=0.6u
X10920 a_9668_11828# cap_shunt_p a_9876_12312# vdd pmos_6p0 w=1.2u l=0.5u
X10921 vss tune_shunt[5] a_9876_51512# vss nmos_6p0 w=0.51u l=0.6u
X10922 vss cap_shunt_n a_14784_23288# vss nmos_6p0 w=0.82u l=0.6u
X10923 a_9668_11828# cap_shunt_p a_9876_12312# vdd pmos_6p0 w=1.2u l=0.5u
X10924 vdd tune_series_gy[3] a_28484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X10925 a_24660_26786# cap_shunt_p a_26376_26724# vss nmos_6p0 w=0.82u l=0.6u
X10926 vss tune_shunt[7] a_21748_23650# vss nmos_6p0 w=0.51u l=0.6u
X10927 vdd a_13564_6647# a_13476_6744# vdd pmos_6p0 w=1.22u l=1u
X10928 a_20740_42104# cap_shunt_p a_21672_42104# vss nmos_6p0 w=0.82u l=0.6u
X10929 vss cap_series_gyp a_7960_4472# vss nmos_6p0 w=0.82u l=0.6u
X10930 a_7168_9176# cap_shunt_p a_5844_9176# vss nmos_6p0 w=0.82u l=0.6u
X10931 vdd a_2140_12919# a_2052_13016# vdd pmos_6p0 w=1.22u l=1u
X10932 a_3620_13396# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10933 a_6740_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10934 a_25572_30644# cap_shunt_p a_25780_31128# vdd pmos_6p0 w=1.2u l=0.5u
X10935 vdd tune_shunt[7] a_16500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X10936 vdd tune_shunt[5] a_3620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X10937 vdd tune_shunt[7] a_24452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X10938 vdd a_5612_33303# a_5524_33400# vdd pmos_6p0 w=1.22u l=1u
X10939 vdd tune_shunt[0] a_28484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X10940 a_14504_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10941 a_12788_20152# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X10942 a_17596_5512# a_17508_5556# vss vss nmos_6p0 w=0.82u l=1u
X10943 a_6740_12312# cap_shunt_p a_8456_12312# vss nmos_6p0 w=0.82u l=0.6u
X10944 vss tune_shunt[7] a_21748_20514# vss nmos_6p0 w=0.51u l=0.6u
X10945 a_17620_47892# cap_shunt_p a_17828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X10946 a_17828_37400# cap_shunt_n a_18760_37400# vss nmos_6p0 w=0.82u l=0.6u
X10947 vdd a_38092_27464# a_38004_27508# vdd pmos_6p0 w=1.22u l=1u
X10948 a_29624_6040# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10949 a_12444_19191# a_12356_19288# vss vss nmos_6p0 w=0.82u l=1u
X10950 a_17828_20152# cap_shunt_p a_19544_20152# vss nmos_6p0 w=0.82u l=0.6u
X10951 a_34844_52552# a_34756_52596# vss vss nmos_6p0 w=0.82u l=1u
X10952 vdd a_19612_55688# a_19524_55732# vdd pmos_6p0 w=1.22u l=1u
X10953 a_27228_42711# a_27140_42808# vss vss nmos_6p0 w=0.82u l=1u
X10954 a_19724_14487# a_19636_14584# vss vss nmos_6p0 w=0.82u l=1u
X10955 a_27888_20152# cap_series_gyp a_25780_20152# vss nmos_6p0 w=0.82u l=0.6u
X10956 vdd tune_shunt[6] a_3620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X10957 a_17828_17016# cap_shunt_p a_17620_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10958 vss tune_series_gygy[4] a_34516_12674# vss nmos_6p0 w=0.51u l=0.6u
X10959 a_7672_13880# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10960 a_9428_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X10961 vdd a_17596_49416# a_17508_49460# vdd pmos_6p0 w=1.22u l=1u
X10962 a_32040_22020# cap_series_gygyn a_31624_22428# vss nmos_6p0 w=0.82u l=0.6u
X10963 a_14504_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X10964 a_17620_44756# cap_shunt_p a_17828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X10965 a_9464_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10966 a_25996_55255# a_25908_55352# vss vss nmos_6p0 w=0.82u l=1u
X10967 vdd a_6508_8215# a_6420_8312# vdd pmos_6p0 w=1.22u l=1u
X10968 vdd a_31820_52552# a_31732_52596# vdd pmos_6p0 w=1.22u l=1u
X10969 a_34188_43672# cap_shunt_gyn a_33920_43734# vss nmos_6p0 w=0.82u l=0.6u
X10970 vdd a_29468_48983# a_29380_49080# vdd pmos_6p0 w=1.22u l=1u
X10971 a_33732_35832# cap_shunt_n a_33524_35348# vdd pmos_6p0 w=1.2u l=0.5u
X10972 vdd tune_series_gy[5] a_18404_11452# vdd pmos_6p0 w=1.2u l=0.5u
X10973 a_11460_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10974 vss cap_shunt_p a_33936_28292# vss nmos_6p0 w=0.82u l=0.6u
X10975 vdd tune_shunt[5] a_16500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X10976 a_9464_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10977 vdd tune_shunt[7] a_6196_22428# vdd pmos_6p0 w=1.2u l=0.5u
X10978 a_31436_6748# cap_series_gygyn a_31624_6748# vdd pmos_6p0 w=1.2u l=0.5u
X10979 a_12444_52552# a_12356_52596# vss vss nmos_6p0 w=0.82u l=1u
X10980 a_6420_13020# cap_shunt_p a_6628_12674# vdd pmos_6p0 w=1.2u l=0.5u
X10981 a_35692_16532# cap_series_gygyn a_35880_16532# vdd pmos_6p0 w=1.2u l=0.5u
X10982 vdd a_5836_7080# a_5748_7124# vdd pmos_6p0 w=1.22u l=1u
X10983 a_15356_13352# a_15268_13396# vss vss nmos_6p0 w=0.82u l=1u
X10984 a_4648_10744# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X10985 vdd a_31372_47848# a_31284_47892# vdd pmos_6p0 w=1.22u l=1u
X10986 vss cap_shunt_p a_33936_25156# vss nmos_6p0 w=0.82u l=0.6u
X10987 vdd tune_shunt[1] a_1716_3612# vdd pmos_6p0 w=1.2u l=0.5u
X10988 a_2500_9884# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10989 a_9332_11452# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X10990 a_35880_19668# cap_series_gygyp a_35692_19668# vdd pmos_6p0 w=1.2u l=0.5u
X10991 vss cap_shunt_n a_11984_37700# vss nmos_6p0 w=0.82u l=0.6u
X10992 a_27676_5079# a_27588_5176# vss vss nmos_6p0 w=0.82u l=1u
X10993 vss cap_shunt_p a_14112_48376# vss nmos_6p0 w=0.82u l=0.6u
X10994 vdd tune_shunt[4] a_17620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X10995 vss tune_shunt[5] a_28692_38968# vss nmos_6p0 w=0.51u l=0.6u
X10996 a_13588_25564# cap_shunt_n a_13796_25218# vdd pmos_6p0 w=1.2u l=0.5u
X10997 vdd tune_shunt[7] a_10452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X10998 a_30616_21236# cap_series_gygyn a_30428_21236# vdd pmos_6p0 w=1.2u l=0.5u
X10999 a_3640_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11000 a_34396_41576# a_34308_41620# vss vss nmos_6p0 w=0.82u l=1u
X11001 a_3172_18100# cap_shunt_p a_3380_18584# vdd pmos_6p0 w=1.2u l=0.5u
X11002 a_10660_4834# cap_series_gyp a_11592_4772# vss nmos_6p0 w=0.82u l=0.6u
X11003 a_28692_9176# cap_series_gyn a_28484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X11004 vdd tune_shunt[6] a_17620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X11005 a_37632_38485# cap_shunt_gyp a_37444_38485# vdd pmos_6p0 w=1.215u l=0.5u
X11006 a_13588_22428# cap_shunt_n a_13796_22082# vdd pmos_6p0 w=1.2u l=0.5u
X11007 a_6532_25940# cap_shunt_n a_6740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X11008 a_18612_9538# cap_series_gyp a_18404_9884# vdd pmos_6p0 w=1.2u l=0.5u
X11009 a_13252_32212# cap_shunt_n a_13460_32696# vdd pmos_6p0 w=1.2u l=0.5u
X11010 a_20740_27992# cap_shunt_n a_22456_27992# vss nmos_6p0 w=0.82u l=0.6u
X11011 a_13796_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11012 vss tune_shunt[3] a_25780_43672# vss nmos_6p0 w=0.51u l=0.6u
X11013 a_6740_53080# cap_shunt_n a_6532_52596# vdd pmos_6p0 w=1.2u l=0.5u
X11014 a_14580_46808# cap_shunt_p a_14372_46324# vdd pmos_6p0 w=1.2u l=0.5u
X11015 a_37652_40536# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X11016 vss cap_shunt_p a_27888_37400# vss nmos_6p0 w=0.82u l=0.6u
X11017 vdd tune_shunt[7] a_10452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X11018 a_28692_6040# cap_shunt_n a_28484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X11019 a_25572_24372# cap_shunt_p a_25780_24856# vdd pmos_6p0 w=1.2u l=0.5u
X11020 vdd tune_series_gy[3] a_25572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X11021 a_5844_11106# cap_shunt_n a_5636_11452# vdd pmos_6p0 w=1.2u l=0.5u
X11022 a_6532_22804# cap_shunt_p a_6740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X11023 a_18612_6402# cap_series_gyn a_18404_6748# vdd pmos_6p0 w=1.2u l=0.5u
X11024 a_34348_8316# cap_series_gygyp a_34536_8316# vdd pmos_6p0 w=1.2u l=0.5u
X11025 vdd a_30812_42711# a_30724_42808# vdd pmos_6p0 w=1.22u l=1u
X11026 vdd tune_series_gy[4] a_15492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X11027 vss cap_series_gygyn a_36624_18884# vss nmos_6p0 w=0.82u l=0.6u
X11028 a_20740_24856# cap_shunt_n a_22456_24856# vss nmos_6p0 w=0.82u l=0.6u
X11029 vss tune_shunt[6] a_14580_43672# vss nmos_6p0 w=0.51u l=0.6u
X11030 vss tune_shunt[5] a_25780_40536# vss nmos_6p0 w=0.51u l=0.6u
X11031 a_7540_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11032 a_13796_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11033 a_13588_34972# cap_shunt_n a_13796_34626# vdd pmos_6p0 w=1.2u l=0.5u
X11034 a_24660_17378# cap_series_gyp a_26376_17316# vss nmos_6p0 w=0.82u l=0.6u
X11035 a_23308_43144# a_23220_43188# vss vss nmos_6p0 w=0.82u l=1u
X11036 vss tune_series_gy[5] a_21748_14242# vss nmos_6p0 w=0.51u l=0.6u
X11037 vdd tune_shunt[6] a_2500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X11038 a_21748_28354# cap_shunt_n a_21540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X11039 a_6740_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11040 a_25572_21236# cap_shunt_p a_25780_21720# vdd pmos_6p0 w=1.2u l=0.5u
X11041 a_27228_36439# a_27140_36536# vss vss nmos_6p0 w=0.82u l=1u
X11042 vss tune_series_gygy[1] a_34516_4834# vss nmos_6p0 w=0.51u l=0.6u
X11043 a_25592_18884# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X11044 vdd tune_shunt[6] a_3620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X11045 a_27104_35832# cap_shunt_p a_25780_35832# vss nmos_6p0 w=0.82u l=0.6u
X11046 vdd a_9980_3511# a_9892_3608# vdd pmos_6p0 w=1.22u l=1u
X11047 a_5844_11106# cap_shunt_n a_6776_11044# vss nmos_6p0 w=0.82u l=0.6u
X11048 vss cap_series_gygyn a_36624_15748# vss nmos_6p0 w=0.82u l=0.6u
X11049 a_9316_50306# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11050 vss tune_shunt[6] a_14580_40536# vss nmos_6p0 w=0.51u l=0.6u
X11051 a_20532_40052# cap_shunt_p a_20740_40536# vdd pmos_6p0 w=1.2u l=0.5u
X11052 a_2708_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11053 a_13588_31836# cap_shunt_n a_13796_31490# vdd pmos_6p0 w=1.2u l=0.5u
X11054 a_23308_40008# a_23220_40052# vss vss nmos_6p0 w=0.82u l=1u
X11055 a_17620_38484# cap_shunt_n a_17828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X11056 a_9464_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11057 vss tune_shunt[7] a_9316_22082# vss nmos_6p0 w=0.51u l=0.6u
X11058 vss tune_series_gy[5] a_21748_11106# vss nmos_6p0 w=0.51u l=0.6u
X11059 vss tune_series_gygy[5] a_35880_22804# vss nmos_6p0 w=0.51u l=0.6u
X11060 a_25996_48983# a_25908_49080# vss vss nmos_6p0 w=0.82u l=1u
X11061 vss tune_shunt_gy[5] a_37632_49080# vss nmos_6p0 w=0.51u l=0.6u
X11062 a_19152_43672# cap_shunt_p a_17828_43672# vss nmos_6p0 w=0.82u l=0.6u
X11063 a_28692_10744# cap_series_gyp a_28484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X11064 a_25592_15748# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X11065 vdd tune_shunt[6] a_3620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11066 a_6292_18584# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11067 a_5544_32696# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11068 a_33732_29560# cap_shunt_p a_33524_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11069 a_1924_6040# cap_shunt_p a_3640_6040# vss nmos_6p0 w=0.82u l=0.6u
X11070 a_27788_50984# a_27700_51028# vss vss nmos_6p0 w=0.82u l=1u
X11071 a_17620_35348# cap_shunt_n a_17828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X11072 a_9464_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11073 vss tune_shunt[5] a_9204_51874# vss nmos_6p0 w=0.51u l=0.6u
X11074 a_9668_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11075 a_19152_40536# cap_shunt_n a_17828_40536# vss nmos_6p0 w=0.82u l=0.6u
X11076 vss cap_shunt_p a_31024_4772# vss nmos_6p0 w=0.82u l=0.6u
X11077 a_31024_34564# cap_shunt_p a_29700_34626# vss nmos_6p0 w=0.82u l=0.6u
X11078 vdd a_36636_53687# a_36548_53784# vdd pmos_6p0 w=1.22u l=1u
X11079 vss cap_series_gyp a_23632_3204# vss nmos_6p0 w=0.82u l=0.6u
X11080 a_31708_53687# a_31620_53784# vss vss nmos_6p0 w=0.82u l=1u
X11081 vdd tune_shunt[7] a_16500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X11082 a_36532_42104# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X11083 a_10452_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11084 vdd tune_shunt[7] a_9332_14588# vdd pmos_6p0 w=1.2u l=0.5u
X11085 a_13588_19292# cap_shunt_p a_13796_18946# vdd pmos_6p0 w=1.2u l=0.5u
X11086 vdd tune_shunt[5] a_20532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X11087 a_9644_35304# a_9556_35348# vss vss nmos_6p0 w=0.82u l=1u
X11088 a_18816_48676# cap_shunt_p a_16708_48738# vss nmos_6p0 w=0.82u l=0.6u
X11089 a_31024_31428# cap_shunt_p a_29700_31490# vss nmos_6p0 w=0.82u l=0.6u
X11090 a_5844_9176# cap_shunt_p a_5636_8692# vdd pmos_6p0 w=1.2u l=0.5u
X11091 a_17828_40536# cap_shunt_n a_17620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X11092 a_31708_50551# a_31620_50648# vss vss nmos_6p0 w=0.82u l=1u
X11093 a_15120_47108# cap_shunt_p a_13796_47170# vss nmos_6p0 w=0.82u l=0.6u
X11094 vdd tune_shunt[6] a_17620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X11095 a_13588_16156# cap_shunt_p a_13796_15810# vdd pmos_6p0 w=1.2u l=0.5u
X11096 vss cap_shunt_p a_4032_45540# vss nmos_6p0 w=0.82u l=0.6u
X11097 vdd a_17260_50551# a_17172_50648# vdd pmos_6p0 w=1.22u l=1u
X11098 vss cap_shunt_n a_11200_53080# vss nmos_6p0 w=0.82u l=0.6u
X11099 a_25100_52119# a_25012_52216# vss vss nmos_6p0 w=0.82u l=1u
X11100 a_12332_50551# a_12244_50648# vss vss nmos_6p0 w=0.82u l=1u
X11101 vdd tune_series_gy[5] a_22436_10260# vdd pmos_6p0 w=1.2u l=0.5u
X11102 a_37652_34264# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X11103 a_24452_42812# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11104 vdd tune_shunt[7] a_17620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11105 a_33732_35832# cap_shunt_n a_33524_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11106 a_10680_8316# cap_series_gyp a_10492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X11107 vdd tune_shunt[5] a_9668_52596# vdd pmos_6p0 w=1.2u l=0.5u
X11108 vss cap_shunt_p a_4032_42404# vss nmos_6p0 w=0.82u l=0.6u
X11109 vdd a_34844_55688# a_34756_55732# vdd pmos_6p0 w=1.22u l=1u
X11110 a_13796_47170# cap_shunt_p a_13588_47516# vdd pmos_6p0 w=1.2u l=0.5u
X11111 a_20740_18584# cap_shunt_p a_22456_18584# vss nmos_6p0 w=0.82u l=0.6u
X11112 a_9316_47170# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11113 a_6420_13020# cap_shunt_p a_6628_12674# vdd pmos_6p0 w=1.2u l=0.5u
X11114 a_13796_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11115 vss tune_shunt[7] a_20740_21720# vss nmos_6p0 w=0.51u l=0.6u
X11116 a_14784_37400# cap_shunt_n a_13460_37400# vss nmos_6p0 w=0.82u l=0.6u
X11117 vss tune_shunt[6] a_25780_34264# vss nmos_6p0 w=0.51u l=0.6u
X11118 a_33524_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11119 a_12780_54120# a_12692_54164# vss vss nmos_6p0 w=0.82u l=1u
X11120 a_6740_43672# cap_shunt_p a_6532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X11121 a_2708_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11122 vdd tune_shunt[6] a_2500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X11123 vdd a_2140_33736# a_2052_33780# vdd pmos_6p0 w=1.22u l=1u
X11124 vdd tune_shunt[7] a_24452_20860# vdd pmos_6p0 w=1.2u l=0.5u
X11125 a_27104_29560# cap_shunt_p a_25780_29560# vss nmos_6p0 w=0.82u l=0.6u
X11126 a_20740_15448# cap_series_gyn a_22456_15448# vss nmos_6p0 w=0.82u l=0.6u
X11127 vss tune_shunt[7] a_25780_31128# vss nmos_6p0 w=0.51u l=0.6u
X11128 a_13588_25564# cap_shunt_n a_13796_25218# vdd pmos_6p0 w=1.2u l=0.5u
X11129 vdd tune_series_gy[4] a_18404_3988# vdd pmos_6p0 w=1.2u l=0.5u
X11130 a_23308_33736# a_23220_33780# vss vss nmos_6p0 w=0.82u l=1u
X11131 a_30616_21236# cap_series_gygyn a_30428_21236# vdd pmos_6p0 w=1.2u l=0.5u
X11132 vdd a_27340_55255# a_27252_55352# vdd pmos_6p0 w=1.22u l=1u
X11133 vdd tune_shunt[7] a_2500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X11134 vdd a_2140_30600# a_2052_30644# vdd pmos_6p0 w=1.22u l=1u
X11135 a_12556_14487# a_12468_14584# vss vss nmos_6p0 w=0.82u l=1u
X11136 a_29700_17378# cap_series_gyp a_29492_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11137 vdd tune_shunt[7] a_3620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11138 a_27104_26424# cap_shunt_p a_25780_26424# vss nmos_6p0 w=0.82u l=0.6u
X11139 a_9540_9538# cap_shunt_p a_11256_9476# vss nmos_6p0 w=0.82u l=0.6u
X11140 a_2708_9538# cap_shunt_n a_4424_9476# vss nmos_6p0 w=0.82u l=0.6u
X11141 a_33920_43189# cap_shunt_gyn a_33920_43734# vdd pmos_6p0 w=1.215u l=0.5u
X11142 a_2708_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11143 a_13588_22428# cap_shunt_n a_13796_22082# vdd pmos_6p0 w=1.2u l=0.5u
X11144 a_27788_44712# a_27700_44756# vss vss nmos_6p0 w=0.82u l=1u
X11145 a_28692_37400# cap_shunt_p a_28484_36916# vdd pmos_6p0 w=1.2u l=0.5u
X11146 a_17620_33780# cap_shunt_n a_17828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X11147 a_23308_30600# a_23220_30644# vss vss nmos_6p0 w=0.82u l=1u
X11148 a_6532_25940# cap_shunt_n a_6740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X11149 vdd a_27340_52119# a_27252_52216# vdd pmos_6p0 w=1.22u l=1u
X11150 a_17620_29076# cap_shunt_n a_17828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X11151 vdd a_6060_38007# a_5972_38104# vdd pmos_6p0 w=1.22u l=1u
X11152 a_19152_34264# cap_shunt_n a_17828_34264# vss nmos_6p0 w=0.82u l=0.6u
X11153 vdd tune_shunt[6] a_9108_47516# vdd pmos_6p0 w=1.2u l=0.5u
X11154 vss tune_shunt_gy[1] a_37632_39672# vss nmos_6p0 w=0.51u l=0.6u
X11155 a_12556_11351# a_12468_11448# vss vss nmos_6p0 w=0.82u l=1u
X11156 a_20532_19668# cap_shunt_p a_20740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X11157 a_6740_53080# cap_shunt_n a_6532_52596# vdd pmos_6p0 w=1.2u l=0.5u
X11158 a_28692_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11159 a_31024_28292# cap_shunt_p a_29700_28354# vss nmos_6p0 w=0.82u l=0.6u
X11160 a_5544_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11161 a_9220_19292# cap_shunt_p a_9428_18946# vdd pmos_6p0 w=1.2u l=0.5u
X11162 a_17620_30644# cap_shunt_n a_17828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X11163 a_6532_22804# cap_shunt_p a_6740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X11164 a_11612_7124# cap_series_gyp a_11800_7124# vdd pmos_6p0 w=1.2u l=0.5u
X11165 a_2500_9884# cap_shunt_n a_2708_9538# vdd pmos_6p0 w=1.2u l=0.5u
X11166 a_19152_31128# cap_shunt_n a_17828_31128# vss nmos_6p0 w=0.82u l=0.6u
X11167 a_21748_44034# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11168 a_9644_29032# a_9556_29076# vss vss nmos_6p0 w=0.82u l=1u
X11169 a_28692_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11170 a_31024_25156# cap_shunt_p a_29700_25218# vss nmos_6p0 w=0.82u l=0.6u
X11171 a_9668_47892# cap_shunt_p a_9876_48376# vdd pmos_6p0 w=1.2u l=0.5u
X11172 vdd tune_shunt[6] a_2500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X11173 a_10548_38968# cap_shunt_n a_10340_38484# vdd pmos_6p0 w=1.2u l=0.5u
X11174 a_21748_28354# cap_shunt_n a_21540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X11175 a_35880_25940# cap_series_gygyp a_36688_26424# vss nmos_6p0 w=0.82u l=0.6u
X11176 a_9644_25896# a_9556_25940# vss vss nmos_6p0 w=0.82u l=1u
X11177 a_7516_54120# a_7428_54164# vss vss nmos_6p0 w=0.82u l=1u
X11178 a_18816_39268# cap_shunt_n a_16708_39330# vss nmos_6p0 w=0.82u l=0.6u
X11179 a_10548_35832# cap_shunt_n a_10340_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11180 vss tune_series_gy[5] a_22644_9176# vss nmos_6p0 w=0.51u l=0.6u
X11181 a_29492_17724# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11182 a_15176_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11183 a_11572_5556# cap_series_gyn a_11780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X11184 a_23980_47848# a_23892_47892# vss vss nmos_6p0 w=0.82u l=1u
X11185 vdd tune_shunt[7] a_12580_16532# vdd pmos_6p0 w=1.2u l=0.5u
X11186 vss cap_shunt_n a_4032_36132# vss nmos_6p0 w=0.82u l=0.6u
X11187 a_24452_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11188 vdd tune_shunt[7] a_17620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11189 a_33732_29560# cap_shunt_p a_33524_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11190 a_25780_6040# cap_series_gyp a_26712_6040# vss nmos_6p0 w=0.82u l=0.6u
X11191 a_36288_39672# cap_shunt_gyn a_36100_39672# vdd pmos_6p0 w=1.215u l=0.5u
X11192 a_35904_24856# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X11193 vdd a_34844_49416# a_34756_49460# vdd pmos_6p0 w=1.22u l=1u
X11194 a_1924_4834# cap_shunt_p a_1716_5180# vdd pmos_6p0 w=1.2u l=0.5u
X11195 vss cap_shunt_p a_18816_18884# vss nmos_6p0 w=0.82u l=0.6u
X11196 vdd a_27004_45847# a_26916_45944# vdd pmos_6p0 w=1.22u l=1u
X11197 a_24452_33404# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11198 a_9332_14588# cap_shunt_p a_9540_14242# vdd pmos_6p0 w=1.2u l=0.5u
X11199 vss cap_shunt_p a_4032_4472# vss nmos_6p0 w=0.82u l=0.6u
X11200 vdd a_15804_14920# a_15716_14964# vdd pmos_6p0 w=1.22u l=1u
X11201 a_3036_52552# a_2948_52596# vss vss nmos_6p0 w=0.82u l=1u
X11202 a_3620_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11203 a_13796_37762# cap_shunt_n a_13588_38108# vdd pmos_6p0 w=1.2u l=0.5u
X11204 a_37420_34871# a_37332_34968# vss vss nmos_6p0 w=0.82u l=1u
X11205 a_21748_29922# cap_shunt_n a_21540_30268# vdd pmos_6p0 w=1.2u l=0.5u
X11206 a_21428_5556# cap_series_gyp a_21636_6040# vdd pmos_6p0 w=1.2u l=0.5u
X11207 vdd a_16364_12919# a_16276_13016# vdd pmos_6p0 w=1.22u l=1u
X11208 a_6740_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11209 vss cap_shunt_p a_18816_15748# vss nmos_6p0 w=0.82u l=0.6u
X11210 a_13588_19292# cap_shunt_p a_13796_18946# vdd pmos_6p0 w=1.2u l=0.5u
X11211 a_16500_49084# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11212 a_4032_48676# cap_shunt_p a_2708_48738# vss nmos_6p0 w=0.82u l=0.6u
X11213 vdd a_27340_48983# a_27252_49080# vdd pmos_6p0 w=1.22u l=1u
X11214 vdd tune_shunt[7] a_2500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X11215 a_32604_13352# a_32516_13396# vss vss nmos_6p0 w=0.82u l=1u
X11216 a_22524_49416# a_22436_49460# vss vss nmos_6p0 w=0.82u l=1u
X11217 a_11460_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11218 a_3248_6040# cap_shunt_p a_1924_6040# vss nmos_6p0 w=0.82u l=0.6u
X11219 vdd a_15804_11784# a_15716_11828# vdd pmos_6p0 w=1.22u l=1u
X11220 a_37420_31735# a_37332_31832# vss vss nmos_6p0 w=0.82u l=1u
X11221 vdd a_2140_24328# a_2052_24372# vdd pmos_6p0 w=1.22u l=1u
X11222 vss cap_series_gyn a_23072_6340# vss nmos_6p0 w=0.82u l=0.6u
X11223 vdd tune_series_gy[5] a_24452_11452# vdd pmos_6p0 w=1.2u l=0.5u
X11224 vdd a_33948_18056# a_33860_18100# vdd pmos_6p0 w=1.22u l=1u
X11225 a_17828_46808# cap_shunt_n a_17620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X11226 a_10452_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11227 a_21748_37762# cap_shunt_n a_22680_37700# vss nmos_6p0 w=0.82u l=0.6u
X11228 a_13588_16156# cap_shunt_p a_13796_15810# vdd pmos_6p0 w=1.2u l=0.5u
X11229 a_32604_10216# a_32516_10260# vss vss nmos_6p0 w=0.82u l=1u
X11230 vss cap_shunt_n a_12656_35832# vss nmos_6p0 w=0.82u l=0.6u
X11231 vss tune_shunt[7] a_16708_26786# vss nmos_6p0 w=0.51u l=0.6u
X11232 vdd tune_series_gy[5] a_22436_10260# vdd pmos_6p0 w=1.2u l=0.5u
X11233 a_23240_3204# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X11234 vdd a_2140_21192# a_2052_21236# vdd pmos_6p0 w=1.22u l=1u
X11235 vdd a_19388_52552# a_19300_52596# vdd pmos_6p0 w=1.22u l=1u
X11236 vdd a_28124_34871# a_28036_34968# vdd pmos_6p0 w=1.22u l=1u
X11237 a_27104_17016# cap_series_gyp a_25780_17016# vss nmos_6p0 w=0.82u l=0.6u
X11238 a_21540_42812# cap_shunt_n a_21748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X11239 a_19524_13396# cap_series_gyn a_19732_13880# vdd pmos_6p0 w=1.2u l=0.5u
X11240 a_4760_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11241 a_34844_38440# a_34756_38484# vss vss nmos_6p0 w=0.82u l=1u
X11242 a_28692_27992# cap_shunt_p a_28484_27508# vdd pmos_6p0 w=1.2u l=0.5u
X11243 a_17620_24372# cap_shunt_n a_17828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X11244 a_13796_47170# cap_shunt_p a_13588_47516# vdd pmos_6p0 w=1.2u l=0.5u
X11245 a_9876_13880# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11246 a_28692_18584# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11247 a_6740_43672# cap_shunt_p a_6532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X11248 vdd tune_shunt[6] a_2500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X11249 a_35448_12612# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X11250 a_17620_21236# cap_shunt_p a_17828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X11251 a_17620_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11252 a_9876_10744# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11253 vss tune_shunt[7] a_25780_21720# vss nmos_6p0 w=0.51u l=0.6u
X11254 a_12768_29860# cap_shunt_n a_10660_29922# vss nmos_6p0 w=0.82u l=0.6u
X11255 a_12892_19191# a_12804_19288# vss vss nmos_6p0 w=0.82u l=1u
X11256 a_7748_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11257 a_27676_42711# a_27588_42808# vss vss nmos_6p0 w=0.82u l=1u
X11258 a_34516_4834# cap_series_gygyp a_34308_5180# vdd pmos_6p0 w=1.2u l=0.5u
X11259 a_28692_15448# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11260 vdd a_33500_40008# a_33412_40052# vdd pmos_6p0 w=1.22u l=1u
X11261 a_10548_29560# cap_shunt_n a_10340_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11262 vdd tune_shunt[7] a_2500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X11263 a_35880_16532# cap_series_gygyn a_36688_17016# vss nmos_6p0 w=0.82u l=0.6u
X11264 a_17828_37400# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11265 a_29700_17378# cap_series_gyp a_29492_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11266 a_10680_8316# cap_series_gyp a_10492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X11267 a_12768_26724# cap_shunt_n a_10660_26786# vss nmos_6p0 w=0.82u l=0.6u
X11268 a_4816_43972# cap_shunt_p a_2708_44034# vss nmos_6p0 w=0.82u l=0.6u
X11269 a_25780_38968# cap_shunt_p a_27496_38968# vss nmos_6p0 w=0.82u l=0.6u
X11270 a_35904_18584# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X11271 a_28692_37400# cap_shunt_p a_28484_36916# vdd pmos_6p0 w=1.2u l=0.5u
X11272 vdd tune_shunt[7] a_6532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X11273 vdd tune_shunt[7] a_13252_33780# vdd pmos_6p0 w=1.2u l=0.5u
X11274 vdd tune_shunt[7] a_3172_16532# vdd pmos_6p0 w=1.2u l=0.5u
X11275 vdd tune_shunt[6] a_3620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X11276 a_20532_19668# cap_shunt_p a_20740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X11277 a_7404_55255# a_7316_55352# vss vss nmos_6p0 w=0.82u l=1u
X11278 a_8064_32696# cap_shunt_n a_6740_32696# vss nmos_6p0 w=0.82u l=0.6u
X11279 a_6508_30167# a_6420_30264# vss vss nmos_6p0 w=0.82u l=1u
X11280 a_15176_23288# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11281 a_24452_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11282 a_35880_5556# tune_series_gygy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X11283 vdd a_2588_52552# a_2500_52596# vdd pmos_6p0 w=1.22u l=1u
X11284 a_12892_52552# a_12804_52596# vss vss nmos_6p0 w=0.82u l=1u
X11285 a_4816_40836# cap_shunt_p a_2708_40898# vss nmos_6p0 w=0.82u l=0.6u
X11286 vdd a_23308_36872# a_23220_36916# vdd pmos_6p0 w=1.22u l=1u
X11287 a_35904_15448# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X11288 a_9220_19292# cap_shunt_p a_9428_18946# vdd pmos_6p0 w=1.2u l=0.5u
X11289 a_37420_28599# a_37332_28696# vss vss nmos_6p0 w=0.82u l=1u
X11290 vss cap_shunt_n a_31808_37700# vss nmos_6p0 w=0.82u l=0.6u
X11291 vdd tune_shunt[7] a_13252_30644# vdd pmos_6p0 w=1.2u l=0.5u
X11292 a_13796_29922# cap_shunt_n a_13588_30268# vdd pmos_6p0 w=1.2u l=0.5u
X11293 a_24660_6402# cap_series_gyn a_25592_6340# vss nmos_6p0 w=0.82u l=0.6u
X11294 vdd tune_series_gy[4] a_18404_3988# vdd pmos_6p0 w=1.2u l=0.5u
X11295 a_10660_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11296 vdd tune_shunt[7] a_3620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X11297 a_6508_27031# a_6420_27128# vss vss nmos_6p0 w=0.82u l=1u
X11298 vss cap_shunt_gyn a_35756_42104# vss nmos_6p0 w=0.82u l=0.6u
X11299 a_10548_38968# cap_shunt_n a_10340_38484# vdd pmos_6p0 w=1.2u l=0.5u
X11300 a_37420_25463# a_37332_25560# vss vss nmos_6p0 w=0.82u l=1u
X11301 vss tune_shunt[6] a_3828_37400# vss nmos_6p0 w=0.51u l=0.6u
X11302 a_10452_36540# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11303 vss cap_shunt_n a_9856_32996# vss nmos_6p0 w=0.82u l=0.6u
X11304 a_14460_6647# a_14372_6744# vss vss nmos_6p0 w=0.82u l=1u
X11305 vss cap_shunt_p a_22064_21720# vss nmos_6p0 w=0.82u l=0.6u
X11306 a_4032_39268# cap_shunt_n a_2708_39330# vss nmos_6p0 w=0.82u l=0.6u
X11307 a_32632_11452# cap_series_gyp a_32444_11452# vdd pmos_6p0 w=1.2u l=0.5u
X11308 a_31808_14180# cap_series_gyp a_29700_14242# vss nmos_6p0 w=0.82u l=0.6u
X11309 a_37980_43144# a_37892_43188# vss vss nmos_6p0 w=0.82u l=1u
X11310 a_32404_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11311 vdd tune_series_gygy[4] a_35692_10260# vdd pmos_6p0 w=1.2u l=0.5u
X11312 a_10548_35832# cap_shunt_n a_10340_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11313 vss cap_shunt_n a_12656_29560# vss nmos_6p0 w=0.82u l=0.6u
X11314 vss tune_shunt[2] a_1924_6402# vss nmos_6p0 w=0.51u l=0.6u
X11315 a_17640_47108# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11316 vdd a_28124_28599# a_28036_28696# vdd pmos_6p0 w=1.22u l=1u
X11317 a_2500_50652# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11318 a_21540_36540# cap_shunt_n a_21748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X11319 a_10452_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11320 a_34516_12674# cap_series_gygyp a_36232_12612# vss nmos_6p0 w=0.82u l=0.6u
X11321 a_6516_20514# cap_shunt_p a_6308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X11322 a_31808_11044# cap_series_gyp a_29700_11106# vss nmos_6p0 w=0.82u l=0.6u
X11323 vss tune_shunt[7] a_10548_32696# vss nmos_6p0 w=0.51u l=0.6u
X11324 vss cap_shunt_n a_12656_26424# vss nmos_6p0 w=0.82u l=0.6u
X11325 vss tune_shunt[7] a_16708_17378# vss nmos_6p0 w=0.51u l=0.6u
X11326 a_21540_33404# cap_shunt_n a_21748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X11327 a_24660_23650# cap_shunt_p a_24452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X11328 vss tune_shunt[7] a_13796_31490# vss nmos_6p0 w=0.51u l=0.6u
X11329 a_11872_27992# cap_shunt_n a_10548_27992# vss nmos_6p0 w=0.82u l=0.6u
X11330 a_13796_37762# cap_shunt_n a_13588_38108# vdd pmos_6p0 w=1.2u l=0.5u
X11331 a_20172_33303# a_20084_33400# vss vss nmos_6p0 w=0.82u l=1u
X11332 a_30408_32696# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11333 vdd a_3932_55255# a_3844_55352# vdd pmos_6p0 w=1.22u l=1u
X11334 a_23756_43144# a_23668_43188# vss vss nmos_6p0 w=0.82u l=1u
X11335 vss tune_shunt[6] a_7748_40898# vss nmos_6p0 w=0.51u l=0.6u
X11336 a_18940_7080# a_18852_7124# vss vss nmos_6p0 w=0.82u l=1u
X11337 vss cap_shunt_p a_26768_39268# vss nmos_6p0 w=0.82u l=0.6u
X11338 vdd a_6060_55688# a_5972_55732# vdd pmos_6p0 w=1.22u l=1u
X11339 a_27676_36439# a_27588_36536# vss vss nmos_6p0 w=0.82u l=1u
X11340 vss cap_shunt_p a_11984_13880# vss nmos_6p0 w=0.82u l=0.6u
X11341 a_10808_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11342 vdd tune_shunt[7] a_2500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X11343 a_11872_24856# cap_shunt_n a_10548_24856# vss nmos_6p0 w=0.82u l=0.6u
X11344 vss tune_series_gy[5] a_25780_12312# vss nmos_6p0 w=0.51u l=0.6u
X11345 vdd a_3932_52119# a_3844_52216# vdd pmos_6p0 w=1.22u l=1u
X11346 a_23756_40008# a_23668_40052# vss vss nmos_6p0 w=0.82u l=1u
X11347 vdd tune_series_gy[5] a_21540_9884# vdd pmos_6p0 w=1.2u l=0.5u
X11348 a_18940_49416# a_18852_49460# vss vss nmos_6p0 w=0.82u l=1u
X11349 vss cap_shunt_p a_11984_10744# vss nmos_6p0 w=0.82u l=0.6u
X11350 vdd a_35292_13352# a_35204_13396# vdd pmos_6p0 w=1.22u l=1u
X11351 a_4940_3944# a_4852_3988# vss vss nmos_6p0 w=0.82u l=1u
X11352 vdd a_3036_55688# a_2948_55732# vdd pmos_6p0 w=1.22u l=1u
X11353 a_28484_40052# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11354 a_14692_6040# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X11355 vdd a_33164_17623# a_33076_17720# vdd pmos_6p0 w=1.22u l=1u
X11356 a_25780_20152# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11357 vdd tune_shunt[6] a_29492_34972# vdd pmos_6p0 w=1.2u l=0.5u
X11358 vss tune_shunt[6] a_2708_45602# vss nmos_6p0 w=0.51u l=0.6u
X11359 a_21540_42812# cap_shunt_n a_21748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X11360 a_14392_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11361 vdd tune_series_gy[4] a_21540_6748# vdd pmos_6p0 w=1.2u l=0.5u
X11362 vss tune_shunt[5] a_9204_51874# vss nmos_6p0 w=0.51u l=0.6u
X11363 a_4816_34564# cap_shunt_n a_2708_34626# vss nmos_6p0 w=0.82u l=0.6u
X11364 vdd a_32604_7080# a_32516_7124# vdd pmos_6p0 w=1.22u l=1u
X11365 vdd a_18940_10216# a_18852_10260# vdd pmos_6p0 w=1.22u l=1u
X11366 a_28692_27992# cap_shunt_p a_28484_27508# vdd pmos_6p0 w=1.2u l=0.5u
X11367 a_6760_3988# cap_series_gyp a_6572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X11368 vdd tune_shunt[7] a_13252_24372# vdd pmos_6p0 w=1.2u l=0.5u
X11369 a_29532_16156# cap_series_gyn a_29720_16156# vdd pmos_6p0 w=1.2u l=0.5u
X11370 vdd tune_shunt[7] a_3620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X11371 a_8064_23288# cap_shunt_p a_6740_23288# vss nmos_6p0 w=0.82u l=0.6u
X11372 a_18404_13020# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11373 vdd tune_shunt[5] a_29492_31836# vdd pmos_6p0 w=1.2u l=0.5u
X11374 a_6404_47170# cap_shunt_p a_8120_47108# vss nmos_6p0 w=0.82u l=0.6u
X11375 vdd a_23308_27464# a_23220_27508# vdd pmos_6p0 w=1.22u l=1u
X11376 a_36688_4472# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X11377 vdd a_2588_43144# a_2500_43188# vdd pmos_6p0 w=1.22u l=1u
X11378 vdd a_35180_34871# a_35092_34968# vdd pmos_6p0 w=1.22u l=1u
X11379 a_4816_31428# cap_shunt_p a_2708_31490# vss nmos_6p0 w=0.82u l=0.6u
X11380 a_32612_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11381 a_18404_9884# cap_series_gyp a_18612_9538# vdd pmos_6p0 w=1.2u l=0.5u
X11382 a_21748_20514# cap_shunt_p a_21540_20860# vdd pmos_6p0 w=1.2u l=0.5u
X11383 vdd tune_shunt[7] a_13252_21236# vdd pmos_6p0 w=1.2u l=0.5u
X11384 vss cap_shunt_p a_11648_15748# vss nmos_6p0 w=0.82u l=0.6u
X11385 vss cap_shunt_p a_8400_17016# vss nmos_6p0 w=0.82u l=0.6u
X11386 vdd tune_shunt[5] a_3620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X11387 a_11612_8692# cap_series_gyp a_11800_8692# vdd pmos_6p0 w=1.2u l=0.5u
X11388 a_7168_11044# cap_shunt_n a_5844_11106# vss nmos_6p0 w=0.82u l=0.6u
X11389 vdd a_20172_48983# a_20084_49080# vdd pmos_6p0 w=1.22u l=1u
X11390 a_13720_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11391 a_10548_29560# cap_shunt_n a_10340_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11392 a_33500_22760# a_33412_22804# vss vss nmos_6p0 w=0.82u l=1u
X11393 a_28236_55255# a_28148_55352# vss vss nmos_6p0 w=0.82u l=1u
X11394 a_14580_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11395 a_25780_42104# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11396 vdd tune_shunt[4] a_33524_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11397 a_18404_6748# cap_series_gyn a_18612_6402# vdd pmos_6p0 w=1.2u l=0.5u
X11398 a_7616_18584# cap_shunt_p a_6292_18584# vss nmos_6p0 w=0.82u l=0.6u
X11399 a_10452_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11400 vss cap_shunt_p a_9856_23588# vss nmos_6p0 w=0.82u l=0.6u
X11401 vdd a_16252_19624# a_16164_19668# vdd pmos_6p0 w=1.22u l=1u
X11402 a_2500_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11403 a_12780_50551# a_12692_50648# vss vss nmos_6p0 w=0.82u l=1u
X11404 a_6420_13020# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11405 a_19936_46808# cap_shunt_n a_17828_46808# vss nmos_6p0 w=0.82u l=0.6u
X11406 vss cap_series_gyp a_7176_4472# vss nmos_6p0 w=0.82u l=0.6u
X11407 a_19524_10260# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11408 vss tune_shunt[4] a_29700_39330# vss nmos_6p0 w=0.51u l=0.6u
X11409 a_14580_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11410 a_3828_42104# cap_shunt_p a_3620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X11411 a_9540_14242# cap_shunt_p a_11256_14180# vss nmos_6p0 w=0.82u l=0.6u
X11412 a_20532_19668# cap_shunt_p a_20740_20152# vdd pmos_6p0 w=1.2u l=0.5u
X11413 a_11200_49944# cap_shunt_p a_9876_49944# vss nmos_6p0 w=0.82u l=0.6u
X11414 vdd a_28124_19191# a_28036_19288# vdd pmos_6p0 w=1.22u l=1u
X11415 a_2500_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11416 a_21540_27132# cap_shunt_n a_21748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X11417 vss tune_shunt[7] a_10548_23288# vss nmos_6p0 w=0.51u l=0.6u
X11418 a_11884_22327# a_11796_22424# vss vss nmos_6p0 w=0.82u l=1u
X11419 a_35880_7124# cap_series_gygyp a_35692_7124# vdd pmos_6p0 w=1.2u l=0.5u
X11420 vss cap_shunt_p a_11424_48676# vss nmos_6p0 w=0.82u l=0.6u
X11421 a_21540_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11422 a_13796_29922# cap_shunt_n a_13588_30268# vdd pmos_6p0 w=1.2u l=0.5u
X11423 a_10660_6402# cap_series_gyn a_10452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X11424 a_9540_11106# cap_shunt_p a_11256_11044# vss nmos_6p0 w=0.82u l=0.6u
X11425 vdd a_33612_16055# a_33524_16152# vdd pmos_6p0 w=1.22u l=1u
X11426 a_11460_44756# cap_shunt_n a_11668_45240# vdd pmos_6p0 w=1.2u l=0.5u
X11427 a_24660_14242# cap_series_gyn a_24452_14588# vdd pmos_6p0 w=1.2u l=0.5u
X11428 a_30616_19668# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11429 vdd a_2140_41143# a_2052_41240# vdd pmos_6p0 w=1.22u l=1u
X11430 vdd a_34060_39575# a_33972_39672# vdd pmos_6p0 w=1.22u l=1u
X11431 vss tune_shunt[7] a_13796_22082# vss nmos_6p0 w=0.51u l=0.6u
X11432 a_5152_20152# cap_shunt_p a_3828_20152# vss nmos_6p0 w=0.82u l=0.6u
X11433 a_20172_23895# a_20084_23992# vss vss nmos_6p0 w=0.82u l=1u
X11434 a_30408_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11435 vss tune_series_gy[4] a_15700_9538# vss nmos_6p0 w=0.51u l=0.6u
X11436 a_9876_49944# cap_shunt_p a_9668_49460# vdd pmos_6p0 w=1.2u l=0.5u
X11437 a_23756_33736# a_23668_33780# vss vss nmos_6p0 w=0.82u l=1u
X11438 vdd tune_shunt[5] a_12580_49460# vdd pmos_6p0 w=1.2u l=0.5u
X11439 a_7748_45602# cap_shunt_p a_7540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X11440 vdd a_37644_32168# a_37556_32212# vdd pmos_6p0 w=1.22u l=1u
X11441 a_15904_22020# cap_shunt_n a_13796_22082# vss nmos_6p0 w=0.82u l=0.6u
X11442 vdd a_33612_12919# a_33524_13016# vdd pmos_6p0 w=1.22u l=1u
X11443 a_32632_11452# cap_series_gyp a_32444_11452# vdd pmos_6p0 w=1.2u l=0.5u
X11444 vdd tune_series_gygy[4] a_35692_10260# vdd pmos_6p0 w=1.2u l=0.5u
X11445 a_16700_11784# a_16612_11828# vss vss nmos_6p0 w=0.82u l=1u
X11446 a_34844_41143# a_34756_41240# vss vss nmos_6p0 w=0.82u l=1u
X11447 a_28692_6040# cap_shunt_n a_30408_6040# vss nmos_6p0 w=0.82u l=0.6u
X11448 a_9876_17016# cap_shunt_p a_9668_16532# vdd pmos_6p0 w=1.2u l=0.5u
X11449 vss tune_shunt[6] a_2708_39330# vss nmos_6p0 w=0.51u l=0.6u
X11450 a_21540_36540# cap_shunt_n a_21748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X11451 a_23756_30600# a_23668_30644# vss vss nmos_6p0 w=0.82u l=1u
X11452 a_9332_9884# cap_shunt_p a_9540_9538# vdd pmos_6p0 w=1.2u l=0.5u
X11453 a_4816_28292# cap_shunt_n a_2708_28354# vss nmos_6p0 w=0.82u l=0.6u
X11454 a_2500_9884# cap_shunt_n a_2708_9538# vdd pmos_6p0 w=1.2u l=0.5u
X11455 a_6516_20514# cap_shunt_p a_6308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X11456 a_5040_10744# cap_shunt_n a_2932_10744# vss nmos_6p0 w=0.82u l=0.6u
X11457 vdd a_3036_46280# a_2948_46324# vdd pmos_6p0 w=1.22u l=1u
X11458 a_17828_20152# cap_shunt_p a_17620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X11459 vdd a_36188_3511# a_36100_3608# vdd pmos_6p0 w=1.22u l=1u
X11460 a_37644_27464# a_37556_27508# vss vss nmos_6p0 w=0.82u l=1u
X11461 a_33948_8648# a_33860_8692# vss vss nmos_6p0 w=0.82u l=1u
X11462 a_17828_42104# cap_shunt_n a_17620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X11463 a_21540_33404# cap_shunt_n a_21748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X11464 vdd tune_shunt[7] a_29492_25564# vdd pmos_6p0 w=1.2u l=0.5u
X11465 a_24660_23650# cap_shunt_p a_24452_23996# vdd pmos_6p0 w=1.2u l=0.5u
X11466 vdd a_36636_52552# a_36548_52596# vdd pmos_6p0 w=1.22u l=1u
X11467 a_4816_25156# cap_shunt_p a_2708_25218# vss nmos_6p0 w=0.82u l=0.6u
X11468 vdd a_13564_55255# a_13476_55352# vdd pmos_6p0 w=1.22u l=1u
X11469 vdd a_35180_28599# a_35092_28696# vdd pmos_6p0 w=1.22u l=1u
X11470 a_1924_3266# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X11471 a_25572_7124# cap_series_gyn a_25780_7608# vdd pmos_6p0 w=1.2u l=0.5u
X11472 a_15492_8316# cap_series_gyn a_15700_7970# vdd pmos_6p0 w=1.2u l=0.5u
X11473 vdd tune_shunt[7] a_20532_18100# vdd pmos_6p0 w=1.2u l=0.5u
X11474 a_13588_49084# cap_shunt_n a_13796_48738# vdd pmos_6p0 w=1.2u l=0.5u
X11475 a_28236_48983# a_28148_49080# vss vss nmos_6p0 w=0.82u l=1u
X11476 vdd tune_shunt[7] a_33524_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11477 a_35692_13396# cap_series_gygyn a_35880_13396# vdd pmos_6p0 w=1.2u l=0.5u
X11478 vdd a_13564_52119# a_13476_52216# vdd pmos_6p0 w=1.22u l=1u
X11479 a_6532_41620# cap_shunt_n a_6740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X11480 a_21748_11106# cap_series_gyn a_21540_11452# vdd pmos_6p0 w=1.2u l=0.5u
X11481 a_9332_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11482 a_7964_54120# a_7876_54164# vss vss nmos_6p0 w=0.82u l=1u
X11483 vdd a_16700_53687# a_16612_53784# vdd pmos_6p0 w=1.22u l=1u
X11484 a_15492_5180# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11485 a_9668_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11486 vdd tune_shunt[7] a_29492_28700# vdd pmos_6p0 w=1.2u l=0.5u
X11487 vdd a_14236_52552# a_14148_52596# vdd pmos_6p0 w=1.22u l=1u
X11488 a_3036_38440# a_2948_38484# vss vss nmos_6p0 w=0.82u l=1u
X11489 a_29720_16156# cap_series_gyn a_30528_15748# vss nmos_6p0 w=0.82u l=0.6u
X11490 a_3640_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11491 a_6760_7124# cap_series_gyp a_6572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X11492 a_26768_12612# cap_series_gyn a_24660_12674# vss nmos_6p0 w=0.82u l=0.6u
X11493 vdd a_10988_44712# a_10900_44756# vdd pmos_6p0 w=1.22u l=1u
X11494 vss cap_shunt_n a_5152_37400# vss nmos_6p0 w=0.82u l=0.6u
X11495 a_6532_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11496 a_21428_5556# cap_series_gyp a_21636_6040# vdd pmos_6p0 w=1.2u l=0.5u
X11497 a_13588_50652# cap_shunt_p a_13796_50306# vdd pmos_6p0 w=1.2u l=0.5u
X11498 vdd a_27452_45847# a_27364_45944# vdd pmos_6p0 w=1.22u l=1u
X11499 vss tune_shunt[6] a_24660_37762# vss nmos_6p0 w=0.51u l=0.6u
X11500 a_20740_37400# cap_shunt_n a_20532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X11501 vss cap_shunt_n a_8848_35832# vss nmos_6p0 w=0.82u l=0.6u
X11502 a_34480_46325# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X11503 a_3640_42404# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11504 a_14372_40052# cap_shunt_n a_14580_40536# vdd pmos_6p0 w=1.2u l=0.5u
X11505 a_3828_32696# cap_shunt_p a_3620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X11506 a_31624_20860# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11507 a_3484_52552# a_3396_52596# vss vss nmos_6p0 w=0.82u l=1u
X11508 a_24204_36872# a_24116_36916# vss vss nmos_6p0 w=0.82u l=1u
X11509 a_14012_8215# a_13924_8312# vss vss nmos_6p0 w=0.82u l=1u
X11510 a_9108_49084# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11511 a_23084_55688# a_22996_55732# vss vss nmos_6p0 w=0.82u l=1u
X11512 a_13384_45240# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11513 vss tune_shunt[6] a_24660_34626# vss nmos_6p0 w=0.51u l=0.6u
X11514 vss tune_shunt[4] a_2708_12674# vss nmos_6p0 w=0.51u l=0.6u
X11515 a_21540_14588# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11516 a_11592_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11517 vdd a_27340_54120# a_27252_54164# vdd pmos_6p0 w=1.22u l=1u
X11518 a_1716_3988# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11519 a_22972_49416# a_22884_49460# vss vss nmos_6p0 w=0.82u l=1u
X11520 a_7748_39330# cap_shunt_n a_7540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X11521 a_13384_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11522 a_24452_39676# cap_shunt_p a_24660_39330# vdd pmos_6p0 w=1.2u l=0.5u
X11523 vss tune_shunt[3] a_5844_10744# vss nmos_6p0 w=0.51u l=0.6u
X11524 a_35880_13396# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11525 a_16500_45948# cap_shunt_p a_16708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X11526 a_19524_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11527 a_11984_20152# cap_shunt_p a_9876_20152# vss nmos_6p0 w=0.82u l=0.6u
X11528 vdd a_27340_50984# a_27252_51028# vdd pmos_6p0 w=1.22u l=1u
X11529 vss cap_shunt_p a_10640_22020# vss nmos_6p0 w=0.82u l=0.6u
X11530 a_2724_11828# cap_shunt_n a_2932_12312# vdd pmos_6p0 w=1.2u l=0.5u
X11531 a_6292_18946# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11532 vdd a_24316_54120# a_24228_54164# vdd pmos_6p0 w=1.22u l=1u
X11533 a_24660_42466# cap_shunt_n a_26376_42404# vss nmos_6p0 w=0.82u l=0.6u
X11534 vss cap_shunt_p a_27552_3204# vss nmos_6p0 w=0.82u l=0.6u
X11535 vdd a_28572_34871# a_28484_34968# vdd pmos_6p0 w=1.22u l=1u
X11536 a_10548_34264# cap_shunt_n a_10340_33780# vdd pmos_6p0 w=1.2u l=0.5u
X11537 a_35880_10260# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11538 a_15020_54120# a_14932_54164# vss vss nmos_6p0 w=0.82u l=1u
X11539 a_25592_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11540 a_35292_55255# a_35204_55352# vss vss nmos_6p0 w=0.82u l=1u
X11541 a_21540_27132# cap_shunt_n a_21748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X11542 a_29720_13020# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11543 vss tune_shunt[6] a_11668_46808# vss nmos_6p0 w=0.51u l=0.6u
X11544 vdd a_24316_50984# a_24228_51028# vdd pmos_6p0 w=1.22u l=1u
X11545 a_37632_47512# cap_shunt_gyp a_37444_47512# vdd pmos_6p0 w=1.215u l=0.5u
X11546 vss cap_shunt_p a_27104_35832# vss nmos_6p0 w=0.82u l=0.6u
X11547 a_10548_31128# cap_shunt_n a_10340_30644# vdd pmos_6p0 w=1.2u l=0.5u
X11548 a_4032_7908# cap_shunt_n a_1924_7970# vss nmos_6p0 w=0.82u l=0.6u
X11549 a_35448_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11550 a_25572_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11551 a_25592_40836# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11552 a_17828_32696# cap_shunt_n a_17620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X11553 a_24660_14242# cap_series_gyn a_24452_14588# vdd pmos_6p0 w=1.2u l=0.5u
X11554 a_18940_52119# a_18852_52216# vss vss nmos_6p0 w=0.82u l=1u
X11555 a_9876_53080# cap_shunt_n a_11592_53080# vss nmos_6p0 w=0.82u l=0.6u
X11556 a_9876_49944# cap_shunt_p a_9668_49460# vdd pmos_6p0 w=1.2u l=0.5u
X11557 a_12788_13880# cap_shunt_p a_14504_13880# vss nmos_6p0 w=0.82u l=0.6u
X11558 a_7748_45602# cap_shunt_p a_7540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X11559 a_25572_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11560 a_29492_28700# cap_shunt_p a_29700_28354# vdd pmos_6p0 w=1.2u l=0.5u
X11561 vss tune_series_gy[4] a_29720_16156# vss nmos_6p0 w=0.51u l=0.6u
X11562 a_6532_32212# cap_shunt_n a_6740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X11563 a_17148_53687# a_17060_53784# vss vss nmos_6p0 w=0.82u l=1u
X11564 vdd a_23308_47415# a_23220_47512# vdd pmos_6p0 w=1.22u l=1u
X11565 vdd a_36188_38440# a_36100_38484# vdd pmos_6p0 w=1.22u l=1u
X11566 a_13588_44380# cap_shunt_n a_13796_44034# vdd pmos_6p0 w=1.2u l=0.5u
X11567 a_6508_5079# a_6420_5176# vss vss nmos_6p0 w=0.82u l=1u
X11568 a_11668_46808# cap_shunt_n a_12600_46808# vss nmos_6p0 w=0.82u l=0.6u
X11569 vdd tune_shunt[6] a_10452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X11570 a_9856_37700# cap_shunt_n a_7748_37762# vss nmos_6p0 w=0.82u l=0.6u
X11571 vss cap_shunt_n a_34720_32996# vss nmos_6p0 w=0.82u l=0.6u
X11572 vss cap_shunt_n a_8848_29560# vss nmos_6p0 w=0.82u l=0.6u
X11573 a_14484_7124# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11574 a_7768_5180# cap_series_gyn a_8576_4772# vss nmos_6p0 w=0.82u l=0.6u
X11575 a_7852_55255# a_7764_55352# vss vss nmos_6p0 w=0.82u l=1u
X11576 a_7540_23996# cap_shunt_p a_7748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X11577 a_3640_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11578 a_6956_30167# a_6868_30264# vss vss nmos_6p0 w=0.82u l=1u
X11579 vdd a_23756_36872# a_23668_36916# vdd pmos_6p0 w=1.22u l=1u
X11580 a_19276_22327# a_19188_22424# vss vss nmos_6p0 w=0.82u l=1u
X11581 vdd tune_shunt[4] a_32404_36540# vdd pmos_6p0 w=1.2u l=0.5u
X11582 a_6532_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11583 a_15512_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11584 a_13588_41244# cap_shunt_n a_13796_40898# vdd pmos_6p0 w=1.2u l=0.5u
X11585 vss tune_shunt[7] a_6740_32696# vss nmos_6p0 w=0.51u l=0.6u
X11586 vdd tune_shunt[7] a_9668_18100# vdd pmos_6p0 w=1.2u l=0.5u
X11587 vss cap_shunt_n a_8848_26424# vss nmos_6p0 w=0.82u l=0.6u
X11588 vdd tune_shunt[6] a_10452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X11589 vss tune_shunt[7] a_24660_28354# vss nmos_6p0 w=0.51u l=0.6u
X11590 a_20740_27992# cap_shunt_n a_20532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X11591 vss cap_shunt_p a_23856_22020# vss nmos_6p0 w=0.82u l=0.6u
X11592 a_37420_47848# a_37332_47892# vss vss nmos_6p0 w=0.82u l=1u
X11593 a_2140_47415# a_2052_47512# vss vss nmos_6p0 w=0.82u l=1u
X11594 vdd a_35628_36439# a_35540_36536# vdd pmos_6p0 w=1.22u l=1u
X11595 a_6956_27031# a_6868_27128# vss vss nmos_6p0 w=0.82u l=1u
X11596 a_6532_13396# cap_shunt_p a_6740_13880# vdd pmos_6p0 w=1.2u l=0.5u
X11597 a_6516_20514# cap_shunt_p a_7448_20452# vss nmos_6p0 w=0.82u l=0.6u
X11598 a_4828_55255# a_4740_55352# vss vss nmos_6p0 w=0.82u l=1u
X11599 a_9540_9538# cap_shunt_p a_10472_9476# vss nmos_6p0 w=0.82u l=0.6u
X11600 vdd tune_shunt[4] a_32404_33404# vdd pmos_6p0 w=1.2u l=0.5u
X11601 a_25780_7608# cap_series_gyn a_27496_7608# vss nmos_6p0 w=0.82u l=0.6u
X11602 a_8412_10216# a_8324_10260# vss vss nmos_6p0 w=0.82u l=1u
X11603 a_17596_54120# a_17508_54164# vss vss nmos_6p0 w=0.82u l=1u
X11604 a_6532_41620# cap_shunt_n a_6740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X11605 a_16500_39676# cap_shunt_n a_16708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X11606 a_9668_21236# cap_shunt_p a_9876_21720# vdd pmos_6p0 w=1.2u l=0.5u
X11607 a_35040_43734# cap_shunt_gyp a_35040_43189# vdd pmos_6p0 w=1.215u l=0.5u
X11608 vss tune_shunt[7] a_24660_25218# vss nmos_6p0 w=0.51u l=0.6u
X11609 vdd a_31708_3944# a_31620_3988# vdd pmos_6p0 w=1.22u l=1u
X11610 a_9668_21236# cap_shunt_p a_9876_21720# vdd pmos_6p0 w=1.2u l=0.5u
X11611 a_20740_43672# cap_shunt_n a_22456_43672# vss nmos_6p0 w=0.82u l=0.6u
X11612 a_11612_7124# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11613 a_2708_17378# cap_shunt_p a_2500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11614 a_24452_13020# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11615 a_24660_36194# cap_shunt_p a_26376_36132# vss nmos_6p0 w=0.82u l=0.6u
X11616 a_23072_20452# cap_shunt_p a_21748_20514# vss nmos_6p0 w=0.82u l=0.6u
X11617 vdd tune_shunt[4] a_33524_33780# vdd pmos_6p0 w=1.2u l=0.5u
X11618 vdd a_28572_28599# a_28484_28696# vdd pmos_6p0 w=1.22u l=1u
X11619 a_29492_11452# cap_series_gyp a_29700_11106# vdd pmos_6p0 w=1.2u l=0.5u
X11620 a_25572_40052# cap_shunt_n a_25780_40536# vdd pmos_6p0 w=1.2u l=0.5u
X11621 a_24752_12312# cap_series_gyn a_22644_12312# vss nmos_6p0 w=0.82u l=0.6u
X11622 a_20740_40536# cap_shunt_p a_22456_40536# vss nmos_6p0 w=0.82u l=0.6u
X11623 a_34516_17378# cap_series_gygyn a_34308_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11624 vdd a_33500_19624# a_33412_19668# vdd pmos_6p0 w=1.22u l=1u
X11625 a_13588_50652# cap_shunt_p a_13796_50306# vdd pmos_6p0 w=1.2u l=0.5u
X11626 a_13496_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X11627 a_20740_37400# cap_shunt_n a_20532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X11628 vss cap_shunt_p a_27104_29560# vss nmos_6p0 w=0.82u l=0.6u
X11629 a_10548_24856# cap_shunt_n a_10340_24372# vdd pmos_6p0 w=1.2u l=0.5u
X11630 a_10452_5180# cap_series_gyp a_10660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X11631 vdd tune_shunt[4] a_33524_30644# vdd pmos_6p0 w=1.2u l=0.5u
X11632 a_35448_29560# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11633 a_14372_40052# cap_shunt_n a_14580_40536# vdd pmos_6p0 w=1.2u l=0.5u
X11634 a_25572_3988# cap_shunt_p a_25780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X11635 a_25592_34564# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11636 a_2708_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11637 vss tune_series_gygy[5] a_34516_22082# vss nmos_6p0 w=0.51u l=0.6u
X11638 vdd tune_shunt[7] a_6532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X11639 a_3828_15448# cap_shunt_p a_3620_14964# vdd pmos_6p0 w=1.2u l=0.5u
X11640 a_6292_50306# cap_shunt_p a_7224_50244# vss nmos_6p0 w=0.82u l=0.6u
X11641 vss cap_shunt_p a_27104_26424# vss nmos_6p0 w=0.82u l=0.6u
X11642 vdd a_20732_53687# a_20644_53784# vdd pmos_6p0 w=1.22u l=1u
X11643 a_21748_9538# cap_series_gyp a_21540_9884# vdd pmos_6p0 w=1.2u l=0.5u
X11644 a_17620_18100# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11645 vdd a_6956_8215# a_6868_8312# vdd pmos_6p0 w=1.22u l=1u
X11646 a_25572_16532# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11647 a_20532_44756# cap_shunt_n a_20740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X11648 a_7748_39330# cap_shunt_n a_7540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X11649 a_32824_20452# cap_series_gygyn a_31624_20860# vss nmos_6p0 w=0.82u l=0.6u
X11650 a_25592_31428# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11651 a_7672_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11652 a_31260_36872# a_31172_36916# vss vss nmos_6p0 w=0.82u l=1u
X11653 vdd tune_shunt[7] a_6532_11828# vdd pmos_6p0 w=1.2u l=0.5u
X11654 a_5612_20759# a_5524_20856# vss vss nmos_6p0 w=0.82u l=1u
X11655 a_16500_45948# cap_shunt_p a_16708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X11656 a_21748_6402# cap_series_gyn a_21540_6748# vdd pmos_6p0 w=1.2u l=0.5u
X11657 vdd a_3484_55688# a_3396_55732# vdd pmos_6p0 w=1.22u l=1u
X11658 a_6060_44279# a_5972_44376# vss vss nmos_6p0 w=0.82u l=1u
X11659 a_36384_43972# tune_shunt_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X11660 a_37868_38007# a_37780_38104# vss vss nmos_6p0 w=0.82u l=1u
X11661 vss tune_shunt[7] a_17828_20152# vss nmos_6p0 w=0.51u l=0.6u
X11662 vss cap_shunt_n a_22848_38968# vss nmos_6p0 w=0.82u l=0.6u
X11663 a_4424_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11664 a_6060_41143# a_5972_41240# vss vss nmos_6p0 w=0.82u l=1u
X11665 a_36384_40836# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11666 a_5936_35832# cap_shunt_n a_3828_35832# vss nmos_6p0 w=0.82u l=0.6u
X11667 a_16708_23650# cap_shunt_n a_16500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X11668 a_15356_19624# a_15268_19668# vss vss nmos_6p0 w=0.82u l=1u
X11669 vdd a_31372_54120# a_31284_54164# vdd pmos_6p0 w=1.22u l=1u
X11670 a_37532_52552# a_37444_52596# vss vss nmos_6p0 w=0.82u l=1u
X11671 vdd a_23756_27464# a_23668_27508# vdd pmos_6p0 w=1.22u l=1u
X11672 vdd tune_shunt[7] a_32404_27132# vdd pmos_6p0 w=1.2u l=0.5u
X11673 a_4424_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11674 a_15512_23588# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11675 a_6084_18100# cap_shunt_p a_6292_18584# vdd pmos_6p0 w=1.2u l=0.5u
X11676 vss tune_shunt[7] a_6740_23288# vss nmos_6p0 w=0.51u l=0.6u
X11677 a_10988_3944# a_10900_3988# vss vss nmos_6p0 w=0.82u l=1u
X11678 vss cap_series_gyn a_16800_9176# vss nmos_6p0 w=0.82u l=0.6u
X11679 vdd a_30812_55255# a_30724_55352# vdd pmos_6p0 w=1.22u l=1u
X11680 vdd a_35628_27031# a_35540_27128# vdd pmos_6p0 w=1.22u l=1u
X11681 a_28684_55255# a_28596_55352# vss vss nmos_6p0 w=0.82u l=1u
X11682 vdd a_31372_50984# a_31284_51028# vdd pmos_6p0 w=1.22u l=1u
X11683 a_9876_49944# cap_shunt_p a_9668_49460# vdd pmos_6p0 w=1.2u l=0.5u
X11684 vss cap_shunt_p a_18816_43972# vss nmos_6p0 w=0.82u l=0.6u
X11685 vss tune_series_gy[5] a_28692_13880# vss nmos_6p0 w=0.51u l=0.6u
X11686 a_23072_14180# cap_series_gyn a_21748_14242# vss nmos_6p0 w=0.82u l=0.6u
X11687 a_16016_4472# cap_series_gyp a_14692_4472# vss nmos_6p0 w=0.82u l=0.6u
X11688 a_6532_32212# cap_shunt_n a_6740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X11689 a_24660_7970# cap_series_gyp a_24452_8316# vdd pmos_6p0 w=1.2u l=0.5u
X11690 vdd a_30812_52119# a_30724_52216# vdd pmos_6p0 w=1.22u l=1u
X11691 a_8456_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11692 a_24660_7970# cap_series_gyp a_26376_7908# vss nmos_6p0 w=0.82u l=0.6u
X11693 a_20740_34264# cap_shunt_n a_22456_34264# vss nmos_6p0 w=0.82u l=0.6u
X11694 a_19732_7608# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11695 a_15132_52552# a_15044_52596# vss vss nmos_6p0 w=0.82u l=1u
X11696 vss cap_shunt_n a_18816_40836# vss nmos_6p0 w=0.82u l=0.6u
X11697 a_13588_44380# cap_shunt_n a_13796_44034# vdd pmos_6p0 w=1.2u l=0.5u
X11698 vss tune_shunt[7] a_16708_31490# vss nmos_6p0 w=0.51u l=0.6u
X11699 vdd tune_series_gygy[0] a_31436_6748# vdd pmos_6p0 w=1.2u l=0.5u
X11700 a_12108_16055# a_12020_16152# vss vss nmos_6p0 w=0.82u l=1u
X11701 vdd a_19724_47415# a_19636_47512# vdd pmos_6p0 w=1.22u l=1u
X11702 a_2708_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11703 vss tune_shunt[3] a_5844_9538# vss nmos_6p0 w=0.51u l=0.6u
X11704 vss tune_series_gy[4] a_28692_10744# vss nmos_6p0 w=0.51u l=0.6u
X11705 a_23072_11044# cap_series_gyn a_21748_11106# vss nmos_6p0 w=0.82u l=0.6u
X11706 a_35840_12612# cap_series_gygyp a_34516_12674# vss nmos_6p0 w=0.82u l=0.6u
X11707 a_18044_13352# a_17956_13396# vss vss nmos_6p0 w=0.82u l=1u
X11708 vss tune_shunt[7] a_6628_14242# vss nmos_6p0 w=0.51u l=0.6u
X11709 vdd a_28572_19191# a_28484_19288# vdd pmos_6p0 w=1.22u l=1u
X11710 a_6740_37400# cap_shunt_n a_7672_37400# vss nmos_6p0 w=0.82u l=0.6u
X11711 a_29700_36194# cap_shunt_n a_29492_36540# vdd pmos_6p0 w=1.2u l=0.5u
X11712 vss cap_shunt_p a_7168_10744# vss nmos_6p0 w=0.82u l=0.6u
X11713 a_35264_45540# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11714 a_25592_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11715 a_20740_31128# cap_shunt_n a_22456_31128# vss nmos_6p0 w=0.82u l=0.6u
X11716 a_1692_38007# a_1604_38104# vss vss nmos_6p0 w=0.82u l=1u
X11717 a_2708_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11718 vdd a_3932_54120# a_3844_54164# vdd pmos_6p0 w=1.22u l=1u
X11719 vdd a_30364_47415# a_30276_47512# vdd pmos_6p0 w=1.22u l=1u
X11720 a_13588_41244# cap_shunt_n a_13796_40898# vdd pmos_6p0 w=1.2u l=0.5u
X11721 a_34516_4834# cap_series_gygyp a_35448_4772# vss nmos_6p0 w=0.82u l=0.6u
X11722 a_20740_27992# cap_shunt_n a_20532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X11723 a_18044_10216# a_17956_10260# vss vss nmos_6p0 w=0.82u l=1u
X11724 a_30616_19668# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11725 a_21672_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11726 a_7768_8316# cap_series_gyn a_7580_8316# vdd pmos_6p0 w=1.2u l=0.5u
X11727 a_35880_10260# cap_series_gygyp a_35692_10260# vdd pmos_6p0 w=1.2u l=0.5u
X11728 a_20532_38484# cap_shunt_n a_20740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X11729 a_32632_14588# cap_series_gyp a_32656_14180# vss nmos_6p0 w=0.82u l=0.6u
X11730 a_12580_14964# cap_shunt_p a_12788_15448# vdd pmos_6p0 w=1.2u l=0.5u
X11731 a_35264_42404# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11732 a_29700_33058# cap_shunt_p a_29492_33404# vdd pmos_6p0 w=1.2u l=0.5u
X11733 a_25592_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11734 a_12376_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X11735 a_18404_3988# cap_series_gyp a_18612_4472# vdd pmos_6p0 w=1.2u l=0.5u
X11736 a_15904_45240# cap_shunt_p a_14580_45240# vss nmos_6p0 w=0.82u l=0.6u
X11737 a_27104_42104# cap_shunt_n a_25780_42104# vss nmos_6p0 w=0.82u l=0.6u
X11738 a_25780_9176# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11739 a_11772_52119# a_11684_52216# vss vss nmos_6p0 w=0.82u l=1u
X11740 a_32268_39575# a_32180_39672# vss vss nmos_6p0 w=0.82u l=1u
X11741 a_2708_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11742 a_6532_41620# cap_shunt_n a_6740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X11743 a_16500_39676# cap_shunt_n a_16708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X11744 a_5612_14487# a_5524_14584# vss vss nmos_6p0 w=0.82u l=1u
X11745 vss cap_series_gyp a_27104_17016# vss nmos_6p0 w=0.82u l=0.6u
X11746 a_2708_17378# cap_shunt_p a_2500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11747 a_6292_51512# cap_shunt_p a_6084_51028# vdd pmos_6p0 w=1.2u l=0.5u
X11748 vdd a_10092_43144# a_10004_43188# vdd pmos_6p0 w=1.22u l=1u
X11749 a_32632_11452# cap_series_gyp a_32656_11044# vss nmos_6p0 w=0.82u l=0.6u
X11750 a_20532_35348# cap_shunt_n a_20740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X11751 a_12580_11828# cap_shunt_p a_12788_12312# vdd pmos_6p0 w=1.2u l=0.5u
X11752 a_15904_42104# cap_shunt_n a_14580_42104# vss nmos_6p0 w=0.82u l=0.6u
X11753 vdd a_27228_31735# a_27140_31832# vdd pmos_6p0 w=1.22u l=1u
X11754 a_10808_51512# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11755 a_13252_36916# cap_shunt_n a_13460_37400# vdd pmos_6p0 w=1.2u l=0.5u
X11756 a_29492_11452# cap_series_gyp a_29700_11106# vdd pmos_6p0 w=1.2u l=0.5u
X11757 a_21748_33058# cap_shunt_n a_23464_32996# vss nmos_6p0 w=0.82u l=0.6u
X11758 a_13588_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11759 vdd a_33500_42711# a_33412_42808# vdd pmos_6p0 w=1.22u l=1u
X11760 a_3620_36916# cap_shunt_n a_3828_37400# vdd pmos_6p0 w=1.2u l=0.5u
X11761 a_6060_34871# a_5972_34968# vss vss nmos_6p0 w=0.82u l=1u
X11762 a_5936_29560# cap_shunt_n a_3828_29560# vss nmos_6p0 w=0.82u l=0.6u
X11763 a_22644_7608# cap_series_gyp a_22436_7124# vdd pmos_6p0 w=1.2u l=0.5u
X11764 a_34516_17378# cap_series_gygyn a_34308_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11765 a_9644_44712# a_9556_44756# vss vss nmos_6p0 w=0.82u l=1u
X11766 vdd tune_shunt[6] a_6532_47892# vdd pmos_6p0 w=1.2u l=0.5u
X11767 a_28692_40536# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11768 a_6084_52220# cap_shunt_p a_6292_51874# vdd pmos_6p0 w=1.2u l=0.5u
X11769 a_19544_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11770 a_29492_36540# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11771 vss cap_series_gyn a_30136_12612# vss nmos_6p0 w=0.82u l=0.6u
X11772 vdd a_31708_13352# a_31620_13396# vdd pmos_6p0 w=1.22u l=1u
X11773 vdd a_9868_53687# a_9780_53784# vdd pmos_6p0 w=1.22u l=1u
X11774 a_5936_26424# cap_shunt_p a_3828_26424# vss nmos_6p0 w=0.82u l=0.6u
X11775 vdd a_37420_9783# a_37332_9880# vdd pmos_6p0 w=1.22u l=1u
X11776 a_16708_14242# cap_shunt_p a_16500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X11777 a_28692_35832# cap_shunt_p a_29624_35832# vss nmos_6p0 w=0.82u l=0.6u
X11778 a_6060_31735# a_5972_31832# vss vss nmos_6p0 w=0.82u l=1u
X11779 vdd a_2588_18056# a_2500_18100# vdd pmos_6p0 w=1.22u l=1u
X11780 a_9644_41576# a_9556_41620# vss vss nmos_6p0 w=0.82u l=1u
X11781 vss cap_shunt_p a_30016_37400# vss nmos_6p0 w=0.82u l=0.6u
X11782 vdd a_30812_48983# a_30724_49080# vdd pmos_6p0 w=1.22u l=1u
X11783 a_7728_47108# cap_shunt_p a_6404_47170# vss nmos_6p0 w=0.82u l=0.6u
X11784 a_32464_46870# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11785 vdd tune_shunt[6] a_6532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X11786 a_35188_43972# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X11787 a_29492_33404# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11788 a_28684_48983# a_28596_49080# vss vss nmos_6p0 w=0.82u l=1u
X11789 a_20532_44756# cap_shunt_n a_20740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X11790 a_2708_29922# cap_shunt_n a_3640_29860# vss nmos_6p0 w=0.82u l=0.6u
X11791 vdd a_37420_6647# a_37332_6744# vdd pmos_6p0 w=1.22u l=1u
X11792 vdd a_10988_55255# a_10900_55352# vdd pmos_6p0 w=1.22u l=1u
X11793 vdd a_36188_55255# a_36100_55352# vdd pmos_6p0 w=1.22u l=1u
X11794 vdd a_13452_3511# a_13364_3608# vdd pmos_6p0 w=1.22u l=1u
X11795 a_37420_53687# a_37332_53784# vss vss nmos_6p0 w=0.82u l=1u
X11796 vdd tune_shunt[3] a_25572_43188# vdd pmos_6p0 w=1.2u l=0.5u
X11797 vss cap_shunt_n a_8064_32696# vss nmos_6p0 w=0.82u l=0.6u
X11798 a_34308_22428# cap_series_gygyp a_34516_22082# vdd pmos_6p0 w=1.2u l=0.5u
X11799 a_35488_42166# cap_shunt_gyn a_35488_41621# vdd pmos_6p0 w=1.215u l=0.5u
X11800 a_5636_9884# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11801 a_31436_20860# cap_series_gygyn a_31624_20860# vdd pmos_6p0 w=1.2u l=0.5u
X11802 vdd a_14684_52552# a_14596_52596# vdd pmos_6p0 w=1.22u l=1u
X11803 vss cap_shunt_p a_8400_51512# vss nmos_6p0 w=0.82u l=0.6u
X11804 vss cap_shunt_n a_18816_34564# vss nmos_6p0 w=0.82u l=0.6u
X11805 a_16708_17378# cap_shunt_p a_16500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X11806 a_2708_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11807 a_2708_26786# cap_shunt_p a_3640_26724# vss nmos_6p0 w=0.82u l=0.6u
X11808 vdd a_37420_3511# a_37332_3608# vdd pmos_6p0 w=1.22u l=1u
X11809 a_7748_39330# cap_shunt_n a_8680_39268# vss nmos_6p0 w=0.82u l=0.6u
X11810 a_2500_34972# cap_shunt_n a_2708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X11811 a_30800_32696# cap_shunt_p a_28692_32696# vss nmos_6p0 w=0.82u l=0.6u
X11812 vdd a_36188_52119# a_36100_52216# vdd pmos_6p0 w=1.22u l=1u
X11813 a_11668_43672# cap_shunt_n a_11460_43188# vdd pmos_6p0 w=1.2u l=0.5u
X11814 a_15568_35832# cap_shunt_n a_13460_35832# vss nmos_6p0 w=0.82u l=0.6u
X11815 vdd a_29468_8215# a_29380_8312# vdd pmos_6p0 w=1.22u l=1u
X11816 vss tune_shunt[7] a_9540_9538# vss nmos_6p0 w=0.51u l=0.6u
X11817 a_20740_46808# cap_shunt_p a_21672_46808# vss nmos_6p0 w=0.82u l=0.6u
X11818 vss cap_shunt_n a_18816_31428# vss nmos_6p0 w=0.82u l=0.6u
X11819 a_17828_27992# cap_shunt_n a_19544_27992# vss nmos_6p0 w=0.82u l=0.6u
X11820 a_27888_27992# cap_shunt_p a_25780_27992# vss nmos_6p0 w=0.82u l=0.6u
X11821 vss tune_shunt[7] a_16708_22082# vss nmos_6p0 w=0.51u l=0.6u
X11822 a_31624_20860# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11823 vdd a_19724_38007# a_19636_38104# vdd pmos_6p0 w=1.22u l=1u
X11824 a_24652_36872# a_24564_36916# vss vss nmos_6p0 w=0.82u l=1u
X11825 a_2500_31836# cap_shunt_p a_2708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X11826 vdd a_2140_40008# a_2052_40052# vdd pmos_6p0 w=1.22u l=1u
X11827 a_29700_26786# cap_shunt_p a_29492_27132# vdd pmos_6p0 w=1.2u l=0.5u
X11828 a_35880_8692# cap_series_gygyn a_35692_8692# vdd pmos_6p0 w=1.2u l=0.5u
X11829 a_11032_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11830 a_6084_18100# cap_shunt_p a_6292_18584# vdd pmos_6p0 w=1.2u l=0.5u
X11831 a_17828_24856# cap_shunt_n a_19544_24856# vss nmos_6p0 w=0.82u l=0.6u
X11832 a_27888_24856# cap_shunt_p a_25780_24856# vss nmos_6p0 w=0.82u l=0.6u
X11833 a_19724_19191# a_19636_19288# vss vss nmos_6p0 w=0.82u l=1u
X11834 a_21672_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11835 vdd a_8748_55255# a_8660_55352# vdd pmos_6p0 w=1.22u l=1u
X11836 vss tune_shunt[6] a_16708_42466# vss nmos_6p0 w=0.51u l=0.6u
X11837 a_20532_29076# cap_shunt_n a_20740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X11838 a_11572_5556# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11839 a_35880_5556# cap_series_gygyn a_35692_5556# vdd pmos_6p0 w=1.2u l=0.5u
X11840 vdd a_27228_25463# a_27140_25560# vdd pmos_6p0 w=1.22u l=1u
X11841 a_17596_7080# a_17508_7124# vss vss nmos_6p0 w=0.82u l=1u
X11842 a_35880_8692# cap_series_gygyn a_36688_9176# vss nmos_6p0 w=0.82u l=0.6u
X11843 a_10660_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11844 a_29624_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X11845 a_30364_19191# a_30276_19288# vss vss nmos_6p0 w=0.82u l=1u
X11846 a_34844_54120# a_34756_54164# vss vss nmos_6p0 w=0.82u l=1u
X11847 a_17620_40052# cap_shunt_n a_17828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X11848 a_6532_32212# cap_shunt_n a_6740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X11849 vss tune_shunt[1] a_25444_3266# vss nmos_6p0 w=0.51u l=0.6u
X11850 vdd a_24764_54120# a_24676_54164# vdd pmos_6p0 w=1.22u l=1u
X11851 a_19724_16055# a_19636_16152# vss vss nmos_6p0 w=0.82u l=1u
X11852 a_35040_44757# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X11853 a_10548_37400# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11854 a_6060_28599# a_5972_28696# vss vss nmos_6p0 w=0.82u l=1u
X11855 a_7560_14180# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11856 vss cap_shunt_p a_8512_47108# vss nmos_6p0 w=0.82u l=0.6u
X11857 a_28692_34264# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11858 a_35904_4472# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X11859 vdd a_27228_22327# a_27140_22424# vdd pmos_6p0 w=1.22u l=1u
X11860 a_10660_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11861 a_13252_27508# cap_shunt_n a_13460_27992# vdd pmos_6p0 w=1.2u l=0.5u
X11862 a_29720_13020# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X11863 vss cap_shunt_n a_13776_43672# vss nmos_6p0 w=0.82u l=0.6u
X11864 a_2140_32168# a_2052_32212# vss vss nmos_6p0 w=0.82u l=1u
X11865 a_21748_23650# cap_shunt_p a_23464_23588# vss nmos_6p0 w=0.82u l=0.6u
X11866 vdd tune_series_gy[3] a_21316_3988# vdd pmos_6p0 w=1.2u l=0.5u
X11867 vdd a_24764_50984# a_24676_51028# vdd pmos_6p0 w=1.22u l=1u
X11868 a_29700_36194# cap_shunt_n a_29492_36540# vdd pmos_6p0 w=1.2u l=0.5u
X11869 a_33948_25896# a_33860_25940# vss vss nmos_6p0 w=0.82u l=1u
X11870 vss cap_shunt_n a_10528_51812# vss nmos_6p0 w=0.82u l=0.6u
X11871 vdd tune_shunt[6] a_21540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X11872 a_28692_29560# cap_shunt_p a_29624_29560# vss nmos_6p0 w=0.82u l=0.6u
X11873 a_3620_27508# cap_shunt_n a_3828_27992# vdd pmos_6p0 w=1.2u l=0.5u
X11874 a_6060_25463# a_5972_25560# vss vss nmos_6p0 w=0.82u l=1u
X11875 a_7560_11044# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X11876 a_34396_49416# a_34308_49460# vss vss nmos_6p0 w=0.82u l=1u
X11877 a_12768_45540# cap_shunt_n a_10660_45602# vss nmos_6p0 w=0.82u l=0.6u
X11878 a_4312_49944# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11879 a_7748_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11880 vdd tune_shunt[6] a_6532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X11881 a_28692_31128# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X11882 a_34308_19292# cap_series_gygyn a_34516_18946# vdd pmos_6p0 w=1.2u l=0.5u
X11883 vss cap_shunt_p a_19152_20152# vss nmos_6p0 w=0.82u l=0.6u
X11884 a_29492_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11885 vss cap_shunt_n a_13776_40536# vss nmos_6p0 w=0.82u l=0.6u
X11886 a_9876_21720# cap_shunt_p a_10808_21720# vss nmos_6p0 w=0.82u l=0.6u
X11887 a_20532_38484# cap_shunt_n a_20740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X11888 a_29700_33058# cap_shunt_p a_29492_33404# vdd pmos_6p0 w=1.2u l=0.5u
X11889 a_12580_14964# cap_shunt_p a_12788_15448# vdd pmos_6p0 w=1.2u l=0.5u
X11890 vdd tune_shunt[7] a_21540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X11891 a_28692_26424# cap_shunt_p a_29624_26424# vss nmos_6p0 w=0.82u l=0.6u
X11892 a_12768_42404# cap_shunt_n a_10660_42466# vss nmos_6p0 w=0.82u l=0.6u
X11893 vdd tune_shunt[6] a_6532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X11894 vdd a_34396_10216# a_34308_10260# vdd pmos_6p0 w=1.22u l=1u
X11895 a_34308_16156# cap_series_gygyn a_34516_15810# vdd pmos_6p0 w=1.2u l=0.5u
X11896 a_9668_51028# cap_shunt_n a_9876_51512# vdd pmos_6p0 w=1.2u l=0.5u
X11897 vss cap_shunt_n a_18816_28292# vss nmos_6p0 w=0.82u l=0.6u
X11898 a_20532_35348# cap_shunt_n a_20740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X11899 a_12580_11828# cap_shunt_p a_12788_12312# vdd pmos_6p0 w=1.2u l=0.5u
X11900 a_21540_13020# cap_series_gyn a_21748_12674# vdd pmos_6p0 w=1.2u l=0.5u
X11901 a_17596_53687# a_17508_53784# vss vss nmos_6p0 w=0.82u l=1u
X11902 a_6508_45847# a_6420_45944# vss vss nmos_6p0 w=0.82u l=1u
X11903 vss tune_shunt[6] a_9876_49944# vss nmos_6p0 w=0.51u l=0.6u
X11904 vdd a_23756_47415# a_23668_47512# vdd pmos_6p0 w=1.22u l=1u
X11905 a_36384_41240# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X11906 a_13252_36916# cap_shunt_n a_13460_37400# vdd pmos_6p0 w=1.2u l=0.5u
X11907 a_29492_11452# cap_series_gyp a_29700_11106# vdd pmos_6p0 w=1.2u l=0.5u
X11908 a_15568_29560# cap_shunt_n a_13460_29560# vss nmos_6p0 w=0.82u l=0.6u
X11909 vss cap_shunt_p a_8064_23288# vss nmos_6p0 w=0.82u l=0.6u
X11910 vdd a_16252_47848# a_16164_47892# vdd pmos_6p0 w=1.22u l=1u
X11911 a_9316_47170# cap_shunt_p a_9108_47516# vdd pmos_6p0 w=1.2u l=0.5u
X11912 a_29492_39676# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11913 a_35880_13396# cap_series_gygyn a_35904_13880# vss nmos_6p0 w=0.82u l=0.6u
X11914 a_7748_34626# cap_shunt_n a_7540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X11915 vss cap_shunt_n a_18816_25156# vss nmos_6p0 w=0.82u l=0.6u
X11916 a_6532_13396# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11917 vdd a_24428_47848# a_24340_47892# vdd pmos_6p0 w=1.22u l=1u
X11918 a_34308_5180# tune_series_gygy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11919 a_6508_42711# a_6420_42808# vss vss nmos_6p0 w=0.82u l=1u
X11920 a_2500_25564# cap_shunt_p a_2708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X11921 a_2708_17378# cap_shunt_p a_3640_17316# vss nmos_6p0 w=0.82u l=0.6u
X11922 a_36384_47108# cap_shunt_gyp a_36384_47512# vdd pmos_6p0 w=1.215u l=0.5u
X11923 a_30800_23288# cap_shunt_p a_28692_23288# vss nmos_6p0 w=0.82u l=0.6u
X11924 a_6084_52220# cap_shunt_p a_6292_51874# vdd pmos_6p0 w=1.2u l=0.5u
X11925 a_21540_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11926 a_15568_26424# cap_shunt_n a_13460_26424# vss nmos_6p0 w=0.82u l=0.6u
X11927 vdd a_4940_8215# a_4852_8312# vdd pmos_6p0 w=1.22u l=1u
X11928 a_12788_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11929 vss cap_shunt_p a_31024_29860# vss nmos_6p0 w=0.82u l=0.6u
X11930 a_35880_10260# cap_series_gygyp a_35904_10744# vss nmos_6p0 w=0.82u l=0.6u
X11931 a_7748_31490# cap_shunt_n a_7540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X11932 a_17828_18584# cap_shunt_p a_19544_18584# vss nmos_6p0 w=0.82u l=0.6u
X11933 vss tune_shunt[7] a_21748_18946# vss nmos_6p0 w=0.51u l=0.6u
X11934 vss tune_series_gygy[1] a_31624_8316# vss nmos_6p0 w=0.51u l=0.6u
X11935 a_2500_22428# cap_shunt_p a_2708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X11936 a_8860_10216# a_8772_10260# vss vss nmos_6p0 w=0.82u l=1u
X11937 a_27888_18584# cap_series_gyn a_25780_18584# vss nmos_6p0 w=0.82u l=0.6u
X11938 vss tune_shunt[7] a_16708_36194# vss nmos_6p0 w=0.51u l=0.6u
X11939 a_20532_44756# cap_shunt_n a_20740_45240# vdd pmos_6p0 w=1.2u l=0.5u
X11940 a_27496_6040# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X11941 a_12788_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11942 vdd a_28124_44279# a_28036_44376# vdd pmos_6p0 w=1.22u l=1u
X11943 vss cap_shunt_p a_31024_26724# vss nmos_6p0 w=0.82u l=0.6u
X11944 a_17828_15448# cap_shunt_p a_19544_15448# vss nmos_6p0 w=0.82u l=0.6u
X11945 vdd a_15356_16488# a_15268_16532# vdd pmos_6p0 w=1.22u l=1u
X11946 a_2500_28700# cap_shunt_n a_2708_28354# vdd pmos_6p0 w=1.2u l=0.5u
X11947 a_9108_22428# cap_shunt_p a_9316_22082# vdd pmos_6p0 w=1.2u l=0.5u
X11948 a_4760_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X11949 a_34308_22428# cap_series_gygyp a_34516_22082# vdd pmos_6p0 w=1.2u l=0.5u
X11950 a_27888_15448# cap_series_gyp a_25780_15448# vss nmos_6p0 w=0.82u l=0.6u
X11951 a_28692_15448# cap_series_gyn a_28484_14964# vdd pmos_6p0 w=1.2u l=0.5u
X11952 a_31436_20860# cap_series_gygyn a_31624_20860# vdd pmos_6p0 w=1.2u l=0.5u
X11953 a_11324_55688# a_11236_55732# vss vss nmos_6p0 w=0.82u l=1u
X11954 vss tune_shunt[7] a_16708_33058# vss nmos_6p0 w=0.51u l=0.6u
X11955 a_16708_47170# cap_shunt_n a_16500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X11956 vdd a_10540_41576# a_10452_41620# vdd pmos_6p0 w=1.22u l=1u
X11957 a_6404_22082# cap_shunt_p a_6196_22428# vdd pmos_6p0 w=1.2u l=0.5u
X11958 vdd a_27228_16055# a_27140_16152# vdd pmos_6p0 w=1.22u l=1u
X11959 a_2500_34972# cap_shunt_n a_2708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X11960 a_11668_43672# cap_shunt_n a_11460_43188# vdd pmos_6p0 w=1.2u l=0.5u
X11961 a_10660_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11962 a_9668_10260# cap_shunt_p a_9876_10744# vdd pmos_6p0 w=1.2u l=0.5u
X11963 a_7540_38108# cap_shunt_n a_7748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X11964 a_35448_22020# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X11965 vdd a_6060_6647# a_5972_6744# vdd pmos_6p0 w=1.22u l=1u
X11966 vss cap_shunt_gyn a_36428_45240# vss nmos_6p0 w=0.82u l=0.6u
X11967 a_35736_9476# cap_series_gygyn a_34536_9884# vss nmos_6p0 w=0.82u l=0.6u
X11968 a_28692_12312# cap_series_gyn a_28484_11828# vdd pmos_6p0 w=1.2u l=0.5u
X11969 a_9876_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11970 a_7748_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X11971 a_1924_7608# cap_shunt_n a_3640_7608# vss nmos_6p0 w=0.82u l=0.6u
X11972 a_32156_11784# a_32068_11828# vss vss nmos_6p0 w=0.82u l=1u
X11973 vdd a_27228_12919# a_27140_13016# vdd pmos_6p0 w=1.22u l=1u
X11974 a_17828_48376# cap_shunt_p a_17620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X11975 a_2500_31836# cap_shunt_p a_2708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X11976 a_10660_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X11977 a_2140_22760# a_2052_22804# vss vss nmos_6p0 w=0.82u l=1u
X11978 a_29700_26786# cap_shunt_p a_29492_27132# vdd pmos_6p0 w=1.2u l=0.5u
X11979 a_33948_16488# a_33860_16532# vss vss nmos_6p0 w=0.82u l=1u
X11980 a_9540_14242# cap_shunt_p a_9332_14588# vdd pmos_6p0 w=1.2u l=0.5u
X11981 a_30616_19668# cap_series_gygyn a_30428_19668# vdd pmos_6p0 w=1.2u l=0.5u
X11982 a_12768_36132# cap_shunt_n a_10660_36194# vss nmos_6p0 w=0.82u l=0.6u
X11983 vdd tune_shunt[5] a_21540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X11984 vdd tune_shunt[7] a_6532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X11985 a_17828_45240# cap_shunt_p a_17620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X11986 a_31708_55255# a_31620_55352# vss vss nmos_6p0 w=0.82u l=1u
X11987 a_9876_12312# cap_shunt_p a_10808_12312# vss nmos_6p0 w=0.82u l=0.6u
X11988 a_20532_29076# cap_shunt_n a_20740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X11989 a_27228_9783# a_27140_9880# vss vss nmos_6p0 w=0.82u l=1u
X11990 vdd tune_shunt[7] a_21540_22428# vdd pmos_6p0 w=1.2u l=0.5u
X11991 a_28692_17016# cap_series_gyn a_29624_17016# vss nmos_6p0 w=0.82u l=0.6u
X11992 a_4816_50244# cap_shunt_n a_2708_50306# vss nmos_6p0 w=0.82u l=0.6u
X11993 vdd a_23308_46280# a_23220_46324# vdd pmos_6p0 w=1.22u l=1u
X11994 a_12332_55255# a_12244_55352# vss vss nmos_6p0 w=0.82u l=1u
X11995 a_37652_38968# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X11996 a_9668_47892# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X11997 a_29916_22327# a_29828_22424# vss vss nmos_6p0 w=0.82u l=1u
X11998 vdd tune_shunt[6] a_3620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X11999 a_34412_48676# cap_shunt_gyn a_34144_48676# vss nmos_6p0 w=0.82u l=0.6u
X12000 a_6508_36439# a_6420_36536# vss vss nmos_6p0 w=0.82u l=1u
X12001 a_1716_3988# cap_shunt_p a_1924_4472# vdd pmos_6p0 w=1.2u l=0.5u
X12002 a_2500_19292# cap_shunt_p a_2708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X12003 a_16500_34972# cap_shunt_n a_16708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X12004 a_13252_27508# cap_shunt_n a_13460_27992# vdd pmos_6p0 w=1.2u l=0.5u
X12005 vdd tune_series_gy[5] a_22436_11828# vdd pmos_6p0 w=1.2u l=0.5u
X12006 a_13796_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12007 vdd a_32156_53687# a_32068_53784# vdd pmos_6p0 w=1.22u l=1u
X12008 vss tune_shunt[6] a_25780_38968# vss nmos_6p0 w=0.51u l=0.6u
X12009 vss cap_shunt_p a_15120_47108# vss nmos_6p0 w=0.82u l=0.6u
X12010 a_24660_28354# cap_shunt_n a_24452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X12011 a_7748_25218# cap_shunt_n a_7540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X12012 a_30016_6040# cap_shunt_n a_28692_6040# vss nmos_6p0 w=0.82u l=0.6u
X12013 a_18424_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12014 vss tune_series_gy[1] a_6760_5556# vss nmos_6p0 w=0.51u l=0.6u
X12015 a_25572_19668# cap_series_gyp a_25780_20152# vdd pmos_6p0 w=1.2u l=0.5u
X12016 a_37980_52552# a_37892_52596# vss vss nmos_6p0 w=0.82u l=1u
X12017 a_2500_16156# cap_shunt_p a_2708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X12018 a_34308_19292# cap_series_gygyn a_34516_18946# vdd pmos_6p0 w=1.2u l=0.5u
X12019 a_16500_31836# cap_shunt_n a_16708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X12020 vss tune_shunt[2] a_1924_6402# vss nmos_6p0 w=0.51u l=0.6u
X12021 a_22644_9176# cap_series_gyp a_22436_8692# vdd pmos_6p0 w=1.2u l=0.5u
X12022 a_9316_48738# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12023 vdd a_32156_50551# a_32068_50648# vdd pmos_6p0 w=1.22u l=1u
X12024 vss cap_shunt_gyp a_34412_43972# vss nmos_6p0 w=0.82u l=0.6u
X12025 a_20532_38484# cap_shunt_n a_20740_38968# vdd pmos_6p0 w=1.2u l=0.5u
X12026 a_24360_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12027 a_23308_38440# a_23220_38484# vss vss nmos_6p0 w=0.82u l=1u
X12028 vdd a_37420_23895# a_37332_23992# vdd pmos_6p0 w=1.22u l=1u
X12029 a_34516_22082# cap_series_gygyp a_36232_22020# vss nmos_6p0 w=0.82u l=0.6u
X12030 vss tune_shunt[7] a_10660_23650# vss nmos_6p0 w=0.51u l=0.6u
X12031 a_34308_16156# cap_series_gygyn a_34516_15810# vdd pmos_6p0 w=1.2u l=0.5u
X12032 a_2708_47170# cap_shunt_p a_2500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X12033 a_20740_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12034 a_3828_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12035 a_20532_35348# cap_shunt_n a_20740_35832# vdd pmos_6p0 w=1.2u l=0.5u
X12036 vss cap_series_gyp a_31024_17316# vss nmos_6p0 w=0.82u l=0.6u
X12037 a_27788_49416# a_27700_49460# vss vss nmos_6p0 w=0.82u l=1u
X12038 vdd a_37420_20759# a_37332_20856# vdd pmos_6p0 w=1.22u l=1u
X12039 vdd tune_shunt[5] a_6084_49084# vdd pmos_6p0 w=1.2u l=0.5u
X12040 vdd a_5276_52552# a_5188_52596# vdd pmos_6p0 w=1.22u l=1u
X12041 a_19152_38968# cap_shunt_n a_17828_38968# vss nmos_6p0 w=0.82u l=0.6u
X12042 a_35840_35832# cap_shunt_n a_33732_35832# vss nmos_6p0 w=0.82u l=0.6u
X12043 vss tune_series_gy[4] a_21636_6040# vss nmos_6p0 w=0.51u l=0.6u
X12044 vdd tune_shunt[7] a_6420_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12045 a_34308_20860# cap_series_gygyp a_34516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X12046 a_15580_52552# a_15492_52596# vss vss nmos_6p0 w=0.82u l=1u
X12047 a_26376_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12048 a_12556_16055# a_12468_16152# vss vss nmos_6p0 w=0.82u l=1u
X12049 a_9316_47170# cap_shunt_p a_9108_47516# vdd pmos_6p0 w=1.2u l=0.5u
X12050 a_3620_13396# cap_shunt_n a_3828_13880# vdd pmos_6p0 w=1.2u l=0.5u
X12051 a_18492_13352# a_18404_13396# vss vss nmos_6p0 w=0.82u l=1u
X12052 a_16708_37762# cap_shunt_n a_16500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X12053 a_27788_46280# a_27700_46324# vss vss nmos_6p0 w=0.82u l=1u
X12054 a_24660_29922# cap_shunt_n a_24452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X12055 a_2500_25564# cap_shunt_p a_2708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X12056 a_6196_47516# cap_shunt_p a_6404_47170# vdd pmos_6p0 w=1.2u l=0.5u
X12057 a_11872_34264# cap_shunt_n a_10548_34264# vss nmos_6p0 w=0.82u l=0.6u
X12058 a_26376_3204# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12059 a_33524_32212# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12060 vdd tune_shunt[7] a_21540_19292# vdd pmos_6p0 w=1.2u l=0.5u
X12061 vss tune_shunt_gy[2] a_37632_41621# vss nmos_6p0 w=0.51u l=0.6u
X12062 a_23464_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12063 a_18492_10216# a_18404_10260# vss vss nmos_6p0 w=0.82u l=1u
X12064 vdd a_20732_52552# a_20644_52596# vdd pmos_6p0 w=1.22u l=1u
X12065 a_10660_44034# cap_shunt_n a_11592_43972# vss nmos_6p0 w=0.82u l=0.6u
X12066 vss cap_shunt_p a_11984_20152# vss nmos_6p0 w=0.82u l=0.6u
X12067 a_2500_22428# cap_shunt_p a_2708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X12068 a_31708_48983# a_31620_49080# vss vss nmos_6p0 w=0.82u l=1u
X12069 a_17828_38968# cap_shunt_n a_17620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X12070 a_11872_31128# cap_shunt_n a_10548_31128# vss nmos_6p0 w=0.82u l=0.6u
X12071 vss tune_series_gygy[4] a_35880_36916# vss nmos_6p0 w=0.51u l=0.6u
X12072 vdd tune_series_gy[5] a_21540_16156# vdd pmos_6p0 w=1.2u l=0.5u
X12073 a_33292_47108# cap_shunt_gyn a_33024_47108# vss nmos_6p0 w=0.82u l=0.6u
X12074 a_7768_5180# cap_series_gyn a_7792_4772# vss nmos_6p0 w=0.82u l=0.6u
X12075 a_12332_48983# a_12244_49080# vss vss nmos_6p0 w=0.82u l=1u
X12076 a_10660_40898# cap_shunt_n a_11592_40836# vss nmos_6p0 w=0.82u l=0.6u
X12077 vdd a_32604_25896# a_32516_25940# vdd pmos_6p0 w=1.22u l=1u
X12078 a_9108_22428# cap_shunt_p a_9316_22082# vdd pmos_6p0 w=1.2u l=0.5u
X12079 a_17828_35832# cap_shunt_n a_17620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X12080 a_31436_20860# cap_series_gygyn a_31624_20860# vdd pmos_6p0 w=1.2u l=0.5u
X12081 vdd a_27676_31735# a_27588_31832# vdd pmos_6p0 w=1.22u l=1u
X12082 a_24660_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12083 vdd tune_shunt[3] a_2724_8692# vdd pmos_6p0 w=1.2u l=0.5u
X12084 a_16708_47170# cap_shunt_n a_16500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X12085 a_34396_52119# a_34308_52216# vss vss nmos_6p0 w=0.82u l=1u
X12086 vss cap_shunt_p a_11200_48376# vss nmos_6p0 w=0.82u l=0.6u
X12087 a_13460_27992# cap_shunt_n a_14392_27992# vss nmos_6p0 w=0.82u l=0.6u
X12088 vdd a_32604_22760# a_32516_22804# vdd pmos_6p0 w=1.22u l=1u
X12089 a_10864_12612# cap_shunt_p a_9540_12674# vss nmos_6p0 w=0.82u l=0.6u
X12090 a_32612_36194# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12091 a_16708_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12092 a_24660_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12093 a_25780_7608# cap_series_gyn a_26712_7608# vss nmos_6p0 w=0.82u l=0.6u
X12094 a_1692_13352# a_1604_13396# vss vss nmos_6p0 w=0.82u l=1u
X12095 a_16500_25564# cap_shunt_n a_16708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X12096 a_13460_24856# cap_shunt_n a_14392_24856# vss nmos_6p0 w=0.82u l=0.6u
X12097 a_5844_3266# cap_shunt_n a_5636_3612# vdd pmos_6p0 w=1.2u l=0.5u
X12098 a_32612_33058# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12099 a_1924_6402# cap_shunt_n a_1716_6748# vdd pmos_6p0 w=1.2u l=0.5u
X12100 a_11572_3988# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12101 vss cap_shunt_p a_4816_20452# vss nmos_6p0 w=0.82u l=0.6u
X12102 vdd tune_series_gygy[5] a_30428_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12103 vdd a_32156_44279# a_32068_44376# vdd pmos_6p0 w=1.22u l=1u
X12104 a_28692_12312# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12105 a_30616_19668# cap_series_gygyn a_30428_19668# vdd pmos_6p0 w=1.2u l=0.5u
X12106 a_1716_3612# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12107 a_18424_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12108 a_32604_8648# a_32516_8692# vss vss nmos_6p0 w=0.82u l=1u
X12109 a_1692_10216# a_1604_10260# vss vss nmos_6p0 w=0.82u l=1u
X12110 a_3036_54120# a_2948_54164# vss vss nmos_6p0 w=0.82u l=1u
X12111 a_29492_5180# cap_shunt_p a_29700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X12112 a_37196_35304# a_37108_35348# vss vss nmos_6p0 w=0.82u l=1u
X12113 a_16500_22428# cap_shunt_n a_16708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X12114 a_20740_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12115 a_20532_29076# cap_shunt_n a_20740_29560# vdd pmos_6p0 w=1.2u l=0.5u
X12116 a_3828_13880# cap_shunt_n a_5544_13880# vss nmos_6p0 w=0.82u l=0.6u
X12117 a_7168_9476# cap_shunt_p a_5844_9538# vss nmos_6p0 w=0.82u l=0.6u
X12118 a_13588_13020# cap_shunt_p a_13796_12674# vdd pmos_6p0 w=1.2u l=0.5u
X12119 vdd a_37420_14487# a_37332_14584# vdd pmos_6p0 w=1.22u l=1u
X12120 a_35840_29560# cap_shunt_p a_33732_29560# vss nmos_6p0 w=0.82u l=0.6u
X12121 a_12712_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12122 a_3248_7608# cap_shunt_n a_1924_7608# vss nmos_6p0 w=0.82u l=0.6u
X12123 vss tune_shunt[7] a_2708_31490# vss nmos_6p0 w=0.51u l=0.6u
X12124 a_10660_28354# cap_shunt_n a_10452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X12125 vss cap_series_gyp a_23072_7908# vss nmos_6p0 w=0.82u l=0.6u
X12126 a_2708_37762# cap_shunt_n a_2500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X12127 a_7560_9176# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12128 a_27496_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12129 a_20740_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12130 a_3828_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12131 a_6572_3988# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12132 vss tune_series_gy[4] a_25780_9176# vss nmos_6p0 w=0.51u l=0.6u
X12133 vdd a_37420_11351# a_37332_11448# vdd pmos_6p0 w=1.22u l=1u
X12134 a_2500_19292# cap_shunt_p a_2708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X12135 a_34844_53687# a_34756_53784# vss vss nmos_6p0 w=0.82u l=1u
X12136 a_22412_47415# a_22324_47512# vss vss nmos_6p0 w=0.82u l=1u
X12137 a_7540_28700# cap_shunt_n a_7748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X12138 a_25572_7124# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12139 vdd tune_series_gygy[3] a_35692_8692# vdd pmos_6p0 w=1.2u l=0.5u
X12140 vdd tune_series_gy[5] a_22436_11828# vdd pmos_6p0 w=1.2u l=0.5u
X12141 a_21540_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12142 a_34536_8316# cap_series_gygyp a_34348_8316# vdd pmos_6p0 w=1.2u l=0.5u
X12143 a_2708_42466# cap_shunt_p a_2500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X12144 a_13460_38968# cap_shunt_n a_13252_38484# vdd pmos_6p0 w=1.2u l=0.5u
X12145 a_24660_28354# cap_shunt_n a_24452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X12146 a_15492_8316# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12147 vdd a_33500_47848# a_33412_47892# vdd pmos_6p0 w=1.22u l=1u
X12148 vdd a_31932_43144# a_31844_43188# vdd pmos_6p0 w=1.22u l=1u
X12149 a_1716_5180# cap_shunt_p a_1924_4834# vdd pmos_6p0 w=1.2u l=0.5u
X12150 a_2500_16156# cap_shunt_p a_2708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X12151 a_34844_50551# a_34756_50648# vss vss nmos_6p0 w=0.82u l=1u
X12152 a_32612_29922# cap_shunt_p a_33544_29860# vss nmos_6p0 w=0.82u l=0.6u
X12153 a_11572_5556# cap_series_gyn a_11780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X12154 vdd tune_series_gygy[2] a_35692_5556# vdd pmos_6p0 w=1.2u l=0.5u
X12155 vss cap_shunt_p a_23072_20452# vss nmos_6p0 w=0.82u l=0.6u
X12156 a_13460_35832# cap_shunt_n a_13252_35348# vdd pmos_6p0 w=1.2u l=0.5u
X12157 a_10660_34626# cap_shunt_n a_11592_34564# vss nmos_6p0 w=0.82u l=0.6u
X12158 a_12788_17016# cap_shunt_p a_12580_16532# vdd pmos_6p0 w=1.2u l=0.5u
X12159 a_35692_18100# cap_series_gygyn a_35880_18100# vdd pmos_6p0 w=1.2u l=0.5u
X12160 vss cap_series_gygyp a_37080_21720# vss nmos_6p0 w=0.82u l=0.6u
X12161 a_17828_29560# cap_shunt_n a_17620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X12162 vdd a_16028_33736# a_15940_33780# vdd pmos_6p0 w=1.22u l=1u
X12163 a_32612_26786# cap_shunt_p a_33544_26724# vss nmos_6p0 w=0.82u l=0.6u
X12164 vdd a_27676_25463# a_27588_25560# vdd pmos_6p0 w=1.22u l=1u
X12165 vdd a_25548_53687# a_25460_53784# vdd pmos_6p0 w=1.22u l=1u
X12166 a_10660_31490# cap_shunt_n a_11592_31428# vss nmos_6p0 w=0.82u l=0.6u
X12167 vdd tune_shunt[5] a_6084_49084# vdd pmos_6p0 w=1.2u l=0.5u
X12168 a_10548_37400# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12169 vdd tune_shunt[7] a_6420_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12170 vdd a_32604_16488# a_32516_16532# vdd pmos_6p0 w=1.22u l=1u
X12171 a_34308_20860# cap_series_gygyp a_34516_20514# vdd pmos_6p0 w=1.2u l=0.5u
X12172 a_9316_47170# cap_shunt_p a_9108_47516# vdd pmos_6p0 w=1.2u l=0.5u
X12173 vdd a_16028_30600# a_15940_30644# vdd pmos_6p0 w=1.22u l=1u
X12174 vdd a_27676_22327# a_27588_22424# vdd pmos_6p0 w=1.22u l=1u
X12175 a_24660_14242# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12176 vdd a_25548_50551# a_25460_50648# vdd pmos_6p0 w=1.22u l=1u
X12177 a_25572_41620# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12178 a_16708_37762# cap_shunt_n a_16500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X12179 a_24660_29922# cap_shunt_n a_24452_30268# vdd pmos_6p0 w=1.2u l=0.5u
X12180 a_22644_9176# cap_series_gyp a_22436_8692# vdd pmos_6p0 w=1.2u l=0.5u
X12181 a_16500_19292# cap_shunt_p a_16708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X12182 a_37652_43972# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12183 a_16708_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12184 vss cap_shunt_n a_4816_14180# vss nmos_6p0 w=0.82u l=0.6u
X12185 a_14012_52119# a_13924_52216# vss vss nmos_6p0 w=0.82u l=1u
X12186 a_24660_11106# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12187 vss cap_shunt_gyp a_36988_48376# vss nmos_6p0 w=0.82u l=0.6u
X12188 a_14372_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12189 a_37644_30600# a_37556_30644# vss vss nmos_6p0 w=0.82u l=1u
X12190 a_35880_7124# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X12191 a_16708_22082# cap_shunt_n a_18424_22020# vss nmos_6p0 w=0.82u l=0.6u
X12192 a_19936_4472# cap_series_gyp a_18612_4472# vss nmos_6p0 w=0.82u l=0.6u
X12193 a_28484_13396# cap_series_gyp a_28692_13880# vdd pmos_6p0 w=1.2u l=0.5u
X12194 a_3036_47848# a_2948_47892# vss vss nmos_6p0 w=0.82u l=1u
X12195 a_10452_42812# cap_shunt_n a_10660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X12196 a_37196_29032# a_37108_29076# vss vss nmos_6p0 w=0.82u l=1u
X12197 a_26768_22020# cap_shunt_p a_24660_22082# vss nmos_6p0 w=0.82u l=0.6u
X12198 vss cap_shunt_p a_11648_9476# vss nmos_6p0 w=0.82u l=0.6u
X12199 a_16500_16156# cap_shunt_p a_16708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X12200 vdd a_10988_54120# a_10900_54164# vdd pmos_6p0 w=1.22u l=1u
X12201 a_37652_40836# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12202 a_24660_7970# cap_series_gyp a_25592_7908# vss nmos_6p0 w=0.82u l=0.6u
X12203 vss cap_shunt_n a_4816_11044# vss nmos_6p0 w=0.82u l=0.6u
X12204 vdd a_36188_54120# a_36100_54164# vdd pmos_6p0 w=1.22u l=1u
X12205 a_6532_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12206 a_4424_43972# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12207 a_5636_8692# cap_shunt_p a_5844_9176# vdd pmos_6p0 w=1.2u l=0.5u
X12208 a_22644_10744# cap_series_gyp a_22436_10260# vdd pmos_6p0 w=1.2u l=0.5u
X12209 vdd tune_series_gygy[4] a_35692_14964# vdd pmos_6p0 w=1.2u l=0.5u
X12210 a_20740_46808# cap_shunt_p a_20532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X12211 vss cap_shunt_p a_8848_45240# vss nmos_6p0 w=0.82u l=0.6u
X12212 vdd tune_series_gy[4] a_25572_18100# vdd pmos_6p0 w=1.2u l=0.5u
X12213 vdd a_2140_19624# a_2052_19668# vdd pmos_6p0 w=1.22u l=1u
X12214 a_6956_45847# a_6868_45944# vss vss nmos_6p0 w=0.82u l=1u
X12215 a_16500_20860# cap_shunt_p a_16708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X12216 vdd tune_shunt[7] a_13588_28700# vdd pmos_6p0 w=1.2u l=0.5u
X12217 a_7580_5180# cap_series_gyn a_7768_5180# vdd pmos_6p0 w=1.2u l=0.5u
X12218 a_14460_8215# a_14372_8312# vss vss nmos_6p0 w=0.82u l=1u
X12219 vdd a_36188_50984# a_36100_51028# vdd pmos_6p0 w=1.22u l=1u
X12220 a_4424_40836# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12221 vdd tune_shunt[7] a_21540_20860# vdd pmos_6p0 w=1.2u l=0.5u
X12222 vdd tune_series_gygy[4] a_35692_11828# vdd pmos_6p0 w=1.2u l=0.5u
X12223 vdd a_16252_55255# a_16164_55352# vdd pmos_6p0 w=1.22u l=1u
X12224 vss tune_shunt[3] a_24660_44034# vss nmos_6p0 w=0.51u l=0.6u
X12225 vss cap_shunt_n a_8848_42104# vss nmos_6p0 w=0.82u l=0.6u
X12226 vss tune_shunt[5] a_2708_22082# vss nmos_6p0 w=0.51u l=0.6u
X12227 vdd a_24876_47848# a_24788_47892# vdd pmos_6p0 w=1.22u l=1u
X12228 a_6956_42711# a_6868_42808# vss vss nmos_6p0 w=0.82u l=1u
X12229 a_27496_12312# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12230 a_17260_12919# a_17172_13016# vss vss nmos_6p0 w=0.82u l=1u
X12231 a_2708_36194# cap_shunt_n a_2500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X12232 a_11592_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12233 a_14692_4472# cap_series_gyp a_14484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X12234 a_20740_17016# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12235 a_18612_11106# cap_series_gyn a_19544_11044# vss nmos_6p0 w=0.82u l=0.6u
X12236 a_17620_19668# cap_shunt_p a_17828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X12237 vdd a_16252_52119# a_16164_52216# vdd pmos_6p0 w=1.22u l=1u
X12238 a_21180_50984# a_21092_51028# vss vss nmos_6p0 w=0.82u l=1u
X12239 a_16708_47170# cap_shunt_n a_17640_47108# vss nmos_6p0 w=0.82u l=0.6u
X12240 vss cap_series_gyn a_23072_14180# vss nmos_6p0 w=0.82u l=0.6u
X12241 vdd tune_series_gygy[5] a_30428_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12242 a_13460_29560# cap_shunt_n a_13252_29076# vdd pmos_6p0 w=1.2u l=0.5u
X12243 a_2708_33058# cap_shunt_p a_2500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X12244 a_35628_33303# a_35540_33400# vss vss nmos_6p0 w=0.82u l=1u
X12245 a_10660_28354# cap_shunt_n a_11592_28292# vss nmos_6p0 w=0.82u l=0.6u
X12246 vdd a_33500_38440# a_33412_38484# vdd pmos_6p0 w=1.22u l=1u
X12247 a_1924_6402# cap_shunt_n a_3640_6340# vss nmos_6p0 w=0.82u l=0.6u
X12248 a_27788_52119# a_27700_52216# vss vss nmos_6p0 w=0.82u l=1u
X12249 vdd a_28572_44279# a_28484_44376# vdd pmos_6p0 w=1.22u l=1u
X12250 a_25780_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12251 a_15700_4834# cap_series_gyn a_15492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X12252 a_35880_19668# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12253 vss cap_series_gyn a_23072_11044# vss nmos_6p0 w=0.82u l=0.6u
X12254 a_11772_55688# a_11684_55732# vss vss nmos_6p0 w=0.82u l=1u
X12255 a_3828_34264# cap_shunt_n a_3620_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12256 a_10660_25218# cap_shunt_n a_11592_25156# vss nmos_6p0 w=0.82u l=0.6u
X12257 a_1924_3266# cap_shunt_n a_3640_3204# vss nmos_6p0 w=0.82u l=0.6u
X12258 vdd tune_shunt[7] a_6532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12259 vss cap_series_gygyp a_37080_12312# vss nmos_6p0 w=0.82u l=0.6u
X12260 a_10660_28354# cap_shunt_n a_10452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X12261 a_25780_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12262 vdd a_27676_16055# a_27588_16152# vdd pmos_6p0 w=1.22u l=1u
X12263 a_25212_45847# a_25124_45944# vss vss nmos_6p0 w=0.82u l=1u
X12264 vdd a_16028_24328# a_15940_24372# vdd pmos_6p0 w=1.22u l=1u
X12265 a_36296_13880# cap_series_gygyn a_35880_13396# vss nmos_6p0 w=0.82u l=0.6u
X12266 a_6172_52552# a_6084_52596# vss vss nmos_6p0 w=0.82u l=1u
X12267 vss tune_shunt[7] a_7748_31490# vss nmos_6p0 w=0.51u l=0.6u
X12268 a_3828_31128# cap_shunt_n a_3620_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12269 a_7540_28700# cap_shunt_n a_7748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X12270 vss cap_shunt_n a_27104_42104# vss nmos_6p0 w=0.82u l=0.6u
X12271 vdd tune_shunt[7] a_6532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12272 a_14692_7608# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12273 a_2708_42466# cap_shunt_p a_2500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X12274 a_13460_38968# cap_shunt_n a_13252_38484# vdd pmos_6p0 w=1.2u l=0.5u
X12275 vdd a_27676_12919# a_27588_13016# vdd pmos_6p0 w=1.22u l=1u
X12276 vdd a_16028_21192# a_15940_21236# vdd pmos_6p0 w=1.22u l=1u
X12277 a_25572_32212# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12278 vss tune_series_gy[5] a_18612_7970# vss nmos_6p0 w=0.51u l=0.6u
X12279 a_9108_49084# cap_shunt_p a_9316_48738# vdd pmos_6p0 w=1.2u l=0.5u
X12280 vss tune_shunt[6] a_12788_48376# vss nmos_6p0 w=0.51u l=0.6u
X12281 a_10452_36540# cap_shunt_n a_10660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X12282 a_36296_10744# cap_series_gygyp a_35880_10260# vss nmos_6p0 w=0.82u l=0.6u
X12283 vdd a_18940_11784# a_18852_11828# vdd pmos_6p0 w=1.22u l=1u
X12284 a_13588_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12285 a_25984_37700# cap_shunt_p a_24660_37762# vss nmos_6p0 w=0.82u l=0.6u
X12286 a_32404_28700# cap_shunt_p a_32612_28354# vdd pmos_6p0 w=1.2u l=0.5u
X12287 a_13460_35832# cap_shunt_n a_13252_35348# vdd pmos_6p0 w=1.2u l=0.5u
X12288 a_6956_5079# a_6868_5176# vss vss nmos_6p0 w=0.82u l=1u
X12289 a_9428_17378# cap_shunt_p a_11144_17316# vss nmos_6p0 w=0.82u l=0.6u
X12290 a_12788_20152# cap_shunt_p a_14504_20152# vss nmos_6p0 w=0.82u l=0.6u
X12291 vss tune_series_gy[4] a_18612_4834# vss nmos_6p0 w=0.51u l=0.6u
X12292 a_24092_3944# a_24004_3988# vss vss nmos_6p0 w=0.82u l=1u
X12293 a_22848_20152# cap_shunt_p a_20740_20152# vss nmos_6p0 w=0.82u l=0.6u
X12294 a_10452_33404# cap_shunt_n a_10660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X12295 a_2500_20860# cap_shunt_p a_2708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X12296 vdd tune_shunt[5] a_9668_52596# vdd pmos_6p0 w=1.2u l=0.5u
X12297 vdd tune_series_gy[4] a_25572_10260# vdd pmos_6p0 w=1.2u l=0.5u
X12298 a_12788_17016# cap_shunt_p a_12580_16532# vdd pmos_6p0 w=1.2u l=0.5u
X12299 a_20740_15448# cap_series_gyn a_20532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X12300 vdd a_23756_46280# a_23668_46324# vdd pmos_6p0 w=1.22u l=1u
X12301 a_16500_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12302 a_9532_55688# a_9444_55732# vss vss nmos_6p0 w=0.82u l=1u
X12303 a_12780_55255# a_12692_55352# vss vss nmos_6p0 w=0.82u l=1u
X12304 vdd a_5612_8215# a_5524_8312# vdd pmos_6p0 w=1.22u l=1u
X12305 a_4424_34564# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12306 a_11780_6040# cap_series_gyn a_11572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X12307 vss tune_shunt[7] a_12788_13880# vss nmos_6p0 w=0.51u l=0.6u
X12308 a_14580_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12309 a_7540_30268# cap_shunt_n a_7748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X12310 a_6956_36439# a_6868_36536# vss vss nmos_6p0 w=0.82u l=1u
X12311 a_2500_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12312 a_16500_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12313 vdd tune_series_gy[5] a_21540_11452# vdd pmos_6p0 w=1.2u l=0.5u
X12314 a_12788_48376# cap_shunt_p a_13720_48376# vss nmos_6p0 w=0.82u l=0.6u
X12315 a_4424_31428# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12316 a_5152_27992# cap_shunt_n a_3828_27992# vss nmos_6p0 w=0.82u l=0.6u
X12317 a_19524_11828# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12318 a_6508_55688# a_6420_55732# vss vss nmos_6p0 w=0.82u l=1u
X12319 vdd a_4940_7080# a_4852_7124# vdd pmos_6p0 w=1.22u l=1u
X12320 a_13340_10216# a_13252_10260# vss vss nmos_6p0 w=0.82u l=1u
X12321 a_16500_49084# cap_shunt_p a_16708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X12322 a_33732_32696# cap_shunt_n a_35448_32696# vss nmos_6p0 w=0.82u l=0.6u
X12323 a_32380_41576# a_32292_41620# vss vss nmos_6p0 w=0.82u l=1u
X12324 a_15904_29860# cap_shunt_n a_13796_29922# vss nmos_6p0 w=0.82u l=0.6u
X12325 a_9540_15810# cap_shunt_p a_11256_15748# vss nmos_6p0 w=0.82u l=0.6u
X12326 a_2708_26786# cap_shunt_p a_2500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X12327 a_11460_41620# cap_shunt_n a_11668_42104# vdd pmos_6p0 w=1.2u l=0.5u
X12328 vss cap_shunt_n a_8960_53380# vss nmos_6p0 w=0.82u l=0.6u
X12329 vdd a_2140_45847# a_2052_45944# vdd pmos_6p0 w=1.22u l=1u
X12330 a_16708_42466# cap_shunt_n a_16500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X12331 a_30632_29860# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12332 vss tune_shunt[7] a_13796_26786# vss nmos_6p0 w=0.51u l=0.6u
X12333 a_35880_8692# cap_series_gygyn a_35904_9176# vss nmos_6p0 w=0.82u l=0.6u
X12334 a_28484_13396# cap_series_gyp a_28692_13880# vdd pmos_6p0 w=1.2u l=0.5u
X12335 a_10452_42812# cap_shunt_n a_10660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X12336 a_5152_24856# cap_shunt_p a_3828_24856# vss nmos_6p0 w=0.82u l=0.6u
X12337 a_12580_19668# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12338 a_7224_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12339 a_23756_38440# a_23668_38484# vss vss nmos_6p0 w=0.82u l=1u
X12340 a_15904_26724# cap_shunt_n a_13796_26786# vss nmos_6p0 w=0.82u l=0.6u
X12341 a_28484_10260# cap_series_gyp a_28692_10744# vdd pmos_6p0 w=1.2u l=0.5u
X12342 a_2588_35304# a_2500_35348# vss vss nmos_6p0 w=0.82u l=1u
X12343 a_22644_10744# cap_series_gyp a_22436_10260# vdd pmos_6p0 w=1.2u l=0.5u
X12344 vdd tune_series_gygy[4] a_35692_14964# vdd pmos_6p0 w=1.2u l=0.5u
X12345 vdd a_2140_42711# a_2052_42808# vdd pmos_6p0 w=1.22u l=1u
X12346 a_28484_38484# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12347 a_30632_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12348 a_20740_46808# cap_shunt_p a_20532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X12349 vdd tune_series_gygy[5] a_34308_23996# vdd pmos_6p0 w=1.2u l=0.5u
X12350 a_11800_7124# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X12351 a_25780_18584# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12352 a_15624_9176# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12353 a_29700_39330# cap_shunt_p a_31416_39268# vss nmos_6p0 w=0.82u l=0.6u
X12354 a_14692_7608# cap_series_gyp a_14484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X12355 a_6852_53442# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12356 vss cap_shunt_n a_18032_32996# vss nmos_6p0 w=0.82u l=0.6u
X12357 vdd tune_series_gygy[4] a_35692_11828# vdd pmos_6p0 w=1.2u l=0.5u
X12358 a_9876_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12359 a_3828_24856# cap_shunt_p a_3620_24372# vdd pmos_6p0 w=1.2u l=0.5u
X12360 vdd tune_shunt[7] a_6532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X12361 a_28692_7608# cap_series_gyp a_30408_7608# vss nmos_6p0 w=0.82u l=0.6u
X12362 a_28484_35348# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12363 a_26376_32996# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12364 a_25780_15448# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12365 a_19724_44279# a_19636_44376# vss vss nmos_6p0 w=0.82u l=1u
X12366 vss tune_series_gy[3] a_18388_3266# vss nmos_6p0 w=0.51u l=0.6u
X12367 a_11256_9476# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12368 a_2708_36194# cap_shunt_n a_2500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X12369 vss tune_shunt[6] a_21748_40898# vss nmos_6p0 w=0.51u l=0.6u
X12370 a_17620_43188# cap_shunt_p a_17828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X12371 a_13588_36540# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12372 vdd tune_shunt[7] a_6532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12373 a_3828_21720# cap_shunt_p a_3620_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12374 a_30364_44279# a_30276_44376# vss vss nmos_6p0 w=0.82u l=1u
X12375 vdd tune_shunt[5] a_3620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X12376 a_19724_41143# a_19636_41240# vss vss nmos_6p0 w=0.82u l=1u
X12377 a_13460_29560# cap_shunt_n a_13252_29076# vdd pmos_6p0 w=1.2u l=0.5u
X12378 a_6060_53687# a_5972_53784# vss vss nmos_6p0 w=0.82u l=1u
X12379 a_2708_33058# cap_shunt_p a_2500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X12380 vdd tune_shunt[5] a_6084_49460# vdd pmos_6p0 w=1.2u l=0.5u
X12381 a_33732_32696# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12382 a_10452_27132# cap_shunt_n a_10660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X12383 a_25572_8692# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12384 a_22064_35832# cap_shunt_n a_20740_35832# vss nmos_6p0 w=0.82u l=0.6u
X12385 a_34308_5180# cap_series_gygyp a_34516_4834# vdd pmos_6p0 w=1.2u l=0.5u
X12386 a_9332_16156# cap_shunt_p a_9540_15810# vdd pmos_6p0 w=1.2u l=0.5u
X12387 vdd a_36300_33736# a_36212_33780# vdd pmos_6p0 w=1.22u l=1u
X12388 a_13588_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12389 vdd tune_shunt[7] a_16500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X12390 a_34536_9884# cap_series_gygyn a_34348_9884# vdd pmos_6p0 w=1.2u l=0.5u
X12391 a_15492_9884# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12392 a_24660_20514# cap_shunt_p a_25592_20452# vss nmos_6p0 w=0.82u l=0.6u
X12393 a_30364_41143# a_30276_41240# vss vss nmos_6p0 w=0.82u l=1u
X12394 a_33948_50984# a_33860_51028# vss vss nmos_6p0 w=0.82u l=1u
X12395 a_12780_48983# a_12692_49080# vss vss nmos_6p0 w=0.82u l=1u
X12396 a_13460_34264# cap_shunt_n a_13252_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12397 a_4424_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12398 a_36384_50244# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12399 a_5936_45240# cap_shunt_p a_3828_45240# vss nmos_6p0 w=0.82u l=0.6u
X12400 a_3380_17016# cap_shunt_p a_3172_16532# vdd pmos_6p0 w=1.2u l=0.5u
X12401 vdd a_16700_18056# a_16612_18100# vdd pmos_6p0 w=1.22u l=1u
X12402 a_3036_53687# a_2948_53784# vss vss nmos_6p0 w=0.82u l=1u
X12403 vss cap_shunt_p a_4032_4772# vss nmos_6p0 w=0.82u l=0.6u
X12404 a_28484_3988# cap_series_gyp a_28692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X12405 vdd a_12444_20759# a_12356_20856# vdd pmos_6p0 w=1.22u l=1u
X12406 vdd a_20284_55255# a_20196_55352# vdd pmos_6p0 w=1.22u l=1u
X12407 a_25572_5556# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12408 a_2500_11452# cap_shunt_n a_2708_11106# vdd pmos_6p0 w=1.2u l=0.5u
X12409 a_2500_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12410 vdd a_36300_30600# a_36212_30644# vdd pmos_6p0 w=1.22u l=1u
X12411 a_16500_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12412 a_15492_6748# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12413 a_34536_6748# cap_series_gygyp a_34348_6748# vdd pmos_6p0 w=1.2u l=0.5u
X12414 a_13460_31128# cap_shunt_n a_13252_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12415 a_4424_25156# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12416 a_5936_42104# cap_shunt_p a_3828_42104# vss nmos_6p0 w=0.82u l=0.6u
X12417 a_16708_29922# cap_shunt_n a_16500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X12418 a_3248_6340# cap_shunt_n a_1924_6402# vss nmos_6p0 w=0.82u l=0.6u
X12419 vdd a_20284_52119# a_20196_52216# vdd pmos_6p0 w=1.22u l=1u
X12420 a_14372_44756# cap_shunt_p a_14580_45240# vdd pmos_6p0 w=1.2u l=0.5u
X12421 a_3828_37400# cap_shunt_n a_3620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X12422 a_16500_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12423 vdd a_2140_39575# a_2052_39672# vdd pmos_6p0 w=1.22u l=1u
X12424 a_16708_36194# cap_shunt_n a_16500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X12425 a_3640_6040# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12426 a_26712_6040# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12427 a_11536_20452# cap_shunt_p a_9428_20514# vss nmos_6p0 w=0.82u l=0.6u
X12428 a_9108_49084# cap_shunt_p a_9316_48738# vdd pmos_6p0 w=1.2u l=0.5u
X12429 a_14728_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12430 a_10452_36540# cap_shunt_n a_10660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X12431 a_2708_45602# cap_shunt_p a_3640_45540# vss nmos_6p0 w=0.82u l=0.6u
X12432 a_3248_3204# cap_shunt_n a_1924_3266# vss nmos_6p0 w=0.82u l=0.6u
X12433 a_32404_28700# cap_shunt_p a_32612_28354# vdd pmos_6p0 w=1.2u l=0.5u
X12434 a_3484_54120# a_3396_54164# vss vss nmos_6p0 w=0.82u l=1u
X12435 a_2588_29032# a_2500_29076# vss vss nmos_6p0 w=0.82u l=1u
X12436 a_20620_22327# a_20532_22424# vss vss nmos_6p0 w=0.82u l=1u
X12437 vdd a_2140_36439# a_2052_36536# vdd pmos_6p0 w=1.22u l=1u
X12438 a_16708_33058# cap_shunt_n a_16500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X12439 a_3620_14964# cap_shunt_p a_3828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X12440 vss tune_shunt[7] a_13796_17378# vss nmos_6p0 w=0.51u l=0.6u
X12441 a_13384_46808# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12442 a_10452_33404# cap_shunt_n a_10660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X12443 a_5152_15448# cap_shunt_p a_3828_15448# vss nmos_6p0 w=0.82u l=0.6u
X12444 a_2500_50652# cap_shunt_n a_2708_50306# vdd pmos_6p0 w=1.2u l=0.5u
X12445 a_2708_42466# cap_shunt_p a_3640_42404# vss nmos_6p0 w=0.82u l=0.6u
X12446 a_35840_22020# cap_series_gygyp a_34516_22082# vss nmos_6p0 w=0.82u l=0.6u
X12447 a_29244_19624# a_29156_19668# vss vss nmos_6p0 w=0.82u l=1u
X12448 a_19164_55688# a_19076_55732# vss vss nmos_6p0 w=0.82u l=1u
X12449 vdd tune_shunt[5] a_6644_53788# vdd pmos_6p0 w=1.2u l=0.5u
X12450 a_32716_9783# a_32628_9880# vss vss nmos_6p0 w=0.82u l=1u
X12451 vdd a_37644_27464# a_37556_27508# vdd pmos_6p0 w=1.22u l=1u
X12452 a_34952_9476# cap_series_gygyn a_34536_9884# vss nmos_6p0 w=0.82u l=0.6u
X12453 a_15904_17316# cap_shunt_p a_13796_17378# vss nmos_6p0 w=0.82u l=0.6u
X12454 a_2588_25896# a_2500_25940# vss vss nmos_6p0 w=0.82u l=1u
X12455 vdd tune_shunt[7] a_13588_20860# vdd pmos_6p0 w=1.2u l=0.5u
X12456 a_17828_43672# cap_shunt_p a_19544_43672# vss nmos_6p0 w=0.82u l=0.6u
X12457 a_6740_35832# cap_shunt_n a_8456_35832# vss nmos_6p0 w=0.82u l=0.6u
X12458 a_5636_10260# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12459 a_9108_50652# cap_shunt_p a_9316_50306# vdd pmos_6p0 w=1.2u l=0.5u
X12460 a_28484_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12461 a_25572_7124# cap_series_gyn a_25780_7608# vdd pmos_6p0 w=1.2u l=0.5u
X12462 a_30632_17316# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12463 a_27888_43672# cap_shunt_p a_25780_43672# vss nmos_6p0 w=0.82u l=0.6u
X12464 a_15492_8316# cap_series_gyn a_15700_7970# vdd pmos_6p0 w=1.2u l=0.5u
X12465 a_22860_47415# a_22772_47512# vss vss nmos_6p0 w=0.82u l=1u
X12466 vss cap_shunt_p a_5936_32696# vss nmos_6p0 w=0.82u l=0.6u
X12467 vdd tune_series_gy[3] a_21316_3612# vdd pmos_6p0 w=1.2u l=0.5u
X12468 a_17828_40536# cap_shunt_n a_19544_40536# vss nmos_6p0 w=0.82u l=0.6u
X12469 vss cap_shunt_n a_18032_23588# vss nmos_6p0 w=0.82u l=0.6u
X12470 a_16500_49084# cap_shunt_p a_16708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X12471 a_30016_12312# cap_series_gyn a_28692_12312# vss nmos_6p0 w=0.82u l=0.6u
X12472 a_32444_14588# cap_series_gyp a_32632_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12473 a_16688_43672# cap_shunt_n a_14580_43672# vss nmos_6p0 w=0.82u l=0.6u
X12474 a_27888_40536# cap_shunt_n a_25780_40536# vss nmos_6p0 w=0.82u l=0.6u
X12475 a_19724_34871# a_19636_34968# vss vss nmos_6p0 w=0.82u l=1u
X12476 a_26376_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12477 vss cap_series_gygyp a_36624_4772# vss nmos_6p0 w=0.82u l=0.6u
X12478 vdd a_33500_55255# a_33412_55352# vdd pmos_6p0 w=1.22u l=1u
X12479 a_17828_37400# cap_shunt_n a_17620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X12480 a_2708_26786# cap_shunt_p a_2500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X12481 a_11460_41620# cap_shunt_n a_11668_42104# vdd pmos_6p0 w=1.2u l=0.5u
X12482 a_32404_30268# cap_shunt_p a_32612_29922# vdd pmos_6p0 w=1.2u l=0.5u
X12483 a_10340_3612# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12484 vdd a_28124_8215# a_28036_8312# vdd pmos_6p0 w=1.22u l=1u
X12485 a_28484_13396# cap_series_gyp a_28692_13880# vdd pmos_6p0 w=1.2u l=0.5u
X12486 a_10452_42812# cap_shunt_n a_10660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X12487 vdd a_27228_41143# a_27140_41240# vdd pmos_6p0 w=1.22u l=1u
X12488 a_22064_29560# cap_shunt_n a_20740_29560# vss nmos_6p0 w=0.82u l=0.6u
X12489 a_22644_7608# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12490 a_24660_14242# cap_series_gyn a_25592_14180# vss nmos_6p0 w=0.82u l=0.6u
X12491 a_13588_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12492 a_34308_20860# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12493 a_16688_40536# cap_shunt_n a_14580_40536# vss nmos_6p0 w=0.82u l=0.6u
X12494 vdd a_8860_17623# a_8772_17720# vdd pmos_6p0 w=1.22u l=1u
X12495 vdd a_33500_52119# a_33412_52216# vdd pmos_6p0 w=1.22u l=1u
X12496 vdd a_30924_47848# a_30836_47892# vdd pmos_6p0 w=1.22u l=1u
X12497 a_3620_46324# cap_shunt_p a_3828_46808# vdd pmos_6p0 w=1.2u l=0.5u
X12498 a_13460_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12499 a_19724_31735# a_19636_31832# vss vss nmos_6p0 w=0.82u l=1u
X12500 a_31624_8316# cap_series_gygyn a_31436_8316# vdd pmos_6p0 w=1.2u l=0.5u
X12501 a_6532_36916# cap_shunt_n a_6740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X12502 vdd a_16476_33736# a_16388_33780# vdd pmos_6p0 w=1.22u l=1u
X12503 a_17620_14964# cap_shunt_p a_17828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X12504 vdd a_25996_53687# a_25908_53784# vdd pmos_6p0 w=1.22u l=1u
X12505 a_10340_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12506 a_19276_30167# a_19188_30264# vss vss nmos_6p0 w=0.82u l=1u
X12507 a_22064_26424# cap_shunt_n a_20740_26424# vss nmos_6p0 w=0.82u l=0.6u
X12508 a_24660_11106# cap_series_gyp a_25592_11044# vss nmos_6p0 w=0.82u l=0.6u
X12509 vdd tune_shunt[7] a_16500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12510 a_13796_47170# cap_shunt_p a_15512_47108# vss nmos_6p0 w=0.82u l=0.6u
X12511 a_9540_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12512 a_16500_19292# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12513 a_33948_41576# a_33860_41620# vss vss nmos_6p0 w=0.82u l=1u
X12514 a_35692_36916# cap_series_gygyp a_35880_36916# vdd pmos_6p0 w=1.2u l=0.5u
X12515 a_13460_24856# cap_shunt_n a_13252_24372# vdd pmos_6p0 w=1.2u l=0.5u
X12516 vss cap_shunt_n a_23856_29860# vss nmos_6p0 w=0.82u l=0.6u
X12517 vdd a_16476_30600# a_16388_30644# vdd pmos_6p0 w=1.22u l=1u
X12518 vdd a_6620_54120# a_6532_54164# vdd pmos_6p0 w=1.22u l=1u
X12519 vdd a_25996_50551# a_25908_50648# vdd pmos_6p0 w=1.22u l=1u
X12520 vdd tune_shunt_gy[6] a_37444_50648# vdd pmos_6p0 w=1.215u l=0.5u
X12521 a_10340_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12522 a_19276_27031# a_19188_27128# vss vss nmos_6p0 w=0.82u l=1u
X12523 a_31624_19292# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12524 a_17148_55255# a_17060_55352# vss vss nmos_6p0 w=0.82u l=1u
X12525 a_9540_11106# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12526 a_16500_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12527 a_13588_45948# cap_shunt_p a_13796_45602# vdd pmos_6p0 w=1.2u l=0.5u
X12528 a_11668_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12529 a_13460_21720# cap_shunt_n a_13252_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12530 vdd tune_shunt[6] a_10452_45948# vdd pmos_6p0 w=1.2u l=0.5u
X12531 vss cap_shunt_n a_23856_26724# vss nmos_6p0 w=0.82u l=0.6u
X12532 a_14460_52119# a_14372_52216# vss vss nmos_6p0 w=0.82u l=1u
X12533 a_3828_27992# cap_shunt_n a_3620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X12534 a_18516_5556# cap_series_gyn a_18724_6040# vdd pmos_6p0 w=1.2u l=0.5u
X12535 a_9540_12674# cap_shunt_p a_9332_13020# vdd pmos_6p0 w=1.2u l=0.5u
X12536 a_25780_13880# cap_series_gyn a_25572_13396# vdd pmos_6p0 w=1.2u l=0.5u
X12537 vdd tune_shunt[5] a_6084_49460# vdd pmos_6p0 w=1.2u l=0.5u
X12538 a_11668_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12539 a_16708_26786# cap_shunt_n a_16500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X12540 a_1924_4472# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X12541 a_2708_36194# cap_shunt_n a_3640_36132# vss nmos_6p0 w=0.82u l=0.6u
X12542 a_10452_27132# cap_shunt_n a_10660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X12543 a_7580_5180# cap_series_gyn a_7768_5180# vdd pmos_6p0 w=1.2u l=0.5u
X12544 a_2500_44380# cap_shunt_p a_2708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X12545 a_11984_18584# cap_shunt_p a_9876_18584# vss nmos_6p0 w=0.82u l=0.6u
X12546 vdd tune_shunt[7] a_16500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X12547 a_11800_8692# cap_series_gyp a_11612_8692# vdd pmos_6p0 w=1.2u l=0.5u
X12548 a_10452_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12549 a_25592_6340# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12550 a_13460_34264# cap_shunt_n a_13252_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12551 a_24452_17724# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12552 vss tune_shunt[6] a_21748_37762# vss nmos_6p0 w=0.51u l=0.6u
X12553 a_6740_29560# cap_shunt_n a_8456_29560# vss nmos_6p0 w=0.82u l=0.6u
X12554 vdd a_2140_27031# a_2052_27128# vdd pmos_6p0 w=1.22u l=1u
X12555 a_14692_4472# cap_series_gyp a_14484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X12556 a_2500_41244# cap_shunt_p a_2708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X12557 a_17024_9476# cap_series_gyn a_15700_9538# vss nmos_6p0 w=0.82u l=0.6u
X12558 a_11984_15448# cap_shunt_p a_9876_15448# vss nmos_6p0 w=0.82u l=0.6u
X12559 a_15120_32996# cap_shunt_n a_13796_33058# vss nmos_6p0 w=0.82u l=0.6u
X12560 a_18760_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12561 vdd a_5612_47415# a_5524_47512# vdd pmos_6p0 w=1.22u l=1u
X12562 a_13460_31128# cap_shunt_n a_13252_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12563 vss tune_shunt[6] a_21748_34626# vss nmos_6p0 w=0.51u l=0.6u
X12564 a_6740_26424# cap_shunt_n a_8456_26424# vss nmos_6p0 w=0.82u l=0.6u
X12565 a_2588_16488# a_2500_16532# vss vss nmos_6p0 w=0.82u l=1u
X12566 a_17828_34264# cap_shunt_n a_19544_34264# vss nmos_6p0 w=0.82u l=0.6u
X12567 a_14372_44756# cap_shunt_p a_14580_45240# vdd pmos_6p0 w=1.2u l=0.5u
X12568 a_27888_34264# cap_shunt_p a_25780_34264# vss nmos_6p0 w=0.82u l=0.6u
X12569 vdd a_33500_48983# a_33412_49080# vdd pmos_6p0 w=1.22u l=1u
X12570 a_28692_34264# cap_shunt_p a_28484_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12571 a_19724_28599# a_19636_28696# vss vss nmos_6p0 w=0.82u l=1u
X12572 a_36652_43972# cap_shunt_gyp a_36384_43972# vss nmos_6p0 w=0.82u l=0.6u
X12573 vss cap_shunt_p a_5936_23288# vss nmos_6p0 w=0.82u l=0.6u
X12574 a_7672_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12575 a_10452_36540# cap_shunt_n a_10660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X12576 a_4940_5079# a_4852_5176# vss vss nmos_6p0 w=0.82u l=1u
X12577 vss cap_shunt_n a_15568_21720# vss nmos_6p0 w=0.82u l=0.6u
X12578 a_12788_49944# cap_shunt_n a_12580_49460# vdd pmos_6p0 w=1.2u l=0.5u
X12579 a_10452_6748# cap_series_gyn a_10660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X12580 a_17828_31128# cap_shunt_n a_19544_31128# vss nmos_6p0 w=0.82u l=0.6u
X12581 vss tune_shunt[1] a_25444_3266# vss nmos_6p0 w=0.51u l=0.6u
X12582 a_27888_31128# cap_shunt_p a_25780_31128# vss nmos_6p0 w=0.82u l=0.6u
X12583 a_28692_31128# cap_shunt_n a_28484_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12584 vss tune_shunt[7] a_17828_27992# vss nmos_6p0 w=0.51u l=0.6u
X12585 a_19724_25463# a_19636_25560# vss vss nmos_6p0 w=0.82u l=1u
X12586 a_36652_40836# cap_shunt_gyp a_36384_40836# vss nmos_6p0 w=0.82u l=0.6u
X12587 a_17828_27992# cap_shunt_n a_17620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X12588 vss cap_series_gyn a_27888_13880# vss nmos_6p0 w=0.82u l=0.6u
X12589 a_29700_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12590 a_7672_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12591 a_9876_48376# cap_shunt_p a_11592_48376# vss nmos_6p0 w=0.82u l=0.6u
X12592 a_10452_33404# cap_shunt_n a_10660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X12593 a_5844_9538# cap_shunt_p a_5636_9884# vdd pmos_6p0 w=1.2u l=0.5u
X12594 vdd a_25548_52552# a_25460_52596# vdd pmos_6p0 w=1.22u l=1u
X12595 a_2500_50652# cap_shunt_n a_2708_50306# vdd pmos_6p0 w=1.2u l=0.5u
X12596 a_10660_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12597 vss tune_shunt[7] a_17828_24856# vss nmos_6p0 w=0.51u l=0.6u
X12598 a_12580_18100# cap_shunt_p a_12788_18584# vdd pmos_6p0 w=1.2u l=0.5u
X12599 vdd tune_shunt[5] a_21540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X12600 a_13460_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12601 vss cap_series_gyn a_27888_10744# vss nmos_6p0 w=0.82u l=0.6u
X12602 a_25660_45847# a_25572_45944# vss vss nmos_6p0 w=0.82u l=1u
X12603 vdd a_16476_24328# a_16388_24372# vdd pmos_6p0 w=1.22u l=1u
X12604 vss tune_series_gy[3] a_28692_9176# vss nmos_6p0 w=0.51u l=0.6u
X12605 a_5844_9176# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X12606 a_2724_10260# cap_shunt_n a_2932_10744# vdd pmos_6p0 w=1.2u l=0.5u
X12607 a_9108_50652# cap_shunt_p a_9316_50306# vdd pmos_6p0 w=1.2u l=0.5u
X12608 a_6532_27508# cap_shunt_n a_6740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X12609 a_10340_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12610 a_1716_3612# cap_shunt_n a_1924_3266# vdd pmos_6p0 w=1.2u l=0.5u
X12611 vdd tune_shunt_gy[3] a_37444_44376# vdd pmos_6p0 w=1.215u l=0.5u
X12612 a_37080_4472# cap_series_gygyp a_35880_3988# vss nmos_6p0 w=0.82u l=0.6u
X12613 a_34844_3944# a_34756_3988# vss vss nmos_6p0 w=0.82u l=1u
X12614 a_22064_17016# cap_shunt_p a_20740_17016# vss nmos_6p0 w=0.82u l=0.6u
X12615 vss cap_shunt_p a_8400_17316# vss nmos_6p0 w=0.82u l=0.6u
X12616 a_33440_14180# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12617 vdd a_16812_50551# a_16724_50648# vdd pmos_6p0 w=1.22u l=1u
X12618 a_13588_39676# cap_shunt_n a_13796_39330# vdd pmos_6p0 w=1.2u l=0.5u
X12619 vdd tune_shunt[6] a_21540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X12620 vdd tune_shunt[6] a_10452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X12621 a_34396_55688# a_34308_55732# vss vss nmos_6p0 w=0.82u l=1u
X12622 vdd a_16476_21192# a_16388_21236# vdd pmos_6p0 w=1.22u l=1u
X12623 vdd a_6060_23895# a_5972_23992# vdd pmos_6p0 w=1.22u l=1u
X12624 a_19276_17623# a_19188_17720# vss vss nmos_6p0 w=0.82u l=1u
X12625 a_7616_18884# cap_shunt_p a_6292_18946# vss nmos_6p0 w=0.82u l=0.6u
X12626 a_32444_14588# cap_series_gyp a_32632_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12627 vdd a_37868_17623# a_37780_17720# vdd pmos_6p0 w=1.22u l=1u
X12628 a_2500_20860# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12629 a_25780_7608# cap_series_gyn a_25572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X12630 a_35692_13396# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12631 a_32404_30268# cap_shunt_p a_32612_29922# vdd pmos_6p0 w=1.2u l=0.5u
X12632 a_34348_8316# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12633 a_33440_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12634 a_15700_7970# cap_series_gyn a_15492_8316# vdd pmos_6p0 w=1.2u l=0.5u
X12635 vss cap_shunt_p a_23856_17316# vss nmos_6p0 w=0.82u l=0.6u
X12636 a_9668_19668# cap_shunt_p a_9876_20152# vdd pmos_6p0 w=1.2u l=0.5u
X12637 a_9668_19668# cap_shunt_p a_9876_20152# vdd pmos_6p0 w=1.2u l=0.5u
X12638 vss tune_shunt[7] a_20740_21720# vss nmos_6p0 w=0.51u l=0.6u
X12639 a_2932_12312# cap_shunt_n a_3864_12312# vss nmos_6p0 w=0.82u l=0.6u
X12640 a_13796_37762# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12641 a_18032_22020# cap_shunt_n a_16708_22082# vss nmos_6p0 w=0.82u l=0.6u
X12642 a_28692_4472# tune_series_gy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X12643 a_24452_13020# cap_series_gyn a_24660_12674# vdd pmos_6p0 w=1.2u l=0.5u
X12644 a_7616_15748# cap_shunt_p a_6292_15810# vss nmos_6p0 w=0.82u l=0.6u
X12645 a_37532_54120# a_37444_54164# vss vss nmos_6p0 w=0.82u l=1u
X12646 a_35532_45540# cap_shunt_gyp a_35264_45540# vss nmos_6p0 w=0.82u l=0.6u
X12647 a_7748_44034# cap_shunt_p a_7540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X12648 vdd a_30588_41576# a_30500_41620# vdd pmos_6p0 w=1.22u l=1u
X12649 a_20532_25940# cap_shunt_n a_20740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X12650 a_23072_18884# cap_shunt_p a_21748_18946# vss nmos_6p0 w=0.82u l=0.6u
X12651 a_25572_38484# cap_shunt_p a_25780_38968# vdd pmos_6p0 w=1.2u l=0.5u
X12652 vdd a_17596_13352# a_17508_13396# vdd pmos_6p0 w=1.22u l=1u
X12653 a_6532_36916# cap_shunt_n a_6740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X12654 a_9980_55688# a_9892_55732# vss vss nmos_6p0 w=0.82u l=1u
X12655 vdd tune_shunt[7] a_16500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12656 a_20740_38968# cap_shunt_n a_22456_38968# vss nmos_6p0 w=0.82u l=0.6u
X12657 a_13796_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12658 a_6572_7124# cap_series_gyp a_6760_7124# vdd pmos_6p0 w=1.2u l=0.5u
X12659 a_36232_4772# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X12660 a_35532_42404# cap_shunt_gyn a_35264_42404# vss nmos_6p0 w=0.82u l=0.6u
X12661 a_13460_24856# cap_shunt_n a_13252_24372# vdd pmos_6p0 w=1.2u l=0.5u
X12662 a_35880_19668# cap_series_gygyp a_35904_20152# vss nmos_6p0 w=0.82u l=0.6u
X12663 a_7748_40898# cap_shunt_n a_7540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X12664 vss tune_shunt[7] a_21748_28354# vss nmos_6p0 w=0.51u l=0.6u
X12665 a_20532_22804# cap_shunt_p a_20740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X12666 a_23072_15748# cap_series_gyn a_21748_15810# vss nmos_6p0 w=0.82u l=0.6u
X12667 a_25572_35348# cap_shunt_p a_25780_35832# vdd pmos_6p0 w=1.2u l=0.5u
X12668 vss cap_series_gygyp a_37080_4472# vss nmos_6p0 w=0.82u l=0.6u
X12669 a_6740_15448# cap_shunt_p a_6532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X12670 a_6956_55688# a_6868_55732# vss vss nmos_6p0 w=0.82u l=1u
X12671 a_7748_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12672 a_31820_50984# a_31732_51028# vss vss nmos_6p0 w=0.82u l=1u
X12673 vdd a_5612_38007# a_5524_38104# vdd pmos_6p0 w=1.22u l=1u
X12674 a_15120_23588# cap_shunt_n a_13796_23650# vss nmos_6p0 w=0.82u l=0.6u
X12675 a_13588_45948# cap_shunt_p a_13796_45602# vdd pmos_6p0 w=1.2u l=0.5u
X12676 vss cap_shunt_n a_31024_36132# vss nmos_6p0 w=0.82u l=0.6u
X12677 a_13460_21720# cap_shunt_n a_13252_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12678 a_6292_48738# cap_shunt_p a_7224_48676# vss nmos_6p0 w=0.82u l=0.6u
X12679 vss tune_shunt[5] a_21748_25218# vss nmos_6p0 w=0.51u l=0.6u
X12680 a_7176_4472# cap_series_gyp a_6760_3988# vss nmos_6p0 w=0.82u l=0.6u
X12681 a_6084_17724# cap_shunt_p a_6292_17378# vdd pmos_6p0 w=1.2u l=0.5u
X12682 vdd a_13228_54120# a_13140_54164# vdd pmos_6p0 w=1.22u l=1u
X12683 a_35880_14964# cap_series_gygyn a_35692_14964# vdd pmos_6p0 w=1.2u l=0.5u
X12684 a_32824_18884# cap_series_gygyn a_31624_19292# vss nmos_6p0 w=0.82u l=0.6u
X12685 a_28692_24856# cap_shunt_p a_28484_24372# vdd pmos_6p0 w=1.2u l=0.5u
X12686 a_6740_12312# cap_shunt_p a_6532_11828# vdd pmos_6p0 w=1.2u l=0.5u
X12687 a_3380_49944# cap_shunt_p a_3172_49460# vdd pmos_6p0 w=1.2u l=0.5u
X12688 a_25780_13880# cap_series_gyn a_25572_13396# vdd pmos_6p0 w=1.2u l=0.5u
X12689 vss tune_series_gygy[5] a_34516_17378# vss nmos_6p0 w=0.51u l=0.6u
X12690 a_10452_27132# cap_shunt_n a_10660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X12691 vss cap_series_gygyp a_35840_12612# vss nmos_6p0 w=0.82u l=0.6u
X12692 a_5612_19191# a_5524_19288# vss vss nmos_6p0 w=0.82u l=1u
X12693 a_30028_52552# a_29940_52596# vss vss nmos_6p0 w=0.82u l=1u
X12694 a_2500_44380# cap_shunt_p a_2708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X12695 a_9464_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12696 a_13796_23650# cap_shunt_n a_13588_23996# vdd pmos_6p0 w=1.2u l=0.5u
X12697 vdd a_26444_47415# a_26356_47512# vdd pmos_6p0 w=1.22u l=1u
X12698 a_35880_11828# cap_series_gygyp a_35692_11828# vdd pmos_6p0 w=1.2u l=0.5u
X12699 vdd a_1692_17623# a_1604_17720# vdd pmos_6p0 w=1.22u l=1u
X12700 vss tune_shunt[7] a_17828_18584# vss nmos_6p0 w=0.51u l=0.6u
X12701 a_15904_46808# cap_shunt_p a_14580_46808# vss nmos_6p0 w=0.82u l=0.6u
X12702 vss tune_series_gygy[0] a_35880_3988# vss nmos_6p0 w=0.51u l=0.6u
X12703 a_7672_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12704 a_5612_16055# a_5524_16152# vss vss nmos_6p0 w=0.82u l=1u
X12705 a_2500_41244# cap_shunt_p a_2708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X12706 vdd a_10988_7080# a_10900_7124# vdd pmos_6p0 w=1.22u l=1u
X12707 vss tune_shunt[7] a_17828_15448# vss nmos_6p0 w=0.51u l=0.6u
X12708 a_15356_18056# a_15268_18100# vss vss nmos_6p0 w=0.82u l=1u
X12709 a_18516_5556# cap_series_gyn a_18724_6040# vdd pmos_6p0 w=1.2u l=0.5u
X12710 a_30408_6040# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12711 vdd tune_shunt[2] a_1716_8316# vdd pmos_6p0 w=1.2u l=0.5u
X12712 a_27676_9783# a_27588_9880# vss vss nmos_6p0 w=0.82u l=1u
X12713 a_9332_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12714 a_25212_55688# a_25124_55732# vss vss nmos_6p0 w=0.82u l=1u
X12715 a_10540_43144# a_10452_43188# vss vss nmos_6p0 w=0.82u l=1u
X12716 a_29720_9884# cap_series_gyn a_29744_9476# vss nmos_6p0 w=0.82u l=0.6u
X12717 a_9644_46280# a_9556_46324# vss vss nmos_6p0 w=0.82u l=1u
X12718 a_15356_14920# a_15268_14964# vss vss nmos_6p0 w=0.82u l=1u
X12719 a_2500_11452# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12720 vdd a_6060_14487# a_5972_14584# vdd pmos_6p0 w=1.22u l=1u
X12721 vdd tune_series_gy[5] a_19524_13396# vdd pmos_6p0 w=1.2u l=0.5u
X12722 a_36688_23288# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X12723 a_10540_40008# a_10452_40052# vss vss nmos_6p0 w=0.82u l=1u
X12724 vss cap_series_gyp a_20720_4472# vss nmos_6p0 w=0.82u l=0.6u
X12725 a_10752_17316# cap_shunt_p a_9428_17378# vss nmos_6p0 w=0.82u l=0.6u
X12726 a_16500_44380# cap_shunt_p a_16708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X12727 a_11800_8692# cap_series_gyp a_12608_9176# vss nmos_6p0 w=0.82u l=0.6u
X12728 vss tune_shunt[6] a_20740_35832# vss nmos_6p0 w=0.51u l=0.6u
X12729 a_13796_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12730 a_3484_53687# a_3396_53784# vss vss nmos_6p0 w=0.82u l=1u
X12731 vdd a_12892_20759# a_12804_20856# vdd pmos_6p0 w=1.22u l=1u
X12732 a_11312_51812# cap_shunt_n a_9204_51874# vss nmos_6p0 w=0.82u l=0.6u
X12733 a_20532_16532# cap_shunt_p a_20740_17016# vdd pmos_6p0 w=1.2u l=0.5u
X12734 a_32612_36194# cap_shunt_n a_32404_36540# vdd pmos_6p0 w=1.2u l=0.5u
X12735 a_25572_29076# cap_shunt_p a_25780_29560# vdd pmos_6p0 w=1.2u l=0.5u
X12736 a_6532_27508# cap_shunt_n a_6740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X12737 a_37420_55255# a_37332_55352# vss vss nmos_6p0 w=0.82u l=1u
X12738 vdd a_2140_47848# a_2052_47892# vdd pmos_6p0 w=1.22u l=1u
X12739 vdd tune_shunt[6] a_24452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X12740 a_36524_30167# a_36436_30264# vss vss nmos_6p0 w=0.82u l=1u
X12741 a_16500_41244# cap_shunt_n a_16708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X12742 a_13796_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12743 a_11592_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12744 a_13588_39676# cap_shunt_n a_13796_39330# vdd pmos_6p0 w=1.2u l=0.5u
X12745 a_9668_51028# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12746 vss tune_shunt[7] a_16708_26786# vss nmos_6p0 w=0.51u l=0.6u
X12747 a_21748_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12748 vdd tune_shunt[5] a_2500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X12749 a_32612_33058# cap_shunt_n a_32404_33404# vdd pmos_6p0 w=1.2u l=0.5u
X12750 vdd a_2140_44712# a_2052_44756# vdd pmos_6p0 w=1.22u l=1u
X12751 a_37632_40053# cap_shunt_gyn a_37652_40536# vss nmos_6p0 w=0.82u l=0.6u
X12752 a_25780_32696# cap_shunt_p a_26712_32696# vss nmos_6p0 w=0.82u l=0.6u
X12753 vdd tune_shunt[7] a_24452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X12754 a_18404_11452# cap_series_gyn a_18612_11106# vdd pmos_6p0 w=1.2u l=0.5u
X12755 a_32444_14588# cap_series_gyp a_32632_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12756 a_6516_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12757 vdd a_6508_31735# a_6420_31832# vdd pmos_6p0 w=1.22u l=1u
X12758 a_36524_27031# a_36436_27128# vss vss nmos_6p0 w=0.82u l=1u
X12759 a_20740_45240# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12760 a_35056_32696# cap_shunt_n a_33732_32696# vss nmos_6p0 w=0.82u l=0.6u
X12761 a_5844_3266# cap_shunt_n a_7560_3204# vss nmos_6p0 w=0.82u l=0.6u
X12762 a_17620_47892# cap_shunt_p a_17828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X12763 vdd a_37420_30167# a_37332_30264# vdd pmos_6p0 w=1.22u l=1u
X12764 a_19152_48376# cap_shunt_p a_17828_48376# vss nmos_6p0 w=0.82u l=0.6u
X12765 a_3828_26424# cap_shunt_p a_3620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X12766 a_24452_13020# cap_series_gyn a_24660_12674# vdd pmos_6p0 w=1.2u l=0.5u
X12767 a_33732_34264# cap_shunt_n a_33524_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12768 vdd a_14908_8215# a_14820_8312# vdd pmos_6p0 w=1.22u l=1u
X12769 a_10808_49944# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12770 a_6196_47516# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12771 a_20740_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12772 a_29692_19624# a_29604_19668# vss vss nmos_6p0 w=0.82u l=1u
X12773 vss tune_shunt[5] a_6292_15810# vss nmos_6p0 w=0.51u l=0.6u
X12774 a_17620_44756# cap_shunt_p a_17828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X12775 a_6532_36916# cap_shunt_n a_6740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X12776 a_13796_14242# cap_shunt_p a_13588_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12777 a_3828_23288# cap_shunt_p a_3620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X12778 vdd a_20844_50551# a_20756_50648# vdd pmos_6p0 w=1.22u l=1u
X12779 a_33732_31128# cap_shunt_n a_33524_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12780 a_28692_38968# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12781 a_17828_37400# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12782 a_12656_32696# cap_shunt_n a_10548_32696# vss nmos_6p0 w=0.82u l=0.6u
X12783 vss cap_shunt_n a_19152_27992# vss nmos_6p0 w=0.82u l=0.6u
X12784 a_31024_39268# cap_shunt_p a_29700_39330# vss nmos_6p0 w=0.82u l=0.6u
X12785 a_16588_55688# a_16500_55732# vss vss nmos_6p0 w=0.82u l=1u
X12786 a_17640_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12787 vdd tune_series_gy[5] a_19524_7124# vdd pmos_6p0 w=1.2u l=0.5u
X12788 vss tune_series_gy[5] a_21748_15810# vss nmos_6p0 w=0.51u l=0.6u
X12789 a_17620_18100# cap_shunt_p a_17828_18584# vdd pmos_6p0 w=1.2u l=0.5u
X12790 vss cap_shunt_n a_19152_24856# vss nmos_6p0 w=0.82u l=0.6u
X12791 a_9876_51512# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12792 a_27552_3204# cap_shunt_p a_25444_3266# vss nmos_6p0 w=0.82u l=0.6u
X12793 a_6084_17724# cap_shunt_p a_6292_17378# vdd pmos_6p0 w=1.2u l=0.5u
X12794 a_6292_50306# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12795 a_17620_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12796 a_29492_5180# tune_shunt[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12797 a_25780_43672# cap_shunt_p a_25572_43188# vdd pmos_6p0 w=1.2u l=0.5u
X12798 vdd a_27676_41143# a_27588_41240# vdd pmos_6p0 w=1.22u l=1u
X12799 a_3380_49944# cap_shunt_p a_3172_49460# vdd pmos_6p0 w=1.2u l=0.5u
X12800 vdd a_34396_14920# a_34308_14964# vdd pmos_6p0 w=1.22u l=1u
X12801 a_13796_23650# cap_shunt_n a_13588_23996# vdd pmos_6p0 w=1.2u l=0.5u
X12802 vdd a_32604_32168# a_32516_32212# vdd pmos_6p0 w=1.22u l=1u
X12803 vss tune_shunt[7] a_20740_29560# vss nmos_6p0 w=0.51u l=0.6u
X12804 a_35692_8692# cap_series_gygyn a_35880_8692# vdd pmos_6p0 w=1.2u l=0.5u
X12805 vss cap_shunt_p a_8400_49944# vss nmos_6p0 w=0.82u l=0.6u
X12806 a_17828_26424# cap_shunt_n a_17620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X12807 a_21540_17724# cap_shunt_p a_21748_17378# vdd pmos_6p0 w=1.2u l=0.5u
X12808 vdd a_33052_55688# a_32964_55732# vdd pmos_6p0 w=1.22u l=1u
X12809 vdd a_20284_54120# a_20196_54164# vdd pmos_6p0 w=1.22u l=1u
X12810 a_26444_52552# a_26356_52596# vss vss nmos_6p0 w=0.82u l=1u
X12811 a_14580_43672# cap_shunt_n a_14372_43188# vdd pmos_6p0 w=1.2u l=0.5u
X12812 vss tune_shunt[6] a_3828_37400# vss nmos_6p0 w=0.51u l=0.6u
X12813 vss cap_shunt_p a_4032_47108# vss nmos_6p0 w=0.82u l=0.6u
X12814 a_36384_45944# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X12815 vdd a_34396_11784# a_34308_11828# vdd pmos_6p0 w=1.22u l=1u
X12816 vdd tune_shunt[7] a_9668_18100# vdd pmos_6p0 w=1.2u l=0.5u
X12817 a_13460_34264# cap_shunt_n a_14392_34264# vss nmos_6p0 w=0.82u l=0.6u
X12818 vss tune_shunt[7] a_20740_26424# vss nmos_6p0 w=0.51u l=0.6u
X12819 a_35692_5556# cap_series_gygyn a_35880_5556# vdd pmos_6p0 w=1.2u l=0.5u
X12820 vdd a_35292_3511# a_35204_3608# vdd pmos_6p0 w=1.22u l=1u
X12821 a_2708_12674# cap_shunt_n a_2500_13020# vdd pmos_6p0 w=1.2u l=0.5u
X12822 a_3380_17016# cap_shunt_p a_4312_17016# vss nmos_6p0 w=0.82u l=0.6u
X12823 a_17828_23288# cap_shunt_n a_17620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X12824 vss cap_series_gyn a_30800_12312# vss nmos_6p0 w=0.82u l=0.6u
X12825 a_31624_19292# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X12826 a_17596_55255# a_17508_55352# vss vss nmos_6p0 w=0.82u l=1u
X12827 vdd a_20284_50984# a_20196_51028# vdd pmos_6p0 w=1.22u l=1u
X12828 a_36384_42808# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X12829 vss cap_shunt_p a_25984_37700# vss nmos_6p0 w=0.82u l=0.6u
X12830 a_32604_27464# a_32516_27508# vss vss nmos_6p0 w=0.82u l=1u
X12831 a_32612_26786# cap_shunt_p a_32404_27132# vdd pmos_6p0 w=1.2u l=0.5u
X12832 vdd a_30028_55688# a_29940_55732# vdd pmos_6p0 w=1.22u l=1u
X12833 vdd a_23420_52552# a_23332_52596# vdd pmos_6p0 w=1.22u l=1u
X12834 a_11668_45240# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12835 a_34328_37700# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12836 vdd tune_shunt[7] a_24452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X12837 a_1692_19624# a_1604_19668# vss vss nmos_6p0 w=0.82u l=1u
X12838 vdd a_2140_38440# a_2052_38484# vdd pmos_6p0 w=1.22u l=1u
X12839 a_37632_33781# cap_shunt_gyn a_37652_34264# vss nmos_6p0 w=0.82u l=0.6u
X12840 a_13460_31128# cap_shunt_n a_14392_31128# vss nmos_6p0 w=0.82u l=0.6u
X12841 vdd a_6508_25463# a_6420_25560# vdd pmos_6p0 w=1.22u l=1u
X12842 a_11592_12312# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12843 a_31808_34564# cap_shunt_p a_29700_34626# vss nmos_6p0 w=0.82u l=0.6u
X12844 a_8576_4772# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12845 vss tune_shunt[7] a_16708_17378# vss nmos_6p0 w=0.51u l=0.6u
X12846 vdd tune_shunt[6] a_2500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X12847 a_32604_24328# a_32516_24372# vss vss nmos_6p0 w=0.82u l=1u
X12848 a_11668_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12849 vdd tune_shunt[7] a_24452_22428# vdd pmos_6p0 w=1.2u l=0.5u
X12850 vdd a_30364_8215# a_30276_8312# vdd pmos_6p0 w=1.22u l=1u
X12851 vdd a_2140_35304# a_2052_35348# vdd pmos_6p0 w=1.22u l=1u
X12852 a_25780_23288# cap_shunt_p a_26712_23288# vss nmos_6p0 w=0.82u l=0.6u
X12853 a_3828_37400# cap_shunt_n a_4760_37400# vss nmos_6p0 w=0.82u l=0.6u
X12854 a_3828_20152# cap_shunt_p a_5544_20152# vss nmos_6p0 w=0.82u l=0.6u
X12855 a_12580_47892# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12856 a_17620_38484# cap_shunt_n a_17828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X12857 a_31808_31428# cap_shunt_p a_29700_31490# vss nmos_6p0 w=0.82u l=0.6u
X12858 vdd a_5612_55688# a_5524_55732# vdd pmos_6p0 w=1.22u l=1u
X12859 vdd tune_shunt[7] a_24452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X12860 a_27496_7608# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12861 a_10472_9476# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X12862 a_7540_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12863 a_24452_8316# cap_series_gyp a_24660_7970# vdd pmos_6p0 w=1.2u l=0.5u
X12864 a_6532_27508# cap_shunt_n a_6740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X12865 a_9668_14964# cap_shunt_p a_9876_15448# vdd pmos_6p0 w=1.2u l=0.5u
X12866 a_17620_35348# cap_shunt_n a_17828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X12867 vdd a_34844_13352# a_34756_13396# vdd pmos_6p0 w=1.22u l=1u
X12868 vss tune_shunt[4] a_3828_13880# vss nmos_6p0 w=0.51u l=0.6u
X12869 vss tune_shunt[6] a_25780_35832# vss nmos_6p0 w=0.51u l=0.6u
X12870 vdd a_32716_17623# a_32628_17720# vdd pmos_6p0 w=1.22u l=1u
X12871 vss cap_shunt_p a_19152_18584# vss nmos_6p0 w=0.82u l=0.6u
X12872 a_7540_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12873 a_12656_23288# cap_shunt_n a_10548_23288# vss nmos_6p0 w=0.82u l=0.6u
X12874 a_9220_20860# cap_shunt_p a_9428_20514# vdd pmos_6p0 w=1.2u l=0.5u
X12875 vdd a_33500_54120# a_33412_54164# vdd pmos_6p0 w=1.22u l=1u
X12876 a_35264_47512# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X12877 a_35600_46870# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12878 vdd tune_shunt[5] a_2500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X12879 vdd tune_shunt_gy[2] a_37444_41621# vdd pmos_6p0 w=1.215u l=0.5u
X12880 a_1924_6040# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X12881 a_20328_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12882 a_11780_4472# cap_series_gyp a_11572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X12883 a_9668_11828# cap_shunt_p a_9876_12312# vdd pmos_6p0 w=1.2u l=0.5u
X12884 a_25780_43672# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X12885 a_17640_23588# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12886 a_18404_11452# cap_series_gyn a_18612_11106# vdd pmos_6p0 w=1.2u l=0.5u
X12887 a_32612_36194# cap_shunt_n a_33544_36132# vss nmos_6p0 w=0.82u l=0.6u
X12888 a_10660_33058# cap_shunt_n a_12376_32996# vss nmos_6p0 w=0.82u l=0.6u
X12889 a_7580_8316# cap_series_gyn a_7768_8316# vdd pmos_6p0 w=1.2u l=0.5u
X12890 vss cap_shunt_p a_19152_15448# vss nmos_6p0 w=0.82u l=0.6u
X12891 vdd a_33500_50984# a_33412_51028# vdd pmos_6p0 w=1.22u l=1u
X12892 vdd a_8860_16488# a_8772_16532# vdd pmos_6p0 w=1.22u l=1u
X12893 a_24452_13020# cap_series_gyn a_24660_12674# vdd pmos_6p0 w=1.2u l=0.5u
X12894 vdd tune_shunt[5] a_3620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X12895 a_25780_40536# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X12896 a_6572_5556# cap_series_gyp a_6760_5556# vdd pmos_6p0 w=1.2u l=0.5u
X12897 a_6292_18946# cap_shunt_p a_6084_19292# vdd pmos_6p0 w=1.2u l=0.5u
X12898 vdd a_25996_52552# a_25908_52596# vdd pmos_6p0 w=1.22u l=1u
X12899 a_6196_47516# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12900 vdd tune_series_gy[4] a_18516_5556# vdd pmos_6p0 w=1.2u l=0.5u
X12901 a_13796_14242# cap_shunt_p a_13588_14588# vdd pmos_6p0 w=1.2u l=0.5u
X12902 a_25100_47415# a_25012_47512# vss vss nmos_6p0 w=0.82u l=1u
X12903 vdd tune_shunt[6] a_3620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X12904 a_6292_15810# cap_shunt_p a_6084_16156# vdd pmos_6p0 w=1.2u l=0.5u
X12905 a_17828_17016# cap_shunt_p a_17620_16532# vdd pmos_6p0 w=1.2u l=0.5u
X12906 a_24452_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12907 vdd a_30028_49416# a_29940_49460# vdd pmos_6p0 w=1.22u l=1u
X12908 a_32404_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12909 vdd a_15804_19624# a_15716_19668# vdd pmos_6p0 w=1.22u l=1u
X12910 vdd tune_series_gy[4] a_24452_19292# vdd pmos_6p0 w=1.2u l=0.5u
X12911 a_20740_34264# cap_shunt_n a_20532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X12912 a_37652_50244# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12913 vss tune_shunt[4] a_20740_17016# vss nmos_6p0 w=0.51u l=0.6u
X12914 a_19388_50984# a_19300_51028# vss vss nmos_6p0 w=0.82u l=1u
X12915 vss cap_shunt_n a_22064_35832# vss nmos_6p0 w=0.82u l=0.6u
X12916 a_6760_5556# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X12917 a_31808_28292# cap_shunt_p a_29700_28354# vss nmos_6p0 w=0.82u l=0.6u
X12918 vdd tune_series_gygy[5] a_35692_24372# vdd pmos_6p0 w=1.2u l=0.5u
X12919 a_19732_13880# cap_series_gyn a_20664_13880# vss nmos_6p0 w=0.82u l=0.6u
X12920 vdd a_32156_18056# a_32068_18100# vdd pmos_6p0 w=1.22u l=1u
X12921 a_32604_18056# a_32516_18100# vss vss nmos_6p0 w=0.82u l=1u
X12922 vdd a_30028_46280# a_29940_46324# vdd pmos_6p0 w=1.22u l=1u
X12923 a_20532_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12924 a_22680_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X12925 a_11460_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12926 vdd a_2140_29032# a_2052_29076# vdd pmos_6p0 w=1.22u l=1u
X12927 vdd tune_series_gy[5] a_24452_16156# vdd pmos_6p0 w=1.2u l=0.5u
X12928 a_16028_32168# a_15940_32212# vss vss nmos_6p0 w=0.82u l=1u
X12929 a_20740_31128# cap_shunt_n a_20532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X12930 a_25780_43672# cap_shunt_p a_25572_43188# vdd pmos_6p0 w=1.2u l=0.5u
X12931 vdd tune_series_gy[4] a_28484_18100# vdd pmos_6p0 w=1.2u l=0.5u
X12932 vdd a_28236_53687# a_28148_53784# vdd pmos_6p0 w=1.22u l=1u
X12933 a_30016_7608# cap_series_gyp a_28692_7608# vss nmos_6p0 w=0.82u l=0.6u
X12934 a_23308_53687# a_23220_53784# vss vss nmos_6p0 w=0.82u l=1u
X12935 a_4424_50244# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X12936 a_31808_25156# cap_shunt_p a_29700_25218# vss nmos_6p0 w=0.82u l=0.6u
X12937 vss tune_series_gy[2] a_6760_7124# vss nmos_6p0 w=0.51u l=0.6u
X12938 a_37980_54120# a_37892_54164# vss vss nmos_6p0 w=0.82u l=1u
X12939 a_10548_3266# cap_series_gyn a_10340_3612# vdd pmos_6p0 w=1.2u l=0.5u
X12940 a_19732_10744# cap_series_gyn a_20664_10744# vss nmos_6p0 w=0.82u l=0.6u
X12941 a_32604_14920# a_32516_14964# vss vss nmos_6p0 w=0.82u l=1u
X12942 vdd tune_series_gygy[5] a_35692_21236# vdd pmos_6p0 w=1.2u l=0.5u
X12943 a_20532_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12944 a_6572_7124# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12945 vdd a_33612_39575# a_33524_39672# vdd pmos_6p0 w=1.22u l=1u
X12946 vss tune_shunt[7] a_13460_37400# vss nmos_6p0 w=0.51u l=0.6u
X12947 a_2932_12312# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X12948 a_14580_43672# cap_shunt_n a_14372_43188# vdd pmos_6p0 w=1.2u l=0.5u
X12949 a_35292_21192# a_35204_21236# vss vss nmos_6p0 w=0.82u l=1u
X12950 vdd a_28236_50551# a_28148_50648# vdd pmos_6p0 w=1.22u l=1u
X12951 a_12108_53687# a_12020_53784# vss vss nmos_6p0 w=0.82u l=1u
X12952 a_23308_50551# a_23220_50648# vss vss nmos_6p0 w=0.82u l=1u
X12953 a_5152_43672# cap_shunt_p a_3828_43672# vss nmos_6p0 w=0.82u l=0.6u
X12954 a_17620_29076# cap_shunt_n a_17828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X12955 a_5612_5079# a_5524_5176# vss vss nmos_6p0 w=0.82u l=1u
X12956 vdd tune_series_gy[0] a_29196_3612# vdd pmos_6p0 w=1.2u l=0.5u
X12957 vss tune_shunt[7] a_25780_29560# vss nmos_6p0 w=0.51u l=0.6u
X12958 a_10660_6402# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X12959 a_9876_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12960 a_22848_4472# cap_series_gyn a_21524_4472# vss nmos_6p0 w=0.82u l=0.6u
X12961 a_15904_45540# cap_shunt_p a_13796_45602# vss nmos_6p0 w=0.82u l=0.6u
X12962 a_7540_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12963 vss tune_shunt[6] a_13796_42466# vss nmos_6p0 w=0.51u l=0.6u
X12964 a_11872_38968# cap_shunt_n a_10548_38968# vss nmos_6p0 w=0.82u l=0.6u
X12965 vdd a_10092_8648# a_10004_8692# vdd pmos_6p0 w=1.22u l=1u
X12966 a_5152_40536# cap_shunt_n a_3828_40536# vss nmos_6p0 w=0.82u l=0.6u
X12967 vss tune_shunt[7] a_25780_26424# vss nmos_6p0 w=0.51u l=0.6u
X12968 a_26376_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X12969 a_9876_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12970 a_35448_17316# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X12971 a_13588_13020# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X12972 vdd a_13676_54120# a_13588_54164# vdd pmos_6p0 w=1.22u l=1u
X12973 a_35692_25940# cap_series_gygyp a_35880_25940# vdd pmos_6p0 w=1.2u l=0.5u
X12974 a_19836_52552# a_19748_52596# vss vss nmos_6p0 w=0.82u l=1u
X12975 a_15904_42404# cap_shunt_n a_13796_42466# vss nmos_6p0 w=0.82u l=0.6u
X12976 a_2588_50984# a_2500_51028# vss vss nmos_6p0 w=0.82u l=1u
X12977 vdd a_1692_25896# a_1604_25940# vdd pmos_6p0 w=1.22u l=1u
X12978 vdd tune_shunt[6] a_2500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X12979 vss cap_shunt_n a_35840_35832# vss nmos_6p0 w=0.82u l=0.6u
X12980 vdd a_10092_5512# a_10004_5556# vdd pmos_6p0 w=1.22u l=1u
X12981 vss cap_series_gyn a_29800_3204# vss nmos_6p0 w=0.82u l=0.6u
X12982 a_20740_21720# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X12983 a_25780_34264# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X12984 a_14692_4472# cap_series_gyp a_16408_4472# vss nmos_6p0 w=0.82u l=0.6u
X12985 a_1692_8648# a_1604_8692# vss vss nmos_6p0 w=0.82u l=1u
X12986 a_4256_12312# cap_shunt_n a_2932_12312# vss nmos_6p0 w=0.82u l=0.6u
X12987 a_10660_23650# cap_shunt_n a_12376_23588# vss nmos_6p0 w=0.82u l=0.6u
X12988 a_30476_52552# a_30388_52596# vss vss nmos_6p0 w=0.82u l=1u
X12989 vdd a_26892_47415# a_26804_47512# vdd pmos_6p0 w=1.22u l=1u
X12990 a_35692_22804# cap_series_gygyp a_35880_22804# vdd pmos_6p0 w=1.2u l=0.5u
X12991 vdd a_15244_55688# a_15156_55732# vdd pmos_6p0 w=1.22u l=1u
X12992 a_4816_48676# cap_shunt_p a_2708_48738# vss nmos_6p0 w=0.82u l=0.6u
X12993 vdd tune_shunt[7] a_13252_38484# vdd pmos_6p0 w=1.2u l=0.5u
X12994 vdd a_1692_22760# a_1604_22804# vdd pmos_6p0 w=1.22u l=1u
X12995 a_32464_44757# cap_shunt_gyp a_32464_45302# vdd pmos_6p0 w=1.215u l=0.5u
X12996 a_3828_40536# cap_shunt_n a_3620_40052# vdd pmos_6p0 w=1.2u l=0.5u
X12997 vdd tune_series_gy[1] a_7580_5180# vdd pmos_6p0 w=1.2u l=0.5u
X12998 vdd tune_shunt[6] a_6532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X12999 vdd tune_shunt[6] a_3620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X13000 a_25780_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13001 a_5096_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13002 vdd a_17820_3511# a_17732_3608# vdd pmos_6p0 w=1.22u l=1u
X13003 vdd tune_series_gygy[4] a_34308_13020# vdd pmos_6p0 w=1.2u l=0.5u
X13004 a_28124_12919# a_28036_13016# vss vss nmos_6p0 w=0.82u l=1u
X13005 a_36296_20152# cap_series_gygyp a_35880_19668# vss nmos_6p0 w=0.82u l=0.6u
X13006 a_21748_34626# cap_shunt_p a_21540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X13007 vdd tune_shunt[7] a_13252_35348# vdd pmos_6p0 w=1.2u l=0.5u
X13008 vss tune_series_gy[0] a_28692_4472# vss nmos_6p0 w=0.51u l=0.6u
X13009 vdd tune_shunt[6] a_3620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X13010 vss cap_shunt_n a_22064_29560# vss nmos_6p0 w=0.82u l=0.6u
X13011 vdd tune_series_gy[4] a_11612_8692# vdd pmos_6p0 w=1.2u l=0.5u
X13012 vdd a_24540_3944# a_24452_3988# vdd pmos_6p0 w=1.22u l=1u
X13013 a_25660_55688# a_25572_55732# vss vss nmos_6p0 w=0.82u l=1u
X13014 a_21748_31490# cap_shunt_n a_21540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X13015 a_20740_24856# cap_shunt_n a_20532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X13016 vss cap_shunt_p a_8400_51812# vss nmos_6p0 w=0.82u l=0.6u
X13017 a_16500_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13018 vss cap_shunt_n a_22064_26424# vss nmos_6p0 w=0.82u l=0.6u
X13019 a_29700_33058# cap_shunt_p a_30632_32996# vss nmos_6p0 w=0.82u l=0.6u
X13020 a_20532_16532# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13021 vss tune_series_gygy[2] a_35880_5556# vss nmos_6p0 w=0.51u l=0.6u
X13022 a_8848_21720# cap_shunt_p a_6740_21720# vss nmos_6p0 w=0.82u l=0.6u
X13023 a_6292_18946# cap_shunt_p a_6084_19292# vdd pmos_6p0 w=1.2u l=0.5u
X13024 a_22636_55688# a_22548_55732# vss vss nmos_6p0 w=0.82u l=1u
X13025 a_10452_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13026 a_16028_22760# a_15940_22804# vss vss nmos_6p0 w=0.82u l=1u
X13027 a_20740_21720# cap_shunt_p a_20532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X13028 a_16500_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13029 a_26712_37400# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13030 vss tune_shunt[4] a_2708_12674# vss nmos_6p0 w=0.51u l=0.6u
X13031 a_34516_17378# cap_series_gygyn a_36232_17316# vss nmos_6p0 w=0.82u l=0.6u
X13032 a_13588_17724# cap_shunt_p a_13796_17378# vdd pmos_6p0 w=1.2u l=0.5u
X13033 a_21748_7970# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13034 vss tune_shunt[5] a_12788_20152# vss nmos_6p0 w=0.51u l=0.6u
X13035 vdd a_14012_9783# a_13924_9880# vdd pmos_6p0 w=1.22u l=1u
X13036 a_6292_15810# cap_shunt_p a_6084_16156# vdd pmos_6p0 w=1.2u l=0.5u
X13037 vss tune_shunt[3] a_5844_10744# vss nmos_6p0 w=0.51u l=0.6u
X13038 a_21540_38108# cap_shunt_n a_21748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X13039 a_3620_33780# cap_shunt_n a_3828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X13040 a_35292_11784# a_35204_11828# vss vss nmos_6p0 w=0.82u l=1u
X13041 vdd a_2140_55255# a_2052_55352# vdd pmos_6p0 w=1.22u l=1u
X13042 vss tune_shunt[7] a_13796_36194# vss nmos_6p0 w=0.51u l=0.6u
X13043 vss tune_series_gy[3] a_29720_9884# vss nmos_6p0 w=0.51u l=0.6u
X13044 a_5152_34264# cap_shunt_n a_3828_34264# vss nmos_6p0 w=0.82u l=0.6u
X13045 a_33524_32212# cap_shunt_n a_33732_32696# vdd pmos_6p0 w=1.2u l=0.5u
X13046 a_21748_4834# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13047 vdd a_14012_6647# a_13924_6744# vdd pmos_6p0 w=1.22u l=1u
X13048 vdd a_26444_49416# a_26356_49460# vdd pmos_6p0 w=1.22u l=1u
X13049 a_15904_36132# cap_shunt_n a_13796_36194# vss nmos_6p0 w=0.82u l=0.6u
X13050 vss cap_shunt_p a_11984_18584# vss nmos_6p0 w=0.82u l=0.6u
X13051 a_24452_42812# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13052 a_2588_44712# a_2500_44756# vss vss nmos_6p0 w=0.82u l=1u
X13053 a_3620_30644# cap_shunt_n a_3828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X13054 vss cap_shunt_p a_35840_29560# vss nmos_6p0 w=0.82u l=0.6u
X13055 vdd tune_series_gygy[5] a_35692_24372# vdd pmos_6p0 w=1.2u l=0.5u
X13056 a_34844_55255# a_34756_55352# vss vss nmos_6p0 w=0.82u l=1u
X13057 vdd a_2140_52119# a_2052_52216# vdd pmos_6p0 w=1.22u l=1u
X13058 a_30632_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13059 vss tune_shunt[7] a_13796_33058# vss nmos_6p0 w=0.51u l=0.6u
X13060 vdd a_6956_31735# a_6868_31832# vdd pmos_6p0 w=1.22u l=1u
X13061 a_11800_7124# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X13062 a_5152_31128# cap_shunt_n a_3828_31128# vss nmos_6p0 w=0.82u l=0.6u
X13063 a_14112_12312# cap_shunt_p a_12788_12312# vss nmos_6p0 w=0.82u l=0.6u
X13064 vss cap_series_gygyp a_36296_37400# vss nmos_6p0 w=0.82u l=0.6u
X13065 vss tune_series_gy[5] a_25780_17016# vss nmos_6p0 w=0.51u l=0.6u
X13066 a_33524_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13067 a_18044_5512# a_17956_5556# vss vss nmos_6p0 w=0.82u l=1u
X13068 vss cap_shunt_n a_5152_13880# vss nmos_6p0 w=0.82u l=0.6u
X13069 vdd tune_series_gy[4] a_28484_18100# vdd pmos_6p0 w=1.2u l=0.5u
X13070 vdd a_26444_46280# a_26356_46324# vdd pmos_6p0 w=1.22u l=1u
X13071 vss cap_shunt_p a_11984_15448# vss nmos_6p0 w=0.82u l=0.6u
X13072 a_35692_16532# cap_series_gygyn a_35880_16532# vdd pmos_6p0 w=1.2u l=0.5u
X13073 vss tune_shunt[4] a_33732_32696# vss nmos_6p0 w=0.51u l=0.6u
X13074 a_5636_3612# cap_shunt_n a_5844_3266# vdd pmos_6p0 w=1.2u l=0.5u
X13075 a_2588_41576# a_2500_41620# vss vss nmos_6p0 w=0.82u l=1u
X13076 a_1716_6748# cap_shunt_n a_1924_6402# vdd pmos_6p0 w=1.2u l=0.5u
X13077 vdd a_1692_16488# a_1604_16532# vdd pmos_6p0 w=1.22u l=1u
X13078 vdd tune_series_gygy[5] a_35692_21236# vdd pmos_6p0 w=1.2u l=0.5u
X13079 a_2140_33303# a_2052_33400# vss vss nmos_6p0 w=0.82u l=1u
X13080 vdd tune_shunt[4] a_29492_39676# vdd pmos_6p0 w=1.2u l=0.5u
X13081 a_4816_39268# cap_shunt_n a_2708_39330# vss nmos_6p0 w=0.82u l=0.6u
X13082 vdd tune_shunt[7] a_13252_29076# vdd pmos_6p0 w=1.2u l=0.5u
X13083 vss cap_shunt_p a_15904_12612# vss nmos_6p0 w=0.82u l=0.6u
X13084 vdd a_35292_53687# a_35204_53784# vdd pmos_6p0 w=1.22u l=1u
X13085 a_30364_53687# a_30276_53784# vss vss nmos_6p0 w=0.82u l=1u
X13086 a_24660_18946# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13087 vdd tune_shunt[7] a_3620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X13088 a_29700_17378# cap_series_gyp a_29492_17724# vdd pmos_6p0 w=1.2u l=0.5u
X13089 a_16708_29922# cap_shunt_n a_18424_29860# vss nmos_6p0 w=0.82u l=0.6u
X13090 a_28692_4472# cap_series_gyp a_28484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X13091 vdd tune_series_gy[2] a_6572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X13092 a_36688_9176# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X13093 a_17620_33780# cap_shunt_n a_17828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X13094 a_26768_29860# cap_shunt_n a_24660_29922# vss nmos_6p0 w=0.82u l=0.6u
X13095 a_16708_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13096 a_21748_25218# cap_shunt_n a_21540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X13097 a_29492_5180# cap_shunt_p a_29700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X13098 vdd tune_series_gygy[5] a_30428_19668# vdd pmos_6p0 w=1.2u l=0.5u
X13099 a_22064_45240# cap_shunt_n a_20740_45240# vss nmos_6p0 w=0.82u l=0.6u
X13100 vss cap_shunt_p a_4816_18884# vss nmos_6p0 w=0.82u l=0.6u
X13101 vdd a_35292_50551# a_35204_50648# vdd pmos_6p0 w=1.22u l=1u
X13102 a_30364_50551# a_30276_50648# vss vss nmos_6p0 w=0.82u l=1u
X13103 vss tune_shunt[7] a_6516_20514# vss nmos_6p0 w=0.51u l=0.6u
X13104 a_16708_26786# cap_shunt_n a_18424_26724# vss nmos_6p0 w=0.82u l=0.6u
X13105 vdd tune_shunt[1] a_25236_3612# vdd pmos_6p0 w=1.2u l=0.5u
X13106 a_26768_26724# cap_shunt_p a_24660_26786# vss nmos_6p0 w=0.82u l=0.6u
X13107 a_19276_45847# a_19188_45944# vss vss nmos_6p0 w=0.82u l=1u
X13108 a_17620_30644# cap_shunt_n a_17828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X13109 a_21748_22082# cap_shunt_p a_21540_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13110 a_28124_5079# a_28036_5176# vss vss nmos_6p0 w=0.82u l=1u
X13111 a_22064_42104# cap_shunt_p a_20740_42104# vss nmos_6p0 w=0.82u l=0.6u
X13112 vss tune_shunt[7] a_6740_32696# vss nmos_6p0 w=0.51u l=0.6u
X13113 vss cap_shunt_p a_4816_15748# vss nmos_6p0 w=0.82u l=0.6u
X13114 a_2500_49084# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13115 vdd tune_shunt[7] a_16500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X13116 a_9876_13880# cap_shunt_p a_9668_13396# vdd pmos_6p0 w=1.2u l=0.5u
X13117 vdd tune_shunt[7] a_12580_13396# vdd pmos_6p0 w=1.2u l=0.5u
X13118 vss cap_shunt_p a_22064_17016# vss nmos_6p0 w=0.82u l=0.6u
X13119 a_9668_47892# cap_shunt_p a_9876_48376# vdd pmos_6p0 w=1.2u l=0.5u
X13120 a_9668_47892# cap_shunt_p a_9876_48376# vdd pmos_6p0 w=1.2u l=0.5u
X13121 vss cap_shunt_p a_23856_45540# vss nmos_6p0 w=0.82u l=0.6u
X13122 a_29700_23650# cap_shunt_p a_30632_23588# vss nmos_6p0 w=0.82u l=0.6u
X13123 vdd a_3036_13352# a_2948_13396# vdd pmos_6p0 w=1.22u l=1u
X13124 a_21748_28354# cap_shunt_n a_21540_28700# vdd pmos_6p0 w=1.2u l=0.5u
X13125 vss cap_series_gygyp a_36296_4472# vss nmos_6p0 w=0.82u l=0.6u
X13126 a_26892_52552# a_26804_52596# vss vss nmos_6p0 w=0.82u l=1u
X13127 a_3828_46808# cap_shunt_p a_3620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X13128 a_19276_42711# a_19188_42808# vss vss nmos_6p0 w=0.82u l=1u
X13129 a_8848_12312# cap_shunt_p a_6740_12312# vss nmos_6p0 w=0.82u l=0.6u
X13130 vdd a_2140_48983# a_2052_49080# vdd pmos_6p0 w=1.22u l=1u
X13131 a_22644_12312# cap_series_gyn a_22436_11828# vdd pmos_6p0 w=1.2u l=0.5u
X13132 a_24660_40898# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13133 vss cap_shunt_p a_8848_46808# vss nmos_6p0 w=0.82u l=0.6u
X13134 vss tune_shunt[7] a_2708_26786# vss nmos_6p0 w=0.51u l=0.6u
X13135 a_9108_22428# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13136 a_34516_12674# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13137 vss cap_shunt_n a_23856_42404# vss nmos_6p0 w=0.82u l=0.6u
X13138 vdd a_30476_55688# a_30388_55732# vdd pmos_6p0 w=1.22u l=1u
X13139 a_23868_52552# a_23780_52596# vss vss nmos_6p0 w=0.82u l=1u
X13140 a_7580_6748# cap_series_gyp a_7768_6748# vdd pmos_6p0 w=1.2u l=0.5u
X13141 a_24452_36540# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13142 a_36160_45302# cap_shunt_gyn a_36160_44757# vdd pmos_6p0 w=1.215u l=0.5u
X13143 a_23072_43972# cap_shunt_n a_21748_44034# vss nmos_6p0 w=0.82u l=0.6u
X13144 a_29492_34972# cap_shunt_p a_29700_34626# vdd pmos_6p0 w=1.2u l=0.5u
X13145 vdd a_6956_25463# a_6868_25560# vdd pmos_6p0 w=1.22u l=1u
X13146 a_3620_24372# cap_shunt_p a_3828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X13147 a_21748_15810# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13148 vdd a_4828_53687# a_4740_53784# vdd pmos_6p0 w=1.22u l=1u
X13149 a_36300_32168# a_36212_32212# vss vss nmos_6p0 w=0.82u l=1u
X13150 vss cap_shunt_p a_23072_18884# vss nmos_6p0 w=0.82u l=0.6u
X13151 a_22436_8692# cap_series_gyp a_22644_9176# vdd pmos_6p0 w=1.2u l=0.5u
X13152 a_33052_41143# a_32964_41240# vss vss nmos_6p0 w=0.82u l=1u
X13153 a_25780_9176# cap_series_gyp a_25572_8692# vdd pmos_6p0 w=1.2u l=0.5u
X13154 a_36624_20452# cap_series_gygyp a_34516_20514# vss nmos_6p0 w=0.82u l=0.6u
X13155 a_36636_50984# a_36548_51028# vss vss nmos_6p0 w=0.82u l=1u
X13156 a_24452_33404# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13157 a_16700_16488# a_16612_16532# vss vss nmos_6p0 w=0.82u l=1u
X13158 a_34144_45944# cap_shunt_gyn a_34144_45540# vdd pmos_6p0 w=1.215u l=0.5u
X13159 a_6740_45240# cap_shunt_p a_8456_45240# vss nmos_6p0 w=0.82u l=0.6u
X13160 a_23072_40836# cap_shunt_p a_21748_40898# vss nmos_6p0 w=0.82u l=0.6u
X13161 a_29492_31836# cap_shunt_p a_29700_31490# vdd pmos_6p0 w=1.2u l=0.5u
X13162 a_15700_9538# cap_series_gyn a_15492_9884# vdd pmos_6p0 w=1.2u l=0.5u
X13163 a_3620_21236# cap_shunt_p a_3828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X13164 a_3620_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13165 a_35880_24372# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13166 vss cap_series_gyn a_17808_4772# vss nmos_6p0 w=0.82u l=0.6u
X13167 vss cap_series_gyn a_23072_15748# vss nmos_6p0 w=0.82u l=0.6u
X13168 a_6292_18946# cap_shunt_p a_6084_19292# vdd pmos_6p0 w=1.2u l=0.5u
X13169 vss tune_shunt[7] a_10548_27992# vss nmos_6p0 w=0.51u l=0.6u
X13170 a_6628_14242# cap_shunt_p a_6420_14588# vdd pmos_6p0 w=1.2u l=0.5u
X13171 vdd tune_shunt[5] a_20532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X13172 a_19524_7124# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13173 a_25780_6040# cap_series_gyp a_25572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X13174 a_1924_7970# cap_shunt_n a_3640_7908# vss nmos_6p0 w=0.82u l=0.6u
X13175 a_14504_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13176 a_12376_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13177 a_34144_42808# cap_shunt_gyn a_34144_42404# vdd pmos_6p0 w=1.215u l=0.5u
X13178 a_6740_42104# cap_shunt_n a_8456_42104# vss nmos_6p0 w=0.82u l=0.6u
X13179 a_3828_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13180 a_2140_23895# a_2052_23992# vss vss nmos_6p0 w=0.82u l=1u
X13181 a_15700_6402# cap_series_gyp a_15492_6748# vdd pmos_6p0 w=1.2u l=0.5u
X13182 vdd tune_shunt[0] a_29492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X13183 a_6292_15810# cap_shunt_p a_6084_16156# vdd pmos_6p0 w=1.2u l=0.5u
X13184 vdd a_20396_47848# a_20308_47892# vdd pmos_6p0 w=1.22u l=1u
X13185 a_17828_46808# cap_shunt_n a_17620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X13186 a_7672_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13187 a_21540_38108# cap_shunt_n a_21748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X13188 vss tune_shunt[7] a_10548_24856# vss nmos_6p0 w=0.51u l=0.6u
X13189 vdd a_28572_8215# a_28484_8312# vdd pmos_6p0 w=1.22u l=1u
X13190 a_22644_7608# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13191 a_21056_9176# cap_series_gyp a_19732_9176# vss nmos_6p0 w=0.82u l=0.6u
X13192 a_14236_50984# a_14148_51028# vss vss nmos_6p0 w=0.82u l=1u
X13193 a_5612_44279# a_5524_44376# vss vss nmos_6p0 w=0.82u l=1u
X13194 a_33524_32212# cap_shunt_n a_33732_32696# vdd pmos_6p0 w=1.2u l=0.5u
X13195 vdd tune_shunt[7] a_13252_25940# vdd pmos_6p0 w=1.2u l=0.5u
X13196 a_21748_18946# cap_shunt_p a_21540_19292# vdd pmos_6p0 w=1.2u l=0.5u
X13197 vss tune_shunt[7] a_17828_20152# vss nmos_6p0 w=0.51u l=0.6u
X13198 a_37080_23288# cap_series_gygyp a_35880_22804# vss nmos_6p0 w=0.82u l=0.6u
X13199 vss tune_shunt[6] a_17828_43672# vss nmos_6p0 w=0.51u l=0.6u
X13200 a_25572_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13201 a_22848_27992# cap_shunt_n a_20740_27992# vss nmos_6p0 w=0.82u l=0.6u
X13202 vss cap_shunt_n a_19936_37400# vss nmos_6p0 w=0.82u l=0.6u
X13203 a_21540_8316# cap_series_gyp a_21748_7970# vdd pmos_6p0 w=1.2u l=0.5u
X13204 vdd a_35292_8648# a_35204_8692# vdd pmos_6p0 w=1.22u l=1u
X13205 a_6172_54120# a_6084_54164# vss vss nmos_6p0 w=0.82u l=1u
X13206 a_7672_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13207 a_6532_46324# cap_shunt_p a_6740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X13208 a_17620_24372# cap_shunt_n a_17828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X13209 a_5612_41143# a_5524_41240# vss vss nmos_6p0 w=0.82u l=1u
X13210 vdd tune_shunt[7] a_13252_22804# vdd pmos_6p0 w=1.2u l=0.5u
X13211 a_21748_15810# cap_series_gyn a_21540_16156# vdd pmos_6p0 w=1.2u l=0.5u
X13212 a_16708_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13213 a_11800_8692# cap_series_gyp a_11824_9176# vss nmos_6p0 w=0.82u l=0.6u
X13214 a_28484_7124# cap_series_gyp a_28692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X13215 a_25780_18584# cap_series_gyn a_25572_18100# vdd pmos_6p0 w=1.2u l=0.5u
X13216 a_7748_44034# cap_shunt_p a_9464_43972# vss nmos_6p0 w=0.82u l=0.6u
X13217 vss tune_shunt[6] a_17828_40536# vss nmos_6p0 w=0.51u l=0.6u
X13218 a_10548_27992# cap_shunt_n a_11480_27992# vss nmos_6p0 w=0.82u l=0.6u
X13219 a_22848_24856# cap_shunt_n a_20740_24856# vss nmos_6p0 w=0.82u l=0.6u
X13220 vdd a_30924_54120# a_30836_54164# vdd pmos_6p0 w=1.22u l=1u
X13221 vdd a_35292_5512# a_35204_5556# vdd pmos_6p0 w=1.22u l=1u
X13222 a_21540_5180# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13223 a_18404_8316# cap_series_gyp a_18612_7970# vdd pmos_6p0 w=1.2u l=0.5u
X13224 a_16708_17378# cap_shunt_p a_18424_17316# vss nmos_6p0 w=0.82u l=0.6u
X13225 vdd tune_series_gy[5] a_25572_14964# vdd pmos_6p0 w=1.2u l=0.5u
X13226 a_26768_17316# cap_series_gyp a_24660_17378# vss nmos_6p0 w=0.82u l=0.6u
X13227 vdd a_29244_41576# a_29156_41620# vdd pmos_6p0 w=1.22u l=1u
X13228 a_13796_28354# cap_shunt_n a_13588_28700# vdd pmos_6p0 w=1.2u l=0.5u
X13229 a_21748_20514# cap_shunt_p a_21540_20860# vdd pmos_6p0 w=1.2u l=0.5u
X13230 a_17620_21236# cap_shunt_p a_17828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X13231 a_19276_36439# a_19188_36536# vss vss nmos_6p0 w=0.82u l=1u
X13232 vss tune_shunt[7] a_6740_23288# vss nmos_6p0 w=0.51u l=0.6u
X13233 a_35880_7124# cap_series_gygyp a_35692_7124# vdd pmos_6p0 w=1.2u l=0.5u
X13234 vdd a_19836_49416# a_19748_49460# vdd pmos_6p0 w=1.22u l=1u
X13235 a_7748_40898# cap_shunt_n a_9464_40836# vss nmos_6p0 w=0.82u l=0.6u
X13236 a_10548_24856# cap_shunt_n a_11480_24856# vss nmos_6p0 w=0.82u l=0.6u
X13237 vdd a_30924_50984# a_30836_51028# vdd pmos_6p0 w=1.22u l=1u
X13238 a_33024_47512# cap_shunt_gyn a_33024_47108# vdd pmos_6p0 w=1.215u l=0.5u
X13239 a_3640_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13240 vss cap_shunt_n a_23856_36132# vss nmos_6p0 w=0.82u l=0.6u
X13241 a_5636_8692# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13242 vdd tune_series_gy[5] a_25572_11828# vdd pmos_6p0 w=1.2u l=0.5u
X13243 a_17828_20152# cap_shunt_p a_18760_20152# vss nmos_6p0 w=0.82u l=0.6u
X13244 vdd a_30476_49416# a_30388_49460# vdd pmos_6p0 w=1.22u l=1u
X13245 a_36428_43672# cap_shunt_gyn a_36160_43734# vss nmos_6p0 w=0.82u l=0.6u
X13246 a_10548_37400# cap_shunt_n a_12264_37400# vss nmos_6p0 w=0.82u l=0.6u
X13247 a_35880_22804# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13248 a_29700_17378# cap_series_gyp a_29492_17724# vdd pmos_6p0 w=1.2u l=0.5u
X13249 a_5844_3266# cap_shunt_n a_6776_3204# vss nmos_6p0 w=0.82u l=0.6u
X13250 a_8736_12612# cap_shunt_p a_6628_12674# vss nmos_6p0 w=0.82u l=0.6u
X13251 vss tune_shunt[5] a_6292_18584# vss nmos_6p0 w=0.51u l=0.6u
X13252 a_31260_13352# a_31172_13396# vss vss nmos_6p0 w=0.82u l=1u
X13253 vdd tune_series_gygy[5] a_30428_19668# vdd pmos_6p0 w=1.2u l=0.5u
X13254 a_21180_49416# a_21092_49460# vss vss nmos_6p0 w=0.82u l=1u
X13255 vss tune_shunt[7] a_2708_17378# vss nmos_6p0 w=0.51u l=0.6u
X13256 a_10548_3266# cap_series_gyn a_10340_3612# vdd pmos_6p0 w=1.2u l=0.5u
X13257 a_33500_3944# a_33412_3988# vss vss nmos_6p0 w=0.82u l=1u
X13258 vdd a_30476_46280# a_30388_46324# vdd pmos_6p0 w=1.22u l=1u
X13259 a_3380_51512# cap_shunt_n a_4312_51512# vss nmos_6p0 w=0.82u l=0.6u
X13260 a_24452_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13261 vdd tune_shunt[7] a_17620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X13262 a_23072_34564# cap_shunt_p a_21748_34626# vss nmos_6p0 w=0.82u l=0.6u
X13263 a_20532_41620# cap_shunt_p a_20740_42104# vdd pmos_6p0 w=1.2u l=0.5u
X13264 a_16476_32168# a_16388_32212# vss vss nmos_6p0 w=0.82u l=1u
X13265 a_29492_25564# cap_shunt_p a_29700_25218# vdd pmos_6p0 w=1.2u l=0.5u
X13266 a_35880_18100# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13267 a_11480_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13268 a_31260_10216# a_31172_10260# vss vss nmos_6p0 w=0.82u l=1u
X13269 a_19732_13880# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13270 a_6292_17016# cap_shunt_p a_6084_16532# vdd pmos_6p0 w=1.2u l=0.5u
X13271 vdd a_28684_53687# a_28596_53784# vdd pmos_6p0 w=1.22u l=1u
X13272 a_23756_53687# a_23668_53784# vss vss nmos_6p0 w=0.82u l=1u
X13273 a_6740_34264# cap_shunt_n a_6532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X13274 vdd tune_shunt[7] a_16500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X13275 a_29700_4834# cap_shunt_p a_29492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X13276 a_28484_14964# cap_series_gyn a_28692_15448# vdd pmos_6p0 w=1.2u l=0.5u
X13277 a_13796_50306# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13278 a_10452_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13279 a_9876_13880# cap_shunt_p a_9668_13396# vdd pmos_6p0 w=1.2u l=0.5u
X13280 vdd tune_shunt[7] a_17620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X13281 vss tune_shunt[5] a_21748_44034# vss nmos_6p0 w=0.51u l=0.6u
X13282 a_10548_38968# cap_shunt_n a_10340_38484# vdd pmos_6p0 w=1.2u l=0.5u
X13283 a_23072_31428# cap_shunt_n a_21748_31490# vss nmos_6p0 w=0.82u l=0.6u
X13284 a_1924_7608# cap_shunt_n a_1716_7124# vdd pmos_6p0 w=1.2u l=0.5u
X13285 a_19732_10744# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13286 a_35880_14964# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13287 a_12556_53687# a_12468_53784# vss vss nmos_6p0 w=0.82u l=1u
X13288 vdd a_28684_50551# a_28596_50648# vdd pmos_6p0 w=1.22u l=1u
X13289 a_23756_50551# a_23668_50648# vss vss nmos_6p0 w=0.82u l=1u
X13290 vdd a_12108_14487# a_12020_14584# vdd pmos_6p0 w=1.22u l=1u
X13291 a_6740_31128# cap_shunt_n a_6532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X13292 a_28484_11828# cap_series_gyn a_28692_12312# vdd pmos_6p0 w=1.2u l=0.5u
X13293 a_22644_12312# cap_series_gyn a_22436_11828# vdd pmos_6p0 w=1.2u l=0.5u
X13294 a_10548_35832# cap_shunt_n a_10340_35348# vdd pmos_6p0 w=1.2u l=0.5u
X13295 vss cap_shunt_n a_35056_32696# vss nmos_6p0 w=0.82u l=0.6u
X13296 a_9668_49460# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13297 vdd tune_series_gy[4] a_14484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X13298 a_28692_40536# cap_shunt_p a_28484_40052# vdd pmos_6p0 w=1.2u l=0.5u
X13299 vdd tune_series_gy[4] a_14484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X13300 vss tune_series_gy[5] a_15720_11452# vss nmos_6p0 w=0.51u l=0.6u
X13301 vdd a_12108_11351# a_12020_11448# vdd pmos_6p0 w=1.22u l=1u
X13302 a_36652_50244# cap_shunt_gyp a_36384_50244# vss nmos_6p0 w=0.82u l=0.6u
X13303 vss cap_shunt_gyp a_35868_49944# vss nmos_6p0 w=0.82u l=0.6u
X13304 a_29700_39330# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13305 a_29492_34972# cap_shunt_p a_29700_34626# vdd pmos_6p0 w=1.2u l=0.5u
X13306 a_7672_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13307 a_5612_34871# a_5524_34968# vss vss nmos_6p0 w=0.82u l=1u
X13308 vss tune_shunt[7] a_7748_26786# vss nmos_6p0 w=0.51u l=0.6u
X13309 a_32612_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13310 vss tune_series_gy[4] a_18724_6040# vss nmos_6p0 w=0.51u l=0.6u
X13311 a_35692_18100# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13312 a_12788_18584# cap_shunt_p a_14504_18584# vss nmos_6p0 w=0.82u l=0.6u
X13313 a_25572_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13314 vss tune_shunt[7] a_17828_34264# vss nmos_6p0 w=0.51u l=0.6u
X13315 vdd a_1692_33303# a_1604_33400# vdd pmos_6p0 w=1.22u l=1u
X13316 vdd tune_series_gy[3] a_14484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X13317 vdd tune_series_gy[4] a_29532_16156# vdd pmos_6p0 w=1.2u l=0.5u
X13318 a_22848_18584# cap_shunt_p a_20740_18584# vss nmos_6p0 w=0.82u l=0.6u
X13319 vss cap_shunt_gyp a_35868_46808# vss nmos_6p0 w=0.82u l=0.6u
X13320 a_18612_12674# cap_series_gyn a_18404_13020# vdd pmos_6p0 w=1.2u l=0.5u
X13321 vss cap_series_gyp a_27888_20152# vss nmos_6p0 w=0.82u l=0.6u
X13322 a_29492_31836# cap_shunt_p a_29700_31490# vdd pmos_6p0 w=1.2u l=0.5u
X13323 a_7672_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13324 vdd a_19724_23895# a_19636_23992# vdd pmos_6p0 w=1.22u l=1u
X13325 a_5612_31735# a_5524_31832# vss vss nmos_6p0 w=0.82u l=1u
X13326 a_6740_13880# cap_shunt_p a_7672_13880# vss nmos_6p0 w=0.82u l=0.6u
X13327 vdd a_15692_55688# a_15604_55732# vdd pmos_6p0 w=1.22u l=1u
X13328 a_35040_43734# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13329 a_12788_15448# cap_shunt_p a_14504_15448# vss nmos_6p0 w=0.82u l=0.6u
X13330 a_6060_55255# a_5972_55352# vss vss nmos_6p0 w=0.82u l=1u
X13331 a_13588_49084# cap_shunt_n a_13796_48738# vdd pmos_6p0 w=1.2u l=0.5u
X13332 a_7748_34626# cap_shunt_n a_9464_34564# vss nmos_6p0 w=0.82u l=0.6u
X13333 vss tune_shunt[7] a_17828_31128# vss nmos_6p0 w=0.51u l=0.6u
X13334 a_22848_15448# cap_series_gyn a_20740_15448# vss nmos_6p0 w=0.82u l=0.6u
X13335 a_34720_37700# cap_shunt_p a_32612_37762# vss nmos_6p0 w=0.82u l=0.6u
X13336 vdd a_19724_20759# a_19636_20856# vdd pmos_6p0 w=1.22u l=1u
X13337 a_21748_11106# cap_series_gyn a_21540_11452# vdd pmos_6p0 w=1.2u l=0.5u
X13338 a_10660_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13339 a_28572_12919# a_28484_13016# vss vss nmos_6p0 w=0.82u l=1u
X13340 vdd a_12668_55688# a_12580_55732# vdd pmos_6p0 w=1.22u l=1u
X13341 a_5936_46808# cap_shunt_p a_3828_46808# vss nmos_6p0 w=0.82u l=0.6u
X13342 a_7792_4772# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13343 vdd tune_series_gy[3] a_18180_3612# vdd pmos_6p0 w=1.2u l=0.5u
X13344 a_3036_55255# a_2948_55352# vss vss nmos_6p0 w=0.82u l=1u
X13345 a_7748_31490# cap_shunt_n a_9464_31428# vss nmos_6p0 w=0.82u l=0.6u
X13346 vdd a_30364_20759# a_30276_20856# vdd pmos_6p0 w=1.22u l=1u
X13347 vdd tune_shunt[6] a_7540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X13348 a_20620_30167# a_20532_30264# vss vss nmos_6p0 w=0.82u l=1u
X13349 a_19732_10744# cap_series_gyn a_19524_10260# vdd pmos_6p0 w=1.2u l=0.5u
X13350 a_13796_47170# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13351 vdd a_6060_30167# a_5972_30264# vdd pmos_6p0 w=1.22u l=1u
X13352 vdd tune_shunt[3] a_32404_38108# vdd pmos_6p0 w=1.2u l=0.5u
X13353 a_8680_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13354 a_6292_50306# cap_shunt_p a_6084_50652# vdd pmos_6p0 w=1.2u l=0.5u
X13355 a_21540_42812# cap_shunt_n a_21748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X13356 a_23072_28292# cap_shunt_n a_21748_28354# vss nmos_6p0 w=0.82u l=0.6u
X13357 vss tune_shunt[7] a_28692_27992# vss nmos_6p0 w=0.51u l=0.6u
X13358 a_24660_4834# cap_series_gyp a_24452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X13359 a_3248_7908# cap_shunt_n a_1924_7970# vss nmos_6p0 w=0.82u l=0.6u
X13360 a_6532_46324# cap_shunt_p a_6740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X13361 a_11480_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13362 vdd a_28236_52552# a_28148_52596# vdd pmos_6p0 w=1.22u l=1u
X13363 a_7560_9476# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13364 a_13796_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13365 a_20620_27031# a_20532_27128# vss vss nmos_6p0 w=0.82u l=1u
X13366 a_25780_18584# cap_series_gyn a_25572_18100# vdd pmos_6p0 w=1.2u l=0.5u
X13367 a_34516_23650# cap_series_gygyp a_34308_23996# vdd pmos_6p0 w=1.2u l=0.5u
X13368 a_3640_7608# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13369 a_26712_7608# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13370 vdd tune_shunt[7] a_17620_16532# vdd pmos_6p0 w=1.2u l=0.5u
X13371 a_20532_32212# cap_shunt_n a_20740_32696# vdd pmos_6p0 w=1.2u l=0.5u
X13372 a_23072_25156# cap_shunt_n a_21748_25218# vss nmos_6p0 w=0.82u l=0.6u
X13373 vss tune_shunt[7] a_28692_24856# vss nmos_6p0 w=0.51u l=0.6u
X13374 a_16476_22760# a_16388_22804# vss vss nmos_6p0 w=0.82u l=1u
X13375 a_13796_28354# cap_shunt_n a_13588_28700# vdd pmos_6p0 w=1.2u l=0.5u
X13376 a_11480_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13377 a_21748_20514# cap_shunt_p a_21540_20860# vdd pmos_6p0 w=1.2u l=0.5u
X13378 a_6740_24856# cap_shunt_p a_6532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X13379 a_5388_3944# a_5300_3988# vss vss nmos_6p0 w=0.82u l=1u
X13380 vdd a_19500_50551# a_19412_50648# vdd pmos_6p0 w=1.22u l=1u
X13381 vss tune_shunt[6] a_16708_42466# vss nmos_6p0 w=0.51u l=0.6u
X13382 vss cap_series_gyp a_30016_13880# vss nmos_6p0 w=0.82u l=0.6u
X13383 vdd tune_shunt[4] a_33524_35348# vdd pmos_6p0 w=1.2u l=0.5u
X13384 a_10548_29560# cap_shunt_n a_10340_29076# vdd pmos_6p0 w=1.2u l=0.5u
X13385 vss tune_shunt[7] a_7748_29922# vss nmos_6p0 w=0.51u l=0.6u
X13386 a_35880_24372# cap_series_gygyp a_35692_24372# vdd pmos_6p0 w=1.2u l=0.5u
X13387 a_33920_45302# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13388 a_25592_39268# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13389 a_2932_10744# cap_shunt_n a_2724_10260# vdd pmos_6p0 w=1.2u l=0.5u
X13390 a_6740_21720# cap_shunt_p a_6532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X13391 a_30588_43144# a_30500_43188# vss vss nmos_6p0 w=0.82u l=1u
X13392 a_6420_13020# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13393 a_5612_28599# a_5524_28696# vss vss nmos_6p0 w=0.82u l=1u
X13394 a_18612_11106# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13395 a_3828_20152# cap_shunt_p a_3620_19668# vdd pmos_6p0 w=1.2u l=0.5u
X13396 vss cap_series_gygyp a_35840_22020# vss nmos_6p0 w=0.82u l=0.6u
X13397 vss cap_series_gyn a_30136_9476# vss nmos_6p0 w=0.82u l=0.6u
X13398 vss cap_series_gyp a_30016_10744# vss nmos_6p0 w=0.82u l=0.6u
X13399 a_20328_11044# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13400 vdd tune_shunt[7] a_6532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X13401 vdd a_26892_49416# a_26804_49460# vdd pmos_6p0 w=1.22u l=1u
X13402 a_10248_47108# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13403 a_35880_21236# cap_series_gygyp a_35692_21236# vdd pmos_6p0 w=1.2u l=0.5u
X13404 a_3828_42104# cap_shunt_p a_3620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X13405 a_18724_6040# cap_series_gyn a_18516_5556# vdd pmos_6p0 w=1.2u l=0.5u
X13406 a_30500_45944# cap_shunt_gyn a_30688_45944# vdd pmos_6p0 w=1.215u l=0.5u
X13407 a_29492_25564# cap_shunt_p a_29700_25218# vdd pmos_6p0 w=1.2u l=0.5u
X13408 a_24660_18946# cap_series_gyn a_25592_18884# vss nmos_6p0 w=0.82u l=0.6u
X13409 a_36076_38007# a_35988_38104# vss vss nmos_6p0 w=0.82u l=1u
X13410 a_5612_25463# a_5524_25560# vss vss nmos_6p0 w=0.82u l=1u
X13411 a_21540_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13412 a_33948_49416# a_33860_49460# vss vss nmos_6p0 w=0.82u l=1u
X13413 vdd a_26892_46280# a_26804_46324# vdd pmos_6p0 w=1.22u l=1u
X13414 a_13796_29922# cap_shunt_n a_13588_30268# vdd pmos_6p0 w=1.2u l=0.5u
X13415 vss cap_series_gyp a_13104_4472# vss nmos_6p0 w=0.82u l=0.6u
X13416 a_6292_17016# cap_shunt_p a_6084_16532# vdd pmos_6p0 w=1.2u l=0.5u
X13417 vdd a_23868_49416# a_23780_49460# vdd pmos_6p0 w=1.22u l=1u
X13418 a_36384_48676# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13419 a_15492_5180# cap_series_gyn a_15700_4834# vdd pmos_6p0 w=1.2u l=0.5u
X13420 a_7748_28354# cap_shunt_n a_9464_28292# vss nmos_6p0 w=0.82u l=0.6u
X13421 a_9876_13880# cap_shunt_p a_9668_13396# vdd pmos_6p0 w=1.2u l=0.5u
X13422 vss cap_shunt_p a_19152_43672# vss nmos_6p0 w=0.82u l=0.6u
X13423 a_14908_5079# a_14820_5176# vss vss nmos_6p0 w=0.82u l=1u
X13424 vss cap_shunt_p a_7952_9176# vss nmos_6p0 w=0.82u l=0.6u
X13425 vdd a_27228_42711# a_27140_42808# vdd pmos_6p0 w=1.22u l=1u
X13426 a_2708_12674# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13427 vdd a_19724_14487# a_19636_14584# vdd pmos_6p0 w=1.22u l=1u
X13428 a_24660_15810# cap_series_gyn a_25592_15748# vss nmos_6p0 w=0.82u l=0.6u
X13429 a_17620_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13430 a_36160_43189# cap_shunt_gyn a_36160_43734# vdd pmos_6p0 w=1.215u l=0.5u
X13431 vdd tune_shunt[5] a_12580_49460# vdd pmos_6p0 w=1.2u l=0.5u
X13432 a_13796_37762# cap_shunt_n a_14728_37700# vss nmos_6p0 w=0.82u l=0.6u
X13433 vdd a_33948_10216# a_33860_10260# vdd pmos_6p0 w=1.22u l=1u
X13434 a_2708_12674# cap_shunt_n a_4424_12612# vss nmos_6p0 w=0.82u l=0.6u
X13435 a_7748_25218# cap_shunt_n a_9464_25156# vss nmos_6p0 w=0.82u l=0.6u
X13436 a_19936_4772# cap_series_gyp a_18612_4834# vss nmos_6p0 w=0.82u l=0.6u
X13437 vss cap_shunt_n a_19152_40536# vss nmos_6p0 w=0.82u l=0.6u
X13438 a_29624_12312# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13439 vdd tune_shunt[6] a_7540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X13440 a_17620_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13441 vdd tune_series_gy[4] a_14484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X13442 a_11536_18884# cap_shunt_p a_9428_18946# vss nmos_6p0 w=0.82u l=0.6u
X13443 a_21540_36540# cap_shunt_n a_21748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X13444 a_29492_34972# cap_shunt_p a_29700_34626# vdd pmos_6p0 w=1.2u l=0.5u
X13445 a_6516_20514# cap_shunt_p a_6308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X13446 vdd a_15804_47848# a_15716_47892# vdd pmos_6p0 w=1.22u l=1u
X13447 vdd tune_series_gy[5] a_18404_8316# vdd pmos_6p0 w=1.2u l=0.5u
X13448 a_7540_23996# cap_shunt_p a_7748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X13449 a_10988_8648# a_10900_8692# vss vss nmos_6p0 w=0.82u l=1u
X13450 vdd tune_shunt[7] a_7540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X13451 a_29916_52119# a_29828_52216# vss vss nmos_6p0 w=0.82u l=1u
X13452 vss tune_shunt[5] a_20740_45240# vss nmos_6p0 w=0.51u l=0.6u
X13453 a_8680_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13454 vss tune_shunt[7] a_9876_13880# vss nmos_6p0 w=0.51u l=0.6u
X13455 vss cap_shunt_p a_18816_48676# vss nmos_6p0 w=0.82u l=0.6u
X13456 a_11668_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13457 a_17828_42104# cap_shunt_n a_17620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X13458 vdd tune_series_gy[4] a_29532_16156# vdd pmos_6p0 w=1.2u l=0.5u
X13459 a_21540_33404# cap_shunt_n a_21748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X13460 a_14260_3612# cap_series_gyn a_14468_3266# vdd pmos_6p0 w=1.2u l=0.5u
X13461 a_16016_9176# cap_series_gyn a_14692_9176# vss nmos_6p0 w=0.82u l=0.6u
X13462 vss tune_series_gy[4] a_28692_18584# vss nmos_6p0 w=0.51u l=0.6u
X13463 a_29492_31836# cap_shunt_p a_29700_31490# vdd pmos_6p0 w=1.2u l=0.5u
X13464 vdd tune_shunt[3] a_24452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X13465 a_20620_17623# a_20532_17720# vss vss nmos_6p0 w=0.82u l=1u
X13466 a_13900_55688# a_13812_55732# vss vss nmos_6p0 w=0.82u l=1u
X13467 a_9316_47170# cap_shunt_p a_11032_47108# vss nmos_6p0 w=0.82u l=0.6u
X13468 a_10092_44712# a_10004_44756# vss vss nmos_6p0 w=0.82u l=1u
X13469 vss tune_shunt[6] a_20740_42104# vss nmos_6p0 w=0.51u l=0.6u
X13470 vss tune_shunt[7] a_9876_10744# vss nmos_6p0 w=0.51u l=0.6u
X13471 a_13588_49084# cap_shunt_n a_13796_48738# vdd pmos_6p0 w=1.2u l=0.5u
X13472 vss tune_shunt[7] a_16708_36194# vss nmos_6p0 w=0.51u l=0.6u
X13473 vdd tune_shunt[7] a_33524_29076# vdd pmos_6p0 w=1.2u l=0.5u
X13474 a_7580_6748# cap_series_gyp a_7768_6748# vdd pmos_6p0 w=1.2u l=0.5u
X13475 a_2500_45948# cap_shunt_p a_2708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X13476 vss tune_series_gy[4] a_28692_15448# vss nmos_6p0 w=0.51u l=0.6u
X13477 a_35840_17316# cap_series_gygyn a_34516_17378# vss nmos_6p0 w=0.82u l=0.6u
X13478 a_21748_11106# cap_series_gyn a_21540_11452# vdd pmos_6p0 w=1.2u l=0.5u
X13479 vdd a_2140_54120# a_2052_54164# vdd pmos_6p0 w=1.22u l=1u
X13480 vdd tune_shunt[5] a_24452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X13481 a_36524_36439# a_36436_36536# vss vss nmos_6p0 w=0.82u l=1u
X13482 a_25592_7908# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X13483 vdd a_6508_41143# a_6420_41240# vdd pmos_6p0 w=1.22u l=1u
X13484 a_15700_7970# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13485 a_10092_41576# a_10004_41620# vss vss nmos_6p0 w=0.82u l=1u
X13486 a_17828_38968# cap_shunt_n a_19544_38968# vss nmos_6p0 w=0.82u l=0.6u
X13487 a_10548_26424# cap_shunt_n a_10340_25940# vdd pmos_6p0 w=1.2u l=0.5u
X13488 a_27888_38968# cap_shunt_p a_25780_38968# vss nmos_6p0 w=0.82u l=0.6u
X13489 vss tune_shunt[7] a_16708_33058# vss nmos_6p0 w=0.51u l=0.6u
X13490 a_32604_40008# a_32516_40052# vss vss nmos_6p0 w=0.82u l=1u
X13491 vss cap_shunt_n a_14784_37400# vss nmos_6p0 w=0.82u l=0.6u
X13492 vdd a_2140_50984# a_2052_51028# vdd pmos_6p0 w=1.22u l=1u
X13493 a_29700_37762# cap_shunt_n a_29492_38108# vdd pmos_6p0 w=1.2u l=0.5u
X13494 a_14692_4472# cap_series_gyp a_15624_4472# vss nmos_6p0 w=0.82u l=0.6u
X13495 vss cap_series_gyp a_16136_11044# vss nmos_6p0 w=0.82u l=0.6u
X13496 a_12580_19668# cap_shunt_p a_12788_20152# vdd pmos_6p0 w=1.2u l=0.5u
X13497 a_6292_50306# cap_shunt_p a_6084_50652# vdd pmos_6p0 w=1.2u l=0.5u
X13498 a_35264_47108# tune_shunt_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13499 vdd a_27228_39575# a_27140_39672# vdd pmos_6p0 w=1.22u l=1u
X13500 a_15700_4834# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X13501 a_10548_23288# cap_shunt_n a_10340_22804# vdd pmos_6p0 w=1.2u l=0.5u
X13502 a_6532_46324# cap_shunt_p a_6740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X13503 vss cap_shunt_n a_15120_32996# vss nmos_6p0 w=0.82u l=0.6u
X13504 a_3828_32696# cap_shunt_p a_3620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X13505 a_5844_9538# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X13506 a_31708_11784# a_31620_11828# vss vss nmos_6p0 w=0.82u l=1u
X13507 a_6740_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13508 a_34516_23650# cap_series_gygyp a_34308_23996# vdd pmos_6p0 w=1.2u l=0.5u
X13509 vdd a_27228_36439# a_27140_36536# vdd pmos_6p0 w=1.22u l=1u
X13510 vss tune_shunt[6] a_10660_40898# vss nmos_6p0 w=0.51u l=0.6u
X13511 a_32156_35304# a_32068_35348# vss vss nmos_6p0 w=0.82u l=1u
X13512 vdd tune_shunt[0] a_29492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X13513 a_21540_14588# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13514 a_6060_39575# a_5972_39672# vss vss nmos_6p0 w=0.82u l=1u
X13515 vdd a_35292_52552# a_35204_52596# vdd pmos_6p0 w=1.22u l=1u
X13516 a_31648_6340# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X13517 vss cap_shunt_n a_19152_34264# vss nmos_6p0 w=0.82u l=0.6u
X13518 a_14484_7124# cap_series_gyp a_14692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X13519 a_29720_16156# cap_series_gyn a_29744_15748# vss nmos_6p0 w=0.82u l=0.6u
X13520 a_22456_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13521 vss cap_series_gyp a_11984_4772# vss nmos_6p0 w=0.82u l=0.6u
X13522 vdd tune_shunt[5] a_3172_49460# vdd pmos_6p0 w=1.2u l=0.5u
X13523 a_17620_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13524 vss tune_series_gygy[4] a_34516_12674# vss nmos_6p0 w=0.51u l=0.6u
X13525 a_14684_50984# a_14596_51028# vss vss nmos_6p0 w=0.82u l=1u
X13526 vss tune_shunt[7] a_9428_20514# vss nmos_6p0 w=0.51u l=0.6u
X13527 vdd tune_shunt[4] a_21540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X13528 a_21748_20514# cap_shunt_p a_22680_20452# vss nmos_6p0 w=0.82u l=0.6u
X13529 a_19732_9176# cap_series_gyp a_19524_8692# vdd pmos_6p0 w=1.2u l=0.5u
X13530 a_2724_11828# cap_shunt_n a_2932_12312# vdd pmos_6p0 w=1.2u l=0.5u
X13531 vss cap_shunt_n a_19152_31128# vss nmos_6p0 w=0.82u l=0.6u
X13532 a_18032_29860# cap_shunt_n a_16708_29922# vss nmos_6p0 w=0.82u l=0.6u
X13533 vdd a_34396_24328# a_34308_24372# vdd pmos_6p0 w=1.22u l=1u
X13534 vss tune_series_gy[3] a_21524_3266# vss nmos_6p0 w=0.51u l=0.6u
X13535 a_28692_13880# cap_series_gyp a_28484_13396# vdd pmos_6p0 w=1.2u l=0.5u
X13536 vdd a_32268_52552# a_32180_52596# vdd pmos_6p0 w=1.22u l=1u
X13537 vdd tune_shunt[7] a_7540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X13538 a_22644_12312# cap_series_gyn a_24360_12312# vss nmos_6p0 w=0.82u l=0.6u
X13539 a_29492_38108# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13540 a_17620_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13541 a_29916_45847# a_29828_45944# vss vss nmos_6p0 w=0.82u l=1u
X13542 a_21540_27132# cap_shunt_n a_21748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X13543 a_16708_23650# cap_shunt_n a_16500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X13544 a_23576_13880# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13545 vdd a_31708_53687# a_31620_53784# vdd pmos_6p0 w=1.22u l=1u
X13546 a_29492_25564# cap_shunt_p a_29700_25218# vdd pmos_6p0 w=1.2u l=0.5u
X13547 a_11996_17623# a_11908_17720# vss vss nmos_6p0 w=0.82u l=1u
X13548 a_18032_26724# cap_shunt_n a_16708_26786# vss nmos_6p0 w=0.82u l=0.6u
X13549 a_1924_6040# cap_shunt_p a_1716_5556# vdd pmos_6p0 w=1.2u l=0.5u
X13550 a_24452_17724# cap_series_gyp a_24660_17378# vdd pmos_6p0 w=1.2u l=0.5u
X13551 a_3380_18584# cap_shunt_p a_5096_18584# vss nmos_6p0 w=0.82u l=0.6u
X13552 vdd a_34396_21192# a_34308_21236# vdd pmos_6p0 w=1.22u l=1u
X13553 a_13796_29922# cap_shunt_n a_13588_30268# vdd pmos_6p0 w=1.2u l=0.5u
X13554 a_6292_17016# cap_shunt_p a_6084_16532# vdd pmos_6p0 w=1.2u l=0.5u
X13555 a_25572_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13556 a_32632_14588# cap_series_gyp a_33440_14180# vss nmos_6p0 w=0.82u l=0.6u
X13557 a_29916_42711# a_29828_42808# vss vss nmos_6p0 w=0.82u l=1u
X13558 vss cap_shunt_n a_18816_39268# vss nmos_6p0 w=0.82u l=0.6u
X13559 a_17828_32696# cap_shunt_n a_17620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X13560 a_34348_9884# cap_series_gygyn a_34536_9884# vdd pmos_6p0 w=1.2u l=0.5u
X13561 vdd a_29692_41576# a_29604_41620# vdd pmos_6p0 w=1.22u l=1u
X13562 a_2500_39676# cap_shunt_n a_2708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X13563 a_23576_10744# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X13564 vdd a_31708_50551# a_31620_50648# vdd pmos_6p0 w=1.22u l=1u
X13565 a_13460_32696# cap_shunt_n a_15176_32696# vss nmos_6p0 w=0.82u l=0.6u
X13566 a_16924_21192# a_16836_21236# vss vss nmos_6p0 w=0.82u l=1u
X13567 vdd a_27228_5079# a_27140_5176# vdd pmos_6p0 w=1.22u l=1u
X13568 a_7748_45602# cap_shunt_p a_7540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X13569 a_35880_24372# cap_series_gygyp a_35904_24856# vss nmos_6p0 w=0.82u l=0.6u
X13570 a_25572_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13571 a_31436_22428# cap_series_gygyn a_31624_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13572 a_32632_11452# cap_series_gyp a_33440_11044# vss nmos_6p0 w=0.82u l=0.6u
X13573 a_34348_6748# cap_series_gygyp a_34536_6748# vdd pmos_6p0 w=1.2u l=0.5u
X13574 vdd a_12332_50551# a_12244_50648# vdd pmos_6p0 w=1.22u l=1u
X13575 a_24660_15810# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13576 a_7224_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13577 a_20532_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13578 a_32604_33736# a_32516_33780# vss vss nmos_6p0 w=0.82u l=1u
X13579 a_17828_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13580 a_34144_43972# cap_shunt_gyp a_34144_44376# vdd pmos_6p0 w=1.215u l=0.5u
X13581 vdd a_21740_55688# a_21652_55732# vdd pmos_6p0 w=1.22u l=1u
X13582 vdd a_4828_52552# a_4740_52596# vdd pmos_6p0 w=1.22u l=1u
X13583 a_13588_42812# cap_shunt_n a_13796_42466# vdd pmos_6p0 w=1.2u l=0.5u
X13584 a_6516_20514# cap_shunt_p a_6308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X13585 vdd a_34844_7080# a_34756_7124# vdd pmos_6p0 w=1.22u l=1u
X13586 a_7224_15748# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13587 a_32604_30600# a_32516_30644# vss vss nmos_6p0 w=0.82u l=1u
X13588 a_11424_50244# cap_shunt_p a_9316_50306# vss nmos_6p0 w=0.82u l=0.6u
X13589 a_7540_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13590 a_32156_29032# a_32068_29076# vss vss nmos_6p0 w=0.82u l=1u
X13591 a_6852_53442# cap_shunt_n a_6644_53788# vdd pmos_6p0 w=1.2u l=0.5u
X13592 a_6740_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13593 a_9540_9538# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13594 a_29132_52552# a_29044_52596# vss vss nmos_6p0 w=0.82u l=1u
X13595 a_33612_5079# a_33524_5176# vss vss nmos_6p0 w=0.82u l=1u
X13596 a_5636_10260# cap_shunt_p a_5844_10744# vdd pmos_6p0 w=1.2u l=0.5u
X13597 a_5636_10260# cap_shunt_p a_5844_10744# vdd pmos_6p0 w=1.2u l=0.5u
X13598 vss cap_shunt_n a_15120_23588# vss nmos_6p0 w=0.82u l=0.6u
X13599 vdd tune_shunt[7] a_20532_18100# vdd pmos_6p0 w=1.2u l=0.5u
X13600 vdd a_22412_55255# a_22324_55352# vdd pmos_6p0 w=1.22u l=1u
X13601 a_6740_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13602 a_35904_9176# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X13603 a_7540_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13604 vdd a_27228_27031# a_27140_27128# vdd pmos_6p0 w=1.22u l=1u
X13605 a_32156_25896# a_32068_25940# vss vss nmos_6p0 w=0.82u l=1u
X13606 a_35692_8692# tune_series_gygy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13607 a_30616_19668# cap_series_gygyn a_31424_20152# vss nmos_6p0 w=0.82u l=0.6u
X13608 a_30028_54120# a_29940_54164# vss vss nmos_6p0 w=0.82u l=1u
X13609 a_2500_45948# cap_shunt_p a_2708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X13610 vss tune_series_gygy[4] a_35880_36916# vss nmos_6p0 w=0.51u l=0.6u
X13611 vdd a_12556_14487# a_12468_14584# vdd pmos_6p0 w=1.22u l=1u
X13612 a_9668_21236# cap_shunt_p a_9876_21720# vdd pmos_6p0 w=1.2u l=0.5u
X13613 vss tune_shunt[6] a_14580_45240# vss nmos_6p0 w=0.51u l=0.6u
X13614 vdd tune_series_gy[3] a_28484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X13615 vss tune_shunt[5] a_3828_20152# vss nmos_6p0 w=0.51u l=0.6u
X13616 vss tune_shunt[4] a_25780_42104# vss nmos_6p0 w=0.51u l=0.6u
X13617 vdd tune_shunt[6] a_21540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X13618 vdd tune_series_gy[5] a_18404_8316# vdd pmos_6p0 w=1.2u l=0.5u
X13619 vss cap_shunt_p a_14112_12312# vss nmos_6p0 w=0.82u l=0.6u
X13620 a_21748_14242# cap_series_gyn a_22680_14180# vss nmos_6p0 w=0.82u l=0.6u
X13621 vdd a_22412_52119# a_22324_52216# vdd pmos_6p0 w=1.22u l=1u
X13622 vdd a_1692_41576# a_1604_41620# vdd pmos_6p0 w=1.22u l=1u
X13623 a_32612_34626# cap_shunt_n a_34328_34564# vss nmos_6p0 w=0.82u l=0.6u
X13624 vss tune_shunt[5] a_29700_31490# vss nmos_6p0 w=0.51u l=0.6u
X13625 a_35692_5556# tune_series_gygy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13626 vdd a_12556_11351# a_12468_11448# vdd pmos_6p0 w=1.22u l=1u
X13627 a_33948_52119# a_33860_52216# vss vss nmos_6p0 w=0.82u l=1u
X13628 a_29700_37762# cap_shunt_n a_29492_38108# vdd pmos_6p0 w=1.2u l=0.5u
X13629 a_2708_23650# cap_shunt_p a_2500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X13630 a_12580_19668# cap_shunt_p a_12788_20152# vdd pmos_6p0 w=1.2u l=0.5u
X13631 a_6292_50306# cap_shunt_p a_6084_50652# vdd pmos_6p0 w=1.2u l=0.5u
X13632 vss tune_shunt[6] a_14580_42104# vss nmos_6p0 w=0.51u l=0.6u
X13633 a_25444_3266# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X13634 vdd tune_shunt[3] a_2500_9884# vdd pmos_6p0 w=1.2u l=0.5u
X13635 a_21748_11106# cap_series_gyn a_22680_11044# vss nmos_6p0 w=0.82u l=0.6u
X13636 a_11648_14180# cap_shunt_p a_9540_14242# vss nmos_6p0 w=0.82u l=0.6u
X13637 a_6628_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13638 a_36384_49080# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X13639 vss cap_shunt_n a_12768_29860# vss nmos_6p0 w=0.82u l=0.6u
X13640 a_30408_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X13641 a_29196_3612# cap_series_gyn a_29384_3612# vdd pmos_6p0 w=1.2u l=0.5u
X13642 a_8996_52220# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13643 a_35600_50006# tune_shunt_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13644 a_32612_31490# cap_shunt_n a_34328_31428# vss nmos_6p0 w=0.82u l=0.6u
X13645 a_35880_25940# cap_series_gygyp a_35692_25940# vdd pmos_6p0 w=1.2u l=0.5u
X13646 a_31436_19292# cap_series_gygyn a_31624_19292# vdd pmos_6p0 w=1.2u l=0.5u
X13647 vdd a_8300_55688# a_8212_55732# vdd pmos_6p0 w=1.22u l=1u
X13648 vdd tune_shunt_gy[3] a_34980_44376# vdd pmos_6p0 w=1.215u l=0.5u
X13649 a_16708_14242# cap_shunt_p a_16500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X13650 a_31436_8316# cap_series_gygyn a_31624_8316# vdd pmos_6p0 w=1.2u l=0.5u
X13651 a_11648_11044# cap_shunt_p a_9540_11106# vss nmos_6p0 w=0.82u l=0.6u
X13652 vss tune_series_gygy[5] a_30616_19668# vss nmos_6p0 w=0.51u l=0.6u
X13653 vdd a_31708_44279# a_31620_44376# vdd pmos_6p0 w=1.22u l=1u
X13654 a_35756_42104# cap_shunt_gyn a_35488_42166# vss nmos_6p0 w=0.82u l=0.6u
X13655 a_18032_17316# cap_shunt_p a_16708_17378# vss nmos_6p0 w=0.82u l=0.6u
X13656 vss cap_shunt_n a_12768_26724# vss nmos_6p0 w=0.82u l=0.6u
X13657 vss cap_shunt_p a_4816_43972# vss nmos_6p0 w=0.82u l=0.6u
X13658 a_35880_22804# cap_series_gygyp a_35692_22804# vdd pmos_6p0 w=1.2u l=0.5u
X13659 a_35880_18100# cap_series_gygyn a_35904_18584# vss nmos_6p0 w=0.82u l=0.6u
X13660 a_7748_39330# cap_shunt_n a_7540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X13661 a_28692_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13662 a_3640_6340# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13663 a_8412_11351# a_8324_11448# vss vss nmos_6p0 w=0.82u l=1u
X13664 a_25572_16532# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13665 vss cap_shunt_n a_22064_45240# vss nmos_6p0 w=0.82u l=0.6u
X13666 a_36748_35304# a_36660_35348# vss vss nmos_6p0 w=0.82u l=1u
X13667 a_8860_18056# a_8772_18100# vss vss nmos_6p0 w=0.82u l=1u
X13668 a_13460_23288# cap_shunt_n a_15176_23288# vss nmos_6p0 w=0.82u l=0.6u
X13669 a_16500_45948# cap_shunt_p a_16708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X13670 a_34516_23650# cap_series_gygyp a_35448_23588# vss nmos_6p0 w=0.82u l=0.6u
X13671 a_22680_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13672 a_31820_49416# a_31732_49460# vss vss nmos_6p0 w=0.82u l=1u
X13673 a_3484_55255# a_3396_55352# vss vss nmos_6p0 w=0.82u l=1u
X13674 vss cap_shunt_p a_4816_40836# vss nmos_6p0 w=0.82u l=0.6u
X13675 a_20740_40536# cap_shunt_p a_20532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X13676 vss tune_series_gygy[4] a_35880_13396# vss nmos_6p0 w=0.51u l=0.6u
X13677 a_35880_14964# cap_series_gygyn a_35904_15448# vss nmos_6p0 w=0.82u l=0.6u
X13678 a_13588_36540# cap_shunt_n a_13796_36194# vdd pmos_6p0 w=1.2u l=0.5u
X13679 vss tune_shunt[7] a_2708_31490# vss nmos_6p0 w=0.51u l=0.6u
X13680 a_3640_3204# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13681 vss cap_shunt_p a_22064_42104# vss nmos_6p0 w=0.82u l=0.6u
X13682 vss tune_shunt[6] a_10660_37762# vss nmos_6p0 w=0.51u l=0.6u
X13683 a_28692_13880# cap_series_gyp a_28484_13396# vdd pmos_6p0 w=1.2u l=0.5u
X13684 a_9108_50652# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13685 vdd tune_shunt[6] a_14372_43188# vdd pmos_6p0 w=1.2u l=0.5u
X13686 a_20532_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13687 a_7748_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13688 a_31820_46280# a_31732_46324# vss vss nmos_6p0 w=0.82u l=1u
X13689 vss tune_shunt[7] a_32612_29922# vss nmos_6p0 w=0.51u l=0.6u
X13690 vdd tune_series_gy[4] a_21428_5556# vdd pmos_6p0 w=1.2u l=0.5u
X13691 vdd a_28684_52552# a_28596_52596# vdd pmos_6p0 w=1.22u l=1u
X13692 vdd a_37420_34871# a_37332_34968# vdd pmos_6p0 w=1.22u l=1u
X13693 a_13588_33404# cap_shunt_n a_13796_33058# vdd pmos_6p0 w=1.2u l=0.5u
X13694 a_16708_23650# cap_shunt_n a_16500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X13695 vss tune_series_gygy[4] a_35880_10260# vss nmos_6p0 w=0.51u l=0.6u
X13696 vss tune_shunt[7] a_10660_34626# vss nmos_6p0 w=0.51u l=0.6u
X13697 a_24452_17724# cap_series_gyp a_24660_17378# vdd pmos_6p0 w=1.2u l=0.5u
X13698 vss cap_series_gyp a_31808_14180# vss nmos_6p0 w=0.82u l=0.6u
X13699 vdd a_22412_48983# a_22324_49080# vdd pmos_6p0 w=1.22u l=1u
X13700 a_20740_46808# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13701 a_11612_8692# cap_series_gyp a_11800_8692# vdd pmos_6p0 w=1.2u l=0.5u
X13702 vdd a_10540_46280# a_10452_46324# vdd pmos_6p0 w=1.22u l=1u
X13703 a_32432_22020# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X13704 a_2500_39676# cap_shunt_n a_2708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X13705 a_30028_47848# a_29940_47892# vss vss nmos_6p0 w=0.82u l=1u
X13706 a_21748_4834# cap_series_gyp a_21540_5180# vdd pmos_6p0 w=1.2u l=0.5u
X13707 vss cap_shunt_n a_23072_43972# vss nmos_6p0 w=0.82u l=0.6u
X13708 a_9876_49944# cap_shunt_p a_9668_49460# vdd pmos_6p0 w=1.2u l=0.5u
X13709 a_31436_22428# cap_series_gygyn a_31624_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13710 vss cap_series_gyp a_31808_11044# vss nmos_6p0 w=0.82u l=0.6u
X13711 a_19936_32696# cap_shunt_n a_17828_32696# vss nmos_6p0 w=0.82u l=0.6u
X13712 a_3172_51028# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13713 a_32612_28354# cap_shunt_p a_34328_28292# vss nmos_6p0 w=0.82u l=0.6u
X13714 vss cap_series_gyp a_27104_6040# vss nmos_6p0 w=0.82u l=0.6u
X13715 a_32156_16488# a_32068_16532# vss vss nmos_6p0 w=0.82u l=1u
X13716 vss cap_shunt_p a_23072_40836# vss nmos_6p0 w=0.82u l=0.6u
X13717 vss cap_shunt_n a_11872_27992# vss nmos_6p0 w=0.82u l=0.6u
X13718 a_5544_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13719 a_28692_32696# cap_shunt_p a_30408_32696# vss nmos_6p0 w=0.82u l=0.6u
X13720 a_33612_23895# a_33524_23992# vss vss nmos_6p0 w=0.82u l=1u
X13721 vss cap_series_gyn a_16800_10744# vss nmos_6p0 w=0.82u l=0.6u
X13722 vdd a_1692_32168# a_1604_32212# vdd pmos_6p0 w=1.22u l=1u
X13723 a_32612_25218# cap_shunt_p a_34328_25156# vss nmos_6p0 w=0.82u l=0.6u
X13724 a_24660_37762# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13725 a_29700_36194# cap_shunt_n a_29492_36540# vdd pmos_6p0 w=1.2u l=0.5u
X13726 a_2708_14242# cap_shunt_n a_2500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X13727 a_9876_17016# cap_shunt_p a_10808_17016# vss nmos_6p0 w=0.82u l=0.6u
X13728 vss cap_shunt_n a_11872_24856# vss nmos_6p0 w=0.82u l=0.6u
X13729 vss tune_series_gygy[5] a_31624_20860# vss nmos_6p0 w=0.51u l=0.6u
X13730 a_6852_53442# cap_shunt_n a_6644_53788# vdd pmos_6p0 w=1.2u l=0.5u
X13731 vdd a_32604_36872# a_32516_36916# vdd pmos_6p0 w=1.22u l=1u
X13732 a_28124_22327# a_28036_22424# vss vss nmos_6p0 w=0.82u l=1u
X13733 a_21748_44034# cap_shunt_n a_21540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X13734 a_16708_33058# cap_shunt_n a_17640_32996# vss nmos_6p0 w=0.82u l=0.6u
X13735 a_28692_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13736 a_35880_16532# cap_series_gygyn a_35692_16532# vdd pmos_6p0 w=1.2u l=0.5u
X13737 vdd a_27676_42711# a_27588_42808# vdd pmos_6p0 w=1.22u l=1u
X13738 a_24660_34626# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13739 a_29700_33058# cap_shunt_p a_29492_33404# vdd pmos_6p0 w=1.2u l=0.5u
X13740 a_36748_29032# a_36660_29076# vss vss nmos_6p0 w=0.82u l=1u
X13741 a_16708_45602# cap_shunt_p a_18424_45540# vss nmos_6p0 w=0.82u l=0.6u
X13742 a_1692_27464# a_1604_27508# vss vss nmos_6p0 w=0.82u l=1u
X13743 a_16500_39676# cap_shunt_n a_16708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X13744 a_13460_38968# cap_shunt_n a_14392_38968# vss nmos_6p0 w=0.82u l=0.6u
X13745 a_16708_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13746 a_21748_40898# cap_shunt_p a_21540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X13747 vss cap_shunt_n a_4816_34564# vss nmos_6p0 w=0.82u l=0.6u
X13748 a_2708_17378# cap_shunt_p a_2500_17724# vdd pmos_6p0 w=1.2u l=0.5u
X13749 a_28692_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13750 a_26444_54120# a_26356_54164# vss vss nmos_6p0 w=0.82u l=1u
X13751 vdd a_34396_41143# a_34308_41240# vdd pmos_6p0 w=1.22u l=1u
X13752 a_33164_16055# a_33076_16152# vss vss nmos_6p0 w=0.82u l=1u
X13753 a_21540_13020# cap_series_gyn a_21748_12674# vdd pmos_6p0 w=1.2u l=0.5u
X13754 vdd a_29132_55688# a_29044_55732# vdd pmos_6p0 w=1.22u l=1u
X13755 vdd a_16364_54120# a_16276_54164# vdd pmos_6p0 w=1.22u l=1u
X13756 a_16708_42466# cap_shunt_n a_18424_42404# vss nmos_6p0 w=0.82u l=0.6u
X13757 a_1692_24328# a_1604_24372# vss vss nmos_6p0 w=0.82u l=1u
X13758 a_26768_42404# cap_shunt_n a_24660_42466# vss nmos_6p0 w=0.82u l=0.6u
X13759 a_37632_38485# cap_shunt_gyp a_37652_38968# vss nmos_6p0 w=0.82u l=0.6u
X13760 vss tune_shunt[5] a_6292_18946# vss nmos_6p0 w=0.51u l=0.6u
X13761 vss tune_series_gy[5] a_18612_11106# vss nmos_6p0 w=0.51u l=0.6u
X13762 vss cap_shunt_gyn a_34412_48676# vss nmos_6p0 w=0.82u l=0.6u
X13763 vss cap_shunt_p a_4816_31428# vss nmos_6p0 w=0.82u l=0.6u
X13764 a_3828_27992# cap_shunt_n a_5544_27992# vss nmos_6p0 w=0.82u l=0.6u
X13765 vdd a_15804_55255# a_15716_55352# vdd pmos_6p0 w=1.22u l=1u
X13766 vdd a_37420_28599# a_37332_28696# vdd pmos_6p0 w=1.22u l=1u
X13767 a_13588_27132# cap_shunt_n a_13796_26786# vdd pmos_6p0 w=1.2u l=0.5u
X13768 a_6740_26424# cap_shunt_n a_6532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X13769 vss tune_shunt[5] a_2708_22082# vss nmos_6p0 w=0.51u l=0.6u
X13770 a_14484_8692# cap_series_gyn a_14692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X13771 a_16812_12919# a_16724_13016# vss vss nmos_6p0 w=0.82u l=1u
X13772 a_11668_46808# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13773 vss tune_shunt[7] a_10660_28354# vss nmos_6p0 w=0.51u l=0.6u
X13774 vdd a_26108_55688# a_26020_55732# vdd pmos_6p0 w=1.22u l=1u
X13775 a_8996_52220# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13776 vdd a_14460_9783# a_14372_9880# vdd pmos_6p0 w=1.22u l=1u
X13777 a_31436_19292# cap_series_gygyn a_31624_19292# vdd pmos_6p0 w=1.2u l=0.5u
X13778 a_6532_52596# cap_shunt_n a_6740_53080# vdd pmos_6p0 w=1.2u l=0.5u
X13779 a_27496_35832# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13780 vss cap_shunt_n a_7168_11044# vss nmos_6p0 w=0.82u l=0.6u
X13781 a_3828_24856# cap_shunt_p a_5544_24856# vss nmos_6p0 w=0.82u l=0.6u
X13782 vss tune_shunt[3] a_2932_9176# vss nmos_6p0 w=0.51u l=0.6u
X13783 a_16708_14242# cap_shunt_p a_16500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X13784 vss cap_shunt_p a_7616_18584# vss nmos_6p0 w=0.82u l=0.6u
X13785 vdd a_15804_52119# a_15716_52216# vdd pmos_6p0 w=1.22u l=1u
X13786 a_20732_50984# a_20644_51028# vss vss nmos_6p0 w=0.82u l=1u
X13787 a_6740_23288# cap_shunt_p a_6532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X13788 vss tune_series_gygy[5] a_31624_22428# vss nmos_6p0 w=0.51u l=0.6u
X13789 a_14484_5556# cap_series_gyn a_14692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X13790 a_32156_3944# a_32068_3988# vss vss nmos_6p0 w=0.82u l=1u
X13791 vss tune_shunt[7] a_10660_25218# vss nmos_6p0 w=0.51u l=0.6u
X13792 a_28692_6040# cap_shunt_n a_29624_6040# vss nmos_6p0 w=0.82u l=0.6u
X13793 a_11984_53080# cap_shunt_n a_9876_53080# vss nmos_6p0 w=0.82u l=0.6u
X13794 vss tune_shunt[6] a_2708_42466# vss nmos_6p0 w=0.51u l=0.6u
X13795 vdd a_14460_6647# a_14372_6744# vdd pmos_6p0 w=1.22u l=1u
X13796 a_1924_6402# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X13797 a_14896_13880# cap_shunt_p a_12788_13880# vss nmos_6p0 w=0.82u l=0.6u
X13798 a_36720_49461# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X13799 a_3620_40052# cap_shunt_n a_3828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X13800 vdd a_6956_41143# a_6868_41240# vdd pmos_6p0 w=1.22u l=1u
X13801 a_34308_22428# cap_series_gygyp a_34516_22082# vdd pmos_6p0 w=1.2u l=0.5u
X13802 vss cap_shunt_p a_23072_34564# vss nmos_6p0 w=0.82u l=0.6u
X13803 a_9876_49944# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13804 a_34516_23650# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13805 vdd tune_series_gy[4] a_29492_11452# vdd pmos_6p0 w=1.2u l=0.5u
X13806 a_6292_48738# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13807 a_36720_46325# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X13808 a_19936_23288# cap_shunt_n a_17828_23288# vss nmos_6p0 w=0.82u l=0.6u
X13809 vdd a_27676_39575# a_27588_39672# vdd pmos_6p0 w=1.22u l=1u
X13810 a_5724_52552# a_5636_52596# vss vss nmos_6p0 w=0.82u l=1u
X13811 vss cap_shunt_n a_23072_31428# vss nmos_6p0 w=0.82u l=0.6u
X13812 a_28692_23288# cap_shunt_p a_30408_23288# vss nmos_6p0 w=0.82u l=0.6u
X13813 vss cap_series_gyn a_25984_6340# vss nmos_6p0 w=0.82u l=0.6u
X13814 vss cap_shunt_p a_5152_20152# vss nmos_6p0 w=0.82u l=0.6u
X13815 vdd tune_series_gy[2] a_10452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X13816 vdd tune_shunt[7] a_9668_10260# vdd pmos_6p0 w=1.2u l=0.5u
X13817 a_34516_20514# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13818 a_1924_7608# tune_shunt[2] vss vss nmos_6p0 w=0.51u l=0.6u
X13819 a_24452_17724# cap_series_gyp a_24660_17378# vdd pmos_6p0 w=1.2u l=0.5u
X13820 a_29700_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13821 vss cap_shunt_n a_15904_22020# vss nmos_6p0 w=0.82u l=0.6u
X13822 vdd a_27676_36439# a_27588_36536# vdd pmos_6p0 w=1.22u l=1u
X13823 a_24660_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13824 a_29700_26786# cap_shunt_p a_29492_27132# vdd pmos_6p0 w=1.2u l=0.5u
X13825 a_24204_19624# a_24116_19668# vss vss nmos_6p0 w=0.82u l=1u
X13826 a_6084_18100# cap_shunt_p a_6292_18584# vdd pmos_6p0 w=1.2u l=0.5u
X13827 a_16708_36194# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13828 vdd a_32604_27464# a_32516_27508# vdd pmos_6p0 w=1.22u l=1u
X13829 a_16708_23650# cap_shunt_n a_17640_23588# vss nmos_6p0 w=0.82u l=0.6u
X13830 vss cap_shunt_n a_4816_28292# vss nmos_6p0 w=0.82u l=0.6u
X13831 a_24660_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13832 a_31436_22428# cap_series_gygyn a_31624_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13833 a_16632_4772# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13834 a_26444_47848# a_26356_47892# vss vss nmos_6p0 w=0.82u l=1u
X13835 vss cap_shunt_gyn a_33292_47108# vss nmos_6p0 w=0.82u l=0.6u
X13836 vdd a_33948_3944# a_33860_3988# vdd pmos_6p0 w=1.22u l=1u
X13837 vdd a_29132_49416# a_29044_49460# vdd pmos_6p0 w=1.22u l=1u
X13838 a_22848_43672# cap_shunt_n a_20740_43672# vss nmos_6p0 w=0.82u l=0.6u
X13839 a_16708_36194# cap_shunt_n a_18424_36132# vss nmos_6p0 w=0.82u l=0.6u
X13840 vdd tune_shunt[6] a_25572_33780# vdd pmos_6p0 w=1.2u l=0.5u
X13841 a_4032_12612# cap_shunt_n a_2708_12674# vss nmos_6p0 w=0.82u l=0.6u
X13842 a_1692_18056# a_1604_18100# vss vss nmos_6p0 w=0.82u l=1u
X13843 a_3172_51028# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13844 a_17620_40052# cap_shunt_n a_17828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X13845 a_26768_36132# cap_shunt_p a_24660_36194# vss nmos_6p0 w=0.82u l=0.6u
X13846 a_28572_5079# a_28484_5176# vss vss nmos_6p0 w=0.82u l=1u
X13847 vss tune_shunt[7] a_9428_20514# vss nmos_6p0 w=0.51u l=0.6u
X13848 a_16708_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13849 a_32740_45944# cap_shunt_gyn a_32928_45944# vdd pmos_6p0 w=1.215u l=0.5u
X13850 a_15176_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13851 vss cap_shunt_p a_4816_25156# vss nmos_6p0 w=0.82u l=0.6u
X13852 a_28692_17016# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X13853 a_1716_8316# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13854 vdd a_29132_46280# a_29044_46324# vdd pmos_6p0 w=1.22u l=1u
X13855 a_22848_40536# cap_shunt_p a_20740_40536# vss nmos_6p0 w=0.82u l=0.6u
X13856 vdd tune_shunt[7] a_25572_30644# vdd pmos_6p0 w=1.2u l=0.5u
X13857 a_1692_14920# a_1604_14964# vss vss nmos_6p0 w=0.82u l=1u
X13858 a_16500_34972# cap_shunt_n a_16708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X13859 a_27496_29560# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13860 a_29700_36194# cap_shunt_n a_29492_36540# vdd pmos_6p0 w=1.2u l=0.5u
X13861 a_6760_7124# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X13862 a_31932_41576# a_31844_41620# vss vss nmos_6p0 w=0.82u l=1u
X13863 vdd tune_shunt[6] a_21540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X13864 vdd a_37420_19191# a_37332_19288# vdd pmos_6p0 w=1.22u l=1u
X13865 a_34308_19292# cap_series_gygyn a_34516_18946# vdd pmos_6p0 w=1.2u l=0.5u
X13866 vss tune_shunt[6] a_2708_36194# vss nmos_6p0 w=0.51u l=0.6u
X13867 a_34516_22082# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13868 a_16500_31836# cap_shunt_n a_16708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X13869 a_27496_26424# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13870 a_7616_50244# cap_shunt_p a_6292_50306# vss nmos_6p0 w=0.82u l=0.6u
X13871 a_6532_43188# cap_shunt_p a_6740_43672# vdd pmos_6p0 w=1.2u l=0.5u
X13872 a_29700_33058# cap_shunt_p a_29492_33404# vdd pmos_6p0 w=1.2u l=0.5u
X13873 a_12580_14964# cap_shunt_p a_12788_15448# vdd pmos_6p0 w=1.2u l=0.5u
X13874 a_33052_53687# a_32964_53784# vss vss nmos_6p0 w=0.82u l=1u
X13875 vss cap_series_gyn a_26768_12612# vss nmos_6p0 w=0.82u l=0.6u
X13876 a_3828_15448# cap_shunt_p a_5544_15448# vss nmos_6p0 w=0.82u l=0.6u
X13877 a_23308_55255# a_23220_55352# vss vss nmos_6p0 w=0.82u l=1u
X13878 a_10640_47108# cap_shunt_p a_9316_47170# vss nmos_6p0 w=0.82u l=0.6u
X13879 vdd tune_shunt[7] a_21540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X13880 a_20720_11044# cap_series_gyn a_18612_11106# vss nmos_6p0 w=0.82u l=0.6u
X13881 a_35692_3988# tune_series_gygy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13882 a_34308_16156# cap_series_gygyn a_34516_15810# vdd pmos_6p0 w=1.2u l=0.5u
X13883 a_9668_51028# cap_shunt_n a_9876_51512# vdd pmos_6p0 w=1.2u l=0.5u
X13884 a_9668_51028# cap_shunt_n a_9876_51512# vdd pmos_6p0 w=1.2u l=0.5u
X13885 vdd a_30140_43144# a_30052_43188# vdd pmos_6p0 w=1.22u l=1u
X13886 vss tune_shunt[7] a_2708_33058# vss nmos_6p0 w=0.51u l=0.6u
X13887 vss cap_shunt_n a_23072_28292# vss nmos_6p0 w=0.82u l=0.6u
X13888 vdd a_12780_50551# a_12692_50648# vdd pmos_6p0 w=1.22u l=1u
X13889 a_28484_33780# cap_shunt_p a_28692_34264# vdd pmos_6p0 w=1.2u l=0.5u
X13890 a_2708_47170# cap_shunt_p a_2500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X13891 a_12580_11828# cap_shunt_p a_12788_12312# vdd pmos_6p0 w=1.2u l=0.5u
X13892 a_33052_50551# a_32964_50648# vss vss nmos_6p0 w=0.82u l=1u
X13893 a_21540_8316# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13894 vdd tune_shunt[6] a_17620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X13895 a_29492_11452# cap_series_gyp a_29700_11106# vdd pmos_6p0 w=1.2u l=0.5u
X13896 a_6852_53442# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X13897 a_13588_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13898 vss cap_shunt_n a_23072_25156# vss nmos_6p0 w=0.82u l=0.6u
X13899 vss tune_shunt[7] a_24660_23650# vss nmos_6p0 w=0.51u l=0.6u
X13900 a_11668_45240# cap_shunt_n a_13384_45240# vss nmos_6p0 w=0.82u l=0.6u
X13901 a_28484_30644# cap_shunt_n a_28692_31128# vdd pmos_6p0 w=1.2u l=0.5u
X13902 vdd a_11884_22327# a_11796_22424# vdd pmos_6p0 w=1.22u l=1u
X13903 a_6532_13396# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13904 a_10660_39330# cap_shunt_n a_11592_39268# vss nmos_6p0 w=0.82u l=0.6u
X13905 a_31436_6748# cap_series_gygyn a_31624_6748# vdd pmos_6p0 w=1.2u l=0.5u
X13906 a_3828_48376# cap_shunt_p a_3620_47892# vdd pmos_6p0 w=1.2u l=0.5u
X13907 vss cap_series_gygyp a_37080_26424# vss nmos_6p0 w=0.82u l=0.6u
X13908 a_15744_11044# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X13909 vdd tune_shunt[6] a_6532_47892# vdd pmos_6p0 w=1.2u l=0.5u
X13910 a_6084_52220# cap_shunt_p a_6292_51874# vdd pmos_6p0 w=1.2u l=0.5u
X13911 a_6196_47516# cap_shunt_p a_6404_47170# vdd pmos_6p0 w=1.2u l=0.5u
X13912 a_25780_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13913 a_31436_19292# cap_series_gygyn a_31624_19292# vdd pmos_6p0 w=1.2u l=0.5u
X13914 vdd a_16028_38440# a_15940_38484# vdd pmos_6p0 w=1.22u l=1u
X13915 a_28348_21192# a_28260_21236# vss vss nmos_6p0 w=0.82u l=1u
X13916 a_29580_52552# a_29492_52596# vss vss nmos_6p0 w=0.82u l=1u
X13917 vss tune_shunt[7] a_24660_20514# vss nmos_6p0 w=0.51u l=0.6u
X13918 a_19836_54120# a_19748_54164# vss vss nmos_6p0 w=0.82u l=1u
X13919 a_11668_42104# cap_shunt_n a_13384_42104# vss nmos_6p0 w=0.82u l=0.6u
X13920 a_7672_53080# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13921 vss tune_shunt[7] a_10548_34264# vss nmos_6p0 w=0.51u l=0.6u
X13922 a_14728_32996# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13923 a_3828_45240# cap_shunt_p a_3620_44756# vdd pmos_6p0 w=1.2u l=0.5u
X13924 a_37280_43734# cap_shunt_gyp a_37280_43189# vdd pmos_6p0 w=1.215u l=0.5u
X13925 vdd a_22860_55255# a_22772_55352# vdd pmos_6p0 w=1.22u l=1u
X13926 a_5612_53687# a_5524_53784# vss vss nmos_6p0 w=0.82u l=1u
X13927 vdd tune_shunt[6] a_6532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X13928 a_12600_43672# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13929 vdd a_27676_27031# a_27588_27128# vdd pmos_6p0 w=1.22u l=1u
X13930 a_17372_3511# a_17284_3608# vss vss nmos_6p0 w=0.82u l=1u
X13931 vdd tune_shunt[5] a_3172_18100# vdd pmos_6p0 w=1.2u l=0.5u
X13932 vdd a_16028_35304# a_15940_35348# vdd pmos_6p0 w=1.22u l=1u
X13933 a_30800_6040# cap_shunt_n a_28692_6040# vss nmos_6p0 w=0.82u l=0.6u
X13934 a_30476_54120# a_30388_54164# vss vss nmos_6p0 w=0.82u l=1u
X13935 a_36296_24856# cap_series_gygyp a_35880_24372# vss nmos_6p0 w=0.82u l=0.6u
X13936 vdd tune_series_gygy[5] a_34308_17724# vdd pmos_6p0 w=1.2u l=0.5u
X13937 vss tune_shunt[7] a_10548_31128# vss nmos_6p0 w=0.51u l=0.6u
X13938 a_24660_44034# cap_shunt_p a_25592_43972# vss nmos_6p0 w=0.82u l=0.6u
X13939 vss tune_shunt[6] a_7748_42466# vss nmos_6p0 w=0.51u l=0.6u
X13940 vdd tune_series_gy[2] a_7580_6748# vdd pmos_6p0 w=1.2u l=0.5u
X13941 vdd a_22860_52119# a_22772_52216# vdd pmos_6p0 w=1.22u l=1u
X13942 a_5612_50551# a_5524_50648# vss vss nmos_6p0 w=0.82u l=1u
X13943 a_19388_49416# a_19300_49460# vss vss nmos_6p0 w=0.82u l=1u
X13944 a_37652_48676# cap_shunt_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X13945 vdd tune_shunt[7] a_13252_32212# vdd pmos_6p0 w=1.2u l=0.5u
X13946 a_34308_22428# cap_series_gygyp a_34516_22082# vdd pmos_6p0 w=1.2u l=0.5u
X13947 a_12600_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X13948 a_24204_5512# a_24116_5556# vss vss nmos_6p0 w=0.82u l=1u
X13949 a_14372_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13950 a_22848_34264# cap_shunt_n a_20740_34264# vss nmos_6p0 w=0.82u l=0.6u
X13951 a_6404_22082# cap_shunt_p a_6196_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13952 vdd tune_shunt[7] a_9108_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13953 vss cap_series_gyp a_20720_4772# vss nmos_6p0 w=0.82u l=0.6u
X13954 a_2500_34972# cap_shunt_n a_2708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X13955 vdd tune_shunt[7] a_25572_24372# vdd pmos_6p0 w=1.2u l=0.5u
X13956 a_11668_43672# cap_shunt_n a_11460_43188# vdd pmos_6p0 w=1.2u l=0.5u
X13957 a_24660_40898# cap_shunt_n a_25592_40836# vss nmos_6p0 w=0.82u l=0.6u
X13958 a_22436_7124# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13959 a_6628_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13960 a_8064_37400# cap_shunt_n a_6740_37400# vss nmos_6p0 w=0.82u l=0.6u
X13961 a_31436_8316# tune_series_gygy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13962 a_4424_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X13963 a_10548_34264# cap_shunt_n a_11480_34264# vss nmos_6p0 w=0.82u l=0.6u
X13964 a_22848_31128# cap_shunt_n a_20740_31128# vss nmos_6p0 w=0.82u l=0.6u
X13965 a_13460_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13966 a_9332_11452# cap_shunt_p a_9540_11106# vdd pmos_6p0 w=1.2u l=0.5u
X13967 vdd tune_series_gygy[5] a_35692_19668# vdd pmos_6p0 w=1.2u l=0.5u
X13968 a_37632_44376# cap_shunt_gyp a_37652_43972# vss nmos_6p0 w=0.82u l=0.6u
X13969 a_2500_31836# cap_shunt_p a_2708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X13970 a_16500_25564# cap_shunt_n a_16708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X13971 vdd tune_shunt[7] a_25572_21236# vdd pmos_6p0 w=1.2u l=0.5u
X13972 vss tune_series_gygy[5] a_30616_19668# vss nmos_6p0 w=0.51u l=0.6u
X13973 a_16500_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X13974 a_29700_26786# cap_shunt_p a_29492_27132# vdd pmos_6p0 w=1.2u l=0.5u
X13975 a_23308_48983# a_23220_49080# vss vss nmos_6p0 w=0.82u l=1u
X13976 a_10660_45602# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X13977 vdd tune_shunt[5] a_21540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X13978 a_33048_14180# cap_series_gyp a_32632_14588# vss nmos_6p0 w=0.82u l=0.6u
X13979 vdd a_23084_47848# a_22996_47892# vdd pmos_6p0 w=1.22u l=1u
X13980 a_33500_36872# a_33412_36916# vss vss nmos_6p0 w=0.82u l=1u
X13981 a_6084_18100# cap_shunt_p a_6292_18584# vdd pmos_6p0 w=1.2u l=0.5u
X13982 a_10548_31128# cap_shunt_n a_11480_31128# vss nmos_6p0 w=0.82u l=0.6u
X13983 a_13460_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X13984 a_8860_11351# a_8772_11448# vss vss nmos_6p0 w=0.82u l=1u
X13985 a_37632_41240# cap_shunt_gyp a_37652_40836# vss nmos_6p0 w=0.82u l=0.6u
X13986 vss tune_series_gygy[3] a_35880_7124# vss nmos_6p0 w=0.51u l=0.6u
X13987 a_16500_22428# cap_shunt_n a_16708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X13988 a_20620_45847# a_20532_45944# vss vss nmos_6p0 w=0.82u l=1u
X13989 vss cap_shunt_n a_9856_37700# vss nmos_6p0 w=0.82u l=0.6u
X13990 vdd a_24204_25896# a_24116_25940# vdd pmos_6p0 w=1.22u l=1u
X13991 a_1716_5180# cap_shunt_p a_1924_4834# vdd pmos_6p0 w=1.2u l=0.5u
X13992 a_29720_9884# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X13993 a_27496_17016# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X13994 a_15720_11452# cap_series_gyp a_15532_11452# vdd pmos_6p0 w=1.2u l=0.5u
X13995 a_18716_55688# a_18628_55732# vss vss nmos_6p0 w=0.82u l=1u
X13996 vdd tune_shunt[7] a_21540_22428# vdd pmos_6p0 w=1.2u l=0.5u
X13997 a_33048_11044# cap_series_gyp a_32632_11452# vss nmos_6p0 w=0.82u l=0.6u
X13998 a_34144_49080# cap_shunt_gyn a_34144_48676# vdd pmos_6p0 w=1.215u l=0.5u
X13999 a_5152_38968# cap_shunt_n a_3828_38968# vss nmos_6p0 w=0.82u l=0.6u
X14000 vdd a_19276_31735# a_19188_31832# vdd pmos_6p0 w=1.22u l=1u
X14001 a_16708_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14002 a_6404_47170# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14003 a_29244_43144# a_29156_43188# vss vss nmos_6p0 w=0.82u l=1u
X14004 a_12608_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X14005 a_13796_33058# cap_shunt_n a_15512_32996# vss nmos_6p0 w=0.82u l=0.6u
X14006 a_23856_32996# cap_shunt_n a_21748_33058# vss nmos_6p0 w=0.82u l=0.6u
X14007 a_20620_42711# a_20532_42808# vss vss nmos_6p0 w=0.82u l=1u
X14008 a_2708_37762# cap_shunt_n a_2500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X14009 a_28484_24372# cap_shunt_p a_28692_24856# vdd pmos_6p0 w=1.2u l=0.5u
X14010 vdd a_24204_22760# a_24116_22804# vdd pmos_6p0 w=1.22u l=1u
X14011 vss cap_series_gyn a_13888_6040# vss nmos_6p0 w=0.82u l=0.6u
X14012 a_2588_49416# a_2500_49460# vss vss nmos_6p0 w=0.82u l=1u
X14013 a_37868_20759# a_37780_20856# vss vss nmos_6p0 w=0.82u l=1u
X14014 vdd tune_shunt[7] a_17620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X14015 vss tune_shunt[7] a_10548_37400# vss nmos_6p0 w=0.51u l=0.6u
X14016 a_16708_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14017 vss tune_shunt[4] a_28692_40536# vss nmos_6p0 w=0.51u l=0.6u
X14018 a_10660_34626# cap_shunt_n a_10452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X14019 a_21748_4834# cap_series_gyp a_21540_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14020 vss tune_series_gy[5] a_24660_14242# vss nmos_6p0 w=0.51u l=0.6u
X14021 a_12580_47892# cap_shunt_p a_12788_48376# vdd pmos_6p0 w=1.2u l=0.5u
X14022 a_6740_40536# cap_shunt_n a_6532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X14023 a_24660_28354# cap_shunt_n a_24452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X14024 a_2588_46280# a_2500_46324# vss vss nmos_6p0 w=0.82u l=1u
X14025 a_3828_38968# cap_shunt_n a_3620_38484# vdd pmos_6p0 w=1.2u l=0.5u
X14026 vdd tune_shunt[6] a_6532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X14027 a_30016_35832# cap_shunt_p a_28692_35832# vss nmos_6p0 w=0.82u l=0.6u
X14028 vss cap_series_gygyn a_37080_17016# vss nmos_6p0 w=0.82u l=0.6u
X14029 a_34308_19292# cap_series_gygyn a_34516_18946# vdd pmos_6p0 w=1.2u l=0.5u
X14030 vdd a_22860_48983# a_22772_49080# vdd pmos_6p0 w=1.22u l=1u
X14031 a_20172_38007# a_20084_38104# vss vss nmos_6p0 w=0.82u l=1u
X14032 a_30408_37400# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14033 vss tune_shunt[6] a_7748_45602# vss nmos_6p0 w=0.51u l=0.6u
X14034 vdd a_16028_29032# a_15940_29076# vdd pmos_6p0 w=1.22u l=1u
X14035 a_30476_47848# a_30388_47892# vss vss nmos_6p0 w=0.82u l=1u
X14036 a_10660_31490# cap_shunt_n a_10452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X14037 a_18044_7080# a_17956_7124# vss vss nmos_6p0 w=0.82u l=1u
X14038 vss tune_series_gy[5] a_24660_11106# vss nmos_6p0 w=0.51u l=0.6u
X14039 a_36296_18584# cap_series_gygyn a_35880_18100# vss nmos_6p0 w=0.82u l=0.6u
X14040 a_14728_23588# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14041 vss cap_series_gyn a_24752_12312# vss nmos_6p0 w=0.82u l=0.6u
X14042 vss tune_shunt[6] a_7748_36194# vss nmos_6p0 w=0.51u l=0.6u
X14043 a_3828_35832# cap_shunt_n a_3620_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14044 vdd tune_shunt[6] a_6532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14045 a_34308_16156# cap_series_gygyn a_34516_15810# vdd pmos_6p0 w=1.2u l=0.5u
X14046 a_31032_20152# cap_series_gygyn a_30616_19668# vss nmos_6p0 w=0.82u l=0.6u
X14047 vdd a_32716_5079# a_32628_5176# vdd pmos_6p0 w=1.22u l=1u
X14048 a_8456_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14049 a_2708_47170# cap_shunt_p a_2500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X14050 vdd a_35292_18056# a_35204_18100# vdd pmos_6p0 w=1.22u l=1u
X14051 a_36296_15448# cap_series_gygyn a_35880_14964# vss nmos_6p0 w=0.82u l=0.6u
X14052 a_2708_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14053 a_24660_34626# cap_shunt_p a_25592_34564# vss nmos_6p0 w=0.82u l=0.6u
X14054 a_13720_12312# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14055 a_30364_55255# a_30276_55352# vss vss nmos_6p0 w=0.82u l=1u
X14056 a_13588_47516# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14057 a_37652_39268# cap_shunt_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X14058 vss tune_shunt[7] a_7748_33058# vss nmos_6p0 w=0.51u l=0.6u
X14059 vss cap_series_gyp a_33832_14180# vss nmos_6p0 w=0.82u l=0.6u
X14060 a_33936_34564# cap_shunt_n a_32612_34626# vss nmos_6p0 w=0.82u l=0.6u
X14061 a_11572_3988# cap_series_gyp a_11780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X14062 a_26444_53687# a_26356_53784# vss vss nmos_6p0 w=0.82u l=1u
X14063 a_2500_25564# cap_shunt_p a_2708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X14064 vss tune_series_gy[5] a_18612_9538# vss nmos_6p0 w=0.51u l=0.6u
X14065 a_10452_38108# cap_shunt_n a_10660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X14066 a_6084_52220# cap_shunt_p a_6292_51874# vdd pmos_6p0 w=1.2u l=0.5u
X14067 a_6196_47516# cap_shunt_p a_6404_47170# vdd pmos_6p0 w=1.2u l=0.5u
X14068 a_22064_46808# cap_shunt_p a_20740_46808# vss nmos_6p0 w=0.82u l=0.6u
X14069 a_24660_31490# cap_shunt_p a_25592_31428# vss nmos_6p0 w=0.82u l=0.6u
X14070 vdd a_19724_30167# a_19636_30264# vdd pmos_6p0 w=1.22u l=1u
X14071 a_16500_19292# cap_shunt_p a_16708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X14072 a_20740_20152# cap_shunt_p a_20532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X14073 a_16500_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14074 vss tune_shunt[4] a_29700_23650# vss nmos_6p0 w=0.51u l=0.6u
X14075 vss cap_series_gyp a_33832_11044# vss nmos_6p0 w=0.82u l=0.6u
X14076 a_6740_20152# cap_shunt_p a_7672_20152# vss nmos_6p0 w=0.82u l=0.6u
X14077 a_10660_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14078 a_33936_31428# cap_shunt_n a_32612_31490# vss nmos_6p0 w=0.82u l=0.6u
X14079 a_34664_27992# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14080 a_28572_22327# a_28484_22424# vss vss nmos_6p0 w=0.82u l=1u
X14081 a_26444_50551# a_26356_50648# vss vss nmos_6p0 w=0.82u l=1u
X14082 a_4424_39268# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14083 a_34508_39575# a_34420_39672# vss vss nmos_6p0 w=0.82u l=1u
X14084 a_6760_5556# cap_series_gyp a_6572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X14085 vdd tune_shunt[7] a_21540_19292# vdd pmos_6p0 w=1.2u l=0.5u
X14086 vss tune_shunt[7] a_12788_18584# vss nmos_6p0 w=0.51u l=0.6u
X14087 a_1692_20759# a_1604_20856# vss vss nmos_6p0 w=0.82u l=1u
X14088 a_2500_22428# cap_shunt_p a_2708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X14089 vss cap_shunt_p a_3248_6040# vss nmos_6p0 w=0.82u l=0.6u
X14090 a_16500_16156# cap_shunt_p a_16708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X14091 a_18516_5556# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14092 vdd a_19276_25463# a_19188_25560# vdd pmos_6p0 w=1.22u l=1u
X14093 vdd tune_series_gy[5] a_21540_16156# vdd pmos_6p0 w=1.2u l=0.5u
X14094 vdd a_17148_53687# a_17060_53784# vdd pmos_6p0 w=1.22u l=1u
X14095 vss tune_series_gy[4] a_21636_6040# vss nmos_6p0 w=0.51u l=0.6u
X14096 vss tune_shunt[7] a_12788_15448# vss nmos_6p0 w=0.51u l=0.6u
X14097 a_26892_54120# a_26804_54164# vss vss nmos_6p0 w=0.82u l=1u
X14098 a_24452_42812# cap_shunt_n a_24660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X14099 vdd a_29580_55688# a_29492_55732# vdd pmos_6p0 w=1.22u l=1u
X14100 a_20620_36439# a_20532_36536# vss vss nmos_6p0 w=0.82u l=1u
X14101 a_18612_11106# cap_series_gyn a_18404_11452# vdd pmos_6p0 w=1.2u l=0.5u
X14102 a_31436_20860# cap_series_gygyn a_31624_20860# vdd pmos_6p0 w=1.2u l=0.5u
X14103 a_11460_46324# cap_shunt_n a_11668_46808# vdd pmos_6p0 w=1.2u l=0.5u
X14104 a_28484_7124# cap_series_gyp a_28692_7608# vdd pmos_6p0 w=1.2u l=0.5u
X14105 vdd a_24204_16488# a_24116_16532# vdd pmos_6p0 w=1.22u l=1u
X14106 a_6532_52596# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14107 a_16708_47170# cap_shunt_n a_16500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X14108 a_12264_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14109 a_6404_22082# cap_shunt_p a_6196_22428# vdd pmos_6p0 w=1.2u l=0.5u
X14110 a_37868_14487# a_37780_14584# vss vss nmos_6p0 w=0.82u l=1u
X14111 a_35600_47893# cap_shunt_gyp a_35600_48438# vdd pmos_6p0 w=1.215u l=0.5u
X14112 vdd a_19276_22327# a_19188_22424# vdd pmos_6p0 w=1.22u l=1u
X14113 a_18404_8316# cap_series_gyp a_18612_7970# vdd pmos_6p0 w=1.2u l=0.5u
X14114 a_16708_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14115 vss tune_shunt[6] a_28692_34264# vss nmos_6p0 w=0.51u l=0.6u
X14116 a_33524_27508# cap_shunt_p a_33732_27992# vdd pmos_6p0 w=1.2u l=0.5u
X14117 a_9072_29860# cap_shunt_n a_7748_29922# vss nmos_6p0 w=0.82u l=0.6u
X14118 a_13796_23650# cap_shunt_n a_15512_23588# vss nmos_6p0 w=0.82u l=0.6u
X14119 a_23868_54120# a_23780_54164# vss vss nmos_6p0 w=0.82u l=1u
X14120 a_23856_23588# cap_shunt_p a_21748_23650# vss nmos_6p0 w=0.82u l=0.6u
X14121 vdd tune_shunt[7] a_13588_34972# vdd pmos_6p0 w=1.2u l=0.5u
X14122 vdd a_5836_3944# a_5748_3988# vdd pmos_6p0 w=1.22u l=1u
X14123 vdd a_26556_55688# a_26468_55732# vdd pmos_6p0 w=1.22u l=1u
X14124 a_12264_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14125 a_37868_11351# a_37780_11448# vss vss nmos_6p0 w=0.82u l=1u
X14126 a_9332_11452# cap_shunt_p a_9540_11106# vdd pmos_6p0 w=1.2u l=0.5u
X14127 vdd tune_series_gygy[5] a_35692_19668# vdd pmos_6p0 w=1.2u l=0.5u
X14128 a_27788_47415# a_27700_47512# vss vss nmos_6p0 w=0.82u l=1u
X14129 a_30016_29560# cap_shunt_p a_28692_29560# vss nmos_6p0 w=0.82u l=0.6u
X14130 a_18404_5180# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14131 vss tune_shunt[6] a_7748_39330# vss nmos_6p0 w=0.51u l=0.6u
X14132 vss tune_shunt[5] a_28692_31128# vss nmos_6p0 w=0.51u l=0.6u
X14133 a_21540_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14134 a_19544_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14135 a_9072_26724# cap_shunt_n a_7748_26786# vss nmos_6p0 w=0.82u l=0.6u
X14136 a_10660_25218# cap_shunt_n a_10452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X14137 vss cap_series_gyn a_12768_6340# vss nmos_6p0 w=0.82u l=0.6u
X14138 vdd tune_shunt[7] a_13588_31836# vdd pmos_6p0 w=1.2u l=0.5u
X14139 vss tune_shunt[7] a_17828_27992# vss nmos_6p0 w=0.51u l=0.6u
X14140 vdd a_13788_50984# a_13700_51028# vdd pmos_6p0 w=1.22u l=1u
X14141 a_6740_46808# cap_shunt_p a_8456_46808# vss nmos_6p0 w=0.82u l=0.6u
X14142 a_3828_29560# cap_shunt_n a_3620_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14143 a_20328_4772# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X14144 vdd tune_shunt[7] a_6532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14145 a_30016_26424# cap_shunt_p a_28692_26424# vss nmos_6p0 w=0.82u l=0.6u
X14146 vdd a_16924_52552# a_16836_52596# vdd pmos_6p0 w=1.22u l=1u
X14147 a_19724_48983# a_19636_49080# vss vss nmos_6p0 w=0.82u l=1u
X14148 a_18180_3612# cap_series_gyn a_18388_3266# vdd pmos_6p0 w=1.2u l=0.5u
X14149 a_29196_3612# tune_series_gy[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14150 a_32268_5079# a_32180_5176# vss vss nmos_6p0 w=0.82u l=1u
X14151 a_20720_4472# cap_series_gyp a_18612_4472# vss nmos_6p0 w=0.82u l=0.6u
X14152 a_13588_13020# cap_shunt_p a_13796_12674# vdd pmos_6p0 w=1.2u l=0.5u
X14153 vss tune_shunt[7] a_17828_24856# vss nmos_6p0 w=0.51u l=0.6u
X14154 a_24660_28354# cap_shunt_n a_25592_28292# vss nmos_6p0 w=0.82u l=0.6u
X14155 vss cap_series_gyn a_8968_4772# vss nmos_6p0 w=0.82u l=0.6u
X14156 a_36972_55688# a_36884_55732# vss vss nmos_6p0 w=0.82u l=1u
X14157 a_30364_48983# a_30276_49080# vss vss nmos_6p0 w=0.82u l=1u
X14158 a_33936_28292# cap_shunt_p a_32612_28354# vss nmos_6p0 w=0.82u l=0.6u
X14159 vdd tune_series_gy[2] a_10452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14160 a_8456_23288# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14161 a_2708_37762# cap_shunt_n a_2500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X14162 a_20740_32696# cap_shunt_n a_21672_32696# vss nmos_6p0 w=0.82u l=0.6u
X14163 vdd tune_shunt[1] a_25572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X14164 a_2500_19292# cap_shunt_p a_2708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X14165 vdd a_31260_25896# a_31172_25940# vdd pmos_6p0 w=1.22u l=1u
X14166 a_2708_22082# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14167 a_19524_10260# cap_series_gyn a_19732_10744# vdd pmos_6p0 w=1.2u l=0.5u
X14168 vss cap_shunt_p a_15904_45240# vss nmos_6p0 w=0.82u l=0.6u
X14169 a_24660_25218# cap_shunt_p a_25592_25156# vss nmos_6p0 w=0.82u l=0.6u
X14170 vss tune_series_gy[2] a_7768_8316# vss nmos_6p0 w=0.51u l=0.6u
X14171 a_13588_38108# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14172 a_10660_34626# cap_shunt_n a_10452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X14173 a_21540_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14174 a_31708_5512# a_31620_5556# vss vss nmos_6p0 w=0.82u l=1u
X14175 a_33948_55688# a_33860_55732# vss vss nmos_6p0 w=0.82u l=1u
X14176 a_12580_47892# cap_shunt_p a_12788_48376# vdd pmos_6p0 w=1.2u l=0.5u
X14177 a_13460_38968# cap_shunt_n a_13252_38484# vdd pmos_6p0 w=1.2u l=0.5u
X14178 a_33936_25156# cap_shunt_p a_32612_25218# vss nmos_6p0 w=0.82u l=0.6u
X14179 a_24660_28354# cap_shunt_n a_24452_28700# vdd pmos_6p0 w=1.2u l=0.5u
X14180 vdd a_5612_23895# a_5524_23992# vdd pmos_6p0 w=1.22u l=1u
X14181 a_2708_22082# cap_shunt_p a_4424_22020# vss nmos_6p0 w=0.82u l=0.6u
X14182 a_21540_9884# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14183 a_31416_29860# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14184 a_17828_27992# cap_shunt_n a_18760_27992# vss nmos_6p0 w=0.82u l=0.6u
X14185 vss cap_shunt_n a_4032_9476# vss nmos_6p0 w=0.82u l=0.6u
X14186 a_1692_14487# a_1604_14584# vss vss nmos_6p0 w=0.82u l=1u
X14187 a_2500_16156# cap_shunt_p a_2708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X14188 a_27228_33303# a_27140_33400# vss vss nmos_6p0 w=0.82u l=1u
X14189 vdd a_31260_22760# a_31172_22804# vdd pmos_6p0 w=1.22u l=1u
X14190 vss cap_shunt_n a_15904_42104# vss nmos_6p0 w=0.82u l=0.6u
X14191 vdd a_36300_35304# a_36212_35348# vdd pmos_6p0 w=1.22u l=1u
X14192 vss tune_series_gy[1] a_7768_5180# vss nmos_6p0 w=0.51u l=0.6u
X14193 vss tune_series_gy[5] a_29700_14242# vss nmos_6p0 w=0.51u l=0.6u
X14194 a_24652_19624# a_24564_19668# vss vss nmos_6p0 w=0.82u l=1u
X14195 a_19388_52119# a_19300_52216# vss vss nmos_6p0 w=0.82u l=1u
X14196 a_9876_51512# cap_shunt_n a_10808_51512# vss nmos_6p0 w=0.82u l=0.6u
X14197 a_17620_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14198 a_10660_31490# cap_shunt_n a_10452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X14199 a_13460_35832# cap_shunt_n a_13252_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14200 a_21540_6748# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14201 vdd a_5612_20759# a_5524_20856# vdd pmos_6p0 w=1.22u l=1u
X14202 a_34480_46325# cap_shunt_gyn a_34480_46870# vdd pmos_6p0 w=1.215u l=0.5u
X14203 a_31416_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14204 a_17828_24856# cap_shunt_n a_18760_24856# vss nmos_6p0 w=0.82u l=0.6u
X14205 a_35692_18100# cap_series_gygyn a_35880_18100# vdd pmos_6p0 w=1.2u l=0.5u
X14206 a_26892_47848# a_26804_47892# vss vss nmos_6p0 w=0.82u l=1u
X14207 a_18032_45540# cap_shunt_p a_16708_45602# vss nmos_6p0 w=0.82u l=0.6u
X14208 vdd a_34396_40008# a_34308_40052# vdd pmos_6p0 w=1.22u l=1u
X14209 a_21636_6040# cap_series_gyp a_21428_5556# vdd pmos_6p0 w=1.2u l=0.5u
X14210 a_1692_11351# a_1604_11448# vss vss nmos_6p0 w=0.82u l=1u
X14211 a_2500_20860# cap_shunt_p a_2708_20514# vdd pmos_6p0 w=1.2u l=0.5u
X14212 a_24452_36540# cap_shunt_p a_24660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X14213 vdd a_29580_49416# a_29492_49460# vdd pmos_6p0 w=1.22u l=1u
X14214 vss tune_series_gy[4] a_29700_11106# vss nmos_6p0 w=0.51u l=0.6u
X14215 vdd a_19276_16055# a_19188_16152# vdd pmos_6p0 w=1.22u l=1u
X14216 a_18032_42404# cap_shunt_n a_16708_42466# vss nmos_6p0 w=0.82u l=0.6u
X14217 a_24452_33404# cap_shunt_p a_24660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X14218 a_7540_30268# cap_shunt_n a_7748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X14219 vdd a_29580_46280# a_29492_46324# vdd pmos_6p0 w=1.22u l=1u
X14220 a_3620_13396# cap_shunt_n a_3828_13880# vdd pmos_6p0 w=1.2u l=0.5u
X14221 a_36624_18884# cap_series_gygyn a_34516_18946# vss nmos_6p0 w=0.82u l=0.6u
X14222 a_6532_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14223 a_25572_41620# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14224 a_3620_19668# cap_shunt_p a_3828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X14225 vss tune_shunt[7] a_9876_20152# vss nmos_6p0 w=0.51u l=0.6u
X14226 a_16708_37762# cap_shunt_n a_16500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X14227 a_7748_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14228 a_2708_47170# cap_shunt_p a_3640_47108# vss nmos_6p0 w=0.82u l=0.6u
X14229 a_10452_38108# cap_shunt_n a_10660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X14230 a_20740_43672# cap_shunt_n a_20532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X14231 a_21748_4834# cap_series_gyp a_22680_4772# vss nmos_6p0 w=0.82u l=0.6u
X14232 a_18760_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14233 vdd tune_shunt[7] a_10340_25940# vdd pmos_6p0 w=1.2u l=0.5u
X14234 a_12788_48376# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14235 a_37444_41240# cap_shunt_gyp a_37632_41240# vdd pmos_6p0 w=1.215u l=0.5u
X14236 a_36624_15748# cap_series_gygyn a_34516_15810# vss nmos_6p0 w=0.82u l=0.6u
X14237 vdd a_15356_49416# a_15268_49460# vdd pmos_6p0 w=1.22u l=1u
X14238 a_14372_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14239 vdd tune_shunt[7] a_13588_25564# vdd pmos_6p0 w=1.2u l=0.5u
X14240 a_19524_8692# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14241 a_17828_48376# cap_shunt_p a_19544_48376# vss nmos_6p0 w=0.82u l=0.6u
X14242 a_23756_55255# a_23668_55352# vss vss nmos_6p0 w=0.82u l=1u
X14243 a_19836_53687# a_19748_53784# vss vss nmos_6p0 w=0.82u l=1u
X14244 vdd tune_shunt[7] a_10340_22804# vdd pmos_6p0 w=1.2u l=0.5u
X14245 a_2588_52119# a_2500_52216# vss vss nmos_6p0 w=0.82u l=1u
X14246 vss cap_shunt_n a_15568_35832# vss nmos_6p0 w=0.82u l=0.6u
X14247 vdd tune_shunt[7] a_13588_22428# vdd pmos_6p0 w=1.2u l=0.5u
X14248 vss tune_shunt[7] a_17828_18584# vss nmos_6p0 w=0.51u l=0.6u
X14249 a_10548_32696# cap_shunt_n a_10340_32212# vdd pmos_6p0 w=1.2u l=0.5u
X14250 a_35692_7124# cap_series_gygyp a_35880_7124# vdd pmos_6p0 w=1.2u l=0.5u
X14251 a_1716_5556# tune_shunt[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14252 a_30016_17016# cap_series_gyn a_28692_17016# vss nmos_6p0 w=0.82u l=0.6u
X14253 a_24452_42812# cap_shunt_n a_24660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X14254 a_1692_9783# a_1604_9880# vss vss nmos_6p0 w=0.82u l=1u
X14255 a_9876_53080# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14256 a_19724_39575# a_19636_39672# vss vss nmos_6p0 w=0.82u l=1u
X14257 a_18612_11106# cap_series_gyn a_18404_11452# vdd pmos_6p0 w=1.2u l=0.5u
X14258 a_11460_46324# cap_shunt_n a_11668_46808# vdd pmos_6p0 w=1.2u l=0.5u
X14259 vss cap_shunt_p a_27888_27992# vss nmos_6p0 w=0.82u l=0.6u
X14260 a_7672_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14261 a_6404_22082# cap_shunt_p a_6196_22428# vdd pmos_6p0 w=1.2u l=0.5u
X14262 a_12788_13880# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14263 a_33524_27508# cap_shunt_p a_33732_27992# vdd pmos_6p0 w=1.2u l=0.5u
X14264 vss tune_shunt[7] a_17828_15448# vss nmos_6p0 w=0.51u l=0.6u
X14265 vdd a_36524_31735# a_36436_31832# vdd pmos_6p0 w=1.22u l=1u
X14266 vss tune_shunt[6] a_17828_38968# vss nmos_6p0 w=0.51u l=0.6u
X14267 vss cap_shunt_p a_27888_24856# vss nmos_6p0 w=0.82u l=0.6u
X14268 a_24660_20514# cap_shunt_p a_24452_20860# vdd pmos_6p0 w=1.2u l=0.5u
X14269 vdd a_16476_38440# a_16388_38484# vdd pmos_6p0 w=1.22u l=1u
X14270 a_20740_23288# cap_shunt_p a_21672_23288# vss nmos_6p0 w=0.82u l=0.6u
X14271 vdd a_12444_19191# a_12356_19288# vdd pmos_6p0 w=1.22u l=1u
X14272 a_17620_19668# cap_shunt_p a_17828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X14273 a_28796_21192# a_28708_21236# vss vss nmos_6p0 w=0.82u l=1u
X14274 a_10340_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14275 vdd a_31260_16488# a_31172_16532# vdd pmos_6p0 w=1.22u l=1u
X14276 vdd a_36300_29032# a_36212_29076# vdd pmos_6p0 w=1.22u l=1u
X14277 a_10660_25218# cap_shunt_n a_10452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X14278 a_34308_22428# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14279 vss tune_series_gygy[5] a_34516_22082# vss nmos_6p0 w=0.51u l=0.6u
X14280 vdd a_33500_7080# a_33412_7124# vdd pmos_6p0 w=1.22u l=1u
X14281 vdd a_9644_33736# a_9556_33780# vdd pmos_6p0 w=1.22u l=1u
X14282 a_13460_29560# cap_shunt_n a_13252_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14283 vdd a_5612_14487# a_5524_14584# vdd pmos_6p0 w=1.22u l=1u
X14284 vdd a_16476_35304# a_16388_35348# vdd pmos_6p0 w=1.22u l=1u
X14285 a_17828_18584# cap_shunt_p a_18760_18584# vss nmos_6p0 w=0.82u l=0.6u
X14286 a_10340_35348# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14287 a_2500_34972# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14288 a_32824_6340# cap_series_gygyn a_31624_6748# vss nmos_6p0 w=0.82u l=0.6u
X14289 a_27228_23895# a_27140_23992# vss vss nmos_6p0 w=0.82u l=1u
X14290 a_16408_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X14291 vss tune_shunt[6] a_20740_35832# vss nmos_6p0 w=0.51u l=0.6u
X14292 vdd a_9644_30600# a_9556_30644# vdd pmos_6p0 w=1.22u l=1u
X14293 a_1716_7124# cap_shunt_n a_1924_7608# vdd pmos_6p0 w=1.2u l=0.5u
X14294 a_11780_4472# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X14295 a_2500_11452# cap_shunt_n a_2708_11106# vdd pmos_6p0 w=1.2u l=0.5u
X14296 a_17828_15448# cap_shunt_p a_18760_15448# vss nmos_6p0 w=0.82u l=0.6u
X14297 a_31416_17316# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X14298 vss cap_shunt_n a_12768_45540# vss nmos_6p0 w=0.82u l=0.6u
X14299 a_18032_36132# cap_shunt_n a_16708_36194# vss nmos_6p0 w=0.82u l=0.6u
X14300 vdd a_6060_34871# a_5972_34968# vdd pmos_6p0 w=1.22u l=1u
X14301 a_2500_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14302 a_24452_27132# cap_shunt_p a_24660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X14303 a_10548_3266# cap_series_gyn a_11480_3204# vss nmos_6p0 w=0.82u l=0.6u
X14304 a_3380_49944# cap_shunt_p a_4312_49944# vss nmos_6p0 w=0.82u l=0.6u
X14305 a_24660_9538# cap_series_gyn a_24452_9884# vdd pmos_6p0 w=1.2u l=0.5u
X14306 vss cap_shunt_p a_34720_37700# vss nmos_6p0 w=0.82u l=0.6u
X14307 a_16708_29922# cap_shunt_n a_16500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X14308 a_2500_49084# cap_shunt_p a_2708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X14309 a_7540_28700# cap_shunt_n a_7748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X14310 a_12788_13880# cap_shunt_p a_12580_13396# vdd pmos_6p0 w=1.2u l=0.5u
X14311 a_13796_48738# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14312 a_18760_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14313 vdd a_27676_5079# a_27588_5176# vdd pmos_6p0 w=1.22u l=1u
X14314 a_19732_12312# cap_series_gyn a_19524_11828# vdd pmos_6p0 w=1.2u l=0.5u
X14315 a_2708_42466# cap_shunt_p a_2500_42812# vdd pmos_6p0 w=1.2u l=0.5u
X14316 vss cap_shunt_n a_12768_42404# vss nmos_6p0 w=0.82u l=0.6u
X14317 a_21748_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14318 a_13460_38968# cap_shunt_n a_13252_38484# vdd pmos_6p0 w=1.2u l=0.5u
X14319 a_15512_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14320 a_25572_32212# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14321 vdd tune_shunt[7] a_13588_19292# vdd pmos_6p0 w=1.2u l=0.5u
X14322 vss tune_shunt[6] a_6740_37400# vss nmos_6p0 w=0.51u l=0.6u
X14323 a_20532_36916# cap_shunt_n a_20740_37400# vdd pmos_6p0 w=1.2u l=0.5u
X14324 a_9108_49084# cap_shunt_p a_9316_48738# vdd pmos_6p0 w=1.2u l=0.5u
X14325 a_24660_6402# cap_series_gyn a_24452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X14326 a_11984_43972# cap_shunt_n a_10660_44034# vss nmos_6p0 w=0.82u l=0.6u
X14327 a_23756_48983# a_23668_49080# vss vss nmos_6p0 w=0.82u l=1u
X14328 a_18760_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14329 a_13460_35832# cap_shunt_n a_13252_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14330 vss cap_shunt_n a_15568_29560# vss nmos_6p0 w=0.82u l=0.6u
X14331 vdd tune_shunt[7] a_13588_16156# vdd pmos_6p0 w=1.2u l=0.5u
X14332 vdd a_37420_53687# a_37332_53784# vdd pmos_6p0 w=1.22u l=1u
X14333 a_32268_12919# a_32180_13016# vss vss nmos_6p0 w=0.82u l=1u
X14334 a_25548_50984# a_25460_51028# vss vss nmos_6p0 w=0.82u l=1u
X14335 vdd a_24652_25896# a_24564_25940# vdd pmos_6p0 w=1.22u l=1u
X14336 a_34396_22760# a_34308_22804# vss vss nmos_6p0 w=0.82u l=1u
X14337 a_12788_17016# cap_shunt_p a_12580_16532# vdd pmos_6p0 w=1.2u l=0.5u
X14338 a_11984_40836# cap_shunt_n a_10660_40898# vss nmos_6p0 w=0.82u l=0.6u
X14339 a_24452_36540# cap_shunt_p a_24660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X14340 a_36652_48676# cap_shunt_gyn a_36384_48676# vss nmos_6p0 w=0.82u l=0.6u
X14341 a_28692_38968# cap_shunt_n a_28484_38484# vdd pmos_6p0 w=1.2u l=0.5u
X14342 vss tune_shunt[1] a_5844_3266# vss nmos_6p0 w=0.51u l=0.6u
X14343 a_29692_43144# a_29604_43188# vss vss nmos_6p0 w=0.82u l=1u
X14344 a_7748_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14345 vss tune_shunt[7] a_13460_32696# vss nmos_6p0 w=0.51u l=0.6u
X14346 vss cap_shunt_p a_4032_32996# vss nmos_6p0 w=0.82u l=0.6u
X14347 vss cap_shunt_n a_15568_26424# vss nmos_6p0 w=0.82u l=0.6u
X14348 vdd a_36524_25463# a_36436_25560# vdd pmos_6p0 w=1.22u l=1u
X14349 vdd a_24652_22760# a_24564_22804# vdd pmos_6p0 w=1.22u l=1u
X14350 a_34308_19292# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14351 a_24452_33404# cap_shunt_p a_24660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X14352 a_28692_35832# cap_shunt_p a_28484_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14353 a_14784_27992# cap_shunt_n a_13460_27992# vss nmos_6p0 w=0.82u l=0.6u
X14354 a_2932_12312# cap_shunt_n a_2724_11828# vdd pmos_6p0 w=1.2u l=0.5u
X14355 vss cap_series_gyn a_27888_18584# vss nmos_6p0 w=0.82u l=0.6u
X14356 a_3620_43188# cap_shunt_p a_3828_43672# vdd pmos_6p0 w=1.2u l=0.5u
X14357 vss cap_shunt_n a_11984_53080# vss nmos_6p0 w=0.82u l=0.6u
X14358 a_10452_38108# cap_shunt_n a_10660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X14359 a_25572_8692# cap_series_gyp a_25780_9176# vdd pmos_6p0 w=1.2u l=0.5u
X14360 a_9428_17378# cap_shunt_p a_9220_17724# vdd pmos_6p0 w=1.2u l=0.5u
X14361 vss cap_shunt_gyp a_36652_43972# vss nmos_6p0 w=0.82u l=0.6u
X14362 vdd tune_series_gygy[3] a_34348_9884# vdd pmos_6p0 w=1.2u l=0.5u
X14363 a_15492_9884# cap_series_gyn a_15700_9538# vdd pmos_6p0 w=1.2u l=0.5u
X14364 a_34308_16156# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14365 vdd tune_shunt[7] a_10340_25940# vdd pmos_6p0 w=1.2u l=0.5u
X14366 a_14784_24856# cap_shunt_n a_13460_24856# vss nmos_6p0 w=0.82u l=0.6u
X14367 a_24660_11106# cap_series_gyp a_24452_11452# vdd pmos_6p0 w=1.2u l=0.5u
X14368 vss cap_series_gyp a_27888_15448# vss nmos_6p0 w=0.82u l=0.6u
X14369 vdd a_16476_29032# a_16388_29076# vdd pmos_6p0 w=1.22u l=1u
X14370 vdd tune_shunt[7] a_2500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X14371 vss tune_series_gy[4] a_28692_12312# vss nmos_6p0 w=0.51u l=0.6u
X14372 a_10340_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14373 a_25572_5556# cap_series_gyp a_25780_6040# vdd pmos_6p0 w=1.2u l=0.5u
X14374 a_1716_8316# cap_shunt_n a_1924_7970# vdd pmos_6p0 w=1.2u l=0.5u
X14375 a_34844_8648# a_34756_8692# vss vss nmos_6p0 w=0.82u l=1u
X14376 a_37080_9176# cap_series_gygyn a_35880_8692# vss nmos_6p0 w=0.82u l=0.6u
X14377 vdd a_33948_14920# a_33860_14964# vdd pmos_6p0 w=1.22u l=1u
X14378 vss cap_shunt_gyp a_36652_40836# vss nmos_6p0 w=0.82u l=0.6u
X14379 a_15492_6748# cap_series_gyp a_15700_6402# vdd pmos_6p0 w=1.2u l=0.5u
X14380 vdd tune_series_gygy[2] a_34348_6748# vdd pmos_6p0 w=1.2u l=0.5u
X14381 vdd tune_shunt[7] a_10340_22804# vdd pmos_6p0 w=1.2u l=0.5u
X14382 a_25444_3266# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X14383 vss tune_shunt[7] a_20740_29560# vss nmos_6p0 w=0.51u l=0.6u
X14384 vdd a_9644_24328# a_9556_24372# vdd pmos_6p0 w=1.22u l=1u
X14385 a_22644_10744# cap_series_gyp a_22436_10260# vdd pmos_6p0 w=1.2u l=0.5u
X14386 vdd a_6060_28599# a_5972_28696# vdd pmos_6p0 w=1.22u l=1u
X14387 a_17596_11784# a_17508_11828# vss vss nmos_6p0 w=0.82u l=1u
X14388 a_24452_42812# cap_shunt_n a_24660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X14389 a_2500_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14390 vdd a_33948_11784# a_33860_11828# vdd pmos_6p0 w=1.22u l=1u
X14391 a_10540_54120# a_10452_54164# vss vss nmos_6p0 w=0.82u l=1u
X14392 a_2708_29922# cap_shunt_n a_2500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X14393 vss tune_shunt[7] a_20740_26424# vss nmos_6p0 w=0.51u l=0.6u
X14394 vdd a_5388_7080# a_5300_7124# vdd pmos_6p0 w=1.22u l=1u
X14395 a_21748_7970# cap_series_gyp a_21540_8316# vdd pmos_6p0 w=1.2u l=0.5u
X14396 a_26892_53687# a_26804_53784# vss vss nmos_6p0 w=0.82u l=1u
X14397 vss cap_shunt_n a_12768_36132# vss nmos_6p0 w=0.82u l=0.6u
X14398 a_2500_22428# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14399 a_28692_9176# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X14400 a_2708_36194# cap_shunt_n a_2500_36540# vdd pmos_6p0 w=1.2u l=0.5u
X14401 vss cap_shunt_p a_30800_35832# vss nmos_6p0 w=0.82u l=0.6u
X14402 a_16708_28354# cap_shunt_n a_16500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X14403 a_24660_20514# cap_shunt_p a_24452_20860# vdd pmos_6p0 w=1.2u l=0.5u
X14404 vdd a_25100_55255# a_25012_55352# vdd pmos_6p0 w=1.22u l=1u
X14405 a_1692_43144# a_1604_43188# vss vss nmos_6p0 w=0.82u l=1u
X14406 a_34956_39575# a_34868_39672# vss vss nmos_6p0 w=0.82u l=1u
X14407 a_26892_50551# a_26804_50648# vss vss nmos_6p0 w=0.82u l=1u
X14408 vss tune_shunt[4] a_20740_46808# vss nmos_6p0 w=0.51u l=0.6u
X14409 vss cap_shunt_n a_4816_50244# vss nmos_6p0 w=0.82u l=0.6u
X14410 a_35532_47108# cap_shunt_gyn a_35264_47108# vss nmos_6p0 w=0.82u l=0.6u
X14411 a_2708_33058# cap_shunt_p a_2500_33404# vdd pmos_6p0 w=1.2u l=0.5u
X14412 a_13460_29560# cap_shunt_n a_13252_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14413 vss tune_series_gy[5] a_19732_7608# vss nmos_6p0 w=0.51u l=0.6u
X14414 a_35692_7124# cap_series_gygyp a_35880_7124# vdd pmos_6p0 w=1.2u l=0.5u
X14415 a_23464_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14416 a_25548_44712# a_25460_44756# vss vss nmos_6p0 w=0.82u l=1u
X14417 a_20532_27508# cap_shunt_n a_20740_27992# vdd pmos_6p0 w=1.2u l=0.5u
X14418 vdd a_25100_52119# a_25012_52216# vdd pmos_6p0 w=1.22u l=1u
X14419 a_11984_34564# cap_shunt_n a_10660_34626# vss nmos_6p0 w=0.82u l=0.6u
X14420 vss cap_series_gygyn a_37080_9176# vss nmos_6p0 w=0.82u l=0.6u
X14421 a_35692_10260# cap_series_gygyp a_35880_10260# vdd pmos_6p0 w=1.2u l=0.5u
X14422 a_1692_40008# a_1604_40052# vss vss nmos_6p0 w=0.82u l=1u
X14423 vdd a_6508_45847# a_6420_45944# vdd pmos_6p0 w=1.22u l=1u
X14424 a_7748_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14425 a_18760_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14426 a_6740_20152# cap_shunt_p a_6532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X14427 a_31820_55688# a_31732_55732# vss vss nmos_6p0 w=0.82u l=1u
X14428 vdd a_17596_53687# a_17508_53784# vdd pmos_6p0 w=1.22u l=1u
X14429 a_10092_46280# a_10004_46324# vss vss nmos_6p0 w=0.82u l=1u
X14430 a_36636_52119# a_36548_52216# vss vss nmos_6p0 w=0.82u l=1u
X14431 a_3828_43672# cap_shunt_p a_5544_43672# vss nmos_6p0 w=0.82u l=0.6u
X14432 a_3380_17016# cap_shunt_p a_3172_16532# vdd pmos_6p0 w=1.2u l=0.5u
X14433 vss tune_series_gygy[5] a_35880_19668# vss nmos_6p0 w=0.51u l=0.6u
X14434 a_6740_42104# cap_shunt_n a_6532_41620# vdd pmos_6p0 w=1.2u l=0.5u
X14435 vdd a_24652_16488# a_24564_16532# vdd pmos_6p0 w=1.22u l=1u
X14436 a_35880_19668# cap_series_gygyp a_35692_19668# vdd pmos_6p0 w=1.2u l=0.5u
X14437 vss tune_shunt[6] a_10660_44034# vss nmos_6p0 w=0.51u l=0.6u
X14438 a_11984_31428# cap_shunt_n a_10660_31490# vss nmos_6p0 w=0.82u l=0.6u
X14439 a_24452_27132# cap_shunt_p a_24660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X14440 a_36296_4472# cap_series_gygyp a_35880_3988# vss nmos_6p0 w=0.82u l=0.6u
X14441 a_2500_9884# cap_shunt_n a_2708_9538# vdd pmos_6p0 w=1.2u l=0.5u
X14442 a_28692_29560# cap_shunt_p a_28484_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14443 vdd a_6508_42711# a_6420_42808# vdd pmos_6p0 w=1.22u l=1u
X14444 a_7748_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14445 a_24452_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14446 vss tune_shunt[7] a_13460_23288# vss nmos_6p0 w=0.51u l=0.6u
X14447 vss tune_shunt[4] a_3828_13880# vss nmos_6p0 w=0.51u l=0.6u
X14448 a_3828_40536# cap_shunt_n a_5544_40536# vss nmos_6p0 w=0.82u l=0.6u
X14449 vss cap_shunt_p a_4032_23588# vss nmos_6p0 w=0.82u l=0.6u
X14450 vss cap_series_gygyn a_35840_17316# vss nmos_6p0 w=0.82u l=0.6u
X14451 a_2500_49084# cap_shunt_p a_2708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X14452 a_16708_29922# cap_shunt_n a_16500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X14453 a_3828_37400# cap_shunt_n a_3620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X14454 vss tune_series_gygy[3] a_35880_8692# vss nmos_6p0 w=0.51u l=0.6u
X14455 a_9108_49084# cap_shunt_p a_9316_48738# vdd pmos_6p0 w=1.2u l=0.5u
X14456 a_29720_9884# cap_series_gyn a_29532_9884# vdd pmos_6p0 w=1.2u l=0.5u
X14457 a_2932_12312# cap_shunt_n a_4648_12312# vss nmos_6p0 w=0.82u l=0.6u
X14458 a_12788_49944# cap_shunt_n a_12580_49460# vdd pmos_6p0 w=1.2u l=0.5u
X14459 a_21672_37400# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14460 a_18816_22020# cap_shunt_n a_16708_22082# vss nmos_6p0 w=0.82u l=0.6u
X14461 a_13588_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14462 vss tune_shunt[7] a_21748_29922# vss nmos_6p0 w=0.51u l=0.6u
X14463 a_32404_28700# cap_shunt_p a_32612_28354# vdd pmos_6p0 w=1.2u l=0.5u
X14464 a_19732_12312# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14465 a_21740_47848# a_21652_47892# vss vss nmos_6p0 w=0.82u l=1u
X14466 vss cap_shunt_n a_19152_38968# vss nmos_6p0 w=0.82u l=0.6u
X14467 a_3620_14964# cap_shunt_p a_3828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X14468 vdd tune_shunt[4] a_2500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X14469 a_2500_19292# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14470 a_24452_36540# cap_shunt_p a_24660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X14471 a_17808_4772# cap_series_gyn a_15700_4834# vss nmos_6p0 w=0.82u l=0.6u
X14472 vdd tune_series_gy[4] a_25572_10260# vdd pmos_6p0 w=1.2u l=0.5u
X14473 a_7952_10744# cap_shunt_p a_5844_10744# vss nmos_6p0 w=0.82u l=0.6u
X14474 vss cap_shunt_n a_11872_34264# vss nmos_6p0 w=0.82u l=0.6u
X14475 a_31648_7908# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X14476 a_3828_13880# cap_shunt_n a_4760_13880# vss nmos_6p0 w=0.82u l=0.6u
X14477 vdd tune_shunt[7] a_13588_20860# vdd pmos_6p0 w=1.2u l=0.5u
X14478 a_14484_8692# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14479 a_5636_10260# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14480 a_21748_37762# cap_shunt_n a_23464_37700# vss nmos_6p0 w=0.82u l=0.6u
X14481 a_2500_16156# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14482 a_24452_33404# cap_shunt_p a_24660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X14483 vss cap_shunt_p a_30800_29560# vss nmos_6p0 w=0.82u l=0.6u
X14484 a_24660_44034# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X14485 vdd tune_shunt[6] a_9108_50652# vdd pmos_6p0 w=1.2u l=0.5u
X14486 vdd a_25100_48983# a_25012_49080# vdd pmos_6p0 w=1.22u l=1u
X14487 vss cap_shunt_n a_11872_31128# vss nmos_6p0 w=0.82u l=0.6u
X14488 vss tune_shunt[4] a_20740_17016# vss nmos_6p0 w=0.51u l=0.6u
X14489 a_14484_5556# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14490 a_16500_49084# cap_shunt_p a_16708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X14491 vdd a_31708_18056# a_31620_18100# vdd pmos_6p0 w=1.22u l=1u
X14492 a_17828_37400# cap_shunt_n a_17620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X14493 a_2708_26786# cap_shunt_p a_2500_27132# vdd pmos_6p0 w=1.2u l=0.5u
X14494 a_11460_41620# cap_shunt_n a_11668_42104# vdd pmos_6p0 w=1.2u l=0.5u
X14495 vss cap_shunt_p a_30800_26424# vss nmos_6p0 w=0.82u l=0.6u
X14496 vss cap_shunt_n a_30016_6040# vss nmos_6p0 w=0.82u l=0.6u
X14497 a_27676_33303# a_27588_33400# vss vss nmos_6p0 w=0.82u l=1u
X14498 a_24660_11106# cap_series_gyp a_24452_11452# vdd pmos_6p0 w=1.2u l=0.5u
X14499 a_23464_14180# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X14500 a_10452_42812# cap_shunt_n a_10660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X14501 vdd tune_shunt[7] a_2500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X14502 vdd tune_shunt[6] a_24452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X14503 a_1692_33736# a_1604_33780# vss vss nmos_6p0 w=0.82u l=1u
X14504 a_11984_28292# cap_shunt_n a_10660_28354# vss nmos_6p0 w=0.82u l=0.6u
X14505 a_17828_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14506 vdd a_6508_39575# a_6420_39672# vdd pmos_6p0 w=1.22u l=1u
X14507 a_7748_42466# cap_shunt_n a_7540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X14508 a_2932_12312# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X14509 vss cap_shunt_p a_10864_12612# vss nmos_6p0 w=0.82u l=0.6u
X14510 a_23464_11044# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X14511 a_36232_12612# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X14512 a_32604_38440# a_32516_38484# vss vss nmos_6p0 w=0.82u l=1u
X14513 a_32612_37762# cap_shunt_p a_32404_38108# vdd pmos_6p0 w=1.2u l=0.5u
X14514 vss cap_shunt_n a_8064_37400# vss nmos_6p0 w=0.82u l=0.6u
X14515 a_10340_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14516 a_1692_30600# a_1604_30644# vss vss nmos_6p0 w=0.82u l=1u
X14517 a_11984_25156# cap_shunt_n a_10660_25218# vss nmos_6p0 w=0.82u l=0.6u
X14518 a_17828_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14519 vdd a_29916_22327# a_29828_22424# vdd pmos_6p0 w=1.22u l=1u
X14520 a_4760_21720# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14521 a_34844_21192# a_34756_21236# vss vss nmos_6p0 w=0.82u l=1u
X14522 vdd a_6508_36439# a_6420_36536# vdd pmos_6p0 w=1.22u l=1u
X14523 vss tune_shunt[3] a_2932_9176# vss nmos_6p0 w=0.51u l=0.6u
X14524 a_3828_34264# cap_shunt_n a_5544_34264# vss nmos_6p0 w=0.82u l=0.6u
X14525 vdd a_32604_3944# a_32516_3988# vdd pmos_6p0 w=1.22u l=1u
X14526 a_30800_37400# cap_shunt_p a_28692_37400# vss nmos_6p0 w=0.82u l=0.6u
X14527 a_6740_32696# cap_shunt_n a_6532_32212# vdd pmos_6p0 w=1.2u l=0.5u
X14528 a_18404_13020# cap_series_gyn a_18612_12674# vdd pmos_6p0 w=1.2u l=0.5u
X14529 a_10340_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14530 a_28692_26424# cap_shunt_p a_28484_25940# vdd pmos_6p0 w=1.2u l=0.5u
X14531 a_29384_3612# cap_series_gyn a_29196_3612# vdd pmos_6p0 w=1.2u l=0.5u
X14532 vdd a_18940_8648# a_18852_8692# vdd pmos_6p0 w=1.22u l=1u
X14533 a_16296_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14534 a_19524_8692# cap_series_gyp a_19732_9176# vdd pmos_6p0 w=1.2u l=0.5u
X14535 a_27496_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14536 a_6776_3204# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14537 a_24452_14588# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14538 vdd a_17820_55688# a_17732_55732# vdd pmos_6p0 w=1.22u l=1u
X14539 a_3828_31128# cap_shunt_n a_5544_31128# vss nmos_6p0 w=0.82u l=0.6u
X14540 vss tune_shunt[7] a_3828_27992# vss nmos_6p0 w=0.51u l=0.6u
X14541 a_13588_36540# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14542 a_3828_27992# cap_shunt_n a_3620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X14543 a_28692_23288# cap_shunt_p a_28484_22804# vdd pmos_6p0 w=1.2u l=0.5u
X14544 a_9540_12674# cap_shunt_p a_9332_13020# vdd pmos_6p0 w=1.2u l=0.5u
X14545 a_12444_21192# a_12356_21236# vss vss nmos_6p0 w=0.82u l=1u
X14546 a_16296_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14547 a_33732_35832# cap_shunt_n a_33524_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14548 a_7540_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14549 a_22436_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14550 a_19524_13396# cap_series_gyn a_19732_13880# vdd pmos_6p0 w=1.2u l=0.5u
X14551 a_14896_20152# cap_shunt_p a_12788_20152# vss nmos_6p0 w=0.82u l=0.6u
X14552 a_25780_21720# cap_shunt_p a_27496_21720# vss nmos_6p0 w=0.82u l=0.6u
X14553 a_29132_54120# a_29044_54164# vss vss nmos_6p0 w=0.82u l=1u
X14554 vss tune_shunt[7] a_3828_24856# vss nmos_6p0 w=0.51u l=0.6u
X14555 a_6420_13020# cap_shunt_p a_6628_12674# vdd pmos_6p0 w=1.2u l=0.5u
X14556 a_13588_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14557 a_10452_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14558 vss tune_shunt[7] a_9428_18946# vss nmos_6p0 w=0.51u l=0.6u
X14559 a_21748_18946# cap_shunt_p a_22680_18884# vss nmos_6p0 w=0.82u l=0.6u
X14560 a_24452_27132# cap_shunt_p a_24660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X14561 a_17620_19668# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14562 vss tune_shunt[6] a_14580_46808# vss nmos_6p0 w=0.51u l=0.6u
X14563 a_29700_39330# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X14564 vss tune_series_gygy[3] a_34536_8316# vss nmos_6p0 w=0.51u l=0.6u
X14565 a_14908_11351# a_14820_11448# vss vss nmos_6p0 w=0.82u l=1u
X14566 a_21540_23996# cap_shunt_p a_21748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X14567 a_21748_15810# cap_series_gyn a_22680_15748# vss nmos_6p0 w=0.82u l=0.6u
X14568 vdd a_34396_19624# a_34308_19668# vdd pmos_6p0 w=1.22u l=1u
X14569 a_25572_25940# cap_shunt_p a_25780_26424# vdd pmos_6p0 w=1.2u l=0.5u
X14570 a_28484_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14571 a_35880_3988# cap_series_gygyp a_35692_3988# vdd pmos_6p0 w=1.2u l=0.5u
X14572 a_23420_50984# a_23332_51028# vss vss nmos_6p0 w=0.82u l=1u
X14573 a_2140_36872# a_2052_36916# vss vss nmos_6p0 w=0.82u l=1u
X14574 vdd a_12892_19191# a_12804_19288# vdd pmos_6p0 w=1.22u l=1u
X14575 vdd a_16028_50984# a_15940_51028# vdd pmos_6p0 w=1.22u l=1u
X14576 a_25780_6040# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X14577 a_11648_15748# cap_shunt_p a_9540_15810# vss nmos_6p0 w=0.82u l=0.6u
X14578 a_36384_41240# cap_shunt_gyp a_36384_40836# vdd pmos_6p0 w=1.215u l=0.5u
X14579 a_10452_36540# cap_shunt_n a_10660_36194# vdd pmos_6p0 w=1.2u l=0.5u
X14580 a_22680_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14581 a_4032_22020# cap_shunt_p a_2708_22082# vss nmos_6p0 w=0.82u l=0.6u
X14582 a_12788_49944# cap_shunt_n a_12580_49460# vdd pmos_6p0 w=1.2u l=0.5u
X14583 a_25572_22804# cap_shunt_p a_25780_23288# vdd pmos_6p0 w=1.2u l=0.5u
X14584 a_28484_22804# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14585 vdd tune_series_gy[3] a_32444_11452# vdd pmos_6p0 w=1.2u l=0.5u
X14586 vdd a_28348_43144# a_28260_43188# vdd pmos_6p0 w=1.22u l=1u
X14587 a_32404_28700# cap_shunt_p a_32612_28354# vdd pmos_6p0 w=1.2u l=0.5u
X14588 a_7748_36194# cap_shunt_n a_7540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X14589 a_17828_27992# cap_shunt_n a_17620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X14590 vss cap_series_gyn a_30800_17016# vss nmos_6p0 w=0.82u l=0.6u
X14591 a_27676_23895# a_27588_23992# vss vss nmos_6p0 w=0.82u l=1u
X14592 a_14692_10744# cap_series_gyn a_14484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X14593 a_2500_50652# cap_shunt_n a_2708_50306# vdd pmos_6p0 w=1.2u l=0.5u
X14594 a_35740_40008# a_35652_40052# vss vss nmos_6p0 w=0.82u l=1u
X14595 a_10452_33404# cap_shunt_n a_10660_33058# vdd pmos_6p0 w=1.2u l=0.5u
X14596 a_22680_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14597 vdd tune_shunt[4] a_2500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X14598 vdd tune_shunt[5] a_25572_40052# vdd pmos_6p0 w=1.2u l=0.5u
X14599 a_17828_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14600 a_36720_48438# cap_shunt_gyp a_36720_47893# vdd pmos_6p0 w=1.215u l=0.5u
X14601 a_20740_45240# cap_shunt_n a_20532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X14602 a_16500_44380# cap_shunt_p a_16708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X14603 a_3640_7908# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14604 a_11592_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14605 vss cap_shunt_p a_22064_46808# vss nmos_6p0 w=0.82u l=0.6u
X14606 a_7748_33058# cap_shunt_n a_7540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X14607 vss tune_series_gy[2] a_11780_4472# vss nmos_6p0 w=0.51u l=0.6u
X14608 vdd tune_shunt[5] a_21540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X14609 a_31808_39268# cap_shunt_p a_29700_39330# vss nmos_6p0 w=0.82u l=0.6u
X14610 a_25236_3612# cap_shunt_p a_25444_3266# vdd pmos_6p0 w=1.2u l=0.5u
X14611 a_20532_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14612 a_10340_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14613 a_34844_11784# a_34756_11828# vss vss nmos_6p0 w=0.82u l=1u
X14614 vdd tune_shunt[6] a_14372_40052# vdd pmos_6p0 w=1.2u l=0.5u
X14615 a_17828_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14616 a_11424_48676# cap_shunt_p a_9316_48738# vss nmos_6p0 w=0.82u l=0.6u
X14617 a_16500_41244# cap_shunt_n a_16708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X14618 vdd a_6508_27031# a_6420_27128# vdd pmos_6p0 w=1.22u l=1u
X14619 a_10452_5180# cap_series_gyp a_10660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X14620 vss cap_shunt_p a_26768_22020# vss nmos_6p0 w=0.82u l=0.6u
X14621 vdd tune_shunt[6] a_21540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X14622 a_20740_18584# cap_shunt_p a_20532_18100# vdd pmos_6p0 w=1.2u l=0.5u
X14623 a_25572_3988# cap_shunt_p a_25780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X14624 a_14468_3266# cap_series_gyn a_14260_3612# vdd pmos_6p0 w=1.2u l=0.5u
X14625 a_28692_17016# cap_series_gyn a_28484_16532# vdd pmos_6p0 w=1.2u l=0.5u
X14626 a_33732_29560# cap_shunt_p a_33524_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14627 vdd tune_series_gy[5] a_20532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X14628 a_7540_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14629 a_16700_49416# a_16612_49460# vss vss nmos_6p0 w=0.82u l=1u
X14630 vdd a_24204_41576# a_24116_41620# vdd pmos_6p0 w=1.22u l=1u
X14631 a_29132_47848# a_29044_47892# vss vss nmos_6p0 w=0.82u l=1u
X14632 a_21748_9538# cap_series_gyp a_21540_9884# vdd pmos_6p0 w=1.2u l=0.5u
X14633 a_25780_32696# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14634 a_9668_19668# cap_shunt_p a_9876_20152# vdd pmos_6p0 w=1.2u l=0.5u
X14635 a_13588_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14636 vss cap_series_gyn a_8184_4772# vss nmos_6p0 w=0.82u l=0.6u
X14637 vss tune_shunt[4] a_33732_32696# vss nmos_6p0 w=0.51u l=0.6u
X14638 a_34308_20860# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14639 a_25996_50984# a_25908_51028# vss vss nmos_6p0 w=0.82u l=1u
X14640 a_25984_20452# cap_shunt_p a_24660_20514# vss nmos_6p0 w=0.82u l=0.6u
X14641 a_28484_40052# cap_shunt_p a_28692_40536# vdd pmos_6p0 w=1.2u l=0.5u
X14642 vss cap_shunt_n a_9072_29860# vss nmos_6p0 w=0.82u l=0.6u
X14643 a_9428_17378# cap_shunt_p a_10360_17316# vss nmos_6p0 w=0.82u l=0.6u
X14644 a_14392_21720# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14645 a_21748_6402# cap_series_gyn a_21540_6748# vdd pmos_6p0 w=1.2u l=0.5u
X14646 a_6760_3988# cap_series_gyp a_6572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X14647 a_25780_12312# cap_series_gyp a_27496_12312# vss nmos_6p0 w=0.82u l=0.6u
X14648 a_20740_35832# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14649 vss tune_shunt[7] a_3828_15448# vss nmos_6p0 w=0.51u l=0.6u
X14650 a_35692_8692# cap_series_gygyn a_35880_8692# vdd pmos_6p0 w=1.2u l=0.5u
X14651 a_35692_36916# cap_series_gygyp a_35880_36916# vdd pmos_6p0 w=1.2u l=0.5u
X14652 vss cap_shunt_p a_7952_9476# vss nmos_6p0 w=0.82u l=0.6u
X14653 a_26712_13880# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X14654 vdd a_34844_53687# a_34756_53784# vdd pmos_6p0 w=1.22u l=1u
X14655 a_28124_30167# a_28036_30264# vss vss nmos_6p0 w=0.82u l=1u
X14656 vss cap_shunt_n a_9072_26724# vss nmos_6p0 w=0.82u l=0.6u
X14657 a_8400_18584# cap_shunt_p a_6292_18584# vss nmos_6p0 w=0.82u l=0.6u
X14658 a_35600_48438# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14659 vdd a_1692_36872# a_1604_36916# vdd pmos_6p0 w=1.22u l=1u
X14660 vss cap_series_gyn a_27104_7608# vss nmos_6p0 w=0.82u l=0.6u
X14661 a_18404_13020# cap_series_gyn a_18612_12674# vdd pmos_6p0 w=1.2u l=0.5u
X14662 vss tune_shunt[7] a_29700_26786# vss nmos_6p0 w=0.51u l=0.6u
X14663 vss cap_shunt_p a_11200_21720# vss nmos_6p0 w=0.82u l=0.6u
X14664 a_35600_50006# cap_shunt_gyp a_35600_49461# vdd pmos_6p0 w=1.215u l=0.5u
X14665 vdd tune_shunt[2] a_1716_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14666 a_6740_15448# cap_shunt_p a_6532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X14667 a_35692_5556# cap_series_gygyn a_35880_5556# vdd pmos_6p0 w=1.2u l=0.5u
X14668 a_21540_14588# cap_series_gyn a_21748_14242# vdd pmos_6p0 w=1.2u l=0.5u
X14669 a_26712_10744# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X14670 vdd a_34844_50551# a_34756_50648# vdd pmos_6p0 w=1.22u l=1u
X14671 a_28124_27031# a_28036_27128# vss vss nmos_6p0 w=0.82u l=1u
X14672 a_25572_16532# cap_series_gyp a_25780_17016# vdd pmos_6p0 w=1.2u l=0.5u
X14673 vss tune_shunt[6] a_11668_45240# vss nmos_6p0 w=0.51u l=0.6u
X14674 a_28484_16532# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14675 vss tune_shunt[7] a_13796_23650# vss nmos_6p0 w=0.51u l=0.6u
X14676 a_35600_46870# cap_shunt_gyp a_35600_46325# vdd pmos_6p0 w=1.215u l=0.5u
X14677 a_24652_5512# a_24564_5556# vss vss nmos_6p0 w=0.82u l=1u
X14678 a_6740_12312# cap_shunt_p a_6532_11828# vdd pmos_6p0 w=1.2u l=0.5u
X14679 a_9540_12674# cap_shunt_p a_9332_13020# vdd pmos_6p0 w=1.2u l=0.5u
X14680 a_3380_49944# cap_shunt_p a_3172_49460# vdd pmos_6p0 w=1.2u l=0.5u
X14681 a_19524_13396# cap_series_gyn a_19732_13880# vdd pmos_6p0 w=1.2u l=0.5u
X14682 a_10452_27132# cap_shunt_n a_10660_26786# vdd pmos_6p0 w=1.2u l=0.5u
X14683 a_2500_44380# cap_shunt_p a_2708_44034# vdd pmos_6p0 w=1.2u l=0.5u
X14684 a_30528_15748# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X14685 a_21748_45602# cap_shunt_p a_21540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X14686 vss tune_shunt[6] a_11668_42104# vss nmos_6p0 w=0.51u l=0.6u
X14687 vss cap_series_gygyn a_36296_13880# vss nmos_6p0 w=0.82u l=0.6u
X14688 vss tune_shunt_gy[5] a_32928_45944# vss nmos_6p0 w=0.51u l=0.6u
X14689 a_20740_38968# cap_shunt_n a_20532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X14690 a_7748_26786# cap_shunt_n a_7540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X14691 vss tune_shunt[7] a_13796_20514# vss nmos_6p0 w=0.51u l=0.6u
X14692 a_21540_17724# cap_shunt_p a_21748_17378# vdd pmos_6p0 w=1.2u l=0.5u
X14693 a_35880_5556# tune_series_gygy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X14694 a_22680_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14695 a_2500_41244# cap_shunt_p a_2708_40898# vdd pmos_6p0 w=1.2u l=0.5u
X14696 a_8848_35832# cap_shunt_n a_6740_35832# vss nmos_6p0 w=0.82u l=0.6u
X14697 vss cap_series_gygyp a_36296_10744# vss nmos_6p0 w=0.82u l=0.6u
X14698 a_20740_35832# cap_shunt_n a_20532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X14699 vss tune_shunt[6] a_9316_50306# vss nmos_6p0 w=0.51u l=0.6u
X14700 vss tune_shunt[7] a_2708_26786# vss nmos_6p0 w=0.51u l=0.6u
X14701 a_21540_23996# cap_shunt_p a_21748_23650# vdd pmos_6p0 w=1.2u l=0.5u
X14702 a_25572_25940# cap_shunt_p a_25780_26424# vdd pmos_6p0 w=1.2u l=0.5u
X14703 a_13460_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14704 a_20532_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14705 a_37632_50648# cap_shunt_gyn a_37652_50244# vss nmos_6p0 w=0.82u l=0.6u
X14706 a_21748_15810# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14707 a_3380_17016# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14708 a_1716_5556# cap_shunt_p a_1924_6040# vdd pmos_6p0 w=1.2u l=0.5u
X14709 a_29720_9884# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X14710 a_3620_47892# cap_shunt_p a_3828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X14711 a_35292_25896# a_35204_25940# vss vss nmos_6p0 w=0.82u l=1u
X14712 a_7768_8316# cap_series_gyn a_7580_8316# vdd pmos_6p0 w=1.2u l=0.5u
X14713 vdd tune_shunt[3] a_5636_8692# vdd pmos_6p0 w=1.2u l=0.5u
X14714 a_5152_48376# cap_shunt_p a_3828_48376# vss nmos_6p0 w=0.82u l=0.6u
X14715 a_11884_47415# a_11796_47512# vss vss nmos_6p0 w=0.82u l=1u
X14716 vdd a_19276_41143# a_19188_41240# vdd pmos_6p0 w=1.22u l=1u
X14717 a_32604_41143# a_32516_41240# vss vss nmos_6p0 w=0.82u l=1u
X14718 a_25572_22804# cap_shunt_p a_25780_23288# vdd pmos_6p0 w=1.2u l=0.5u
X14719 a_13460_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14720 a_25984_14180# cap_series_gyn a_24660_14242# vss nmos_6p0 w=0.82u l=0.6u
X14721 a_25996_44712# a_25908_44756# vss vss nmos_6p0 w=0.82u l=1u
X14722 vdd a_24204_32168# a_24116_32212# vdd pmos_6p0 w=1.22u l=1u
X14723 a_9220_19292# cap_shunt_p a_9428_18946# vdd pmos_6p0 w=1.2u l=0.5u
X14724 a_3620_44756# cap_shunt_p a_3828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X14725 vdd tune_series_gygy[1] a_34308_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14726 vdd a_6956_45847# a_6868_45944# vdd pmos_6p0 w=1.22u l=1u
X14727 a_20740_29560# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14728 a_25780_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14729 a_28692_7608# cap_series_gyp a_29624_7608# vss nmos_6p0 w=0.82u l=0.6u
X14730 a_18044_52552# a_17956_52596# vss vss nmos_6p0 w=0.82u l=1u
X14731 a_9072_45540# cap_shunt_p a_7748_45602# vss nmos_6p0 w=0.82u l=0.6u
X14732 a_10660_44034# cap_shunt_n a_10452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X14733 a_3828_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14734 vss cap_shunt_n a_5152_27992# vss nmos_6p0 w=0.82u l=0.6u
X14735 a_25984_11044# cap_series_gyp a_24660_11106# vss nmos_6p0 w=0.82u l=0.6u
X14736 a_15904_47108# cap_shunt_p a_13796_47170# vss nmos_6p0 w=0.82u l=0.6u
X14737 vss tune_shunt[7] a_9540_14242# vss nmos_6p0 w=0.51u l=0.6u
X14738 a_2588_55688# a_2500_55732# vss vss nmos_6p0 w=0.82u l=1u
X14739 vdd tune_shunt[4] a_13588_50652# vdd pmos_6p0 w=1.2u l=0.5u
X14740 a_32612_36194# cap_shunt_n a_32404_36540# vdd pmos_6p0 w=1.2u l=0.5u
X14741 vss cap_shunt_n a_15904_29860# vss nmos_6p0 w=0.82u l=0.6u
X14742 a_14484_3988# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14743 vdd a_6956_42711# a_6868_42808# vdd pmos_6p0 w=1.22u l=1u
X14744 a_3640_32996# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14745 a_20740_26424# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14746 a_9072_42404# cap_shunt_n a_7748_42466# vss nmos_6p0 w=0.82u l=0.6u
X14747 a_24204_27464# a_24116_27508# vss vss nmos_6p0 w=0.82u l=1u
X14748 a_18492_7080# a_18404_7124# vss vss nmos_6p0 w=0.82u l=1u
X14749 vss tune_series_gy[2] a_10660_6402# vss nmos_6p0 w=0.51u l=0.6u
X14750 a_14692_9176# cap_series_gyn a_16408_9176# vss nmos_6p0 w=0.82u l=0.6u
X14751 vss tune_series_gygy[4] a_31624_19292# vss nmos_6p0 w=0.51u l=0.6u
X14752 a_10660_40898# cap_shunt_n a_10452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X14753 vss cap_shunt_p a_5152_24856# vss nmos_6p0 w=0.82u l=0.6u
X14754 a_21524_4472# cap_series_gyn a_22456_4472# vss nmos_6p0 w=0.82u l=0.6u
X14755 vss tune_shunt[7] a_9540_11106# vss nmos_6p0 w=0.51u l=0.6u
X14756 a_19732_13880# cap_series_gyn a_21448_13880# vss nmos_6p0 w=0.82u l=0.6u
X14757 vdd tune_shunt[7] a_9668_14964# vdd pmos_6p0 w=1.2u l=0.5u
X14758 a_3620_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14759 vss tune_shunt[6] a_17828_43672# vss nmos_6p0 w=0.51u l=0.6u
X14760 a_32612_33058# cap_shunt_n a_32404_33404# vdd pmos_6p0 w=1.2u l=0.5u
X14761 vdd a_1692_27464# a_1604_27508# vdd pmos_6p0 w=1.22u l=1u
X14762 vss cap_shunt_n a_15904_26724# vss nmos_6p0 w=0.82u l=0.6u
X14763 vss tune_series_gy[4] a_29700_17378# vss nmos_6p0 w=0.51u l=0.6u
X14764 a_32040_6340# cap_series_gygyn a_31624_6748# vss nmos_6p0 w=0.82u l=0.6u
X14765 vss cap_shunt_p a_11200_12312# vss nmos_6p0 w=0.82u l=0.6u
X14766 a_32444_14588# cap_series_gyp a_32632_14588# vdd pmos_6p0 w=1.2u l=0.5u
X14767 a_5724_54120# a_5636_54164# vss vss nmos_6p0 w=0.82u l=1u
X14768 a_24204_24328# a_24116_24372# vss vss nmos_6p0 w=0.82u l=1u
X14769 vss cap_series_gyp a_25984_7908# vss nmos_6p0 w=0.82u l=0.6u
X14770 a_17620_47892# cap_shunt_p a_17828_48376# vdd pmos_6p0 w=1.2u l=0.5u
X14771 vdd tune_series_gy[2] a_10452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X14772 a_19732_10744# cap_series_gyn a_21448_10744# vss nmos_6p0 w=0.82u l=0.6u
X14773 vdd tune_shunt[7] a_9668_11828# vdd pmos_6p0 w=1.2u l=0.5u
X14774 a_28124_17623# a_28036_17720# vss vss nmos_6p0 w=0.82u l=1u
X14775 a_21748_39330# cap_shunt_p a_21540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X14776 a_3036_21192# a_2948_21236# vss vss nmos_6p0 w=0.82u l=1u
X14777 a_4492_3944# a_4404_3988# vss vss nmos_6p0 w=0.82u l=1u
X14778 vss tune_shunt[6] a_17828_40536# vss nmos_6p0 w=0.51u l=0.6u
X14779 a_3828_26424# cap_shunt_p a_3620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X14780 vss tune_shunt[6] a_9316_47170# vss nmos_6p0 w=0.51u l=0.6u
X14781 a_14580_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14782 vss tune_shunt[7] a_13796_14242# vss nmos_6p0 w=0.51u l=0.6u
X14783 vss tune_series_gy[3] a_28692_9176# vss nmos_6p0 w=0.51u l=0.6u
X14784 a_28484_7124# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14785 a_14484_8692# cap_series_gyn a_14692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X14786 a_16500_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14787 a_24660_33058# cap_shunt_p a_26376_32996# vss nmos_6p0 w=0.82u l=0.6u
X14788 vdd a_25212_45847# a_25124_45944# vdd pmos_6p0 w=1.22u l=1u
X14789 a_17620_44756# cap_shunt_p a_17828_45240# vdd pmos_6p0 w=1.2u l=0.5u
X14790 vdd a_32156_7080# a_32068_7124# vdd pmos_6p0 w=1.22u l=1u
X14791 a_8848_29560# cap_shunt_n a_6740_29560# vss nmos_6p0 w=0.82u l=0.6u
X14792 a_20740_29560# cap_shunt_n a_20532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X14793 a_3828_23288# cap_shunt_p a_3620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X14794 a_16500_49084# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14795 a_14580_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14796 a_14484_5556# cap_series_gyn a_14692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X14797 a_3828_13880# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X14798 a_17828_43672# cap_shunt_p a_18760_43672# vss nmos_6p0 w=0.82u l=0.6u
X14799 a_18612_7970# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14800 a_8848_26424# cap_shunt_n a_6740_26424# vss nmos_6p0 w=0.82u l=0.6u
X14801 vss cap_shunt_p a_11424_22020# vss nmos_6p0 w=0.82u l=0.6u
X14802 a_6740_15448# cap_shunt_p a_6532_14964# vdd pmos_6p0 w=1.2u l=0.5u
X14803 a_7448_20452# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14804 a_20732_49416# a_20644_49460# vss vss nmos_6p0 w=0.82u l=1u
X14805 a_21540_14588# cap_series_gyn a_21748_14242# vdd pmos_6p0 w=1.2u l=0.5u
X14806 vss tune_shunt[7] a_2708_17378# vss nmos_6p0 w=0.51u l=0.6u
X14807 a_34664_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14808 a_28692_4472# tune_series_gy[0] vss vss nmos_6p0 w=0.51u l=0.6u
X14809 a_25572_16532# cap_series_gyp a_25780_17016# vdd pmos_6p0 w=1.2u l=0.5u
X14810 a_17828_40536# cap_shunt_n a_18760_40536# vss nmos_6p0 w=0.82u l=0.6u
X14811 a_35180_30167# a_35092_30264# vss vss nmos_6p0 w=0.82u l=1u
X14812 a_18612_4834# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X14813 a_17620_14964# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14814 a_6740_12312# cap_shunt_p a_6532_11828# vdd pmos_6p0 w=1.2u l=0.5u
X14815 a_25780_43672# cap_shunt_p a_25572_43188# vdd pmos_6p0 w=1.2u l=0.5u
X14816 a_3620_38484# cap_shunt_n a_3828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X14817 a_35292_16488# a_35204_16532# vss vss nmos_6p0 w=0.82u l=1u
X14818 vdd a_6956_39575# a_6868_39672# vdd pmos_6p0 w=1.22u l=1u
X14819 a_34664_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14820 a_21748_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X14821 vdd a_17596_52552# a_17508_52596# vdd pmos_6p0 w=1.22u l=1u
X14822 a_11984_48376# cap_shunt_p a_9876_48376# vss nmos_6p0 w=0.82u l=0.6u
X14823 a_35180_27031# a_35092_27128# vss vss nmos_6p0 w=0.82u l=1u
X14824 a_21748_9538# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14825 a_33052_55255# a_32964_55352# vss vss nmos_6p0 w=0.82u l=1u
X14826 vdd tune_shunt[6] a_13588_44380# vdd pmos_6p0 w=1.2u l=0.5u
X14827 a_14580_43672# cap_shunt_n a_14372_43188# vdd pmos_6p0 w=1.2u l=0.5u
X14828 a_3620_35348# cap_shunt_n a_3828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X14829 vdd a_6956_36439# a_6868_36536# vdd pmos_6p0 w=1.22u l=1u
X14830 a_12264_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14831 vss cap_series_gygyn a_31032_21720# vss nmos_6p0 w=0.82u l=0.6u
X14832 a_14112_17016# cap_shunt_p a_12788_17016# vss nmos_6p0 w=0.82u l=0.6u
X14833 a_9072_36132# cap_shunt_n a_7748_36194# vss nmos_6p0 w=0.82u l=0.6u
X14834 vss cap_shunt_n a_11984_43972# vss nmos_6p0 w=0.82u l=0.6u
X14835 vss cap_series_gygyn a_35736_9476# vss nmos_6p0 w=0.82u l=0.6u
X14836 a_16700_52119# a_16612_52216# vss vss nmos_6p0 w=0.82u l=1u
X14837 vss cap_shunt_p a_10640_47108# vss nmos_6p0 w=0.82u l=0.6u
X14838 vss cap_series_gyn a_20720_11044# vss nmos_6p0 w=0.82u l=0.6u
X14839 a_34516_18946# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14840 vdd tune_shunt[6] a_13588_41244# vdd pmos_6p0 w=1.2u l=0.5u
X14841 a_32612_26786# cap_shunt_p a_32404_27132# vdd pmos_6p0 w=1.2u l=0.5u
X14842 a_25572_25940# cap_shunt_p a_25780_26424# vdd pmos_6p0 w=1.2u l=0.5u
X14843 a_12264_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14844 a_3640_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14845 a_21428_5556# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14846 vdd a_20620_31735# a_20532_31832# vdd pmos_6p0 w=1.22u l=1u
X14847 a_3828_13880# cap_shunt_n a_3620_13396# vdd pmos_6p0 w=1.2u l=0.5u
X14848 a_20740_17016# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X14849 a_7224_50244# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14850 a_11668_46808# cap_shunt_n a_13384_46808# vss nmos_6p0 w=0.82u l=0.6u
X14851 vss cap_shunt_p a_5152_15448# vss nmos_6p0 w=0.82u l=0.6u
X14852 a_24204_18056# a_24116_18100# vss vss nmos_6p0 w=0.82u l=1u
X14853 vss cap_shunt_n a_11984_40836# vss nmos_6p0 w=0.82u l=0.6u
X14854 vss tune_shunt[6] a_10548_38968# vss nmos_6p0 w=0.51u l=0.6u
X14855 a_12892_21192# a_12804_21236# vss vss nmos_6p0 w=0.82u l=1u
X14856 vss tune_shunt[7] a_17828_34264# vss nmos_6p0 w=0.51u l=0.6u
X14857 a_25572_22804# cap_shunt_p a_25780_23288# vdd pmos_6p0 w=1.2u l=0.5u
X14858 vss cap_shunt_p a_15904_17316# vss nmos_6p0 w=0.82u l=0.6u
X14859 a_29580_54120# a_29492_54164# vss vss nmos_6p0 w=0.82u l=1u
X14860 a_3172_51028# cap_shunt_n a_3380_51512# vdd pmos_6p0 w=1.2u l=0.5u
X14861 a_37280_45302# tune_shunt_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X14862 vss tune_series_gy[3] a_11800_7124# vss nmos_6p0 w=0.51u l=0.6u
X14863 a_24204_14920# a_24116_14964# vss vss nmos_6p0 w=0.82u l=1u
X14864 vss cap_shunt_p a_27888_43672# vss nmos_6p0 w=0.82u l=0.6u
X14865 vdd tune_shunt[7] a_10452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X14866 vss tune_shunt[7] a_9428_18946# vss nmos_6p0 w=0.51u l=0.6u
X14867 a_17620_38484# cap_shunt_n a_17828_38968# vdd pmos_6p0 w=1.2u l=0.5u
X14868 vdd tune_series_gygy[3] a_35692_7124# vdd pmos_6p0 w=1.2u l=0.5u
X14869 a_11256_12612# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14870 a_6516_20514# cap_shunt_p a_8232_20452# vss nmos_6p0 w=0.82u l=0.6u
X14871 a_5612_55255# a_5524_55352# vss vss nmos_6p0 w=0.82u l=1u
X14872 vdd tune_shunt[7] a_13252_36916# vdd pmos_6p0 w=1.2u l=0.5u
X14873 vss tune_shunt[7] a_17828_31128# vss nmos_6p0 w=0.51u l=0.6u
X14874 vss tune_shunt[3] a_2932_12312# vss nmos_6p0 w=0.51u l=0.6u
X14875 vdd a_18940_55255# a_18852_55352# vdd pmos_6p0 w=1.22u l=1u
X14876 a_10660_44034# cap_shunt_n a_10452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X14877 a_30800_7608# cap_series_gyp a_28692_7608# vss nmos_6p0 w=0.82u l=0.6u
X14878 a_22848_38968# cap_shunt_n a_20740_38968# vss nmos_6p0 w=0.82u l=0.6u
X14879 a_7540_34972# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14880 vss cap_shunt_n a_16688_43672# vss nmos_6p0 w=0.82u l=0.6u
X14881 a_24660_23650# cap_shunt_p a_26376_23588# vss nmos_6p0 w=0.82u l=0.6u
X14882 vss cap_shunt_n a_27888_40536# vss nmos_6p0 w=0.82u l=0.6u
X14883 a_32612_36194# cap_shunt_n a_32404_36540# vdd pmos_6p0 w=1.2u l=0.5u
X14884 a_17620_35348# cap_shunt_n a_17828_35832# vdd pmos_6p0 w=1.2u l=0.5u
X14885 a_21748_34626# cap_shunt_p a_21540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X14886 vdd tune_shunt[7] a_10452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X14887 a_28124_9783# a_28036_9880# vss vss nmos_6p0 w=0.82u l=1u
X14888 a_11668_40536# cap_shunt_n a_11460_40052# vdd pmos_6p0 w=1.2u l=0.5u
X14889 vdd a_31260_32168# a_31172_32212# vdd pmos_6p0 w=1.22u l=1u
X14890 a_34536_6748# cap_series_gygyp a_34560_6340# vss nmos_6p0 w=0.82u l=0.6u
X14891 vdd a_18940_52119# a_18852_52216# vdd pmos_6p0 w=1.22u l=1u
X14892 a_10660_40898# cap_shunt_n a_10452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X14893 a_32404_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14894 a_18612_4834# cap_series_gyp a_18404_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14895 a_10548_38968# cap_shunt_n a_11480_38968# vss nmos_6p0 w=0.82u l=0.6u
X14896 a_7540_31836# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14897 a_8860_19191# a_8772_19288# vss vss nmos_6p0 w=0.82u l=1u
X14898 vss cap_shunt_n a_16688_40536# vss nmos_6p0 w=0.82u l=0.6u
X14899 vdd a_5612_30167# a_5524_30264# vdd pmos_6p0 w=1.22u l=1u
X14900 a_31416_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14901 a_17828_34264# cap_shunt_n a_18760_34264# vss nmos_6p0 w=0.82u l=0.6u
X14902 a_32612_33058# cap_shunt_n a_32404_33404# vdd pmos_6p0 w=1.2u l=0.5u
X14903 vdd a_6060_53687# a_5972_53784# vdd pmos_6p0 w=1.22u l=1u
X14904 vdd a_16476_50984# a_16388_51028# vdd pmos_6p0 w=1.22u l=1u
X14905 a_7616_48676# cap_shunt_p a_6292_48738# vss nmos_6p0 w=0.82u l=0.6u
X14906 a_21748_31490# cap_shunt_n a_21540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X14907 vss cap_series_gygyn a_36296_9176# vss nmos_6p0 w=0.82u l=0.6u
X14908 a_2500_50652# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14909 a_19276_47415# a_19188_47512# vss vss nmos_6p0 w=0.82u l=1u
X14910 vss tune_series_gy[3] a_25780_6040# vss nmos_6p0 w=0.51u l=0.6u
X14911 vdd tune_series_gygy[1] a_34308_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14912 a_8860_16055# a_8772_16152# vss vss nmos_6p0 w=0.82u l=1u
X14913 a_28484_18100# cap_series_gyp a_28692_18584# vdd pmos_6p0 w=1.2u l=0.5u
X14914 vdd a_28796_43144# a_28708_43188# vdd pmos_6p0 w=1.22u l=1u
X14915 a_31260_27464# a_31172_27508# vss vss nmos_6p0 w=0.82u l=1u
X14916 a_34516_17378# tune_series_gygy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14917 a_22076_52552# a_21988_52596# vss vss nmos_6p0 w=0.82u l=1u
X14918 a_17828_31128# cap_shunt_n a_18760_31128# vss nmos_6p0 w=0.82u l=0.6u
X14919 a_24452_13020# cap_series_gyn a_24660_12674# vdd pmos_6p0 w=1.2u l=0.5u
X14920 a_33052_48983# a_32964_49080# vss vss nmos_6p0 w=0.82u l=1u
X14921 vdd a_6508_5079# a_6420_5176# vdd pmos_6p0 w=1.22u l=1u
X14922 vdd tune_series_gy[5] a_19524_8692# vdd pmos_6p0 w=1.2u l=0.5u
X14923 vdd a_3036_53687# a_2948_53784# vdd pmos_6p0 w=1.22u l=1u
X14924 a_27900_45847# a_27812_45944# vss vss nmos_6p0 w=0.82u l=1u
X14925 a_31436_6748# cap_series_gygyn a_31624_6748# vdd pmos_6p0 w=1.2u l=0.5u
X14926 a_3620_29076# cap_shunt_n a_3828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X14927 a_29492_39676# cap_shunt_p a_29700_39330# vdd pmos_6p0 w=1.2u l=0.5u
X14928 vdd a_37868_8215# a_37780_8312# vdd pmos_6p0 w=1.22u l=1u
X14929 a_31260_24328# a_31172_24372# vss vss nmos_6p0 w=0.82u l=1u
X14930 vss cap_series_gyn a_30584_3204# vss nmos_6p0 w=0.82u l=0.6u
X14931 a_6532_13396# cap_shunt_p a_6740_13880# vdd pmos_6p0 w=1.2u l=0.5u
X14932 a_11460_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14933 a_6740_48376# cap_shunt_p a_6532_47892# vdd pmos_6p0 w=1.2u l=0.5u
X14934 a_18760_45240# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14935 a_1716_6748# cap_shunt_n a_1924_6402# vdd pmos_6p0 w=1.2u l=0.5u
X14936 a_35692_13396# cap_series_gygyn a_35880_13396# vdd pmos_6p0 w=1.2u l=0.5u
X14937 a_24452_38108# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14938 vdd tune_shunt[7] a_17620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X14939 vdd a_6956_27031# a_6868_27128# vdd pmos_6p0 w=1.22u l=1u
X14940 vdd a_20620_25463# a_20532_25560# vdd pmos_6p0 w=1.22u l=1u
X14941 vss cap_series_gyn a_17808_9476# vss nmos_6p0 w=0.82u l=0.6u
X14942 a_21748_9538# cap_series_gyp a_21540_9884# vdd pmos_6p0 w=1.2u l=0.5u
X14943 vss tune_series_gy[4] a_24660_18946# vss nmos_6p0 w=0.51u l=0.6u
X14944 a_6740_45240# cap_shunt_p a_6532_44756# vdd pmos_6p0 w=1.2u l=0.5u
X14945 a_18760_42104# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X14946 vss cap_series_gyp a_23856_4772# vss nmos_6p0 w=0.82u l=0.6u
X14947 vss cap_shunt_n a_11984_34564# vss nmos_6p0 w=0.82u l=0.6u
X14948 vdd tune_shunt[7] a_10340_32212# vdd pmos_6p0 w=1.2u l=0.5u
X14949 vdd a_2588_14920# a_2500_14964# vdd pmos_6p0 w=1.22u l=1u
X14950 a_20532_25940# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14951 a_25572_16532# cap_series_gyp a_25780_17016# vdd pmos_6p0 w=1.2u l=0.5u
X14952 vdd a_24652_41576# a_24564_41620# vdd pmos_6p0 w=1.22u l=1u
X14953 vdd a_20620_22327# a_20532_22424# vdd pmos_6p0 w=1.22u l=1u
X14954 vdd a_37084_40008# a_36996_40052# vdd pmos_6p0 w=1.22u l=1u
X14955 a_21748_6402# cap_series_gyn a_21540_6748# vdd pmos_6p0 w=1.2u l=0.5u
X14956 a_29580_47848# a_29492_47892# vss vss nmos_6p0 w=0.82u l=1u
X14957 a_34144_43972# tune_shunt_gy[6] vss vss nmos_6p0 w=0.51u l=0.6u
X14958 vdd a_32828_41576# a_32740_41620# vdd pmos_6p0 w=1.22u l=1u
X14959 a_7672_48376# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14960 a_25780_43672# cap_shunt_p a_25572_43188# vdd pmos_6p0 w=1.2u l=0.5u
X14961 a_35628_38007# a_35540_38104# vss vss nmos_6p0 w=0.82u l=1u
X14962 vss cap_shunt_n a_11984_31428# vss nmos_6p0 w=0.82u l=0.6u
X14963 a_5612_48983# a_5524_49080# vss vss nmos_6p0 w=0.82u l=1u
X14964 vss tune_shunt[7] a_12788_12312# vss nmos_6p0 w=0.51u l=0.6u
X14965 a_20532_22804# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14966 a_18404_13020# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14967 a_29720_13020# cap_series_gyn a_29532_13020# vdd pmos_6p0 w=1.2u l=0.5u
X14968 vss tune_shunt[4] a_17828_48376# vss nmos_6p0 w=0.51u l=0.6u
X14969 vdd a_1692_47415# a_1604_47512# vdd pmos_6p0 w=1.22u l=1u
X14970 vss cap_shunt_p a_22848_21720# vss nmos_6p0 w=0.82u l=0.6u
X14971 a_14580_43672# cap_shunt_n a_14372_43188# vdd pmos_6p0 w=1.2u l=0.5u
X14972 vss cap_shunt_p a_27888_34264# vss nmos_6p0 w=0.82u l=0.6u
X14973 vdd a_20172_17623# a_20084_17720# vdd pmos_6p0 w=1.22u l=1u
X14974 a_17620_29076# cap_shunt_n a_17828_29560# vdd pmos_6p0 w=1.2u l=0.5u
X14975 vdd tune_shunt[7] a_10452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X14976 a_12788_20152# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X14977 a_6740_27992# cap_shunt_n a_7672_27992# vss nmos_6p0 w=0.82u l=0.6u
X14978 vdd tune_shunt[7] a_13252_27508# vdd pmos_6p0 w=1.2u l=0.5u
X14979 a_1924_4834# cap_shunt_p a_1716_5180# vdd pmos_6p0 w=1.2u l=0.5u
X14980 a_28572_30167# a_28484_30264# vss vss nmos_6p0 w=0.82u l=1u
X14981 a_30136_12612# cap_series_gyn a_29720_13020# vss nmos_6p0 w=0.82u l=0.6u
X14982 a_7540_25564# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14983 a_15356_47848# a_15268_47892# vss vss nmos_6p0 w=0.82u l=1u
X14984 a_29624_35832# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X14985 vss cap_shunt_p a_27888_31128# vss nmos_6p0 w=0.82u l=0.6u
X14986 vdd tune_series_gy[4] a_25572_19668# vdd pmos_6p0 w=1.2u l=0.5u
X14987 vdd a_18044_49416# a_17956_49460# vdd pmos_6p0 w=1.22u l=1u
X14988 vdd a_19724_34871# a_19636_34968# vdd pmos_6p0 w=1.22u l=1u
X14989 a_32612_26786# cap_shunt_p a_32404_27132# vdd pmos_6p0 w=1.2u l=0.5u
X14990 a_2500_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X14991 a_21748_25218# cap_shunt_n a_21540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X14992 a_6740_24856# cap_shunt_p a_7672_24856# vss nmos_6p0 w=0.82u l=0.6u
X14993 a_28572_27031# a_28484_27128# vss vss nmos_6p0 w=0.82u l=1u
X14994 a_29700_23650# cap_shunt_p a_29492_23996# vdd pmos_6p0 w=1.2u l=0.5u
X14995 a_19732_9176# cap_series_gyp a_20664_9176# vss nmos_6p0 w=0.82u l=0.6u
X14996 a_26444_55255# a_26356_55352# vss vss nmos_6p0 w=0.82u l=1u
X14997 a_27104_32696# cap_shunt_p a_25780_32696# vss nmos_6p0 w=0.82u l=0.6u
X14998 vss tune_shunt[5] a_20740_45240# vss nmos_6p0 w=0.51u l=0.6u
X14999 vdd a_9644_40008# a_9556_40052# vdd pmos_6p0 w=1.22u l=1u
X15000 vdd a_36076_33303# a_35988_33400# vdd pmos_6p0 w=1.22u l=1u
X15001 vss cap_shunt_p a_7952_10744# vss nmos_6p0 w=0.82u l=0.6u
X15002 a_12788_12312# cap_shunt_p a_13720_12312# vss nmos_6p0 w=0.82u l=0.6u
X15003 vdd a_6060_44279# a_5972_44376# vdd pmos_6p0 w=1.22u l=1u
X15004 a_2500_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15005 a_21748_22082# cap_shunt_p a_21540_22428# vdd pmos_6p0 w=1.2u l=0.5u
X15006 a_3172_51028# cap_shunt_n a_3380_51512# vdd pmos_6p0 w=1.2u l=0.5u
X15007 vdd a_37868_38007# a_37780_38104# vdd pmos_6p0 w=1.22u l=1u
X15008 vss tune_shunt[6] a_20740_42104# vss nmos_6p0 w=0.51u l=0.6u
X15009 a_35344_9476# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X15010 a_31260_18056# a_31172_18100# vss vss nmos_6p0 w=0.82u l=1u
X15011 vss cap_shunt_n a_3248_7608# vss nmos_6p0 w=0.82u l=0.6u
X15012 a_9668_13396# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15013 a_18612_4472# cap_series_gyp a_18404_3988# vdd pmos_6p0 w=1.2u l=0.5u
X15014 a_33500_8648# a_33412_8692# vss vss nmos_6p0 w=0.82u l=1u
X15015 a_37868_19191# a_37780_19288# vss vss nmos_6p0 w=0.82u l=1u
X15016 vss cap_shunt_p a_7616_18884# vss nmos_6p0 w=0.82u l=0.6u
X15017 a_20732_52119# a_20644_52216# vss vss nmos_6p0 w=0.82u l=1u
X15018 vss cap_series_gyn a_12656_3204# vss nmos_6p0 w=0.82u l=0.6u
X15019 a_16708_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15020 a_20532_46324# cap_shunt_p a_20740_46808# vdd pmos_6p0 w=1.2u l=0.5u
X15021 a_23072_39268# cap_shunt_p a_21748_39330# vss nmos_6p0 w=0.82u l=0.6u
X15022 vss tune_shunt[5] a_28692_38968# vss nmos_6p0 w=0.51u l=0.6u
X15023 a_19544_27992# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15024 vss tune_shunt[7] a_9540_9538# vss nmos_6p0 w=0.51u l=0.6u
X15025 a_21748_34626# cap_shunt_p a_21540_34972# vdd pmos_6p0 w=1.2u l=0.5u
X15026 a_31260_14920# a_31172_14964# vss vss nmos_6p0 w=0.82u l=1u
X15027 a_6740_38968# cap_shunt_n a_6532_38484# vdd pmos_6p0 w=1.2u l=0.5u
X15028 a_11592_51512# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15029 vss cap_shunt_n a_11984_28292# vss nmos_6p0 w=0.82u l=0.6u
X15030 a_28484_8692# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15031 a_5844_9176# cap_shunt_p a_5636_8692# vdd pmos_6p0 w=1.2u l=0.5u
X15032 a_9644_32168# a_9556_32212# vss vss nmos_6p0 w=0.82u l=1u
X15033 a_6760_5556# cap_series_gyp a_7568_6040# vss nmos_6p0 w=0.82u l=0.6u
X15034 a_37868_16055# a_37780_16152# vss vss nmos_6p0 w=0.82u l=1u
X15035 vss cap_shunt_p a_7616_15748# vss nmos_6p0 w=0.82u l=0.6u
X15036 vss cap_shunt_p a_30016_27992# vss nmos_6p0 w=0.82u l=0.6u
X15037 vdd tune_shunt[7] a_17620_27508# vdd pmos_6p0 w=1.2u l=0.5u
X15038 a_18404_9884# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15039 a_19544_24856# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15040 vdd a_20620_16055# a_20532_16152# vdd pmos_6p0 w=1.22u l=1u
X15041 a_21748_31490# cap_shunt_n a_21540_31836# vdd pmos_6p0 w=1.2u l=0.5u
X15042 a_29492_23996# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15043 vss tune_shunt[5] a_6292_50306# vss nmos_6p0 w=0.51u l=0.6u
X15044 a_6740_35832# cap_shunt_n a_6532_35348# vdd pmos_6p0 w=1.2u l=0.5u
X15045 vss cap_shunt_n a_11984_25156# vss nmos_6p0 w=0.82u l=0.6u
X15046 a_13796_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15047 a_28484_5556# tune_shunt[0] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15048 vdd a_17596_8648# a_17508_8692# vdd pmos_6p0 w=1.22u l=1u
X15049 a_28484_18100# cap_series_gyp a_28692_18584# vdd pmos_6p0 w=1.2u l=0.5u
X15050 vss cap_shunt_p a_30016_24856# vss nmos_6p0 w=0.82u l=0.6u
X15051 a_18404_6748# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15052 a_20532_16532# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15053 a_31708_35304# a_31620_35348# vss vss nmos_6p0 w=0.82u l=1u
X15054 vdd a_24652_32168# a_24564_32212# vdd pmos_6p0 w=1.22u l=1u
X15055 a_6292_18946# cap_shunt_p a_6084_19292# vdd pmos_6p0 w=1.2u l=0.5u
X15056 vdd tune_shunt[7] a_9332_14588# vdd pmos_6p0 w=1.2u l=0.5u
X15057 a_13588_17724# cap_shunt_p a_13796_17378# vdd pmos_6p0 w=1.2u l=0.5u
X15058 a_18492_52552# a_18404_52596# vss vss nmos_6p0 w=0.82u l=1u
X15059 a_13796_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15060 a_5612_39575# a_5524_39672# vss vss nmos_6p0 w=0.82u l=1u
X15061 a_29492_39676# cap_shunt_p a_29700_39330# vdd pmos_6p0 w=1.2u l=0.5u
X15062 vdd a_17596_5512# a_17508_5556# vdd pmos_6p0 w=1.22u l=1u
X15063 a_6532_13396# cap_shunt_p a_6740_13880# vdd pmos_6p0 w=1.2u l=0.5u
X15064 vdd a_34844_52552# a_34756_52596# vdd pmos_6p0 w=1.22u l=1u
X15065 vdd tune_shunt[7] a_9668_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15066 a_2708_29922# cap_shunt_n a_4424_29860# vss nmos_6p0 w=0.82u l=0.6u
X15067 vdd a_1692_38007# a_1604_38104# vdd pmos_6p0 w=1.22u l=1u
X15068 vdd tune_series_gy[4] a_24452_8316# vdd pmos_6p0 w=1.2u l=0.5u
X15069 a_6292_15810# cap_shunt_p a_6084_16156# vdd pmos_6p0 w=1.2u l=0.5u
X15070 a_14784_34264# cap_shunt_n a_13460_34264# vss nmos_6p0 w=0.82u l=0.6u
X15071 a_3620_33780# cap_shunt_n a_3828_34264# vdd pmos_6p0 w=1.2u l=0.5u
X15072 a_10528_51812# cap_shunt_n a_9204_51874# vss nmos_6p0 w=0.82u l=0.6u
X15073 vss cap_shunt_n a_18032_37700# vss nmos_6p0 w=0.82u l=0.6u
X15074 a_29624_29560# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15075 vdd a_19724_28599# a_19636_28696# vdd pmos_6p0 w=1.22u l=1u
X15076 a_2708_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15077 a_4704_17016# cap_shunt_p a_3380_17016# vss nmos_6p0 w=0.82u l=0.6u
X15078 a_24652_27464# a_24564_27508# vss vss nmos_6p0 w=0.82u l=1u
X15079 a_21748_18946# cap_shunt_p a_21540_19292# vdd pmos_6p0 w=1.2u l=0.5u
X15080 a_17620_47892# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15081 a_26376_37700# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15082 vdd tune_series_gy[2] a_10452_6748# vdd pmos_6p0 w=1.2u l=0.5u
X15083 vdd a_33948_24328# a_33860_24372# vdd pmos_6p0 w=1.22u l=1u
X15084 vdd a_11772_52119# a_11684_52216# vdd pmos_6p0 w=1.22u l=1u
X15085 vss cap_shunt_gyp a_36652_50244# vss nmos_6p0 w=0.82u l=0.6u
X15086 a_26444_48983# a_26356_49080# vss vss nmos_6p0 w=0.82u l=1u
X15087 a_2708_26786# cap_shunt_p a_4424_26724# vss nmos_6p0 w=0.82u l=0.6u
X15088 vss tune_shunt[4] a_21748_45602# vss nmos_6p0 w=0.51u l=0.6u
X15089 a_21748_44034# cap_shunt_n a_22680_43972# vss nmos_6p0 w=0.82u l=0.6u
X15090 a_7748_39330# cap_shunt_n a_9464_39268# vss nmos_6p0 w=0.82u l=0.6u
X15091 vdd tune_shunt[7] a_10340_32212# vdd pmos_6p0 w=1.2u l=0.5u
X15092 a_1692_19191# a_1604_19288# vss vss nmos_6p0 w=0.82u l=1u
X15093 a_14784_31128# cap_shunt_n a_13460_31128# vss nmos_6p0 w=0.82u l=0.6u
X15094 a_3620_30644# cap_shunt_n a_3828_31128# vdd pmos_6p0 w=1.2u l=0.5u
X15095 vss cap_series_gyp a_19936_4472# vss nmos_6p0 w=0.82u l=0.6u
X15096 a_29624_26424# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15097 a_19524_11828# cap_series_gyn a_19732_12312# vdd pmos_6p0 w=1.2u l=0.5u
X15098 vss cap_shunt_p a_15904_46808# vss nmos_6p0 w=0.82u l=0.6u
X15099 vdd tune_shunt[7] a_2500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X15100 a_24652_24328# a_24564_24372# vss vss nmos_6p0 w=0.82u l=1u
X15101 a_21748_15810# cap_series_gyn a_21540_16156# vdd pmos_6p0 w=1.2u l=0.5u
X15102 a_28236_50984# a_28148_51028# vss vss nmos_6p0 w=0.82u l=1u
X15103 a_17620_44756# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15104 a_31708_7080# a_31620_7124# vss vss nmos_6p0 w=0.82u l=1u
X15105 a_6740_15448# cap_shunt_p a_7672_15448# vss nmos_6p0 w=0.82u l=0.6u
X15106 vdd a_12444_52552# a_12356_52596# vdd pmos_6p0 w=1.22u l=1u
X15107 a_29700_14242# cap_series_gyp a_29492_14588# vdd pmos_6p0 w=1.2u l=0.5u
X15108 a_28572_17623# a_28484_17720# vss vss nmos_6p0 w=0.82u l=1u
X15109 vdd a_33948_21192# a_33860_21236# vdd pmos_6p0 w=1.22u l=1u
X15110 a_27104_23288# cap_shunt_p a_25780_23288# vss nmos_6p0 w=0.82u l=0.6u
X15111 a_21748_40898# cap_shunt_p a_22680_40836# vss nmos_6p0 w=0.82u l=0.6u
X15112 a_18724_6040# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X15113 a_31436_20860# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15114 a_1692_16055# a_1604_16152# vss vss nmos_6p0 w=0.82u l=1u
X15115 vdd tune_shunt[7] a_16500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X15116 a_9332_9884# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15117 a_29720_13020# cap_series_gyn a_29532_13020# vdd pmos_6p0 w=1.2u l=0.5u
X15118 vdd tune_shunt[7] a_24452_20860# vdd pmos_6p0 w=1.2u l=0.5u
X15119 a_10548_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15120 a_11612_7124# cap_series_gyp a_11800_7124# vdd pmos_6p0 w=1.2u l=0.5u
X15121 vdd a_25660_45847# a_25572_45944# vdd pmos_6p0 w=1.22u l=1u
X15122 a_28484_8692# cap_series_gyn a_28692_9176# vdd pmos_6p0 w=1.2u l=0.5u
X15123 a_1692_52552# a_1604_52596# vss vss nmos_6p0 w=0.82u l=1u
X15124 a_21292_55688# a_21204_55732# vss vss nmos_6p0 w=0.82u l=1u
X15125 a_10548_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15126 vdd a_7068_54120# a_6980_54164# vdd pmos_6p0 w=1.22u l=1u
X15127 a_28484_5556# cap_shunt_n a_28692_6040# vdd pmos_6p0 w=1.2u l=0.5u
X15128 a_17828_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15129 a_35168_44376# cap_shunt_gyn a_34980_44376# vdd pmos_6p0 w=1.215u l=0.5u
X15130 a_34536_8316# cap_series_gygyp a_34348_8316# vdd pmos_6p0 w=1.2u l=0.5u
X15131 a_19544_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15132 vdd a_29916_41143# a_29828_41240# vdd pmos_6p0 w=1.22u l=1u
X15133 a_21748_25218# cap_shunt_n a_21540_25564# vdd pmos_6p0 w=1.2u l=0.5u
X15134 a_35880_22804# cap_series_gygyp a_36688_23288# vss nmos_6p0 w=0.82u l=0.6u
X15135 a_17828_43672# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15136 a_29700_23650# cap_shunt_p a_29492_23996# vdd pmos_6p0 w=1.2u l=0.5u
X15137 vdd a_6508_55255# a_6420_55352# vdd pmos_6p0 w=1.22u l=1u
X15138 a_37444_45944# cap_shunt_gyn a_37632_45944# vdd pmos_6p0 w=1.215u l=0.5u
X15139 a_6740_29560# cap_shunt_n a_6532_29076# vdd pmos_6p0 w=1.2u l=0.5u
X15140 vss cap_shunt_p a_10752_17316# vss nmos_6p0 w=0.82u l=0.6u
X15141 a_12768_32996# cap_shunt_n a_10660_33058# vss nmos_6p0 w=0.82u l=0.6u
X15142 a_9644_22760# a_9556_22804# vss vss nmos_6p0 w=0.82u l=1u
X15143 vss cap_series_gyp a_30016_18584# vss nmos_6p0 w=0.82u l=0.6u
X15144 a_35264_45540# cap_shunt_gyp a_35264_45944# vdd pmos_6p0 w=1.215u l=0.5u
X15145 a_29492_14588# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15146 a_19544_15448# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15147 vdd a_22524_54120# a_22436_54164# vdd pmos_6p0 w=1.22u l=1u
X15148 vss cap_shunt_n a_11312_51812# vss nmos_6p0 w=0.82u l=0.6u
X15149 a_31708_29032# a_31620_29076# vss vss nmos_6p0 w=0.82u l=1u
X15150 a_21748_22082# cap_shunt_p a_21540_22428# vdd pmos_6p0 w=1.2u l=0.5u
X15151 a_3380_51512# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X15152 a_17828_40536# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15153 vss cap_series_gygyn a_32824_22020# vss nmos_6p0 w=0.82u l=0.6u
X15154 a_37444_42808# cap_shunt_gyn a_37632_42808# vdd pmos_6p0 w=1.215u l=0.5u
X15155 a_29532_9884# cap_series_gyn a_29720_9884# vdd pmos_6p0 w=1.2u l=0.5u
X15156 vdd tune_shunt[7] a_12580_13396# vdd pmos_6p0 w=1.2u l=0.5u
X15157 a_13796_14242# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15158 a_1924_4834# cap_shunt_p a_1716_5180# vdd pmos_6p0 w=1.2u l=0.5u
X15159 a_9668_47892# cap_shunt_p a_9876_48376# vdd pmos_6p0 w=1.2u l=0.5u
X15160 a_10548_37400# cap_shunt_n a_10340_36916# vdd pmos_6p0 w=1.2u l=0.5u
X15161 vss cap_series_gyn a_30016_15448# vss nmos_6p0 w=0.82u l=0.6u
X15162 a_9876_21720# cap_shunt_p a_11592_21720# vss nmos_6p0 w=0.82u l=0.6u
X15163 a_35264_42404# cap_shunt_gyn a_35264_42808# vdd pmos_6p0 w=1.215u l=0.5u
X15164 a_3828_46808# cap_shunt_p a_3620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X15165 a_31708_25896# a_31620_25940# vss vss nmos_6p0 w=0.82u l=1u
X15166 a_19836_55255# a_19748_55352# vss vss nmos_6p0 w=0.82u l=1u
X15167 vdd a_22524_50984# a_22436_51028# vdd pmos_6p0 w=1.22u l=1u
X15168 a_6508_33303# a_6420_33400# vss vss nmos_6p0 w=0.82u l=1u
X15169 a_21428_5556# cap_series_gyp a_21636_6040# vdd pmos_6p0 w=1.2u l=0.5u
X15170 a_24452_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15171 vss tune_shunt[5] a_3828_20152# vss nmos_6p0 w=0.51u l=0.6u
X15172 vdd a_22076_49416# a_21988_49460# vdd pmos_6p0 w=1.22u l=1u
X15173 vss tune_shunt[6] a_3828_43672# vss nmos_6p0 w=0.51u l=0.6u
X15174 vss tune_shunt[6] a_21748_39330# vss nmos_6p0 w=0.51u l=0.6u
X15175 vss cap_shunt_n a_5936_37400# vss nmos_6p0 w=0.82u l=0.6u
X15176 a_14908_9783# a_14820_9880# vss vss nmos_6p0 w=0.82u l=1u
X15177 vss cap_shunt_p a_19152_48376# vss nmos_6p0 w=0.82u l=0.6u
X15178 a_22456_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15179 a_3620_24372# cap_shunt_p a_3828_24856# vdd pmos_6p0 w=1.2u l=0.5u
X15180 a_21540_5180# cap_series_gyp a_21748_4834# vdd pmos_6p0 w=1.2u l=0.5u
X15181 a_30920_15748# cap_series_gyn a_29720_16156# vss nmos_6p0 w=0.82u l=0.6u
X15182 a_2708_17378# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15183 vdd a_8860_49416# a_8772_49460# vdd pmos_6p0 w=1.22u l=1u
X15184 a_32404_34972# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15185 a_2140_8648# a_2052_8692# vss vss nmos_6p0 w=0.82u l=1u
X15186 vdd a_32156_10216# a_32068_10260# vdd pmos_6p0 w=1.22u l=1u
X15187 a_24652_18056# a_24564_18100# vss vss nmos_6p0 w=0.82u l=1u
X15188 vdd a_19724_19191# a_19636_19288# vdd pmos_6p0 w=1.22u l=1u
X15189 vss cap_shunt_p a_25984_20452# vss nmos_6p0 w=0.82u l=0.6u
X15190 a_28236_44712# a_28148_44756# vss vss nmos_6p0 w=0.82u l=1u
X15191 a_17620_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15192 a_31260_3944# a_31172_3988# vss vss nmos_6p0 w=0.82u l=1u
X15193 a_21056_13880# cap_series_gyn a_19732_13880# vss nmos_6p0 w=0.82u l=0.6u
X15194 a_9876_49944# cap_shunt_p a_10808_49944# vss nmos_6p0 w=0.82u l=0.6u
X15195 vss cap_shunt_gyp a_35308_43672# vss nmos_6p0 w=0.82u l=0.6u
X15196 vss tune_shunt[6] a_3828_40536# vss nmos_6p0 w=0.51u l=0.6u
X15197 a_2708_17378# cap_shunt_p a_4424_17316# vss nmos_6p0 w=0.82u l=0.6u
X15198 a_17828_43672# cap_shunt_p a_17620_43188# vdd pmos_6p0 w=1.2u l=0.5u
X15199 a_21748_34626# cap_shunt_p a_22680_34564# vss nmos_6p0 w=0.82u l=0.6u
X15200 a_19936_9476# cap_series_gyp a_18612_9538# vss nmos_6p0 w=0.82u l=0.6u
X15201 vdd tune_series_gy[4] a_28484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15202 a_15356_53687# a_15268_53784# vss vss nmos_6p0 w=0.82u l=1u
X15203 a_28484_18100# cap_series_gyp a_28692_18584# vdd pmos_6p0 w=1.2u l=0.5u
X15204 vdd a_30364_19191# a_30276_19288# vdd pmos_6p0 w=1.22u l=1u
X15205 vdd a_21516_47415# a_21428_47512# vdd pmos_6p0 w=1.22u l=1u
X15206 vdd a_34396_38440# a_34308_38484# vdd pmos_6p0 w=1.22u l=1u
X15207 a_29624_17016# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X15208 a_3620_21236# cap_shunt_p a_3828_21720# vdd pmos_6p0 w=1.2u l=0.5u
X15209 a_32404_31836# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15210 a_5636_8692# cap_shunt_p a_5844_9176# vdd pmos_6p0 w=1.2u l=0.5u
X15211 a_24652_14920# a_24564_14964# vss vss nmos_6p0 w=0.82u l=1u
X15212 a_17620_35348# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15213 vss cap_shunt_n a_12656_32696# vss nmos_6p0 w=0.82u l=0.6u
X15214 a_21056_10744# cap_series_gyn a_19732_10744# vss nmos_6p0 w=0.82u l=0.6u
X15215 a_6292_48738# cap_shunt_p a_6084_49084# vdd pmos_6p0 w=1.2u l=0.5u
X15216 a_13460_37400# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15217 vss tune_shunt[3] a_2932_12312# vss nmos_6p0 w=0.51u l=0.6u
X15218 a_21748_31490# cap_shunt_n a_22680_31428# vss nmos_6p0 w=0.82u l=0.6u
X15219 a_29492_39676# cap_shunt_p a_29700_39330# vdd pmos_6p0 w=1.2u l=0.5u
X15220 a_6740_13880# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15221 a_3828_20152# cap_shunt_p a_4760_20152# vss nmos_6p0 w=0.82u l=0.6u
X15222 a_25572_41620# cap_shunt_n a_25780_42104# vdd pmos_6p0 w=1.2u l=0.5u
X15223 a_32824_7908# cap_series_gygyn a_31624_8316# vss nmos_6p0 w=0.82u l=0.6u
X15224 a_6532_13396# cap_shunt_p a_6740_13880# vdd pmos_6p0 w=1.2u l=0.5u
X15225 vdd tune_shunt[6] a_7540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X15226 vdd tune_series_gy[5] a_24452_11452# vdd pmos_6p0 w=1.2u l=0.5u
X15227 vss tune_shunt[7] a_9876_18584# vss nmos_6p0 w=0.51u l=0.6u
X15228 a_17828_46808# cap_shunt_n a_17620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X15229 a_21540_38108# cap_shunt_n a_21748_37762# vdd pmos_6p0 w=1.2u l=0.5u
X15230 vdd a_37868_55688# a_37780_55732# vdd pmos_6p0 w=1.22u l=1u
X15231 a_22680_45540# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15232 a_16924_35304# a_16836_35348# vss vss nmos_6p0 w=0.82u l=1u
X15233 vss tune_series_gygy[4] a_35880_13396# vss nmos_6p0 w=0.51u l=0.6u
X15234 a_21748_18946# cap_shunt_p a_21540_19292# vdd pmos_6p0 w=1.2u l=0.5u
X15235 a_14372_41620# cap_shunt_n a_14580_42104# vdd pmos_6p0 w=1.2u l=0.5u
X15236 a_37444_39672# cap_shunt_gyp a_37632_39672# vdd pmos_6p0 w=1.215u l=0.5u
X15237 a_25572_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15238 vdd tune_shunt[7] a_3620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X15239 vss tune_shunt[7] a_9876_15448# vss nmos_6p0 w=0.51u l=0.6u
X15240 a_11032_22020# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15241 a_21540_42812# cap_shunt_n a_21748_42466# vdd pmos_6p0 w=1.2u l=0.5u
X15242 a_24660_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15243 a_7748_26786# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15244 vss tune_shunt[7] a_32612_29922# vss nmos_6p0 w=0.51u l=0.6u
X15245 a_17620_25940# cap_shunt_n a_17828_26424# vdd pmos_6p0 w=1.2u l=0.5u
X15246 a_36232_22020# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X15247 a_22680_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15248 vdd tune_shunt[7] a_2500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X15249 a_6572_5556# cap_series_gyp a_6760_5556# vdd pmos_6p0 w=1.2u l=0.5u
X15250 vss tune_series_gygy[4] a_35880_10260# vss nmos_6p0 w=0.51u l=0.6u
X15251 a_21748_15810# cap_series_gyn a_21540_16156# vdd pmos_6p0 w=1.2u l=0.5u
X15252 a_17828_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15253 vdd a_33164_23895# a_33076_23992# vdd pmos_6p0 w=1.22u l=1u
X15254 a_29700_14242# cap_series_gyp a_29492_14588# vdd pmos_6p0 w=1.2u l=0.5u
X15255 a_25780_18584# cap_series_gyn a_25572_18100# vdd pmos_6p0 w=1.2u l=0.5u
X15256 vdd tune_shunt[7] a_3620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X15257 a_13000_9176# cap_series_gyp a_11800_8692# vss nmos_6p0 w=0.82u l=0.6u
X15258 a_12768_23588# cap_shunt_n a_10660_23650# vss nmos_6p0 w=0.82u l=0.6u
X15259 a_31436_20860# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15260 vdd a_3484_53687# a_3396_53784# vdd pmos_6p0 w=1.22u l=1u
X15261 a_17620_22804# cap_shunt_n a_17828_23288# vdd pmos_6p0 w=1.2u l=0.5u
X15262 vdd tune_shunt[7] a_16500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X15263 a_29720_13020# cap_series_gyn a_29532_13020# vdd pmos_6p0 w=1.2u l=0.5u
X15264 vss cap_shunt_gyn a_34188_45240# vss nmos_6p0 w=0.82u l=0.6u
X15265 a_17828_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15266 a_10452_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15267 a_14692_9176# cap_series_gyn a_15624_9176# vss nmos_6p0 w=0.82u l=0.6u
X15268 vdd tune_shunt[7] a_20532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X15269 a_15700_9538# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X15270 a_35292_50984# a_35204_51028# vss vss nmos_6p0 w=0.82u l=1u
X15271 vdd a_27788_47848# a_27700_47892# vdd pmos_6p0 w=1.22u l=1u
X15272 a_10548_27992# cap_shunt_n a_10340_27508# vdd pmos_6p0 w=1.2u l=0.5u
X15273 a_9876_12312# cap_shunt_p a_11592_12312# vss nmos_6p0 w=0.82u l=0.6u
X15274 a_19544_4472# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X15275 a_30640_21720# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X15276 a_9876_48376# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15277 vss cap_shunt_p a_31808_34564# vss nmos_6p0 w=0.82u l=0.6u
X15278 a_31708_16488# a_31620_16532# vss vss nmos_6p0 w=0.82u l=1u
X15279 a_15120_37700# cap_shunt_n a_13796_37762# vss nmos_6p0 w=0.82u l=0.6u
X15280 a_28692_32696# cap_shunt_p a_28484_32212# vdd pmos_6p0 w=1.2u l=0.5u
X15281 vdd tune_shunt[7] a_20532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X15282 a_22456_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15283 a_6508_23895# a_6420_23992# vss vss nmos_6p0 w=0.82u l=1u
X15284 vdd a_27788_44712# a_27700_44756# vdd pmos_6p0 w=1.22u l=1u
X15285 a_11800_7124# cap_series_gyp a_11612_7124# vdd pmos_6p0 w=1.2u l=0.5u
X15286 a_10540_3944# a_10452_3988# vss vss nmos_6p0 w=0.82u l=1u
X15287 vss cap_series_gyn a_25984_14180# vss nmos_6p0 w=0.82u l=0.6u
X15288 a_32268_50984# a_32180_51028# vss vss nmos_6p0 w=0.82u l=1u
X15289 a_7952_3204# cap_shunt_n a_5844_3266# vss nmos_6p0 w=0.82u l=0.6u
X15290 vss tune_shunt[6] a_3828_34264# vss nmos_6p0 w=0.51u l=0.6u
X15291 vss cap_shunt_p a_31808_31428# vss nmos_6p0 w=0.82u l=0.6u
X15292 a_21748_28354# cap_shunt_n a_22680_28292# vss nmos_6p0 w=0.82u l=0.6u
X15293 vdd tune_shunt[7] a_17620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X15294 a_13888_6040# cap_series_gyn a_11780_6040# vss nmos_6p0 w=0.82u l=0.6u
X15295 vss cap_shunt_p a_9072_45540# vss nmos_6p0 w=0.82u l=0.6u
X15296 a_22456_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15297 a_32404_25564# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15298 vdd a_1692_55688# a_1604_55732# vdd pmos_6p0 w=1.22u l=1u
X15299 vss cap_series_gyp a_25984_11044# vss nmos_6p0 w=0.82u l=0.6u
X15300 a_5500_11784# a_5412_11828# vss vss nmos_6p0 w=0.82u l=1u
X15301 a_12580_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15302 a_17620_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15303 vss tune_shunt[1] a_1924_3266# vss nmos_6p0 w=0.51u l=0.6u
X15304 vss tune_series_gygy[5] a_34516_17378# vss nmos_6p0 w=0.51u l=0.6u
X15305 vss tune_shunt[7] a_3828_31128# vss nmos_6p0 w=0.51u l=0.6u
X15306 a_6740_34264# cap_shunt_n a_6532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X15307 a_10452_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15308 vss cap_series_gyp a_13000_9176# vss nmos_6p0 w=0.82u l=0.6u
X15309 a_21748_25218# cap_shunt_n a_22680_25156# vss nmos_6p0 w=0.82u l=0.6u
X15310 vdd tune_shunt[7] a_17620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X15311 vdd a_18940_54120# a_18852_54164# vdd pmos_6p0 w=1.22u l=1u
X15312 vss cap_shunt_n a_9072_42404# vss nmos_6p0 w=0.82u l=0.6u
X15313 a_7840_20452# cap_shunt_p a_6516_20514# vss nmos_6p0 w=0.82u l=0.6u
X15314 vss cap_shunt_n a_12656_23288# vss nmos_6p0 w=0.82u l=0.6u
X15315 a_10452_5180# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15316 vss tune_shunt[7] a_25780_21720# vss nmos_6p0 w=0.51u l=0.6u
X15317 a_6740_31128# cap_shunt_n a_6532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X15318 a_22644_12312# cap_series_gyn a_22436_11828# vdd pmos_6p0 w=1.2u l=0.5u
X15319 vdd a_37868_49416# a_37780_49460# vdd pmos_6p0 w=1.22u l=1u
X15320 a_21540_30268# cap_shunt_n a_21748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X15321 a_35740_52552# a_35652_52596# vss vss nmos_6p0 w=0.82u l=1u
X15322 a_28124_42711# a_28036_42808# vss vss nmos_6p0 w=0.82u l=1u
X15323 a_16924_29032# a_16836_29076# vss vss nmos_6p0 w=0.82u l=1u
X15324 a_32716_16055# a_32628_16152# vss vss nmos_6p0 w=0.82u l=1u
X15325 vdd a_18940_50984# a_18852_51028# vdd pmos_6p0 w=1.22u l=1u
X15326 vdd a_33948_41143# a_33860_41240# vdd pmos_6p0 w=1.22u l=1u
X15327 a_25572_32212# cap_shunt_p a_25780_32696# vdd pmos_6p0 w=1.2u l=0.5u
X15328 a_28484_32212# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15329 vss cap_shunt_n a_3248_6340# vss nmos_6p0 w=0.82u l=0.6u
X15330 a_25572_3988# tune_shunt[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15331 vdd a_15916_54120# a_15828_54164# vdd pmos_6p0 w=1.22u l=1u
X15332 a_35880_36916# cap_series_gygyp a_35692_36916# vdd pmos_6p0 w=1.2u l=0.5u
X15333 a_29916_47415# a_29828_47512# vss vss nmos_6p0 w=0.82u l=1u
X15334 vdd a_18492_49416# a_18404_49460# vdd pmos_6p0 w=1.22u l=1u
X15335 a_21540_36540# cap_shunt_n a_21748_36194# vdd pmos_6p0 w=1.2u l=0.5u
X15336 vss tune_series_gy[5] a_18612_11106# vss nmos_6p0 w=0.51u l=0.6u
X15337 a_16500_42812# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15338 a_23308_21192# a_23220_21236# vss vss nmos_6p0 w=0.82u l=1u
X15339 vdd a_37868_46280# a_37780_46324# vdd pmos_6p0 w=1.22u l=1u
X15340 a_26892_55255# a_26804_55352# vss vss nmos_6p0 w=0.82u l=1u
X15341 a_22680_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15342 a_16924_25896# a_16836_25940# vss vss nmos_6p0 w=0.82u l=1u
X15343 a_32716_52552# a_32628_52596# vss vss nmos_6p0 w=0.82u l=1u
X15344 vss cap_shunt_n a_3248_3204# vss nmos_6p0 w=0.82u l=0.6u
X15345 a_35692_18100# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15346 a_9876_53080# cap_shunt_n a_9668_52596# vdd pmos_6p0 w=1.2u l=0.5u
X15347 a_36688_37400# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X15348 a_25572_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15349 vdd tune_series_gy[4] a_28484_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15350 a_25548_49416# a_25460_49460# vss vss nmos_6p0 w=0.82u l=1u
X15351 a_21540_33404# cap_shunt_n a_21748_33058# vdd pmos_6p0 w=1.2u l=0.5u
X15352 a_18612_4472# cap_series_gyp a_18404_3988# vdd pmos_6p0 w=1.2u l=0.5u
X15353 a_5544_13880# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15354 a_35692_14964# cap_series_gygyn a_35880_14964# vdd pmos_6p0 w=1.2u l=0.5u
X15355 vdd a_3036_52552# a_2948_52596# vdd pmos_6p0 w=1.22u l=1u
X15356 a_17620_16532# cap_shunt_p a_17828_17016# vdd pmos_6p0 w=1.2u l=0.5u
X15357 a_13340_52552# a_13252_52596# vss vss nmos_6p0 w=0.82u l=1u
X15358 a_20532_46324# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15359 a_19152_21720# cap_shunt_p a_17828_21720# vss nmos_6p0 w=0.82u l=0.6u
X15360 a_6292_48738# cap_shunt_p a_6084_49084# vdd pmos_6p0 w=1.2u l=0.5u
X15361 vss tune_series_gygy[5] a_35880_24372# vss nmos_6p0 w=0.51u l=0.6u
X15362 a_16252_13352# a_16164_13396# vss vss nmos_6p0 w=0.82u l=1u
X15363 a_13588_47516# cap_shunt_p a_13796_47170# vdd pmos_6p0 w=1.2u l=0.5u
X15364 vss tune_shunt[6] a_2708_42466# vss nmos_6p0 w=0.51u l=0.6u
X15365 a_25548_46280# a_25460_46324# vss vss nmos_6p0 w=0.82u l=1u
X15366 a_35692_11828# cap_series_gygyp a_35880_11828# vdd pmos_6p0 w=1.2u l=0.5u
X15367 a_25572_41620# cap_shunt_n a_25780_42104# vdd pmos_6p0 w=1.2u l=0.5u
X15368 vss cap_shunt_p a_31808_28292# vss nmos_6p0 w=0.82u l=0.6u
X15369 vdd a_37196_30600# a_37108_30644# vdd pmos_6p0 w=1.22u l=1u
X15370 vdd tune_shunt[5] a_20532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X15371 vdd a_4492_8215# a_4404_8312# vdd pmos_6p0 w=1.22u l=1u
X15372 a_27900_55688# a_27812_55732# vss vss nmos_6p0 w=0.82u l=1u
X15373 a_19948_50551# a_19860_50648# vss vss nmos_6p0 w=0.82u l=1u
X15374 a_18816_29860# cap_shunt_n a_16708_29922# vss nmos_6p0 w=0.82u l=0.6u
X15375 a_10548_26424# cap_shunt_n a_10340_25940# vdd pmos_6p0 w=1.2u l=0.5u
X15376 vss tune_series_gygy[1] a_31624_8316# vss nmos_6p0 w=0.51u l=0.6u
X15377 a_33612_9783# a_33524_9880# vss vss nmos_6p0 w=0.82u l=1u
X15378 a_14372_41620# cap_shunt_n a_14580_42104# vdd pmos_6p0 w=1.2u l=0.5u
X15379 vdd tune_shunt[6] a_7540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X15380 vss cap_shunt_p a_31808_25156# vss nmos_6p0 w=0.82u l=0.6u
X15381 a_33544_29860# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15382 a_20720_4772# cap_series_gyp a_18612_4834# vss nmos_6p0 w=0.82u l=0.6u
X15383 vdd tune_shunt[6] a_29492_34972# vdd pmos_6p0 w=1.2u l=0.5u
X15384 vdd tune_shunt[7] a_20532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X15385 vss cap_shunt_p a_11984_48376# vss nmos_6p0 w=0.82u l=0.6u
X15386 vdd a_1692_49416# a_1604_49460# vdd pmos_6p0 w=1.22u l=1u
X15387 a_18816_26724# cap_shunt_n a_16708_26786# vss nmos_6p0 w=0.82u l=0.6u
X15388 a_10548_23288# cap_shunt_n a_10340_22804# vdd pmos_6p0 w=1.2u l=0.5u
X15389 a_20740_45240# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X15390 vss cap_shunt_p a_5152_43672# vss nmos_6p0 w=0.82u l=0.6u
X15391 a_33544_26724# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15392 a_25780_18584# cap_series_gyn a_25572_18100# vdd pmos_6p0 w=1.2u l=0.5u
X15393 vdd tune_shunt[5] a_29492_31836# vdd pmos_6p0 w=1.2u l=0.5u
X15394 vdd tune_shunt[7] a_17620_16532# vdd pmos_6p0 w=1.2u l=0.5u
X15395 vss cap_shunt_p a_14112_17016# vss nmos_6p0 w=0.82u l=0.6u
X15396 a_32156_52119# a_32068_52216# vss vss nmos_6p0 w=0.82u l=1u
X15397 vss cap_shunt_n a_9072_36132# vss nmos_6p0 w=0.82u l=0.6u
X15398 vdd tune_series_gy[4] a_24452_8316# vdd pmos_6p0 w=1.2u l=0.5u
X15399 a_22456_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15400 vdd a_1692_46280# a_1604_46324# vdd pmos_6p0 w=1.22u l=1u
X15401 vss cap_shunt_p a_15904_45540# vss nmos_6p0 w=0.82u l=0.6u
X15402 a_3620_33780# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15403 a_13796_28354# cap_shunt_n a_13588_28700# vdd pmos_6p0 w=1.2u l=0.5u
X15404 vdd tune_series_gy[5] a_25572_14964# vdd pmos_6p0 w=1.2u l=0.5u
X15405 vss tune_shunt[5] a_29700_36194# vss nmos_6p0 w=0.51u l=0.6u
X15406 a_12768_6340# cap_series_gyn a_10660_6402# vss nmos_6p0 w=0.82u l=0.6u
X15407 a_21748_20514# cap_shunt_p a_21540_20860# vdd pmos_6p0 w=1.2u l=0.5u
X15408 a_20740_42104# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15409 vss cap_shunt_n a_11872_38968# vss nmos_6p0 w=0.82u l=0.6u
X15410 a_6740_24856# cap_shunt_p a_6532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X15411 a_24204_43144# a_24116_43188# vss vss nmos_6p0 w=0.82u l=1u
X15412 vss cap_shunt_n a_5152_40536# vss nmos_6p0 w=0.82u l=0.6u
X15413 a_26712_20152# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X15414 a_28124_36439# a_28036_36536# vss vss nmos_6p0 w=0.82u l=1u
X15415 vss cap_shunt_n a_15904_42404# vss nmos_6p0 w=0.82u l=0.6u
X15416 vss tune_shunt[5] a_24660_40898# vss nmos_6p0 w=0.51u l=0.6u
X15417 a_3620_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15418 vdd tune_series_gy[5] a_25572_11828# vdd pmos_6p0 w=1.2u l=0.5u
X15419 vss tune_shunt[5] a_29700_33058# vss nmos_6p0 w=0.51u l=0.6u
X15420 vss tune_series_gy[5] a_25780_12312# vss nmos_6p0 w=0.51u l=0.6u
X15421 a_2932_10744# cap_shunt_n a_2724_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15422 a_6740_21720# cap_shunt_p a_6532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X15423 a_24204_40008# a_24116_40052# vss vss nmos_6p0 w=0.82u l=1u
X15424 a_16500_36540# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15425 vss cap_shunt_n a_4256_12312# vss nmos_6p0 w=0.82u l=0.6u
X15426 a_26892_48983# a_26804_49080# vss vss nmos_6p0 w=0.82u l=1u
X15427 a_5636_9884# cap_shunt_p a_5844_9538# vdd pmos_6p0 w=1.2u l=0.5u
X15428 a_18424_22020# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15429 vss cap_shunt_p a_4816_48676# vss nmos_6p0 w=0.82u l=0.6u
X15430 a_3828_42104# cap_shunt_p a_3620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X15431 vdd a_34396_55255# a_34308_55352# vdd pmos_6p0 w=1.22u l=1u
X15432 a_23464_18884# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15433 a_28684_50984# a_28596_51028# vss vss nmos_6p0 w=0.82u l=1u
X15434 a_21540_27132# cap_shunt_n a_21748_26786# vdd pmos_6p0 w=1.2u l=0.5u
X15435 vdd a_12892_52552# a_12804_52596# vdd pmos_6p0 w=1.22u l=1u
X15436 a_1692_38440# a_1604_38484# vss vss nmos_6p0 w=0.82u l=1u
X15437 a_16500_33404# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15438 a_9332_9884# cap_shunt_p a_9540_9538# vdd pmos_6p0 w=1.2u l=0.5u
X15439 a_8848_45240# cap_shunt_p a_6740_45240# vss nmos_6p0 w=0.82u l=0.6u
X15440 a_6292_17016# cap_shunt_p a_6084_16532# vdd pmos_6p0 w=1.2u l=0.5u
X15441 vss cap_series_gygyp a_36296_20152# vss nmos_6p0 w=0.82u l=0.6u
X15442 a_6740_34264# cap_shunt_n a_6532_33780# vdd pmos_6p0 w=1.2u l=0.5u
X15443 vss cap_series_gyp a_30016_7608# vss nmos_6p0 w=0.82u l=0.6u
X15444 a_9876_13880# cap_shunt_p a_9668_13396# vdd pmos_6p0 w=1.2u l=0.5u
X15445 vss tune_series_gygy[5] a_35880_18100# vss nmos_6p0 w=0.51u l=0.6u
X15446 vdd a_34396_52119# a_34308_52216# vdd pmos_6p0 w=1.22u l=1u
X15447 vss tune_shunt[6] a_2708_36194# vss nmos_6p0 w=0.51u l=0.6u
X15448 a_23464_15748# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X15449 a_10548_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15450 a_32604_53687# a_32516_53784# vss vss nmos_6p0 w=0.82u l=1u
X15451 vdd a_3036_43144# a_2948_43188# vdd pmos_6p0 w=1.22u l=1u
X15452 a_17620_33780# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15453 a_8848_42104# cap_shunt_n a_6740_42104# vss nmos_6p0 w=0.82u l=0.6u
X15454 a_3828_38968# cap_shunt_n a_5544_38968# vss nmos_6p0 w=0.82u l=0.6u
X15455 a_13588_38108# cap_shunt_n a_13796_37762# vdd pmos_6p0 w=1.2u l=0.5u
X15456 a_6740_31128# cap_shunt_n a_6532_30644# vdd pmos_6p0 w=1.2u l=0.5u
X15457 vss tune_series_gygy[4] a_35880_14964# vss nmos_6p0 w=0.51u l=0.6u
X15458 a_6740_37400# cap_shunt_n a_6532_36916# vdd pmos_6p0 w=1.2u l=0.5u
X15459 vss tune_shunt[7] a_2708_33058# vss nmos_6p0 w=0.51u l=0.6u
X15460 a_21540_30268# cap_shunt_n a_21748_29922# vdd pmos_6p0 w=1.2u l=0.5u
X15461 a_10680_8316# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X15462 a_10548_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15463 vss tune_series_gy[1] a_6760_5556# vss nmos_6p0 w=0.51u l=0.6u
X15464 a_32604_50551# a_32516_50648# vss vss nmos_6p0 w=0.82u l=1u
X15465 a_37632_50648# cap_shunt_gyn a_37444_50648# vdd pmos_6p0 w=1.215u l=0.5u
X15466 vdd tune_shunt[6] a_7540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X15467 a_25572_32212# cap_shunt_p a_25780_32696# vdd pmos_6p0 w=1.2u l=0.5u
X15468 a_19544_11044# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X15469 a_17620_30644# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15470 a_9428_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15471 a_21748_45602# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X15472 a_29492_34972# cap_shunt_p a_29700_34626# vdd pmos_6p0 w=1.2u l=0.5u
X15473 vdd a_6956_55255# a_6868_55352# vdd pmos_6p0 w=1.22u l=1u
X15474 a_25780_37400# cap_shunt_p a_26712_37400# vss nmos_6p0 w=0.82u l=0.6u
X15475 vdd tune_shunt[7] a_7540_33404# vdd pmos_6p0 w=1.2u l=0.5u
X15476 vdd a_23308_53687# a_23220_53784# vdd pmos_6p0 w=1.22u l=1u
X15477 a_16296_46808# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15478 a_25780_10744# cap_series_gyn a_25572_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15479 a_9876_53080# cap_shunt_n a_9668_52596# vdd pmos_6p0 w=1.2u l=0.5u
X15480 vdd tune_shunt[7] a_29492_25564# vdd pmos_6p0 w=1.2u l=0.5u
X15481 vdd a_35740_55688# a_35652_55732# vdd pmos_6p0 w=1.22u l=1u
X15482 vdd a_22972_54120# a_22884_54164# vdd pmos_6p0 w=1.22u l=1u
X15483 a_9856_43972# cap_shunt_p a_7748_44034# vss nmos_6p0 w=0.82u l=0.6u
X15484 a_29492_31836# cap_shunt_p a_29700_31490# vdd pmos_6p0 w=1.2u l=0.5u
X15485 a_18816_17316# cap_shunt_p a_16708_17378# vss nmos_6p0 w=0.82u l=0.6u
X15486 a_12332_22327# a_12244_22424# vss vss nmos_6p0 w=0.82u l=1u
X15487 a_13796_20514# cap_shunt_n a_13588_20860# vdd pmos_6p0 w=1.2u l=0.5u
X15488 vdd a_12108_53687# a_12020_53784# vdd pmos_6p0 w=1.22u l=1u
X15489 vdd a_23308_50551# a_23220_50648# vdd pmos_6p0 w=1.22u l=1u
X15490 a_6292_48738# cap_shunt_p a_6084_49084# vdd pmos_6p0 w=1.2u l=0.5u
X15491 vss cap_shunt_n a_5152_34264# vss nmos_6p0 w=0.82u l=0.6u
X15492 a_32156_42711# a_32068_42808# vss vss nmos_6p0 w=0.82u l=1u
X15493 vdd a_22972_50984# a_22884_51028# vdd pmos_6p0 w=1.22u l=1u
X15494 a_9856_40836# cap_shunt_n a_7748_40898# vss nmos_6p0 w=0.82u l=0.6u
X15495 vss cap_shunt_n a_8848_32696# vss nmos_6p0 w=0.82u l=0.6u
X15496 a_3620_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15497 a_25572_41620# cap_shunt_n a_25780_42104# vdd pmos_6p0 w=1.2u l=0.5u
X15498 vss cap_shunt_n a_15904_36132# vss nmos_6p0 w=0.82u l=0.6u
X15499 a_21748_11106# cap_series_gyn a_21540_11452# vdd pmos_6p0 w=1.2u l=0.5u
X15500 a_6956_33303# a_6868_33400# vss vss nmos_6p0 w=0.82u l=1u
X15501 a_12656_37400# cap_shunt_n a_10548_37400# vss nmos_6p0 w=0.82u l=0.6u
X15502 a_24204_33736# a_24116_33780# vss vss nmos_6p0 w=0.82u l=1u
X15503 a_4032_29860# cap_shunt_n a_2708_29922# vss nmos_6p0 w=0.82u l=0.6u
X15504 a_9644_3944# a_9556_3988# vss vss nmos_6p0 w=0.82u l=1u
X15505 vss cap_shunt_n a_5152_31128# vss nmos_6p0 w=0.82u l=0.6u
X15506 a_10548_26424# cap_shunt_n a_10340_25940# vdd pmos_6p0 w=1.2u l=0.5u
X15507 vdd a_4940_3944# a_4852_3988# vdd pmos_6p0 w=1.22u l=1u
X15508 vdd tune_shunt[7] a_9668_21236# vdd pmos_6p0 w=1.2u l=0.5u
X15509 a_37420_12919# a_37332_13016# vss vss nmos_6p0 w=0.82u l=1u
X15510 a_3620_21236# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15511 a_17640_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15512 a_2708_23650# cap_shunt_p a_2500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X15513 a_36384_45944# cap_shunt_gyp a_36384_45540# vdd pmos_6p0 w=1.215u l=0.5u
X15514 a_29700_37762# cap_shunt_n a_29492_38108# vdd pmos_6p0 w=1.2u l=0.5u
X15515 a_6292_50306# cap_shunt_p a_6084_50652# vdd pmos_6p0 w=1.2u l=0.5u
X15516 a_28684_44712# a_28596_44756# vss vss nmos_6p0 w=0.82u l=1u
X15517 a_24204_30600# a_24116_30644# vss vss nmos_6p0 w=0.82u l=1u
X15518 a_4032_26724# cap_shunt_p a_2708_26786# vss nmos_6p0 w=0.82u l=0.6u
X15519 a_16500_27132# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15520 a_16800_4472# cap_series_gyp a_14692_4472# vss nmos_6p0 w=0.82u l=0.6u
X15521 a_11144_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15522 a_4704_51512# cap_shunt_n a_3380_51512# vss nmos_6p0 w=0.82u l=0.6u
X15523 a_34560_9476# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X15524 a_10548_23288# cap_shunt_n a_10340_22804# vdd pmos_6p0 w=1.2u l=0.5u
X15525 vdd a_21964_47415# a_21876_47512# vdd pmos_6p0 w=1.22u l=1u
X15526 vss cap_shunt_n a_4816_39268# vss nmos_6p0 w=0.82u l=0.6u
X15527 a_3828_32696# cap_shunt_p a_3620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X15528 vss tune_series_gy[5] a_19732_13880# vss nmos_6p0 w=0.51u l=0.6u
X15529 a_34516_23650# cap_series_gygyp a_34308_23996# vdd pmos_6p0 w=1.2u l=0.5u
X15530 a_25780_7608# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X15531 vss cap_series_gyn a_11872_3204# vss nmos_6p0 w=0.82u l=0.6u
X15532 a_9108_49084# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15533 a_16708_47170# cap_shunt_n a_18424_47108# vss nmos_6p0 w=0.82u l=0.6u
X15534 a_36384_42808# cap_shunt_gyn a_36384_42404# vdd pmos_6p0 w=1.215u l=0.5u
X15535 a_13796_28354# cap_shunt_n a_13588_28700# vdd pmos_6p0 w=1.2u l=0.5u
X15536 vdd a_14012_55255# a_13924_55352# vdd pmos_6p0 w=1.22u l=1u
X15537 vdd a_22636_47848# a_22548_47892# vdd pmos_6p0 w=1.22u l=1u
X15538 vss cap_shunt_n a_26768_29860# vss nmos_6p0 w=0.82u l=0.6u
X15539 a_6740_24856# cap_shunt_p a_6532_24372# vdd pmos_6p0 w=1.2u l=0.5u
X15540 a_14692_4472# cap_series_gyp a_14484_3988# vdd pmos_6p0 w=1.2u l=0.5u
X15541 vss tune_series_gy[5] a_19732_10744# vss nmos_6p0 w=0.51u l=0.6u
X15542 a_6760_5556# cap_series_gyp a_6784_6040# vss nmos_6p0 w=0.82u l=0.6u
X15543 a_34516_4834# cap_series_gygyp a_36232_4772# vss nmos_6p0 w=0.82u l=0.6u
X15544 a_37632_44376# cap_shunt_gyp a_37444_44376# vdd pmos_6p0 w=1.215u l=0.5u
X15545 vdd tune_shunt[6] a_14372_44756# vdd pmos_6p0 w=1.2u l=0.5u
X15546 vss cap_shunt_p a_27104_32696# vss nmos_6p0 w=0.82u l=0.6u
X15547 a_3828_20152# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X15548 vdd a_14012_52119# a_13924_52216# vdd pmos_6p0 w=1.22u l=1u
X15549 a_16500_45948# cap_shunt_p a_16708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X15550 a_35448_32696# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15551 a_17620_24372# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15552 vss cap_shunt_p a_26768_26724# vss nmos_6p0 w=0.82u l=0.6u
X15553 a_8412_54120# a_8324_54164# vss vss nmos_6p0 w=0.82u l=1u
X15554 a_6740_21720# cap_shunt_p a_6532_21236# vdd pmos_6p0 w=1.2u l=0.5u
X15555 vdd tune_shunt[4] a_21540_45948# vdd pmos_6p0 w=1.2u l=0.5u
X15556 a_6740_27992# cap_shunt_n a_6532_27508# vdd pmos_6p0 w=1.2u l=0.5u
X15557 a_25548_52119# a_25460_52216# vss vss nmos_6p0 w=0.82u l=1u
X15558 a_21748_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15559 a_29700_31490# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X15560 a_32156_8648# a_32068_8692# vss vss nmos_6p0 w=0.82u l=1u
X15561 vdd tune_shunt[7] a_7540_27132# vdd pmos_6p0 w=1.2u l=0.5u
X15562 a_6292_49944# cap_shunt_p a_6084_49460# vdd pmos_6p0 w=1.2u l=0.5u
X15563 a_2932_9176# cap_shunt_n a_2724_8692# vdd pmos_6p0 w=1.2u l=0.5u
X15564 a_35180_36439# a_35092_36536# vss vss nmos_6p0 w=0.82u l=1u
X15565 a_10452_6748# cap_series_gyn a_10660_6402# vdd pmos_6p0 w=1.2u l=0.5u
X15566 a_17620_21236# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15567 a_35692_10260# tune_series_gygy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15568 a_14896_18584# cap_shunt_p a_12788_18584# vss nmos_6p0 w=0.82u l=0.6u
X15569 a_29492_25564# cap_shunt_p a_29700_25218# vdd pmos_6p0 w=1.2u l=0.5u
X15570 a_10452_23996# cap_shunt_n a_10660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X15571 vss cap_shunt_p a_19936_20152# vss nmos_6p0 w=0.82u l=0.6u
X15572 vss tune_series_gy[4] a_29720_13020# vss nmos_6p0 w=0.51u l=0.6u
X15573 a_9668_16532# cap_shunt_p a_9876_17016# vdd pmos_6p0 w=1.2u l=0.5u
X15574 a_31260_40008# a_31172_40052# vss vss nmos_6p0 w=0.82u l=1u
X15575 vss cap_shunt_p a_23072_39268# vss nmos_6p0 w=0.82u l=0.6u
X15576 vss tune_shunt[6] a_24660_37762# vss nmos_6p0 w=0.51u l=0.6u
X15577 a_10920_51812# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15578 vss tune_series_gy[5] a_21748_7970# vss nmos_6p0 w=0.51u l=0.6u
X15579 a_8064_13880# cap_shunt_p a_6740_13880# vss nmos_6p0 w=0.82u l=0.6u
X15580 a_35264_47512# cap_shunt_gyn a_35264_47108# vdd pmos_6p0 w=1.215u l=0.5u
X15581 vdd a_16700_14920# a_16612_14964# vdd pmos_6p0 w=1.22u l=1u
X15582 a_14896_15448# cap_shunt_p a_12788_15448# vss nmos_6p0 w=0.82u l=0.6u
X15583 vdd a_2588_33736# a_2500_33780# vdd pmos_6p0 w=1.22u l=1u
X15584 a_9856_34564# cap_shunt_n a_7748_34626# vss nmos_6p0 w=0.82u l=0.6u
X15585 vdd a_32716_49416# a_32628_49460# vdd pmos_6p0 w=1.22u l=1u
X15586 vdd a_20620_41143# a_20532_41240# vdd pmos_6p0 w=1.22u l=1u
X15587 a_37868_5079# a_37780_5176# vss vss nmos_6p0 w=0.82u l=1u
X15588 vdd a_17260_12919# a_17172_13016# vdd pmos_6p0 w=1.22u l=1u
X15589 vss tune_shunt[6] a_24660_34626# vss nmos_6p0 w=0.51u l=0.6u
X15590 a_9540_9538# cap_shunt_p a_9332_9884# vdd pmos_6p0 w=1.2u l=0.5u
X15591 vdd a_27788_55255# a_27700_55352# vdd pmos_6p0 w=1.22u l=1u
X15592 vss tune_shunt[7] a_10660_29922# vss nmos_6p0 w=0.51u l=0.6u
X15593 vss tune_series_gy[4] a_21748_4834# vss nmos_6p0 w=0.51u l=0.6u
X15594 a_2708_9538# cap_shunt_n a_2500_9884# vdd pmos_6p0 w=1.2u l=0.5u
X15595 a_23420_49416# a_23332_49460# vss vss nmos_6p0 w=0.82u l=1u
X15596 vdd a_16700_11784# a_16612_11828# vdd pmos_6p0 w=1.22u l=1u
X15597 a_33500_13352# a_33412_13396# vss vss nmos_6p0 w=0.82u l=1u
X15598 vdd a_2588_30600# a_2500_30644# vdd pmos_6p0 w=1.22u l=1u
X15599 a_20532_41620# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15600 a_25572_32212# cap_shunt_p a_25780_32696# vdd pmos_6p0 w=1.2u l=0.5u
X15601 a_9856_31428# cap_shunt_n a_7748_31490# vss nmos_6p0 w=0.82u l=0.6u
X15602 vss cap_shunt_p a_8848_23288# vss nmos_6p0 w=0.82u l=0.6u
X15603 vdd a_34844_18056# a_34756_18100# vdd pmos_6p0 w=1.22u l=1u
X15604 a_6956_23895# a_6868_23992# vss vss nmos_6p0 w=0.82u l=1u
X15605 vss tune_series_gy[3] a_11800_7124# vss nmos_6p0 w=0.51u l=0.6u
X15606 vdd tune_shunt[7] a_32404_30268# vdd pmos_6p0 w=1.2u l=0.5u
X15607 vdd a_27788_52119# a_27700_52216# vdd pmos_6p0 w=1.22u l=1u
X15608 a_13588_42812# cap_shunt_n a_13796_42466# vdd pmos_6p0 w=1.2u l=0.5u
X15609 a_15700_7970# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X15610 vdd tune_shunt[6] a_10452_44380# vdd pmos_6p0 w=1.2u l=0.5u
X15611 vss cap_series_gyp a_21840_9176# vss nmos_6p0 w=0.82u l=0.6u
X15612 a_33500_10216# a_33412_10260# vss vss nmos_6p0 w=0.82u l=1u
X15613 vdd tune_shunt[1] a_5636_3612# vdd pmos_6p0 w=1.2u l=0.5u
X15614 a_29532_9884# cap_series_gyn a_29720_9884# vdd pmos_6p0 w=1.2u l=0.5u
X15615 a_12788_48376# cap_shunt_p a_14504_48376# vss nmos_6p0 w=0.82u l=0.6u
X15616 a_10660_37762# cap_shunt_n a_12376_37700# vss nmos_6p0 w=0.82u l=0.6u
X15617 vdd tune_shunt[2] a_1716_6748# vdd pmos_6p0 w=1.2u l=0.5u
X15618 a_17828_18584# cap_shunt_p a_17620_18100# vdd pmos_6p0 w=1.2u l=0.5u
X15619 a_10540_55255# a_10452_55352# vss vss nmos_6p0 w=0.82u l=1u
X15620 a_16632_9476# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X15621 a_25780_10744# cap_series_gyn a_25572_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15622 a_2708_14242# cap_shunt_n a_2500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X15623 a_9876_53080# cap_shunt_n a_9668_52596# vdd pmos_6p0 w=1.2u l=0.5u
X15624 a_7540_44380# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15625 a_35740_38440# a_35652_38484# vss vss nmos_6p0 w=0.82u l=1u
X15626 vdd tune_shunt[6] a_11460_40052# vdd pmos_6p0 w=1.2u l=0.5u
X15627 a_15700_4834# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X15628 a_4032_17316# cap_shunt_p a_2708_17378# vss nmos_6p0 w=0.82u l=0.6u
X15629 vss tune_shunt[6] a_11668_46808# vss nmos_6p0 w=0.51u l=0.6u
X15630 vdd tune_shunt[6] a_10452_41244# vdd pmos_6p0 w=1.2u l=0.5u
X15631 vdd tune_shunt[6] a_25572_38484# vdd pmos_6p0 w=1.2u l=0.5u
X15632 vdd a_20172_33303# a_20084_33400# vdd pmos_6p0 w=1.22u l=1u
X15633 a_28572_9783# a_28484_9880# vss vss nmos_6p0 w=0.82u l=1u
X15634 a_21748_44034# cap_shunt_n a_21540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X15635 a_13796_20514# cap_shunt_n a_13588_20860# vdd pmos_6p0 w=1.2u l=0.5u
X15636 a_6740_43672# cap_shunt_p a_7672_43672# vss nmos_6p0 w=0.82u l=0.6u
X15637 a_10452_5180# cap_series_gyp a_10660_4834# vdd pmos_6p0 w=1.2u l=0.5u
X15638 a_5636_10260# cap_shunt_p a_5844_10744# vdd pmos_6p0 w=1.2u l=0.5u
X15639 a_1692_44279# a_1604_44376# vss vss nmos_6p0 w=0.82u l=1u
X15640 a_7540_41244# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15641 vdd a_30364_53687# a_30276_53784# vdd pmos_6p0 w=1.22u l=1u
X15642 a_2500_45948# cap_shunt_p a_2708_45602# vdd pmos_6p0 w=1.2u l=0.5u
X15643 a_25572_3988# cap_shunt_p a_25780_4472# vdd pmos_6p0 w=1.2u l=0.5u
X15644 a_16500_39676# cap_shunt_n a_16708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X15645 vdd tune_shunt[6] a_25572_35348# vdd pmos_6p0 w=1.2u l=0.5u
X15646 a_30408_13880# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X15647 a_30140_41576# a_30052_41620# vss vss nmos_6p0 w=0.82u l=1u
X15648 a_21748_40898# cap_shunt_p a_21540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X15649 a_6740_40536# cap_shunt_n a_7672_40536# vss nmos_6p0 w=0.82u l=0.6u
X15650 a_28572_42711# a_28484_42808# vss vss nmos_6p0 w=0.82u l=1u
X15651 vdd tune_shunt[6] a_21540_39676# vdd pmos_6p0 w=1.2u l=0.5u
X15652 a_35880_7124# tune_series_gygy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X15653 a_13460_38968# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15654 vdd tune_shunt[5] a_6084_17724# vdd pmos_6p0 w=1.2u l=0.5u
X15655 vdd a_30364_50551# a_30276_50648# vdd pmos_6p0 w=1.22u l=1u
X15656 a_1692_41143# a_1604_41240# vss vss nmos_6p0 w=0.82u l=1u
X15657 vss cap_shunt_p a_27104_23288# vss nmos_6p0 w=0.82u l=0.6u
X15658 a_30408_10744# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X15659 a_2708_23650# cap_shunt_p a_2500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X15660 vdd a_6956_5079# a_6868_5176# vdd pmos_6p0 w=1.22u l=1u
X15661 a_12580_19668# cap_shunt_p a_12788_20152# vdd pmos_6p0 w=1.2u l=0.5u
X15662 a_23756_21192# a_23668_21236# vss vss nmos_6p0 w=0.82u l=1u
X15663 a_29700_37762# cap_shunt_n a_29492_38108# vdd pmos_6p0 w=1.2u l=0.5u
X15664 a_25572_13396# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15665 vss cap_series_gyp a_26768_17316# vss nmos_6p0 w=0.82u l=0.6u
X15666 vdd a_19276_45847# a_19188_45944# vdd pmos_6p0 w=1.22u l=1u
X15667 a_16708_37762# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15668 a_31260_33736# a_31172_33780# vss vss nmos_6p0 w=0.82u l=1u
X15669 a_13588_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15670 a_25984_18884# cap_series_gyn a_24660_18946# vss nmos_6p0 w=0.82u l=0.6u
X15671 a_8300_55255# a_8212_55352# vss vss nmos_6p0 w=0.82u l=1u
X15672 a_25996_49416# a_25908_49460# vss vss nmos_6p0 w=0.82u l=1u
X15673 a_16028_36872# a_15940_36916# vss vss nmos_6p0 w=0.82u l=1u
X15674 a_35880_25940# cap_series_gygyp a_35692_25940# vdd pmos_6p0 w=1.2u l=0.5u
X15675 a_28484_38484# cap_shunt_n a_28692_38968# vdd pmos_6p0 w=1.2u l=0.5u
X15676 vdd a_24204_36872# a_24116_36916# vdd pmos_6p0 w=1.22u l=1u
X15677 a_10340_33780# cap_shunt_n a_10548_34264# vdd pmos_6p0 w=1.2u l=0.5u
X15678 a_34516_23650# cap_series_gygyp a_34308_23996# vdd pmos_6p0 w=1.2u l=0.5u
X15679 vdd a_3484_52552# a_3396_52596# vdd pmos_6p0 w=1.22u l=1u
X15680 a_37868_34871# a_37780_34968# vss vss nmos_6p0 w=0.82u l=1u
X15681 vdd tune_shunt[5] a_17620_46324# vdd pmos_6p0 w=1.2u l=0.5u
X15682 a_9856_28292# cap_shunt_n a_7748_28354# vss nmos_6p0 w=0.82u l=0.6u
X15683 vdd a_19276_42711# a_19188_42808# vdd pmos_6p0 w=1.22u l=1u
X15684 a_16708_34626# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15685 a_19544_43672# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15686 a_31260_30600# a_31172_30644# vss vss nmos_6p0 w=0.82u l=1u
X15687 vss tune_shunt[7] a_24660_28354# vss nmos_6p0 w=0.51u l=0.6u
X15688 a_25984_15748# cap_series_gyn a_24660_15810# vss nmos_6p0 w=0.82u l=0.6u
X15689 vdd a_27788_48983# a_27700_49080# vdd pmos_6p0 w=1.22u l=1u
X15690 a_25996_46280# a_25908_46324# vss vss nmos_6p0 w=0.82u l=1u
X15691 a_35880_22804# cap_series_gygyp a_35692_22804# vdd pmos_6p0 w=1.2u l=0.5u
X15692 a_28484_35348# cap_shunt_p a_28692_35832# vdd pmos_6p0 w=1.2u l=0.5u
X15693 a_5936_32696# cap_shunt_p a_3828_32696# vss nmos_6p0 w=0.82u l=0.6u
X15694 a_10340_30644# cap_shunt_n a_10548_31128# vdd pmos_6p0 w=1.2u l=0.5u
X15695 vss cap_series_gyp a_11880_7908# vss nmos_6p0 w=0.82u l=0.6u
X15696 a_37868_31735# a_37780_31832# vss vss nmos_6p0 w=0.82u l=1u
X15697 vdd a_2588_24328# a_2500_24372# vdd pmos_6p0 w=1.22u l=1u
X15698 a_4816_12612# cap_shunt_n a_2708_12674# vss nmos_6p0 w=0.82u l=0.6u
X15699 a_9856_25156# cap_shunt_n a_7748_25218# vss nmos_6p0 w=0.82u l=0.6u
X15700 a_18044_54120# a_17956_54164# vss vss nmos_6p0 w=0.82u l=1u
X15701 a_19544_40536# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15702 a_10660_45602# cap_shunt_n a_10452_45948# vdd pmos_6p0 w=1.2u l=0.5u
X15703 vss tune_shunt[7] a_24660_25218# vss nmos_6p0 w=0.51u l=0.6u
X15704 a_13588_36540# cap_shunt_n a_13796_36194# vdd pmos_6p0 w=1.2u l=0.5u
X15705 a_35868_49944# cap_shunt_gyp a_35600_50006# vss nmos_6p0 w=0.82u l=0.6u
X15706 vdd tune_series_gy[5] a_22436_8692# vdd pmos_6p0 w=1.2u l=0.5u
X15707 vdd a_2588_21192# a_2500_21236# vdd pmos_6p0 w=1.22u l=1u
X15708 vss cap_shunt_p a_30016_40536# vss nmos_6p0 w=0.82u l=0.6u
X15709 a_6292_49944# cap_shunt_p a_6084_49460# vdd pmos_6p0 w=1.2u l=0.5u
X15710 a_20532_32212# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15711 a_22436_13396# cap_series_gyn a_22644_13880# vdd pmos_6p0 w=1.2u l=0.5u
X15712 a_9428_20514# cap_shunt_p a_9220_20860# vdd pmos_6p0 w=1.2u l=0.5u
X15713 a_13588_33404# cap_shunt_n a_13796_33058# vdd pmos_6p0 w=1.2u l=0.5u
X15714 a_16708_23650# cap_shunt_n a_16500_23996# vdd pmos_6p0 w=1.2u l=0.5u
X15715 a_2708_33058# cap_shunt_p a_3640_32996# vss nmos_6p0 w=0.82u l=0.6u
X15716 a_10452_23996# cap_shunt_n a_10660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X15717 a_35868_46808# cap_shunt_gyp a_35600_46870# vss nmos_6p0 w=0.82u l=0.6u
X15718 a_32040_7908# cap_series_gygyn a_31624_8316# vss nmos_6p0 w=0.82u l=0.6u
X15719 vss tune_shunt[7] a_13796_18946# vss nmos_6p0 w=0.51u l=0.6u
X15720 vdd tune_series_gygy[0] a_31436_6748# vdd pmos_6p0 w=1.2u l=0.5u
X15721 a_2708_45602# cap_shunt_p a_4424_45540# vss nmos_6p0 w=0.82u l=0.6u
X15722 vss cap_series_gyp a_20720_9476# vss nmos_6p0 w=0.82u l=0.6u
X15723 a_2500_39676# cap_shunt_n a_2708_39330# vdd pmos_6p0 w=1.2u l=0.5u
X15724 vdd tune_shunt[3] a_2724_10260# vdd pmos_6p0 w=1.2u l=0.5u
X15725 a_2708_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15726 vdd tune_shunt[7] a_25572_29076# vdd pmos_6p0 w=1.2u l=0.5u
X15727 vdd a_19724_44279# a_19636_44376# vdd pmos_6p0 w=1.22u l=1u
X15728 a_24652_43144# a_24564_43188# vss vss nmos_6p0 w=0.82u l=1u
X15729 vss tune_shunt[5] a_29700_37762# vss nmos_6p0 w=0.51u l=0.6u
X15730 a_11592_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15731 vss tune_shunt[6] a_9316_48738# vss nmos_6p0 w=0.51u l=0.6u
X15732 a_6740_34264# cap_shunt_n a_7672_34264# vss nmos_6p0 w=0.82u l=0.6u
X15733 a_32828_43144# a_32740_43188# vss vss nmos_6p0 w=0.82u l=1u
X15734 a_28572_36439# a_28484_36536# vss vss nmos_6p0 w=0.82u l=1u
X15735 a_2708_42466# cap_shunt_p a_4424_42404# vss nmos_6p0 w=0.82u l=0.6u
X15736 vdd a_33948_40008# a_33860_40052# vdd pmos_6p0 w=1.22u l=1u
X15737 a_7768_8316# cap_series_gyn a_7580_8316# vdd pmos_6p0 w=1.2u l=0.5u
X15738 vss cap_series_gyn a_21056_13880# vss nmos_6p0 w=0.82u l=0.6u
X15739 a_37632_49080# cap_shunt_gyn a_37652_48676# vss nmos_6p0 w=0.82u l=0.6u
X15740 vdd a_30364_44279# a_30276_44376# vdd pmos_6p0 w=1.22u l=1u
X15741 a_1692_34871# a_1604_34968# vss vss nmos_6p0 w=0.82u l=1u
X15742 a_9332_16156# cap_shunt_p a_9540_15810# vdd pmos_6p0 w=1.2u l=0.5u
X15743 a_18404_3988# cap_series_gyp a_18612_4472# vdd pmos_6p0 w=1.2u l=0.5u
X15744 a_24652_40008# a_24564_40052# vss vss nmos_6p0 w=0.82u l=1u
X15745 vss tune_shunt[6] a_29700_34626# vss nmos_6p0 w=0.51u l=0.6u
X15746 a_11592_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15747 a_6740_31128# cap_shunt_n a_7672_31128# vss nmos_6p0 w=0.82u l=0.6u
X15748 a_29700_29922# cap_shunt_p a_29492_30268# vdd pmos_6p0 w=1.2u l=0.5u
X15749 vdd a_19276_39575# a_19188_39672# vdd pmos_6p0 w=1.22u l=1u
X15750 vss cap_series_gyn a_21056_10744# vss nmos_6p0 w=0.82u l=0.6u
X15751 a_29916_6647# a_29828_6744# vss vss nmos_6p0 w=0.82u l=1u
X15752 a_1692_31735# a_1604_31832# vss vss nmos_6p0 w=0.82u l=1u
X15753 a_2708_14242# cap_shunt_n a_2500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X15754 a_37868_28599# a_37780_28696# vss vss nmos_6p0 w=0.82u l=1u
X15755 a_6852_53442# cap_shunt_n a_6644_53788# vdd pmos_6p0 w=1.2u l=0.5u
X15756 vdd tune_shunt[6] a_11460_40052# vdd pmos_6p0 w=1.2u l=0.5u
X15757 a_29700_37762# cap_shunt_n a_30632_37700# vss nmos_6p0 w=0.82u l=0.6u
X15758 vdd a_19276_36439# a_19188_36536# vdd pmos_6p0 w=1.22u l=1u
X15759 a_16708_28354# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15760 a_22644_7608# cap_series_gyp a_22436_7124# vdd pmos_6p0 w=1.2u l=0.5u
X15761 a_21748_44034# cap_shunt_n a_21540_44380# vdd pmos_6p0 w=1.2u l=0.5u
X15762 a_10660_40898# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15763 a_13588_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15764 vdd tune_series_gy[3] a_11612_7124# vdd pmos_6p0 w=1.2u l=0.5u
X15765 a_5636_10260# cap_shunt_p a_5844_10744# vdd pmos_6p0 w=1.2u l=0.5u
X15766 a_20620_47415# a_20532_47512# vss vss nmos_6p0 w=0.82u l=1u
X15767 a_28484_29076# cap_shunt_p a_28692_29560# vdd pmos_6p0 w=1.2u l=0.5u
X15768 a_10340_24372# cap_shunt_n a_10548_24856# vdd pmos_6p0 w=1.2u l=0.5u
X15769 a_12580_14964# cap_shunt_p a_12788_15448# vdd pmos_6p0 w=1.2u l=0.5u
X15770 a_35880_16532# cap_series_gygyn a_35692_16532# vdd pmos_6p0 w=1.2u l=0.5u
X15771 vdd a_24204_27464# a_24116_27508# vdd pmos_6p0 w=1.22u l=1u
X15772 a_12264_38968# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15773 a_37868_25463# a_37780_25560# vss vss nmos_6p0 w=0.82u l=1u
X15774 a_16708_25218# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15775 vdd tune_shunt[7] a_6308_20860# vdd pmos_6p0 w=1.2u l=0.5u
X15776 a_19544_34264# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15777 vdd a_4492_7080# a_4404_7124# vdd pmos_6p0 w=1.22u l=1u
X15778 a_21748_40898# cap_shunt_p a_21540_41244# vdd pmos_6p0 w=1.2u l=0.5u
X15779 a_10660_39330# cap_shunt_n a_10452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X15780 a_21448_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X15781 a_13104_6040# cap_series_gyn a_11780_6040# vss nmos_6p0 w=0.82u l=0.6u
X15782 a_12580_11828# cap_shunt_p a_12788_12312# vdd pmos_6p0 w=1.2u l=0.5u
X15783 vdd tune_shunt[6] a_13588_45948# vdd pmos_6p0 w=1.2u l=0.5u
X15784 a_5936_23288# cap_shunt_p a_3828_23288# vss nmos_6p0 w=0.82u l=0.6u
X15785 a_10660_4834# cap_series_gyp a_10452_5180# vdd pmos_6p0 w=1.2u l=0.5u
X15786 a_32444_14588# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15787 a_13796_20514# cap_shunt_n a_14728_20452# vss nmos_6p0 w=0.82u l=0.6u
X15788 a_28692_32696# cap_shunt_p a_29624_32696# vss nmos_6p0 w=0.82u l=0.6u
X15789 vdd tune_shunt[5] a_6084_17724# vdd pmos_6p0 w=1.2u l=0.5u
X15790 a_9428_20514# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15791 vss cap_shunt_p a_30016_34264# vss nmos_6p0 w=0.82u l=0.6u
X15792 a_19544_31128# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15793 a_18612_4472# cap_series_gyp a_20328_4472# vss nmos_6p0 w=0.82u l=0.6u
X15794 a_29492_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15795 a_25780_4472# cap_shunt_p a_25572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X15796 vss cap_series_gyp a_12216_9176# vss nmos_6p0 w=0.82u l=0.6u
X15797 a_13588_27132# cap_shunt_n a_13796_26786# vdd pmos_6p0 w=1.2u l=0.5u
X15798 vss tune_shunt[6] a_17828_38968# vss nmos_6p0 w=0.51u l=0.6u
X15799 vdd a_23756_53687# a_23668_53784# vdd pmos_6p0 w=1.22u l=1u
X15800 vss cap_shunt_n a_30016_31128# vss nmos_6p0 w=0.82u l=0.6u
X15801 a_35880_25940# cap_series_gygyp a_35692_25940# vdd pmos_6p0 w=1.2u l=0.5u
X15802 a_5488_18584# cap_shunt_p a_3380_18584# vss nmos_6p0 w=0.82u l=0.6u
X15803 a_12780_22327# a_12692_22424# vss vss nmos_6p0 w=0.82u l=1u
X15804 a_16708_14242# cap_shunt_p a_16500_14588# vdd pmos_6p0 w=1.2u l=0.5u
X15805 a_2708_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15806 a_2708_23650# cap_shunt_p a_3640_23588# vss nmos_6p0 w=0.82u l=0.6u
X15807 a_13720_17016# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15808 vdd a_12556_53687# a_12468_53784# vdd pmos_6p0 w=1.22u l=1u
X15809 vdd a_23756_50551# a_23668_50648# vdd pmos_6p0 w=1.22u l=1u
X15810 a_24660_39330# cap_shunt_p a_25592_39268# vss nmos_6p0 w=0.82u l=0.6u
X15811 a_2140_38007# a_2052_38104# vss vss nmos_6p0 w=0.82u l=1u
X15812 a_15568_32696# cap_shunt_n a_13460_32696# vss nmos_6p0 w=0.82u l=0.6u
X15813 a_35880_22804# cap_series_gygyp a_35692_22804# vdd pmos_6p0 w=1.2u l=0.5u
X15814 a_6572_3988# cap_series_gyp a_6760_3988# vdd pmos_6p0 w=1.2u l=0.5u
X15815 a_2708_36194# cap_shunt_n a_4424_36132# vss nmos_6p0 w=0.82u l=0.6u
X15816 a_2500_13020# tune_shunt[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15817 a_1692_28599# a_1604_28696# vss vss nmos_6p0 w=0.82u l=1u
X15818 a_35880_8692# cap_series_gygyn a_35692_8692# vdd pmos_6p0 w=1.2u l=0.5u
X15819 a_3620_40052# cap_shunt_n a_3828_40536# vdd pmos_6p0 w=1.2u l=0.5u
X15820 a_12220_52119# a_12132_52216# vss vss nmos_6p0 w=0.82u l=1u
X15821 a_11668_45240# cap_shunt_n a_11460_44756# vdd pmos_6p0 w=1.2u l=0.5u
X15822 vdd a_31260_36872# a_31172_36916# vdd pmos_6p0 w=1.22u l=1u
X15823 a_2708_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15824 vss cap_shunt_n a_7168_3204# vss nmos_6p0 w=0.82u l=0.6u
X15825 a_28692_9176# cap_series_gyn a_28484_8692# vdd pmos_6p0 w=1.2u l=0.5u
X15826 vss tune_series_gy[5] a_24660_15810# vss nmos_6p0 w=0.51u l=0.6u
X15827 a_24652_33736# a_24564_33780# vss vss nmos_6p0 w=0.82u l=1u
X15828 vss tune_shunt[7] a_29700_28354# vss nmos_6p0 w=0.51u l=0.6u
X15829 a_36384_50244# cap_shunt_gyp a_36384_50648# vdd pmos_6p0 w=1.215u l=0.5u
X15830 a_10660_45602# cap_shunt_n a_10452_45948# vdd pmos_6p0 w=1.2u l=0.5u
X15831 a_37080_37400# cap_series_gygyp a_35880_36916# vss nmos_6p0 w=0.82u l=0.6u
X15832 a_18612_9538# cap_series_gyp a_18404_9884# vdd pmos_6p0 w=1.2u l=0.5u
X15833 vdd a_5612_34871# a_5524_34968# vdd pmos_6p0 w=1.22u l=1u
X15834 vss cap_shunt_p a_31024_32996# vss nmos_6p0 w=0.82u l=0.6u
X15835 a_37632_41621# cap_shunt_gyp a_37444_41621# vdd pmos_6p0 w=1.215u l=0.5u
X15836 a_35740_41143# a_35652_41240# vss vss nmos_6p0 w=0.82u l=1u
X15837 a_17828_38968# cap_shunt_n a_18760_38968# vss nmos_6p0 w=0.82u l=0.6u
X15838 a_1692_25463# a_1604_25560# vss vss nmos_6p0 w=0.82u l=1u
X15839 a_35880_5556# cap_series_gygyn a_35692_5556# vdd pmos_6p0 w=1.2u l=0.5u
X15840 vdd a_34396_54120# a_34308_54164# vdd pmos_6p0 w=1.22u l=1u
X15841 a_37632_39672# cap_shunt_gyp a_37652_39268# vss nmos_6p0 w=0.82u l=0.6u
X15842 a_2500_34972# cap_shunt_n a_2708_34626# vdd pmos_6p0 w=1.2u l=0.5u
X15843 a_6292_49944# cap_shunt_p a_6084_49460# vdd pmos_6p0 w=1.2u l=0.5u
X15844 a_28692_6040# cap_shunt_n a_28484_5556# vdd pmos_6p0 w=1.2u l=0.5u
X15845 a_34536_8316# cap_series_gygyp a_34560_7908# vss nmos_6p0 w=0.82u l=0.6u
X15846 a_24652_30600# a_24564_30644# vss vss nmos_6p0 w=0.82u l=1u
X15847 vss tune_shunt[7] a_29700_25218# vss nmos_6p0 w=0.51u l=0.6u
X15848 a_18612_6402# cap_series_gyn a_18404_6748# vdd pmos_6p0 w=1.2u l=0.5u
X15849 a_10452_23996# cap_shunt_n a_10660_23650# vdd pmos_6p0 w=1.2u l=0.5u
X15850 vdd a_34396_50984# a_34308_51028# vdd pmos_6p0 w=1.22u l=1u
X15851 a_2500_31836# cap_shunt_p a_2708_31490# vdd pmos_6p0 w=1.2u l=0.5u
X15852 a_36076_14487# a_35988_14584# vss vss nmos_6p0 w=0.82u l=1u
X15853 a_24452_17724# cap_series_gyp a_24660_17378# vdd pmos_6p0 w=1.2u l=0.5u
X15854 vss tune_shunt[6] a_6740_37400# vss nmos_6p0 w=0.51u l=0.6u
X15855 a_23968_9176# cap_series_gyp a_22644_9176# vss nmos_6p0 w=0.82u l=0.6u
X15856 vdd a_37532_52552# a_37444_52596# vdd pmos_6p0 w=1.22u l=1u
X15857 vss tune_series_gy[3] a_25780_7608# vss nmos_6p0 w=0.51u l=0.6u
X15858 a_9876_18584# cap_shunt_p a_9668_18100# vdd pmos_6p0 w=1.2u l=0.5u
X15859 a_10548_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15860 vdd tune_shunt[7] a_12580_18100# vdd pmos_6p0 w=1.2u l=0.5u
X15861 vdd a_14460_55255# a_14372_55352# vdd pmos_6p0 w=1.22u l=1u
X15862 vdd a_19276_27031# a_19188_27128# vdd pmos_6p0 w=1.22u l=1u
X15863 a_22076_54120# a_21988_54164# vss vss nmos_6p0 w=0.82u l=1u
X15864 vdd a_10988_3944# a_10900_3988# vdd pmos_6p0 w=1.22u l=1u
X15865 a_24452_8316# cap_series_gyp a_24660_7970# vdd pmos_6p0 w=1.2u l=0.5u
X15866 a_6292_17016# cap_shunt_p a_7224_17016# vss nmos_6p0 w=0.82u l=0.6u
X15867 a_31816_20152# cap_series_gygyn a_30616_19668# vss nmos_6p0 w=0.82u l=0.6u
X15868 a_16924_50984# a_16836_51028# vss vss nmos_6p0 w=0.82u l=1u
X15869 a_27160_3204# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15870 a_36076_11351# a_35988_11448# vss vss nmos_6p0 w=0.82u l=1u
X15871 a_35880_36916# tune_series_gygy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X15872 a_33948_22760# a_33860_22804# vss vss nmos_6p0 w=0.82u l=1u
X15873 a_31436_22428# cap_series_gygyn a_31624_22428# vdd pmos_6p0 w=1.2u l=0.5u
X15874 vss cap_series_gyn a_22848_4472# vss nmos_6p0 w=0.82u l=0.6u
X15875 a_6420_14588# cap_shunt_p a_6628_14242# vdd pmos_6p0 w=1.2u l=0.5u
X15876 vdd tune_shunt[6] a_3620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X15877 vdd tune_shunt[7] a_13588_39676# vdd pmos_6p0 w=1.2u l=0.5u
X15878 a_15720_11452# cap_series_gyp a_15532_11452# vdd pmos_6p0 w=1.2u l=0.5u
X15879 a_13796_14242# cap_shunt_p a_14728_14180# vss nmos_6p0 w=0.82u l=0.6u
X15880 a_10548_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15881 vdd a_14460_52119# a_14372_52216# vdd pmos_6p0 w=1.22u l=1u
X15882 a_7748_42466# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15883 a_9332_16156# cap_shunt_p a_9540_15810# vdd pmos_6p0 w=1.2u l=0.5u
X15884 vdd a_11436_55255# a_11348_55352# vdd pmos_6p0 w=1.22u l=1u
X15885 a_8860_54120# a_8772_54164# vss vss nmos_6p0 w=0.82u l=1u
X15886 a_7224_48676# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15887 a_14504_12312# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15888 a_17620_41620# cap_shunt_n a_17828_42104# vdd pmos_6p0 w=1.2u l=0.5u
X15889 a_24452_5180# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15890 a_25996_52119# a_25908_52216# vss vss nmos_6p0 w=0.82u l=1u
X15891 a_18760_46808# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15892 vdd tune_shunt[7] a_10340_36916# vdd pmos_6p0 w=1.2u l=0.5u
X15893 a_29700_29922# cap_shunt_p a_29492_30268# vdd pmos_6p0 w=1.2u l=0.5u
X15894 vdd a_15132_52552# a_15044_52596# vdd pmos_6p0 w=1.22u l=1u
X15895 a_33732_32696# cap_shunt_n a_33524_32212# vdd pmos_6p0 w=1.2u l=0.5u
X15896 a_28692_23288# cap_shunt_p a_29624_23288# vss nmos_6p0 w=0.82u l=0.6u
X15897 a_20328_9476# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X15898 a_11984_6340# cap_series_gyn a_10660_6402# vss nmos_6p0 w=0.82u l=0.6u
X15899 a_32268_9783# a_32180_9880# vss vss nmos_6p0 w=0.82u l=1u
X15900 a_8400_18884# cap_shunt_p a_6292_18946# vss nmos_6p0 w=0.82u l=0.6u
X15901 a_4380_52552# a_4292_52596# vss vss nmos_6p0 w=0.82u l=1u
X15902 a_35880_16532# cap_series_gygyn a_35692_16532# vdd pmos_6p0 w=1.2u l=0.5u
X15903 vss cap_shunt_p a_27888_38968# vss nmos_6p0 w=0.82u l=0.6u
X15904 a_24660_34626# cap_shunt_p a_24452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X15905 vss tune_shunt[6] a_28692_35832# vss nmos_6p0 w=0.51u l=0.6u
X15906 vss tune_shunt[7] a_6740_13880# vss nmos_6p0 w=0.51u l=0.6u
X15907 a_8400_15748# cap_shunt_p a_6292_15810# vss nmos_6p0 w=0.82u l=0.6u
X15908 a_22456_45240# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15909 a_8184_4772# cap_series_gyn a_7768_5180# vss nmos_6p0 w=0.82u l=0.6u
X15910 a_36384_43972# cap_shunt_gyp a_36384_44376# vdd pmos_6p0 w=1.215u l=0.5u
X15911 a_10660_39330# cap_shunt_n a_10452_39676# vdd pmos_6p0 w=1.2u l=0.5u
X15912 a_15568_23288# cap_shunt_n a_13460_23288# vss nmos_6p0 w=0.82u l=0.6u
X15913 a_9668_51028# cap_shunt_n a_9876_51512# vdd pmos_6p0 w=1.2u l=0.5u
X15914 a_22436_7124# cap_series_gyp a_22644_7608# vdd pmos_6p0 w=1.2u l=0.5u
X15915 a_33920_43189# tune_shunt_gy[6] vdd vdd pmos_6p0 w=1.215u l=0.5u
X15916 vdd a_5612_28599# a_5524_28696# vdd pmos_6p0 w=1.22u l=1u
X15917 vdd a_4940_5079# a_4852_5176# vdd pmos_6p0 w=1.22u l=1u
X15918 a_24660_31490# cap_shunt_p a_24452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X15919 a_32444_14588# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15920 vss tune_shunt[6] a_6404_47170# vss nmos_6p0 w=0.51u l=0.6u
X15921 vdd tune_shunt[6] a_17620_41620# vdd pmos_6p0 w=1.2u l=0.5u
X15922 a_22456_42104# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15923 a_1924_6402# cap_shunt_n a_1716_6748# vdd pmos_6p0 w=1.2u l=0.5u
X15924 vdd a_31260_27464# a_31172_27508# vdd pmos_6p0 w=1.22u l=1u
X15925 a_29468_20759# a_29380_20856# vss vss nmos_6p0 w=0.82u l=1u
X15926 vdd a_9644_44712# a_9556_44756# vdd pmos_6p0 w=1.22u l=1u
X15927 vss cap_shunt_p a_31024_23588# vss nmos_6p0 w=0.82u l=0.6u
X15928 vdd a_15356_13352# a_15268_13396# vdd pmos_6p0 w=1.22u l=1u
X15929 a_2500_25564# cap_shunt_p a_2708_25218# vdd pmos_6p0 w=1.2u l=0.5u
X15930 a_2500_45948# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15931 a_16500_17724# cap_shunt_p a_16708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X15932 a_31436_19292# cap_series_gygyn a_31624_19292# vdd pmos_6p0 w=1.2u l=0.5u
X15933 a_20740_21720# cap_shunt_p a_22456_21720# vss nmos_6p0 w=0.82u l=0.6u
X15934 a_7768_8316# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X15935 vss tune_shunt[4] a_20740_46808# vss nmos_6p0 w=0.51u l=0.6u
X15936 a_2500_22428# cap_shunt_p a_2708_22082# vdd pmos_6p0 w=1.2u l=0.5u
X15937 a_6740_20152# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15938 a_18032_47108# cap_shunt_n a_16708_47170# vss nmos_6p0 w=0.82u l=0.6u
X15939 a_24452_38108# cap_shunt_p a_24660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X15940 a_37444_49080# cap_shunt_gyn a_37632_49080# vdd pmos_6p0 w=1.215u l=0.5u
X15941 vss cap_series_gygyp a_36624_12612# vss nmos_6p0 w=0.82u l=0.6u
X15942 a_23464_43972# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X15943 a_2708_23650# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15944 a_7768_5180# tune_series_gy[1] vss vss nmos_6p0 w=0.51u l=0.6u
X15945 a_24660_39330# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15946 a_7748_36194# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X15947 a_35264_48676# cap_shunt_gyn a_35264_49080# vdd pmos_6p0 w=1.215u l=0.5u
X15948 a_21748_9538# cap_series_gyp a_22680_9476# vss nmos_6p0 w=0.82u l=0.6u
X15949 vss tune_series_gygy[5] a_35880_19668# vss nmos_6p0 w=0.51u l=0.6u
X15950 vss tune_shunt_gy[3] a_37632_45944# vss nmos_6p0 w=0.51u l=0.6u
X15951 a_22644_13880# cap_series_gyn a_23576_13880# vss nmos_6p0 w=0.82u l=0.6u
X15952 a_20532_25940# cap_shunt_n a_20740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X15953 a_25592_12612# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X15954 a_14372_46324# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15955 vdd tune_shunt[7] a_3620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X15956 a_17620_14964# cap_shunt_p a_17828_15448# vdd pmos_6p0 w=1.2u l=0.5u
X15957 a_23464_40836# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X15958 a_2708_20514# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X15959 a_7748_33058# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15960 a_18044_53687# a_17956_53784# vss vss nmos_6p0 w=0.82u l=1u
X15961 vdd a_24204_47415# a_24116_47512# vdd pmos_6p0 w=1.22u l=1u
X15962 vdd a_37084_38440# a_36996_38484# vdd pmos_6p0 w=1.22u l=1u
X15963 a_17620_32212# cap_shunt_n a_17828_32696# vdd pmos_6p0 w=1.2u l=0.5u
X15964 vss tune_shunt_gy[2] a_37632_42808# vss nmos_6p0 w=0.51u l=0.6u
X15965 a_22644_10744# cap_series_gyp a_23576_10744# vss nmos_6p0 w=0.82u l=0.6u
X15966 vdd tune_shunt[7] a_10340_27508# vdd pmos_6p0 w=1.2u l=0.5u
X15967 a_20532_22804# cap_shunt_p a_20740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X15968 a_6760_7124# cap_series_gyp a_7568_7608# vss nmos_6p0 w=0.82u l=0.6u
X15969 a_16476_36872# a_16388_36916# vss vss nmos_6p0 w=0.82u l=1u
X15970 vdd a_23308_43144# a_23220_43188# vdd pmos_6p0 w=1.22u l=1u
X15971 vdd a_24652_36872# a_24564_36916# vdd pmos_6p0 w=1.22u l=1u
X15972 vdd tune_series_gy[2] a_11572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X15973 vdd tune_shunt[7] a_9332_11452# vdd pmos_6p0 w=1.2u l=0.5u
X15974 a_9876_18584# cap_shunt_p a_9668_18100# vdd pmos_6p0 w=1.2u l=0.5u
X15975 vdd tune_shunt[6] a_20532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X15976 vss tune_shunt[7] a_28692_29560# vss nmos_6p0 w=0.51u l=0.6u
X15977 a_12788_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15978 vss tune_series_gy[4] a_15700_7970# vss nmos_6p0 w=0.51u l=0.6u
X15979 vdd a_27788_54120# a_27700_54164# vdd pmos_6p0 w=1.22u l=1u
X15980 a_18816_45540# cap_shunt_p a_16708_45602# vss nmos_6p0 w=0.82u l=0.6u
X15981 vdd a_36524_36439# a_36436_36536# vdd pmos_6p0 w=1.22u l=1u
X15982 vdd tune_shunt[7] a_9668_14964# vdd pmos_6p0 w=1.2u l=0.5u
X15983 a_6420_14588# cap_shunt_p a_6628_14242# vdd pmos_6p0 w=1.2u l=0.5u
X15984 a_14784_38968# cap_shunt_n a_13460_38968# vss nmos_6p0 w=0.82u l=0.6u
X15985 a_24660_25218# cap_shunt_p a_24452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X15986 a_18492_54120# a_18404_54164# vss vss nmos_6p0 w=0.82u l=1u
X15987 a_15720_11452# cap_series_gyp a_15532_11452# vdd pmos_6p0 w=1.2u l=0.5u
X15988 a_13588_13020# cap_shunt_p a_13796_12674# vdd pmos_6p0 w=1.2u l=0.5u
X15989 vss tune_shunt[7] a_28692_26424# vss nmos_6p0 w=0.51u l=0.6u
X15990 a_4492_5079# a_4404_5176# vss vss nmos_6p0 w=0.82u l=1u
X15991 a_12788_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X15992 vdd tune_shunt[6] a_25572_33780# vdd pmos_6p0 w=1.2u l=0.5u
X15993 vss tune_series_gy[3] a_15700_4834# vss nmos_6p0 w=0.51u l=0.6u
X15994 vdd a_27788_50984# a_27700_51028# vdd pmos_6p0 w=1.22u l=1u
X15995 a_18816_42404# cap_shunt_n a_16708_42466# vss nmos_6p0 w=0.82u l=0.6u
X15996 a_21316_3988# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X15997 vdd tune_shunt[7] a_9668_11828# vdd pmos_6p0 w=1.2u l=0.5u
X15998 vss tune_shunt[1] a_1924_3266# vss nmos_6p0 w=0.51u l=0.6u
X15999 vdd tune_shunt[7] a_10340_36916# vdd pmos_6p0 w=1.2u l=0.5u
X16000 a_10492_8316# tune_series_gy[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16001 vdd a_5612_19191# a_5524_19288# vdd pmos_6p0 w=1.22u l=1u
X16002 vdd a_9644_38440# a_9556_38484# vdd pmos_6p0 w=1.22u l=1u
X16003 vdd tune_shunt[7] a_17620_32212# vdd pmos_6p0 w=1.2u l=0.5u
X16004 a_33732_32696# cap_shunt_n a_33524_32212# vdd pmos_6p0 w=1.2u l=0.5u
X16005 a_7748_29922# cap_shunt_n a_8680_29860# vss nmos_6p0 w=0.82u l=0.6u
X16006 a_24660_22082# cap_shunt_p a_24452_22428# vdd pmos_6p0 w=1.2u l=0.5u
X16007 a_2500_19292# cap_shunt_p a_2708_18946# vdd pmos_6p0 w=1.2u l=0.5u
X16008 a_15468_54120# a_15380_54164# vss vss nmos_6p0 w=0.82u l=1u
X16009 a_2500_39676# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16010 vdd tune_shunt[7] a_25572_30644# vdd pmos_6p0 w=1.2u l=0.5u
X16011 a_10660_34626# cap_shunt_n a_10452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X16012 a_16408_9176# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X16013 a_20740_32696# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16014 a_22456_4472# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X16015 a_6740_40536# cap_shunt_n a_6532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X16016 vdd a_9644_35304# a_9556_35348# vdd pmos_6p0 w=1.22u l=1u
X16017 a_7540_34972# cap_shunt_n a_7748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X16018 a_35840_32696# cap_shunt_n a_33732_32696# vss nmos_6p0 w=0.82u l=0.6u
X16019 a_7748_26786# cap_shunt_n a_8680_26724# vss nmos_6p0 w=0.82u l=0.6u
X16020 a_2500_16156# cap_shunt_p a_2708_15810# vdd pmos_6p0 w=1.2u l=0.5u
X16021 a_8008_18584# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16022 a_34396_3944# a_34308_3988# vss vss nmos_6p0 w=0.82u l=1u
X16023 a_10660_31490# cap_shunt_n a_10452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X16024 a_24660_34626# cap_shunt_p a_24452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X16025 a_17828_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16026 a_11592_49944# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16027 a_7540_31836# cap_shunt_n a_7748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X16028 a_2708_47170# cap_shunt_p a_2500_47516# vdd pmos_6p0 w=1.2u l=0.5u
X16029 a_23464_34564# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16030 a_24660_31490# cap_shunt_p a_24452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X16031 a_17828_24856# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16032 vss cap_series_gyp a_16016_4472# vss nmos_6p0 w=0.82u l=0.6u
X16033 a_29384_3612# cap_series_gyn a_29408_3204# vss nmos_6p0 w=0.82u l=0.6u
X16034 a_2708_14242# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X16035 vdd a_29916_45847# a_29828_45944# vdd pmos_6p0 w=1.22u l=1u
X16036 a_35692_24372# cap_series_gygyp a_35880_24372# vdd pmos_6p0 w=1.2u l=0.5u
X16037 a_1692_54120# a_1604_54164# vss vss nmos_6p0 w=0.82u l=1u
X16038 vss tune_shunt[5] a_6292_48738# vss nmos_6p0 w=0.51u l=0.6u
X16039 vdd a_4380_55688# a_4292_55732# vdd pmos_6p0 w=1.22u l=1u
X16040 a_8680_37700# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16041 a_32612_33058# cap_shunt_n a_33544_32996# vss nmos_6p0 w=0.82u l=0.6u
X16042 a_20532_16532# cap_shunt_p a_20740_17016# vdd pmos_6p0 w=1.2u l=0.5u
X16043 a_17372_55688# a_17284_55732# vss vss nmos_6p0 w=0.82u l=1u
X16044 a_23464_31428# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16045 a_2708_11106# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X16046 a_18612_12674# cap_series_gyn a_20328_12612# vss nmos_6p0 w=0.82u l=0.6u
X16047 a_32268_17623# a_32180_17720# vss vss nmos_6p0 w=0.82u l=1u
X16048 a_5544_20152# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16049 a_6196_47516# cap_shunt_p a_6404_47170# vdd pmos_6p0 w=1.2u l=0.5u
X16050 vdd a_29916_42711# a_29828_42808# vdd pmos_6p0 w=1.22u l=1u
X16051 a_16500_17724# cap_shunt_p a_16708_17378# vdd pmos_6p0 w=1.2u l=0.5u
X16052 a_35692_21236# cap_series_gygyp a_35880_21236# vdd pmos_6p0 w=1.2u l=0.5u
X16053 a_13796_18946# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16054 vss tune_shunt[7] a_3828_27992# vss nmos_6p0 w=0.51u l=0.6u
X16055 a_37868_47848# a_37780_47892# vss vss nmos_6p0 w=0.82u l=1u
X16056 a_16252_19624# a_16164_19668# vss vss nmos_6p0 w=0.82u l=1u
X16057 a_6628_14242# cap_shunt_p a_8344_14180# vss nmos_6p0 w=0.82u l=0.6u
X16058 a_9220_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16059 a_14348_55688# a_14260_55732# vss vss nmos_6p0 w=0.82u l=1u
X16060 vdd a_24652_27464# a_24564_27508# vdd pmos_6p0 w=1.22u l=1u
X16061 a_24452_38108# cap_shunt_p a_24660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X16062 a_6060_12919# a_5972_13016# vss vss nmos_6p0 w=0.82u l=1u
X16063 a_24660_18946# cap_series_gyn a_24452_19292# vdd pmos_6p0 w=1.2u l=0.5u
X16064 vss tune_shunt[7] a_3828_24856# vss nmos_6p0 w=0.51u l=0.6u
X16065 a_1924_6402# cap_shunt_n a_1716_6748# vdd pmos_6p0 w=1.2u l=0.5u
X16066 vdd tune_shunt[7] a_6532_25940# vdd pmos_6p0 w=1.2u l=0.5u
X16067 a_18816_36132# cap_shunt_n a_16708_36194# vss nmos_6p0 w=0.82u l=0.6u
X16068 vdd a_36524_27031# a_36436_27128# vdd pmos_6p0 w=1.22u l=1u
X16069 vss cap_shunt_gyn a_36652_48676# vss nmos_6p0 w=0.82u l=0.6u
X16070 a_10548_32696# cap_shunt_n a_10340_32212# vdd pmos_6p0 w=1.2u l=0.5u
X16071 a_20532_25940# cap_shunt_n a_20740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X16072 a_6532_52596# tune_shunt[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16073 a_33544_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16074 a_21540_9884# cap_series_gyp a_21748_9538# vdd pmos_6p0 w=1.2u l=0.5u
X16075 a_24660_15810# cap_series_gyn a_24452_16156# vdd pmos_6p0 w=1.2u l=0.5u
X16076 a_5844_3266# tune_shunt[1] vss vss nmos_6p0 w=0.51u l=0.6u
X16077 vdd a_32156_14920# a_32068_14964# vdd pmos_6p0 w=1.22u l=1u
X16078 vss tune_series_gy[4] a_28692_17016# vss nmos_6p0 w=0.51u l=0.6u
X16079 a_28236_49416# a_28148_49460# vss vss nmos_6p0 w=0.82u l=1u
X16080 vdd tune_shunt[7] a_6532_22804# vdd pmos_6p0 w=1.2u l=0.5u
X16081 vss cap_shunt_p a_8064_13880# vss nmos_6p0 w=0.82u l=0.6u
X16082 a_35904_21720# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X16083 vdd tune_shunt[7] a_25572_24372# vdd pmos_6p0 w=1.2u l=0.5u
X16084 a_1716_7124# cap_shunt_n a_1924_7608# vdd pmos_6p0 w=1.2u l=0.5u
X16085 a_37196_32168# a_37108_32212# vss vss nmos_6p0 w=0.82u l=1u
X16086 vdd a_33948_19624# a_33860_19668# vdd pmos_6p0 w=1.22u l=1u
X16087 vdd tune_series_gy[4] a_28484_14964# vdd pmos_6p0 w=1.2u l=0.5u
X16088 vdd tune_shunt[7] a_13588_34972# vdd pmos_6p0 w=1.2u l=0.5u
X16089 vdd a_9644_29032# a_9556_29076# vdd pmos_6p0 w=1.22u l=1u
X16090 a_3828_27992# cap_shunt_n a_4760_27992# vss nmos_6p0 w=0.82u l=0.6u
X16091 vdd tune_shunt[7] a_10340_27508# vdd pmos_6p0 w=1.2u l=0.5u
X16092 a_20532_22804# cap_shunt_p a_20740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X16093 a_34144_45944# tune_shunt_gy[5] vdd vdd pmos_6p0 w=1.215u l=0.5u
X16094 a_21540_6748# cap_series_gyn a_21748_6402# vdd pmos_6p0 w=1.2u l=0.5u
X16095 a_9332_11452# cap_shunt_p a_9540_11106# vdd pmos_6p0 w=1.2u l=0.5u
X16096 vdd a_32156_11784# a_32068_11828# vdd pmos_6p0 w=1.22u l=1u
X16097 a_30800_13880# cap_series_gyp a_28692_13880# vss nmos_6p0 w=0.82u l=0.6u
X16098 a_28236_46280# a_28148_46324# vss vss nmos_6p0 w=0.82u l=1u
X16099 a_21540_28700# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16100 a_6572_3988# tune_series_gy[1] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16101 a_3620_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16102 vdd tune_shunt[7] a_25572_21236# vdd pmos_6p0 w=1.2u l=0.5u
X16103 a_10660_25218# cap_shunt_n a_10452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X16104 a_20740_23288# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16105 vdd tune_series_gy[4] a_28484_11828# vdd pmos_6p0 w=1.2u l=0.5u
X16106 vss cap_series_gyn a_30920_15748# vss nmos_6p0 w=0.82u l=0.6u
X16107 a_9876_18584# cap_shunt_p a_9668_18100# vdd pmos_6p0 w=1.2u l=0.5u
X16108 a_15356_55255# a_15268_55352# vss vss nmos_6p0 w=0.82u l=1u
X16109 vdd a_31260_47415# a_31172_47512# vdd pmos_6p0 w=1.22u l=1u
X16110 vdd tune_shunt[7] a_13588_31836# vdd pmos_6p0 w=1.2u l=0.5u
X16111 a_3828_24856# cap_shunt_p a_4760_24856# vss nmos_6p0 w=0.82u l=0.6u
X16112 a_4032_45540# cap_shunt_p a_2708_45602# vss nmos_6p0 w=0.82u l=0.6u
X16113 a_34536_8316# cap_series_gygyp a_34348_8316# vdd pmos_6p0 w=1.2u l=0.5u
X16114 a_34144_42808# tune_shunt_gy[4] vdd vdd pmos_6p0 w=1.215u l=0.5u
X16115 a_7540_25564# cap_shunt_n a_7748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X16116 a_30800_10744# cap_series_gyp a_28692_10744# vss nmos_6p0 w=0.82u l=0.6u
X16117 a_23464_28292# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16118 a_17828_18584# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16119 a_33164_39575# a_33076_39672# vss vss nmos_6p0 w=0.82u l=1u
X16120 a_24660_25218# cap_shunt_p a_24452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X16121 a_15720_11452# cap_series_gyp a_15532_11452# vdd pmos_6p0 w=1.2u l=0.5u
X16122 a_13588_13020# cap_shunt_p a_13796_12674# vdd pmos_6p0 w=1.2u l=0.5u
X16123 a_1692_47848# a_1604_47892# vss vss nmos_6p0 w=0.82u l=1u
X16124 a_4032_42404# cap_shunt_p a_2708_42466# vss nmos_6p0 w=0.82u l=0.6u
X16125 vss tune_shunt[7] a_16708_23650# vss nmos_6p0 w=0.51u l=0.6u
X16126 vss tune_shunt[5] a_6852_53442# vss nmos_6p0 w=0.51u l=0.6u
X16127 a_2708_37762# cap_shunt_n a_2500_38108# vdd pmos_6p0 w=1.2u l=0.5u
X16128 vdd a_28124_31735# a_28036_31832# vdd pmos_6p0 w=1.22u l=1u
X16129 a_17828_15448# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16130 a_13776_45240# cap_shunt_n a_11668_45240# vss nmos_6p0 w=0.82u l=0.6u
X16131 a_23464_25156# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16132 a_24660_22082# cap_shunt_p a_24452_22428# vdd pmos_6p0 w=1.2u l=0.5u
X16133 a_3380_49944# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X16134 a_11984_39268# cap_shunt_n a_10660_39330# vss nmos_6p0 w=0.82u l=0.6u
X16135 a_17828_38968# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X16136 a_4760_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16137 a_7540_28700# cap_shunt_n a_7748_28354# vdd pmos_6p0 w=1.2u l=0.5u
X16138 a_19524_10260# cap_series_gyn a_19732_10744# vdd pmos_6p0 w=1.2u l=0.5u
X16139 a_12788_13880# cap_shunt_p a_12580_13396# vdd pmos_6p0 w=1.2u l=0.5u
X16140 a_10660_34626# cap_shunt_n a_10452_34972# vdd pmos_6p0 w=1.2u l=0.5u
X16141 a_12580_47892# cap_shunt_p a_12788_48376# vdd pmos_6p0 w=1.2u l=0.5u
X16142 vss tune_shunt[7] a_16708_20514# vss nmos_6p0 w=0.51u l=0.6u
X16143 a_3828_48376# cap_shunt_p a_5544_48376# vss nmos_6p0 w=0.82u l=0.6u
X16144 a_6740_40536# cap_shunt_n a_6532_40052# vdd pmos_6p0 w=1.2u l=0.5u
X16145 a_8996_52220# cap_shunt_n a_9204_51874# vdd pmos_6p0 w=1.2u l=0.5u
X16146 a_6740_46808# cap_shunt_p a_6532_46324# vdd pmos_6p0 w=1.2u l=0.5u
X16147 a_13776_42104# cap_shunt_n a_11668_42104# vss nmos_6p0 w=0.82u l=0.6u
X16148 vdd a_37980_52552# a_37892_52596# vdd pmos_6p0 w=1.22u l=1u
X16149 a_7540_34972# cap_shunt_n a_7748_34626# vdd pmos_6p0 w=1.2u l=0.5u
X16150 a_10548_34264# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16151 a_36296_9176# cap_series_gygyn a_35880_8692# vss nmos_6p0 w=0.82u l=0.6u
X16152 vdd a_8412_11351# a_8324_11448# vdd pmos_6p0 w=1.22u l=1u
X16153 vdd a_32604_13352# a_32516_13396# vdd pmos_6p0 w=1.22u l=1u
X16154 a_2140_13352# a_2052_13396# vss vss nmos_6p0 w=0.82u l=1u
X16155 vdd a_31260_7080# a_31172_7124# vdd pmos_6p0 w=1.22u l=1u
X16156 a_17620_40052# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16157 a_10660_31490# cap_shunt_n a_10452_31836# vdd pmos_6p0 w=1.2u l=0.5u
X16158 vss tune_shunt[5] a_3380_18584# vss nmos_6p0 w=0.51u l=0.6u
X16159 vss cap_shunt_n a_26768_42404# vss nmos_6p0 w=0.82u l=0.6u
X16160 a_28692_12312# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X16161 a_7540_31836# cap_shunt_n a_7748_31490# vdd pmos_6p0 w=1.2u l=0.5u
X16162 a_10548_31128# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16163 a_19732_7608# tune_series_gy[5] vss vss nmos_6p0 w=0.51u l=0.6u
X16164 a_2140_10216# a_2052_10260# vss vss nmos_6p0 w=0.82u l=1u
X16165 a_25984_43972# cap_shunt_p a_24660_44034# vss nmos_6p0 w=0.82u l=0.6u
X16166 a_28692_37400# cap_shunt_p a_28484_36916# vdd pmos_6p0 w=1.2u l=0.5u
X16167 a_32404_34972# cap_shunt_n a_32612_34626# vdd pmos_6p0 w=1.2u l=0.5u
X16168 vdd a_11884_55255# a_11796_55352# vdd pmos_6p0 w=1.22u l=1u
X16169 vss tune_shunt[7] a_3828_15448# vss nmos_6p0 w=0.51u l=0.6u
X16170 a_25780_35832# cap_shunt_p a_27496_35832# vss nmos_6p0 w=0.82u l=0.6u
X16171 a_7580_8316# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16172 vss cap_series_gyn a_25984_18884# vss nmos_6p0 w=0.82u l=0.6u
X16173 a_30584_3204# cap_series_gyn a_29384_3612# vss nmos_6p0 w=0.82u l=0.6u
X16174 vdd a_22188_55688# a_22100_55732# vdd pmos_6p0 w=1.22u l=1u
X16175 vdd a_15580_52552# a_15492_52596# vdd pmos_6p0 w=1.22u l=1u
X16176 vss tune_shunt[6] a_3828_38968# vss nmos_6p0 w=0.51u l=0.6u
X16177 a_13588_47516# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16178 a_25984_40836# cap_shunt_n a_24660_40898# vss nmos_6p0 w=0.82u l=0.6u
X16179 a_20532_16532# cap_shunt_p a_20740_17016# vdd pmos_6p0 w=1.2u l=0.5u
X16180 a_6532_43188# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16181 a_32404_31836# cap_shunt_n a_32612_31490# vdd pmos_6p0 w=1.2u l=0.5u
X16182 a_3620_19668# cap_shunt_p a_3828_20152# vdd pmos_6p0 w=1.2u l=0.5u
X16183 a_35904_12312# cap_series_gygyp vss vss nmos_6p0 w=0.82u l=0.6u
X16184 vss cap_series_gyn a_25984_15748# vss nmos_6p0 w=0.82u l=0.6u
X16185 a_17808_9476# cap_series_gyn a_15700_9538# vss nmos_6p0 w=0.82u l=0.6u
X16186 a_30616_21236# cap_series_gygyn a_30640_21720# vss nmos_6p0 w=0.82u l=0.6u
X16187 a_20740_43672# cap_shunt_n a_20532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X16188 vss tune_shunt[7] a_13460_27992# vss nmos_6p0 w=0.51u l=0.6u
X16189 vss cap_shunt_p a_14896_13880# vss nmos_6p0 w=0.82u l=0.6u
X16190 vss cap_shunt_n a_15120_37700# vss nmos_6p0 w=0.82u l=0.6u
X16191 a_23856_4772# cap_series_gyp a_21748_4834# vss nmos_6p0 w=0.82u l=0.6u
X16192 a_6740_37400# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X16193 vdd tune_shunt[7] a_13588_25564# vdd pmos_6p0 w=1.2u l=0.5u
X16194 vss tune_shunt[6] a_10660_45602# vss nmos_6p0 w=0.51u l=0.6u
X16195 a_9220_17724# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16196 a_24452_38108# cap_shunt_p a_24660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X16197 a_37420_22327# a_37332_22424# vss vss nmos_6p0 w=0.82u l=1u
X16198 a_11824_7608# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X16199 vss tune_shunt[7] a_13460_24856# vss nmos_6p0 w=0.51u l=0.6u
X16200 a_2724_8692# tune_shunt[3] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16201 a_29492_17724# tune_series_gy[4] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16202 a_24660_18946# cap_series_gyn a_24452_19292# vdd pmos_6p0 w=1.2u l=0.5u
X16203 a_3828_15448# cap_shunt_p a_4760_15448# vss nmos_6p0 w=0.82u l=0.6u
X16204 a_4032_36132# cap_shunt_n a_2708_36194# vss nmos_6p0 w=0.82u l=0.6u
X16205 vdd tune_shunt[7] a_13588_22428# vdd pmos_6p0 w=1.2u l=0.5u
X16206 a_25572_36916# cap_shunt_p a_25780_37400# vdd pmos_6p0 w=1.2u l=0.5u
X16207 a_28484_36916# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16208 a_10548_32696# cap_shunt_n a_10340_32212# vdd pmos_6p0 w=1.2u l=0.5u
X16209 vdd a_9644_55255# a_9556_55352# vdd pmos_6p0 w=1.22u l=1u
X16210 vss tune_shunt[6] a_6404_47170# vss nmos_6p0 w=0.51u l=0.6u
X16211 a_15904_32996# cap_shunt_n a_13796_33058# vss nmos_6p0 w=0.82u l=0.6u
X16212 a_20532_25940# cap_shunt_n a_20740_26424# vdd pmos_6p0 w=1.2u l=0.5u
X16213 vdd a_28124_25463# a_28036_25560# vdd pmos_6p0 w=1.22u l=1u
X16214 a_10452_6748# tune_series_gy[2] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16215 a_15700_4834# cap_series_gyn a_15492_5180# vdd pmos_6p0 w=1.2u l=0.5u
X16216 a_11460_46324# cap_shunt_n a_11668_46808# vdd pmos_6p0 w=1.2u l=0.5u
X16217 a_2708_29922# cap_shunt_n a_2500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X16218 a_15700_4834# cap_series_gyn a_17416_4772# vss nmos_6p0 w=0.82u l=0.6u
X16219 a_24660_15810# cap_series_gyn a_24452_16156# vdd pmos_6p0 w=1.2u l=0.5u
X16220 a_35740_54120# a_35652_54164# vss vss nmos_6p0 w=0.82u l=1u
X16221 a_30632_32996# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16222 a_28692_18584# cap_series_gyp a_28484_18100# vdd pmos_6p0 w=1.2u l=0.5u
X16223 a_4760_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16224 vss cap_shunt_n a_3248_7908# vss nmos_6p0 w=0.82u l=0.6u
X16225 vss cap_shunt_p a_7840_20452# vss nmos_6p0 w=0.82u l=0.6u
X16226 vss tune_shunt[7] a_16708_14242# vss nmos_6p0 w=0.51u l=0.6u
X16227 vdd tune_series_gy[4] a_28484_14964# vdd pmos_6p0 w=1.2u l=0.5u
X16228 a_16708_28354# cap_shunt_n a_16500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X16229 a_20532_22804# cap_shunt_p a_20740_23288# vdd pmos_6p0 w=1.2u l=0.5u
X16230 vdd a_28124_22327# a_28036_22424# vdd pmos_6p0 w=1.22u l=1u
X16231 a_36232_17316# cap_series_gygyn vss vss nmos_6p0 w=0.82u l=0.6u
X16232 a_24660_20514# cap_shunt_p a_24452_20860# vdd pmos_6p0 w=1.2u l=0.5u
X16233 a_10340_38484# tune_shunt[6] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16234 a_34844_25896# a_34756_25940# vss vss nmos_6p0 w=0.82u l=1u
X16235 vdd a_10540_7080# a_10452_7124# vdd pmos_6p0 w=1.22u l=1u
X16236 a_32716_54120# a_32628_54164# vss vss nmos_6p0 w=0.82u l=1u
X16237 a_4760_26424# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16238 a_20664_9176# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X16239 a_10660_25218# cap_shunt_n a_10452_25564# vdd pmos_6p0 w=1.2u l=0.5u
X16240 vss cap_shunt_p a_26768_36132# vss nmos_6p0 w=0.82u l=0.6u
X16241 a_19732_7608# cap_series_gyp a_19524_7124# vdd pmos_6p0 w=1.2u l=0.5u
X16242 vdd tune_series_gy[4] a_28484_11828# vdd pmos_6p0 w=1.2u l=0.5u
X16243 vdd a_37980_43144# a_37892_43188# vdd pmos_6p0 w=1.22u l=1u
X16244 a_13460_37400# cap_shunt_n a_15176_37400# vss nmos_6p0 w=0.82u l=0.6u
X16245 a_7540_25564# cap_shunt_n a_7748_25218# vdd pmos_6p0 w=1.2u l=0.5u
X16246 a_10340_35348# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16247 a_32612_31490# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X16248 vdd a_11436_54120# a_11348_54164# vdd pmos_6p0 w=1.22u l=1u
X16249 vdd a_11884_48983# a_11796_49080# vdd pmos_6p0 w=1.22u l=1u
X16250 vdd tune_series_gy[1] a_6572_3988# vdd pmos_6p0 w=1.2u l=0.5u
X16251 a_6292_17378# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X16252 a_7784_53380# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16253 a_37868_53687# a_37780_53784# vss vss nmos_6p0 w=0.82u l=1u
X16254 a_25780_29560# cap_shunt_p a_27496_29560# vss nmos_6p0 w=0.82u l=0.6u
X16255 vdd a_35292_10216# a_35204_10260# vdd pmos_6p0 w=1.22u l=1u
X16256 a_14112_49944# cap_shunt_n a_12788_49944# vss nmos_6p0 w=0.82u l=0.6u
X16257 a_32268_49416# a_32180_49460# vss vss nmos_6p0 w=0.82u l=1u
X16258 a_6292_51512# cap_shunt_p a_7224_51512# vss nmos_6p0 w=0.82u l=0.6u
X16259 a_17828_26424# cap_shunt_n a_17620_25940# vdd pmos_6p0 w=1.2u l=0.5u
X16260 vdd tune_series_gy[3] a_25572_7124# vdd pmos_6p0 w=1.2u l=0.5u
X16261 a_28692_27992# cap_shunt_p a_28484_27508# vdd pmos_6p0 w=1.2u l=0.5u
X16262 a_34348_8316# cap_series_gygyp a_34536_8316# vdd pmos_6p0 w=1.2u l=0.5u
X16263 a_25984_34564# cap_shunt_p a_24660_34626# vss nmos_6p0 w=0.82u l=0.6u
X16264 a_32404_25564# cap_shunt_p a_32612_25218# vdd pmos_6p0 w=1.2u l=0.5u
X16265 a_18492_53687# a_18404_53784# vss vss nmos_6p0 w=0.82u l=1u
X16266 vdd a_24652_47415# a_24564_47512# vdd pmos_6p0 w=1.22u l=1u
X16267 a_12656_3204# cap_series_gyn a_10548_3266# vss nmos_6p0 w=0.82u l=0.6u
X16268 a_14392_35832# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16269 a_29532_16156# cap_series_gyn a_29720_16156# vdd pmos_6p0 w=1.2u l=0.5u
X16270 vss cap_shunt_p a_7616_50244# vss nmos_6p0 w=0.82u l=0.6u
X16271 a_25780_26424# cap_shunt_p a_27496_26424# vss nmos_6p0 w=0.82u l=0.6u
X16272 a_10452_30268# cap_shunt_n a_10660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X16273 a_11780_6040# cap_series_gyn a_11572_5556# vdd pmos_6p0 w=1.2u l=0.5u
X16274 a_2932_9176# tune_shunt[3] vss vss nmos_6p0 w=0.51u l=0.6u
X16275 a_12788_13880# cap_shunt_p a_12580_13396# vdd pmos_6p0 w=1.2u l=0.5u
X16276 a_13588_38108# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16277 a_17828_23288# cap_shunt_n a_17620_22804# vdd pmos_6p0 w=1.2u l=0.5u
X16278 a_29532_13020# cap_series_gyn a_29720_13020# vdd pmos_6p0 w=1.2u l=0.5u
X16279 vss tune_shunt[3] a_24660_44034# vss nmos_6p0 w=0.51u l=0.6u
X16280 vdd a_23756_43144# a_23668_43188# vdd pmos_6p0 w=1.22u l=1u
X16281 a_10660_31490# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16282 a_25984_31428# cap_shunt_p a_24660_31490# vss nmos_6p0 w=0.82u l=0.6u
X16283 a_26712_27992# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16284 a_7568_6040# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X16285 a_6420_14588# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16286 vdd tune_shunt[7] a_13588_19292# vdd pmos_6p0 w=1.2u l=0.5u
X16287 vss tune_shunt[6] a_10660_39330# vss nmos_6p0 w=0.51u l=0.6u
X16288 vdd a_5612_5079# a_5524_5176# vdd pmos_6p0 w=1.22u l=1u
X16289 a_8064_20152# cap_shunt_p a_6740_20152# vss nmos_6p0 w=0.82u l=0.6u
X16290 vdd a_2588_40008# a_2500_40052# vdd pmos_6p0 w=1.22u l=1u
X16291 a_20740_46808# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X16292 vdd a_35180_31735# a_35092_31832# vdd pmos_6p0 w=1.22u l=1u
X16293 a_28348_41576# a_28260_41620# vss vss nmos_6p0 w=0.82u l=1u
X16294 vss cap_shunt_p a_11648_12612# vss nmos_6p0 w=0.82u l=0.6u
X16295 vdd tune_shunt[6] a_9108_49084# vdd pmos_6p0 w=1.2u l=0.5u
X16296 a_36384_49080# cap_shunt_gyn a_36384_48676# vdd pmos_6p0 w=1.215u l=0.5u
X16297 a_18424_29860# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16298 a_26712_24856# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16299 vss cap_series_gyp a_19936_4772# vss nmos_6p0 w=0.82u l=0.6u
X16300 vdd tune_shunt[7] a_13588_16156# vdd pmos_6p0 w=1.2u l=0.5u
X16301 a_33500_19624# a_33412_19668# vss vss nmos_6p0 w=0.82u l=1u
X16302 a_28236_52119# a_28148_52216# vss vss nmos_6p0 w=0.82u l=1u
X16303 vss tune_shunt[7] a_13796_37762# vss nmos_6p0 w=0.51u l=0.6u
X16304 vdd tune_shunt[4] a_33524_32212# vdd pmos_6p0 w=1.2u l=0.5u
X16305 a_32404_34972# cap_shunt_n a_32612_34626# vdd pmos_6p0 w=1.2u l=0.5u
X16306 vss tune_series_gygy[3] a_34536_9884# vss nmos_6p0 w=0.51u l=0.6u
X16307 vdd a_16252_16488# a_16164_16532# vdd pmos_6p0 w=1.22u l=1u
X16308 a_25572_27508# cap_shunt_p a_25780_27992# vdd pmos_6p0 w=1.2u l=0.5u
X16309 a_18424_26724# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16310 a_12220_55688# a_12132_55732# vss vss nmos_6p0 w=0.82u l=1u
X16311 a_28484_27508# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16312 vss tune_shunt[7] a_13796_34626# vss nmos_6p0 w=0.51u l=0.6u
X16313 a_2708_28354# cap_shunt_n a_2500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X16314 a_6740_53080# cap_shunt_n a_7672_53080# vss nmos_6p0 w=0.82u l=0.6u
X16315 a_3828_13880# tune_shunt[4] vss vss nmos_6p0 w=0.51u l=0.6u
X16316 a_20532_16532# cap_shunt_p a_20740_17016# vdd pmos_6p0 w=1.2u l=0.5u
X16317 a_32404_31836# cap_shunt_n a_32612_31490# vdd pmos_6p0 w=1.2u l=0.5u
X16318 a_15904_23588# cap_shunt_n a_13796_23650# vss nmos_6p0 w=0.82u l=0.6u
X16319 a_2932_12312# cap_shunt_n a_2724_11828# vdd pmos_6p0 w=1.2u l=0.5u
X16320 vdd a_28124_16055# a_28036_16152# vdd pmos_6p0 w=1.22u l=1u
X16321 a_2588_32168# a_2500_32212# vss vss nmos_6p0 w=0.82u l=1u
X16322 a_1692_53687# a_1604_53784# vss vss nmos_6p0 w=0.82u l=1u
X16323 a_10452_38108# cap_shunt_n a_10660_37762# vdd pmos_6p0 w=1.2u l=0.5u
X16324 a_14692_7608# cap_series_gyp a_14484_7124# vdd pmos_6p0 w=1.2u l=0.5u
X16325 a_30632_23588# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16326 a_16500_49084# cap_shunt_p a_16708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X16327 a_32716_47848# a_32628_47892# vss vss nmos_6p0 w=0.82u l=1u
X16328 a_11592_45540# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16329 a_20740_43672# cap_shunt_n a_20532_43188# vdd pmos_6p0 w=1.2u l=0.5u
X16330 vss cap_series_gygyp a_36296_24856# vss nmos_6p0 w=0.82u l=0.6u
X16331 a_21540_20860# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16332 vss tune_shunt[7] a_7748_31490# vss nmos_6p0 w=0.51u l=0.6u
X16333 a_7748_37762# cap_shunt_n a_7540_38108# vdd pmos_6p0 w=1.2u l=0.5u
X16334 a_11460_41620# cap_shunt_n a_11668_42104# vdd pmos_6p0 w=1.2u l=0.5u
X16335 a_24660_11106# cap_series_gyp a_24452_11452# vdd pmos_6p0 w=1.2u l=0.5u
X16336 vdd a_28124_12919# a_28036_13016# vdd pmos_6p0 w=1.22u l=1u
X16337 a_1692_50551# a_1604_50648# vss vss nmos_6p0 w=0.82u l=1u
X16338 vss tune_shunt[6] a_12788_48376# vss nmos_6p0 w=0.51u l=0.6u
X16339 a_10340_29076# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16340 a_8848_46808# cap_shunt_p a_6740_46808# vss nmos_6p0 w=0.82u l=0.6u
X16341 a_21748_29922# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16342 a_34844_16488# a_34756_16532# vss vss nmos_6p0 w=0.82u l=1u
X16343 a_11592_42404# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16344 vss tune_series_gy[4] a_15700_6402# vss nmos_6p0 w=0.51u l=0.6u
X16345 a_20172_20759# a_20084_20856# vss vss nmos_6p0 w=0.82u l=1u
X16346 a_13460_26424# cap_shunt_n a_13252_25940# vdd pmos_6p0 w=1.2u l=0.5u
X16347 a_7748_42466# cap_shunt_n a_7540_42812# vdd pmos_6p0 w=1.2u l=0.5u
X16348 a_32604_55255# a_32516_55352# vss vss nmos_6p0 w=0.82u l=1u
X16349 a_16708_47170# tune_shunt[5] vss vss nmos_6p0 w=0.51u l=0.6u
X16350 a_25572_36916# cap_shunt_p a_25780_37400# vdd pmos_6p0 w=1.2u l=0.5u
X16351 a_6404_22082# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16352 a_5844_10744# cap_shunt_p a_7560_10744# vss nmos_6p0 w=0.82u l=0.6u
X16353 a_24452_42812# cap_shunt_n a_24660_42466# vdd pmos_6p0 w=1.2u l=0.5u
X16354 a_25984_28292# cap_shunt_n a_24660_28354# vss nmos_6p0 w=0.82u l=0.6u
X16355 vdd tune_shunt[7] a_20532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X16356 vdd a_24204_46280# a_24116_46324# vdd pmos_6p0 w=1.22u l=1u
X16357 a_2708_29922# cap_shunt_n a_2500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X16358 a_14392_29560# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16359 a_13460_23288# cap_shunt_n a_13252_22804# vdd pmos_6p0 w=1.2u l=0.5u
X16360 a_34308_5180# cap_series_gygyp a_34516_4834# vdd pmos_6p0 w=1.2u l=0.5u
X16361 vss tune_series_gy[2] a_6760_7124# vss nmos_6p0 w=0.51u l=0.6u
X16362 a_28692_18584# cap_series_gyp a_28484_18100# vdd pmos_6p0 w=1.2u l=0.5u
X16363 a_16708_44034# tune_shunt[6] vss vss nmos_6p0 w=0.51u l=0.6u
X16364 a_22064_32696# cap_shunt_n a_20740_32696# vss nmos_6p0 w=0.82u l=0.6u
X16365 a_11780_4472# tune_series_gy[2] vss vss nmos_6p0 w=0.51u l=0.6u
X16366 a_17828_17016# cap_shunt_p a_17620_16532# vdd pmos_6p0 w=1.2u l=0.5u
X16367 a_13588_30268# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16368 a_25984_25156# cap_shunt_p a_24660_25218# vss nmos_6p0 w=0.82u l=0.6u
X16369 a_28484_3988# cap_series_gyp a_28692_4472# vdd pmos_6p0 w=1.2u l=0.5u
X16370 a_25780_15448# cap_series_gyp a_25572_14964# vdd pmos_6p0 w=1.2u l=0.5u
X16371 a_16708_28354# cap_shunt_n a_16500_28700# vdd pmos_6p0 w=1.2u l=0.5u
X16372 a_33948_5512# a_33860_5556# vss vss nmos_6p0 w=0.82u l=1u
X16373 a_14392_26424# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16374 a_24660_20514# cap_shunt_p a_24452_20860# vdd pmos_6p0 w=1.2u l=0.5u
X16375 a_4816_22020# cap_shunt_p a_2708_22082# vss nmos_6p0 w=0.82u l=0.6u
X16376 a_25780_17016# cap_series_gyp a_27496_17016# vss nmos_6p0 w=0.82u l=0.6u
X16377 vdd a_23308_18056# a_23220_18100# vdd pmos_6p0 w=1.22u l=1u
X16378 vdd a_35180_25463# a_35092_25560# vdd pmos_6p0 w=1.22u l=1u
X16379 vdd a_33052_53687# a_32964_53784# vdd pmos_6p0 w=1.22u l=1u
X16380 a_19276_33303# a_19188_33400# vss vss nmos_6p0 w=0.82u l=1u
X16381 a_35880_3988# cap_series_gygyp a_35692_3988# vdd pmos_6p0 w=1.2u l=0.5u
X16382 vss cap_shunt_n a_5152_38968# vss nmos_6p0 w=0.82u l=0.6u
X16383 a_34308_22428# tune_series_gygy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16384 vdd tune_series_gy[5] a_18404_11452# vdd pmos_6p0 w=1.2u l=0.5u
X16385 a_25780_12312# cap_series_gyp a_25572_11828# vdd pmos_6p0 w=1.2u l=0.5u
X16386 a_26712_18584# cap_series_gyn vss vss nmos_6p0 w=0.82u l=0.6u
X16387 a_14796_55688# a_14708_55732# vss vss nmos_6p0 w=0.82u l=1u
X16388 a_2140_9783# a_2052_9880# vss vss nmos_6p0 w=0.82u l=1u
X16389 a_31624_6748# cap_series_gygyn a_31648_6340# vss nmos_6p0 w=0.82u l=0.6u
X16390 vss cap_shunt_n a_23856_32996# vss nmos_6p0 w=0.82u l=0.6u
X16391 a_35692_10260# cap_series_gygyp a_35880_10260# vdd pmos_6p0 w=1.2u l=0.5u
X16392 a_9332_13020# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16393 vdd a_33052_50551# a_32964_50648# vdd pmos_6p0 w=1.22u l=1u
X16394 a_24204_38440# a_24116_38484# vss vss nmos_6p0 w=0.82u l=1u
X16395 a_6740_20152# cap_shunt_p a_6532_19668# vdd pmos_6p0 w=1.2u l=0.5u
X16396 a_24660_7970# tune_series_gy[4] vss vss nmos_6p0 w=0.51u l=0.6u
X16397 a_26712_15448# cap_series_gyp vss vss nmos_6p0 w=0.82u l=0.6u
X16398 a_9668_16532# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16399 a_19936_37400# cap_shunt_n a_17828_37400# vss nmos_6p0 w=0.82u l=0.6u
X16400 a_3036_35304# a_2948_35348# vss vss nmos_6p0 w=0.82u l=1u
X16401 a_29720_13020# cap_series_gyn a_30528_12612# vss nmos_6p0 w=0.82u l=0.6u
X16402 vdd a_10988_41576# a_10900_41620# vdd pmos_6p0 w=1.22u l=1u
X16403 vss tune_shunt[7] a_13796_28354# vss nmos_6p0 w=0.51u l=0.6u
X16404 a_32404_25564# cap_shunt_p a_32612_25218# vdd pmos_6p0 w=1.2u l=0.5u
X16405 a_28684_49416# a_28596_49460# vss vss nmos_6p0 w=0.82u l=1u
X16406 a_24452_23996# tune_shunt[7] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16407 a_28692_37400# cap_shunt_p a_30408_37400# vss nmos_6p0 w=0.82u l=0.6u
X16408 a_24660_4834# tune_series_gy[3] vss vss nmos_6p0 w=0.51u l=0.6u
X16409 a_29532_16156# cap_series_gyn a_29720_16156# vdd pmos_6p0 w=1.2u l=0.5u
X16410 vdd a_6172_52552# a_6084_52596# vdd pmos_6p0 w=1.22u l=1u
X16411 a_2500_49084# cap_shunt_p a_2708_48738# vdd pmos_6p0 w=1.2u l=0.5u
X16412 a_16708_29922# cap_shunt_n a_16500_30268# vdd pmos_6p0 w=1.2u l=0.5u
X16413 a_18424_17316# cap_shunt_p vss vss nmos_6p0 w=0.82u l=0.6u
X16414 a_10452_30268# cap_shunt_n a_10660_29922# vdd pmos_6p0 w=1.2u l=0.5u
X16415 a_3828_37400# cap_shunt_n a_3620_36916# vdd pmos_6p0 w=1.2u l=0.5u
X16416 vss cap_series_gygyn a_36296_18584# vss nmos_6p0 w=0.82u l=0.6u
X16417 vss tune_shunt[7] a_13796_25218# vss nmos_6p0 w=0.51u l=0.6u
X16418 vss tune_shunt[7] a_9540_14242# vss nmos_6p0 w=0.51u l=0.6u
X16419 vdd a_5612_53687# a_5524_53784# vdd pmos_6p0 w=1.22u l=1u
X16420 a_28684_46280# a_28596_46324# vss vss nmos_6p0 w=0.82u l=1u
X16421 vss tune_shunt[6] a_21748_40898# vss nmos_6p0 w=0.51u l=0.6u
X16422 a_6740_32696# cap_shunt_n a_8456_32696# vss nmos_6p0 w=0.82u l=0.6u
X16423 a_3828_27992# tune_shunt[7] vss vss nmos_6p0 w=0.51u l=0.6u
X16424 a_2588_22760# a_2500_22804# vss vss nmos_6p0 w=0.82u l=1u
X16425 vdd a_17372_3511# a_17284_3608# vdd pmos_6p0 w=1.22u l=1u
X16426 a_36988_48376# cap_shunt_gyp a_36720_48438# vss nmos_6p0 w=0.82u l=0.6u
X16427 vdd a_20060_55688# a_19972_55732# vdd pmos_6p0 w=1.22u l=1u
X16428 a_16708_37762# cap_shunt_n a_17640_37700# vss nmos_6p0 w=0.82u l=0.6u
X16429 a_1924_4472# cap_shunt_p a_1716_3988# vdd pmos_6p0 w=1.2u l=0.5u
X16430 a_21540_11452# tune_series_gy[5] vdd vdd pmos_6p0 w=1.2u l=0.5u
X16431 a_20172_14487# a_20084_14584# vss vss nmos_6p0 w=0.82u l=1u
X16432 a_11592_36132# cap_shunt_n vss vss nmos_6p0 w=0.82u l=0.6u
X16433 vss cap_series_gygyn a_36296_15448# vss nmos_6p0 w=0.82u l=0.6u
X16434 a_21628_52552# a_21540_52596# vss vss nmos_6p0 w=0.82u l=1u
X16435 vss tune_shunt[7] a_9540_11106# vss nmos_6p0 w=0.51u l=0.6u
X16436 a_7748_36194# cap_shunt_n a_7540_36540# vdd pmos_6p0 w=1.2u l=0.5u
X16437 vdd a_5612_50551# a_5524_50648# vdd pmos_6p0 w=1.22u l=1u
X16438 vdd a_19276_48983# a_19188_49080# vdd pmos_6p0 w=1.22u l=1u
X16439 vdd a_24092_3944# a_24004_3988# vdd pmos_6p0 w=1.22u l=1u
C0 cap_shunt_gyn tune_shunt_gy[6] 2.17fF
C1 vdd tune_series_gy[3] 2.07fF
C2 cap_shunt_gyp tune_shunt_gy[5] 3.00fF
C3 cap_shunt_n tune_shunt[4] 7.76fF
C4 cap_shunt_gyp tune_shunt_gy[6] 4.48fF
C5 tune_shunt[5] cap_shunt_n 8.74fF
C6 vdd cap_shunt_p 38.56fF
C7 cap_shunt_n tune_shunt[6] 14.82fF
C8 tune_shunt[5] tune_shunt[4] 4.81fF
C9 cap_shunt_gyp cap_shunt_gyn 6.72fF
C10 tune_shunt[5] tune_shunt[6] 2.89fF
C11 tune_series_gy[2] tune_shunt[1] 2.48fF
C12 vdd cap_series_gyn 10.50fF
C13 cap_series_gyn tune_series_gy[3] 2.31fF
C14 vdd tune_series_gy[4] 4.39fF
C15 vdd cap_series_gyp 10.42fF
C16 cap_series_gyp tune_series_gy[3] 4.18fF
C17 cap_shunt_p cap_series_gyn 4.36fF
C18 vdd cap_series_gygyn 5.16fF
C19 vdd tune_series_gygy[5] 2.30fF
C20 cap_shunt_p cap_series_gyp 3.19fF
C21 vdd tune_series_gygy[4] 2.09fF
C22 vdd cap_series_gygyp 5.97fF
C23 vdd tune_shunt[7] 24.85fF
C24 tune_series_gy[4] cap_series_gyn 6.71fF
C25 cap_shunt_n tune_shunt[1] 2.19fF
C26 cap_shunt_p tune_shunt[7] 29.11fF
C27 cap_series_gyp cap_series_gyn 17.93fF
C28 vdd tune_shunt[3] 3.53fF
C29 cap_series_gyp tune_series_gy[4] 5.67fF
C30 tune_series_gy[3] tune_shunt[0] 2.74fF
C31 vdd tune_shunt_gy[5] 2.06fF
C32 cap_shunt_p tune_shunt[3] 2.56fF
C33 vdd tune_shunt_gy[6] 2.14fF
C34 cap_series_gyn tune_series_gy[0] 2.38fF
C35 vdd cap_shunt_gyn 4.62fF
C36 vdd cap_shunt_n 39.12fF
C37 vdd tune_shunt[4] 5.62fF
C38 vdd tune_shunt[5] 7.34fF
C39 vdd tune_shunt[6] 12.93fF
C40 tune_series_gygy[4] cap_series_gygyn 4.33fF
C41 cap_shunt_n cap_shunt_p 22.81fF
C42 vdd cap_shunt_gyp 4.36fF
C43 cap_shunt_p tune_shunt[4] 10.85fF
C44 cap_series_gygyp cap_series_gygyn 3.46fF
C45 tune_series_gygy[4] tune_series_gygy[5] 6.30fF
C46 vdd tune_series_gy[5] 4.38fF
C47 tune_shunt[5] cap_shunt_p 8.91fF
C48 cap_shunt_p tune_shunt[6] 13.11fF
C49 cap_series_gyp tune_shunt[0] 2.73fF
C50 cap_shunt_n cap_series_gyn 3.24fF
C51 tune_shunt[2] tune_shunt[1] 2.41fF
C52 cap_shunt_n cap_series_gyp 3.85fF
C53 tune_shunt[0] tune_series_gy[0] 2.50fF
C54 cap_series_gyn tune_series_gy[5] 7.53fF
C55 tune_shunt[5] cap_series_gyp 2.45fF
C56 tune_shunt[3] tune_shunt[7] 4.70fF
C57 tune_shunt[6] cap_series_gyp 3.86fF
C58 cap_series_gyp tune_series_gy[5] 5.17fF
C59 cap_shunt_n tune_shunt[7] 26.33fF
C60 tune_shunt[4] tune_shunt[7] 3.17fF
C61 tune_series_gy[3] tune_shunt[1] 2.13fF
C62 tune_shunt[5] tune_shunt[7] 6.88fF
C63 tune_shunt[6] tune_shunt[7] 2.19fF
C64 cap_shunt_n tune_shunt[3] 4.20fF
C65 cap_shunt_gyn tune_shunt_gy[5] 2.79fF
C66 tune_series_gy[0] vss 3.90fF
C67 tune_shunt[1] vss 6.39fF
C68 tune_shunt[0] vss 3.60fF
C69 tune_series_gy[1] vss 6.42fF
C70 tune_series_gygy[2] vss 3.08fF
C71 tune_series_gygy[0] vss 3.67fF
C72 tune_series_gygy[1] vss 3.22fF
C73 tune_series_gy[2] vss 11.90fF
C74 tune_shunt[2] vss 9.66fF
C75 tune_series_gygy[3] vss 6.06fF
C76 tune_series_gy[3] vss 23.53fF
C77 tune_series_gy[5] vss 45.82fF
C78 cap_series_gyn vss 123.37fF
C79 tune_series_gy[4] vss 45.23fF
C80 cap_series_gyp vss 123.52fF
C81 cap_series_gygyn vss 46.65fF
C82 tune_series_gygy[5] vss 23.26fF
C83 tune_series_gygy[4] vss 12.99fF
C84 cap_series_gygyp vss 47.50fF
C85 tune_shunt[7] vss 266.59fF
C86 tune_shunt_gy[1] vss 2.65fF
C87 tune_shunt_gy[2] vss 2.32fF
C88 tune_shunt[3] vss 18.17fF
C89 tune_shunt_gy[3] vss 4.25fF
C90 tune_shunt_gy[5] vss 8.46fF
C91 tune_shunt_gy[6] vss 8.37fF
C92 cap_shunt_gyn vss 22.70fF
C93 tune_shunt[4] vss 36.00fF
C94 tune_shunt[6] vss 132.42fF
C95 cap_shunt_gyp vss 22.67fF
C96 tune_shunt_gy[4] vss 4.36fF
C97 cap_shunt_p vss 487.66fF
C98 cap_shunt_n vss 490.19fF
C99 tune_shunt[5] vss 67.15fF
C100 vdd vss 3407.22fF
.ends
