* NGSPICE file created from aoi21_flat.ext - technology: gf180mcuC

.subckt aoi21_flat A1 A2 B ZN VDD VSS
X0 VDD B a_36_472# VDD pmos_6p0 w=1.215u l=0.5u
X1 ZN A2 a_36_472# VDD pmos_6p0 w=1.215u l=0.5u
X2 a_36_472# A1 ZN VDD pmos_6p0 w=1.215u l=0.5u
X3 VSS B ZN VSS nmos_6p0 w=0.51u l=0.6u
X4 ZN A1 a_244_68# VSS nmos_6p0 w=0.82u l=0.6u
X5 a_244_68# A2 VSS VSS nmos_6p0 w=0.82u l=0.6u
.ends
