magic
tech gf180mcuC
magscale 1 10
timestamp 1669581515
<< nwell >>
rect -419 1180 -15 2768
rect -419 349 -15 817
<< pwell >>
rect -419 2768 -15 3122
rect -419 819 -16 1180
rect -419 817 -15 819
rect -419 -137 -15 349
<< nmos >>
rect -332 2942 -172 2998
rect -245 904 -189 1064
rect -332 119 -172 175
<< pmos >>
rect -245 1358 -189 2638
rect -245 479 -189 639
<< ndiff >>
rect -332 3073 -172 3086
rect -332 3027 -319 3073
rect -185 3027 -172 3073
rect -332 2998 -172 3027
rect -332 2913 -172 2942
rect -332 2867 -319 2913
rect -185 2867 -172 2913
rect -332 2854 -172 2867
rect -333 1051 -245 1064
rect -333 917 -320 1051
rect -274 917 -245 1051
rect -333 904 -245 917
rect -189 1051 -101 1064
rect -189 917 -160 1051
rect -114 917 -101 1051
rect -189 904 -101 917
rect -332 250 -172 263
rect -332 204 -319 250
rect -185 204 -172 250
rect -332 175 -172 204
rect -332 90 -172 119
rect -332 44 -319 90
rect -185 44 -172 90
rect -332 31 -172 44
<< pdiff >>
rect -333 2625 -245 2638
rect -333 1371 -320 2625
rect -274 1371 -245 2625
rect -333 1358 -245 1371
rect -189 2625 -101 2638
rect -189 1371 -160 2625
rect -114 1371 -101 2625
rect -189 1358 -101 1371
rect -333 626 -245 639
rect -333 492 -320 626
rect -274 492 -245 626
rect -333 479 -245 492
rect -189 626 -101 639
rect -189 492 -160 626
rect -114 492 -101 626
rect -189 479 -101 492
<< ndiffc >>
rect -319 3027 -185 3073
rect -319 2867 -185 2913
rect -320 917 -274 1051
rect -160 917 -114 1051
rect -319 204 -185 250
rect -319 44 -185 90
<< pdiffc >>
rect -320 1371 -274 2625
rect -160 1371 -114 2625
rect -320 492 -274 626
rect -160 492 -114 626
<< psubdiff >>
rect -395 -48 -59 -35
rect -395 -94 -375 -48
rect -79 -94 -59 -48
rect -395 -107 -59 -94
<< psubdiffcont >>
rect -375 -94 -79 -48
<< polysilicon >>
rect -141 2998 -69 3006
rect -376 2942 -332 2998
rect -172 2993 -69 2998
rect -172 2947 -128 2993
rect -82 2947 -69 2993
rect -172 2942 -69 2947
rect -141 2934 -69 2942
rect -253 2728 -181 2741
rect -253 2682 -240 2728
rect -194 2682 -181 2728
rect -253 2669 -181 2682
rect -245 2638 -189 2669
rect -245 1327 -189 1358
rect -253 1314 -181 1327
rect -253 1268 -240 1314
rect -194 1268 -181 1314
rect -253 1255 -181 1268
rect -253 1154 -181 1167
rect -253 1108 -240 1154
rect -194 1108 -181 1154
rect -253 1095 -181 1108
rect -245 1064 -189 1095
rect -245 860 -189 904
rect -253 729 -181 742
rect -253 683 -240 729
rect -194 683 -181 729
rect -253 670 -181 683
rect -245 639 -189 670
rect -245 435 -189 479
rect -141 175 -69 183
rect -376 119 -332 175
rect -172 170 -69 175
rect -172 124 -128 170
rect -82 124 -69 170
rect -172 119 -69 124
rect -141 111 -69 119
<< polycontact >>
rect -128 2947 -82 2993
rect -240 2682 -194 2728
rect -240 1268 -194 1314
rect -240 1108 -194 1154
rect -240 683 -194 729
rect -128 124 -82 170
<< metal1 >>
rect -372 3085 -174 3087
rect -372 3029 -360 3085
rect -304 3073 -252 3085
rect -196 3073 -174 3085
rect -372 3027 -319 3029
rect -185 3027 -174 3073
rect -128 3070 -68 3082
rect -128 3014 -126 3070
rect -70 3014 -68 3070
rect -128 2993 -68 3014
rect -82 2962 -68 2993
rect -330 2867 -319 2913
rect -185 2867 -174 2913
rect -128 2906 -126 2947
rect -70 2906 -68 2962
rect -128 2894 -68 2906
rect -330 2848 -174 2867
rect -330 2788 -8 2848
rect -312 2740 -124 2742
rect -312 2684 -300 2740
rect -244 2728 -192 2740
rect -244 2684 -240 2728
rect -312 2682 -240 2684
rect -194 2684 -192 2728
rect -136 2684 -124 2740
rect -194 2682 -124 2684
rect -320 2625 -114 2636
rect -274 2576 -160 2625
rect -274 2511 -260 2576
rect -262 2455 -260 2511
rect -274 2403 -260 2455
rect -262 2381 -260 2403
rect -262 2347 -160 2381
rect -274 2321 -160 2347
rect -274 2295 -260 2321
rect -262 2239 -260 2295
rect -274 2187 -260 2239
rect -262 2141 -260 2187
rect -262 2131 -160 2141
rect -274 2081 -160 2131
rect -274 2079 -260 2081
rect -262 2023 -260 2079
rect -274 1971 -260 2023
rect -262 1915 -260 1971
rect -274 1901 -260 1915
rect -274 1863 -160 1901
rect -262 1841 -160 1863
rect -262 1807 -260 1841
rect -274 1755 -260 1807
rect -262 1699 -260 1755
rect -274 1661 -260 1699
rect -274 1647 -160 1661
rect -262 1601 -160 1647
rect -262 1591 -260 1601
rect -274 1539 -260 1591
rect -262 1483 -260 1539
rect -274 1420 -260 1483
rect -274 1371 -160 1420
rect -320 1360 -114 1371
rect -312 1312 -240 1314
rect -312 1256 -300 1312
rect -244 1268 -240 1312
rect -194 1312 -124 1314
rect -194 1268 -192 1312
rect -244 1256 -192 1268
rect -136 1256 -124 1312
rect -312 1254 -124 1256
rect -311 1166 -123 1168
rect -311 1110 -299 1166
rect -243 1154 -191 1166
rect -243 1110 -240 1154
rect -311 1108 -240 1110
rect -194 1110 -191 1154
rect -135 1110 -123 1166
rect -194 1108 -123 1110
rect -68 1062 -8 2788
rect -320 1051 -274 1062
rect -320 907 -274 917
rect -426 847 -274 907
rect -160 1051 -8 1062
rect -114 1002 -8 1051
rect -114 917 -105 1002
rect -160 906 -105 917
rect -426 349 -366 847
rect -311 741 -123 743
rect -311 685 -299 741
rect -243 729 -191 741
rect -243 685 -240 729
rect -311 683 -240 685
rect -194 685 -191 729
rect -135 685 -123 741
rect -194 683 -123 685
rect -320 626 -274 637
rect -168 626 -114 637
rect -274 614 -260 626
rect -262 558 -260 614
rect -274 506 -260 558
rect -320 450 -318 492
rect -262 450 -260 506
rect -320 438 -260 450
rect -168 614 -160 626
rect -114 614 -108 626
rect -168 558 -166 614
rect -110 558 -108 614
rect -168 506 -160 558
rect -114 506 -108 558
rect -168 450 -166 506
rect -110 450 -108 506
rect -168 438 -108 450
rect -426 296 -174 349
rect -330 250 -174 296
rect -330 204 -319 250
rect -185 204 -174 250
rect -128 229 -68 241
rect -128 173 -126 229
rect -70 173 -68 229
rect -128 170 -68 173
rect -82 124 -68 170
rect -128 121 -68 124
rect -372 88 -319 90
rect -372 32 -360 88
rect -185 44 -174 90
rect -128 65 -126 121
rect -70 65 -68 121
rect -128 53 -68 65
rect -304 32 -252 44
rect -196 32 -174 44
rect -372 30 -174 32
rect -386 -94 -375 -48
rect -79 -94 -68 -48
<< via1 >>
rect -360 3073 -304 3085
rect -252 3073 -196 3085
rect -360 3029 -319 3073
rect -319 3029 -304 3073
rect -252 3029 -196 3073
rect -126 3014 -70 3070
rect -126 2947 -82 2962
rect -82 2947 -70 2962
rect -126 2906 -70 2947
rect -300 2684 -244 2740
rect -192 2684 -136 2740
rect -318 2455 -274 2511
rect -274 2455 -262 2511
rect -318 2347 -274 2403
rect -274 2347 -262 2403
rect -318 2239 -274 2295
rect -274 2239 -262 2295
rect -318 2131 -274 2187
rect -274 2131 -262 2187
rect -318 2023 -274 2079
rect -274 2023 -262 2079
rect -318 1915 -274 1971
rect -274 1915 -262 1971
rect -318 1807 -274 1863
rect -274 1807 -262 1863
rect -318 1699 -274 1755
rect -274 1699 -262 1755
rect -318 1591 -274 1647
rect -274 1591 -262 1647
rect -318 1483 -274 1539
rect -274 1483 -262 1539
rect -300 1256 -244 1312
rect -192 1256 -136 1312
rect -299 1110 -243 1166
rect -191 1110 -135 1166
rect -299 685 -243 741
rect -191 685 -135 741
rect -318 558 -274 614
rect -274 558 -262 614
rect -318 492 -274 506
rect -274 492 -262 506
rect -318 450 -262 492
rect -166 558 -160 614
rect -160 558 -114 614
rect -114 558 -110 614
rect -166 492 -160 506
rect -160 492 -114 506
rect -114 492 -110 506
rect -166 450 -110 492
rect -126 173 -70 229
rect -360 44 -319 88
rect -319 44 -304 88
rect -252 44 -196 88
rect -126 65 -70 121
rect -360 32 -304 44
rect -252 32 -196 44
<< metal2 >>
rect -372 3085 -184 3147
rect -372 3029 -360 3085
rect -304 3029 -252 3085
rect -196 3029 -184 3085
rect -372 3027 -184 3029
rect -128 3070 -68 3082
rect -128 3014 -126 3070
rect -70 3014 -68 3070
rect -128 3006 -68 3014
rect -128 2962 -56 3006
rect -128 2906 -126 2962
rect -70 2934 -56 2962
rect -70 2906 -68 2934
rect -128 2894 -68 2906
rect -312 2740 -124 2742
rect -312 2684 -300 2740
rect -244 2684 -192 2740
rect -136 2684 -124 2740
rect -312 2682 -124 2684
rect -320 2511 -260 2523
rect -320 2455 -318 2511
rect -262 2455 -260 2511
rect -320 2403 -260 2455
rect -320 2347 -318 2403
rect -262 2347 -260 2403
rect -320 2295 -260 2347
rect -320 2239 -318 2295
rect -262 2239 -260 2295
rect -320 2187 -260 2239
rect -320 2131 -318 2187
rect -262 2131 -260 2187
rect -320 2079 -260 2131
rect -320 2023 -318 2079
rect -262 2023 -260 2079
rect -320 1971 -260 2023
rect -320 1915 -318 1971
rect -262 1915 -260 1971
rect -320 1863 -260 1915
rect -320 1807 -318 1863
rect -262 1807 -260 1863
rect -320 1755 -260 1807
rect -320 1699 -318 1755
rect -262 1699 -260 1755
rect -320 1647 -260 1699
rect -320 1591 -318 1647
rect -262 1591 -260 1647
rect -320 1539 -260 1591
rect -320 1483 -318 1539
rect -262 1483 -260 1539
rect -320 1471 -260 1483
rect -196 1314 -124 2682
rect -312 1312 -124 1314
rect -312 1256 -300 1312
rect -244 1256 -192 1312
rect -136 1256 -124 1312
rect -312 1254 -124 1256
rect -253 1168 -181 1254
rect -311 1166 -123 1168
rect -311 1110 -299 1166
rect -243 1110 -191 1166
rect -135 1110 -123 1166
rect -311 1108 -123 1110
rect -253 743 -181 1108
rect -311 741 -123 743
rect -311 685 -299 741
rect -243 685 -191 741
rect -135 685 -123 741
rect -311 683 -123 685
rect -320 614 -260 626
rect -320 558 -318 614
rect -262 558 -260 614
rect -320 506 -260 558
rect -320 450 -318 506
rect -262 450 -260 506
rect -320 438 -260 450
rect -168 614 -108 626
rect -168 558 -166 614
rect -110 558 -108 614
rect -168 506 -108 558
rect -168 450 -166 506
rect -110 450 -108 506
rect -168 438 -108 450
rect -128 229 -68 241
rect -128 173 -126 229
rect -70 183 -68 229
rect -70 173 -56 183
rect -128 121 -56 173
rect -372 88 -184 90
rect -372 32 -360 88
rect -304 32 -252 88
rect -196 32 -184 88
rect -128 65 -126 121
rect -70 111 -56 121
rect -70 65 -68 111
rect -128 53 -68 65
rect -372 -30 -184 32
<< via2 >>
rect -126 3014 -70 3070
rect -126 2906 -70 2962
rect -318 2131 -262 2187
rect -318 2023 -262 2079
rect -318 1915 -262 1971
rect -318 1807 -262 1863
rect -318 558 -262 614
rect -318 450 -262 506
rect -166 558 -110 614
rect -166 450 -110 506
rect -126 173 -70 229
rect -126 65 -70 121
<< metal3 >>
rect -419 3070 -15 3082
rect -419 3014 -126 3070
rect -70 3014 -15 3070
rect -419 2962 -15 3014
rect -419 2906 -126 2962
rect -70 2906 -15 2962
rect -419 2894 -15 2906
rect -419 2187 -15 2197
rect -419 2131 -318 2187
rect -262 2131 -15 2187
rect -419 2079 -15 2131
rect -419 2023 -318 2079
rect -262 2023 -15 2079
rect -419 1971 -15 2023
rect -419 1915 -318 1971
rect -262 1915 -15 1971
rect -419 1863 -15 1915
rect -419 1807 -318 1863
rect -262 1807 -15 1863
rect -419 1797 -15 1807
rect -426 614 -15 626
rect -426 558 -318 614
rect -262 558 -166 614
rect -110 558 -15 614
rect -426 506 -15 558
rect -426 450 -318 506
rect -262 450 -166 506
rect -110 450 -15 506
rect -426 438 -15 450
rect -419 229 -15 241
rect -419 173 -126 229
rect -70 173 -15 229
rect -419 121 -15 173
rect -419 65 -126 121
rect -70 65 -15 121
rect -419 53 -15 65
rect -373 35 -172 53
<< comment >>
rect -217 706 -216 2742
<< end >>
