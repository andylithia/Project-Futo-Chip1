magic
tech gf180mcuC
magscale 1 10
timestamp 1670231070
<< metal1 >>
rect 111570 6638 111582 6690
rect 111634 6687 111646 6690
rect 112130 6687 112142 6690
rect 111634 6641 112142 6687
rect 111634 6638 111646 6641
rect 112130 6638 112142 6641
rect 112194 6638 112206 6690
rect 1344 6298 159092 6332
rect 1344 6246 40196 6298
rect 40248 6246 40320 6298
rect 40372 6246 40444 6298
rect 40496 6246 40568 6298
rect 40620 6246 40692 6298
rect 40744 6246 40816 6298
rect 40868 6246 40940 6298
rect 40992 6246 41064 6298
rect 41116 6246 79508 6298
rect 79560 6246 79632 6298
rect 79684 6246 79756 6298
rect 79808 6246 79880 6298
rect 79932 6246 80004 6298
rect 80056 6246 80128 6298
rect 80180 6246 80252 6298
rect 80304 6246 80376 6298
rect 80428 6246 118820 6298
rect 118872 6246 118944 6298
rect 118996 6246 119068 6298
rect 119120 6246 119192 6298
rect 119244 6246 119316 6298
rect 119368 6246 119440 6298
rect 119492 6246 119564 6298
rect 119616 6246 119688 6298
rect 119740 6246 158132 6298
rect 158184 6246 158256 6298
rect 158308 6246 158380 6298
rect 158432 6246 158504 6298
rect 158556 6246 158628 6298
rect 158680 6246 158752 6298
rect 158804 6246 158876 6298
rect 158928 6246 159000 6298
rect 159052 6246 159092 6298
rect 1344 6212 159092 6246
rect 10658 5966 10670 6018
rect 10722 5966 10734 6018
rect 2146 5854 2158 5906
rect 2210 5854 2222 5906
rect 8866 5854 8878 5906
rect 8930 5854 8942 5906
rect 9986 5854 9998 5906
rect 10050 5854 10062 5906
rect 13906 5854 13918 5906
rect 13970 5854 13982 5906
rect 17826 5854 17838 5906
rect 17890 5854 17902 5906
rect 21634 5854 21646 5906
rect 21698 5854 21710 5906
rect 25554 5854 25566 5906
rect 25618 5854 25630 5906
rect 29474 5854 29486 5906
rect 29538 5854 29550 5906
rect 33506 5854 33518 5906
rect 33570 5854 33582 5906
rect 37314 5854 37326 5906
rect 37378 5854 37390 5906
rect 41346 5854 41358 5906
rect 41410 5854 41422 5906
rect 45266 5854 45278 5906
rect 45330 5854 45342 5906
rect 49074 5854 49086 5906
rect 49138 5854 49150 5906
rect 52994 5854 53006 5906
rect 53058 5854 53070 5906
rect 57026 5854 57038 5906
rect 57090 5854 57102 5906
rect 60834 5854 60846 5906
rect 60898 5854 60910 5906
rect 64754 5854 64766 5906
rect 64818 5854 64830 5906
rect 68674 5854 68686 5906
rect 68738 5854 68750 5906
rect 72594 5854 72606 5906
rect 72658 5854 72670 5906
rect 76626 5854 76638 5906
rect 76690 5854 76702 5906
rect 80322 5854 80334 5906
rect 80386 5854 80398 5906
rect 84130 5854 84142 5906
rect 84194 5854 84206 5906
rect 90962 5854 90974 5906
rect 91026 5854 91038 5906
rect 94882 5854 94894 5906
rect 94946 5854 94958 5906
rect 98802 5854 98814 5906
rect 98866 5854 98878 5906
rect 102722 5854 102734 5906
rect 102786 5854 102798 5906
rect 103954 5854 103966 5906
rect 104018 5854 104030 5906
rect 110562 5854 110574 5906
rect 110626 5854 110638 5906
rect 114370 5854 114382 5906
rect 114434 5854 114446 5906
rect 115602 5854 115614 5906
rect 115666 5854 115678 5906
rect 119522 5854 119534 5906
rect 119586 5854 119598 5906
rect 120194 5854 120206 5906
rect 120258 5854 120270 5906
rect 123330 5854 123342 5906
rect 123394 5854 123406 5906
rect 127250 5854 127262 5906
rect 127314 5854 127326 5906
rect 131282 5854 131294 5906
rect 131346 5854 131358 5906
rect 135090 5854 135102 5906
rect 135154 5854 135166 5906
rect 139010 5854 139022 5906
rect 139074 5854 139086 5906
rect 145730 5854 145742 5906
rect 145794 5854 145806 5906
rect 2818 5742 2830 5794
rect 2882 5742 2894 5794
rect 4946 5742 4958 5794
rect 5010 5742 5022 5794
rect 5954 5742 5966 5794
rect 6018 5742 6030 5794
rect 8082 5742 8094 5794
rect 8146 5742 8158 5794
rect 12786 5742 12798 5794
rect 12850 5742 12862 5794
rect 14578 5742 14590 5794
rect 14642 5742 14654 5794
rect 16706 5742 16718 5794
rect 16770 5742 16782 5794
rect 18498 5742 18510 5794
rect 18562 5742 18574 5794
rect 20626 5742 20638 5794
rect 20690 5742 20702 5794
rect 22418 5742 22430 5794
rect 22482 5742 22494 5794
rect 24546 5742 24558 5794
rect 24610 5742 24622 5794
rect 26338 5742 26350 5794
rect 26402 5742 26414 5794
rect 28466 5742 28478 5794
rect 28530 5742 28542 5794
rect 30258 5742 30270 5794
rect 30322 5742 30334 5794
rect 32386 5742 32398 5794
rect 32450 5742 32462 5794
rect 34178 5742 34190 5794
rect 34242 5742 34254 5794
rect 36306 5742 36318 5794
rect 36370 5742 36382 5794
rect 38098 5742 38110 5794
rect 38162 5742 38174 5794
rect 40226 5742 40238 5794
rect 40290 5742 40302 5794
rect 42018 5742 42030 5794
rect 42082 5742 42094 5794
rect 44146 5742 44158 5794
rect 44210 5742 44222 5794
rect 45938 5742 45950 5794
rect 46002 5742 46014 5794
rect 48066 5742 48078 5794
rect 48130 5742 48142 5794
rect 49858 5742 49870 5794
rect 49922 5742 49934 5794
rect 51986 5742 51998 5794
rect 52050 5742 52062 5794
rect 53778 5742 53790 5794
rect 53842 5742 53854 5794
rect 55906 5742 55918 5794
rect 55970 5742 55982 5794
rect 57698 5742 57710 5794
rect 57762 5742 57774 5794
rect 59826 5742 59838 5794
rect 59890 5742 59902 5794
rect 61618 5742 61630 5794
rect 61682 5742 61694 5794
rect 63746 5742 63758 5794
rect 63810 5742 63822 5794
rect 65538 5742 65550 5794
rect 65602 5742 65614 5794
rect 67666 5742 67678 5794
rect 67730 5742 67742 5794
rect 69458 5742 69470 5794
rect 69522 5742 69534 5794
rect 71586 5742 71598 5794
rect 71650 5742 71662 5794
rect 73378 5742 73390 5794
rect 73442 5742 73454 5794
rect 75506 5742 75518 5794
rect 75570 5742 75582 5794
rect 77298 5742 77310 5794
rect 77362 5742 77374 5794
rect 79426 5742 79438 5794
rect 79490 5742 79502 5794
rect 80994 5742 81006 5794
rect 81058 5742 81070 5794
rect 83122 5742 83134 5794
rect 83186 5742 83198 5794
rect 84914 5742 84926 5794
rect 84978 5742 84990 5794
rect 87042 5742 87054 5794
rect 87106 5742 87118 5794
rect 88050 5742 88062 5794
rect 88114 5742 88126 5794
rect 90178 5742 90190 5794
rect 90242 5742 90254 5794
rect 91970 5742 91982 5794
rect 92034 5742 92046 5794
rect 94098 5742 94110 5794
rect 94162 5742 94174 5794
rect 95890 5742 95902 5794
rect 95954 5742 95966 5794
rect 98018 5742 98030 5794
rect 98082 5742 98094 5794
rect 99810 5742 99822 5794
rect 99874 5742 99886 5794
rect 101938 5742 101950 5794
rect 102002 5742 102014 5794
rect 104738 5742 104750 5794
rect 104802 5742 104814 5794
rect 106866 5742 106878 5794
rect 106930 5742 106942 5794
rect 107650 5742 107662 5794
rect 107714 5742 107726 5794
rect 109778 5742 109790 5794
rect 109842 5742 109854 5794
rect 111570 5742 111582 5794
rect 111634 5742 111646 5794
rect 113698 5742 113710 5794
rect 113762 5742 113774 5794
rect 116274 5742 116286 5794
rect 116338 5742 116350 5794
rect 118402 5742 118414 5794
rect 118466 5742 118478 5794
rect 122322 5742 122334 5794
rect 122386 5742 122398 5794
rect 124114 5742 124126 5794
rect 124178 5742 124190 5794
rect 126242 5742 126254 5794
rect 126306 5742 126318 5794
rect 128034 5742 128046 5794
rect 128098 5742 128110 5794
rect 130162 5742 130174 5794
rect 130226 5742 130238 5794
rect 131954 5742 131966 5794
rect 132018 5742 132030 5794
rect 134082 5742 134094 5794
rect 134146 5742 134158 5794
rect 135874 5742 135886 5794
rect 135938 5742 135950 5794
rect 138002 5742 138014 5794
rect 138066 5742 138078 5794
rect 139794 5742 139806 5794
rect 139858 5742 139870 5794
rect 141922 5742 141934 5794
rect 141986 5742 141998 5794
rect 142930 5742 142942 5794
rect 142994 5742 143006 5794
rect 145058 5742 145070 5794
rect 145122 5742 145134 5794
rect 1344 5514 158592 5548
rect 1344 5462 20540 5514
rect 20592 5462 20664 5514
rect 20716 5462 20788 5514
rect 20840 5462 20912 5514
rect 20964 5462 21036 5514
rect 21088 5462 21160 5514
rect 21212 5462 21284 5514
rect 21336 5462 21408 5514
rect 21460 5462 59852 5514
rect 59904 5462 59976 5514
rect 60028 5462 60100 5514
rect 60152 5462 60224 5514
rect 60276 5462 60348 5514
rect 60400 5462 60472 5514
rect 60524 5462 60596 5514
rect 60648 5462 60720 5514
rect 60772 5462 99164 5514
rect 99216 5462 99288 5514
rect 99340 5462 99412 5514
rect 99464 5462 99536 5514
rect 99588 5462 99660 5514
rect 99712 5462 99784 5514
rect 99836 5462 99908 5514
rect 99960 5462 100032 5514
rect 100084 5462 138476 5514
rect 138528 5462 138600 5514
rect 138652 5462 138724 5514
rect 138776 5462 138848 5514
rect 138900 5462 138972 5514
rect 139024 5462 139096 5514
rect 139148 5462 139220 5514
rect 139272 5462 139344 5514
rect 139396 5462 158592 5514
rect 1344 5428 158592 5462
rect 2818 5182 2830 5234
rect 2882 5182 2894 5234
rect 4946 5182 4958 5234
rect 5010 5182 5022 5234
rect 9426 5182 9438 5234
rect 9490 5182 9502 5234
rect 10770 5182 10782 5234
rect 10834 5182 10846 5234
rect 12898 5182 12910 5234
rect 12962 5182 12974 5234
rect 14690 5182 14702 5234
rect 14754 5182 14766 5234
rect 16818 5182 16830 5234
rect 16882 5182 16894 5234
rect 20850 5182 20862 5234
rect 20914 5182 20926 5234
rect 23202 5182 23214 5234
rect 23266 5182 23278 5234
rect 25330 5182 25342 5234
rect 25394 5182 25406 5234
rect 28802 5182 28814 5234
rect 28866 5182 28878 5234
rect 33282 5182 33294 5234
rect 33346 5182 33358 5234
rect 34626 5182 34638 5234
rect 34690 5182 34702 5234
rect 36754 5182 36766 5234
rect 36818 5182 36830 5234
rect 39106 5182 39118 5234
rect 39170 5182 39182 5234
rect 41234 5182 41246 5234
rect 41298 5182 41310 5234
rect 42578 5182 42590 5234
rect 42642 5182 42654 5234
rect 44706 5182 44718 5234
rect 44770 5182 44782 5234
rect 49186 5182 49198 5234
rect 49250 5182 49262 5234
rect 50530 5182 50542 5234
rect 50594 5182 50606 5234
rect 52658 5182 52670 5234
rect 52722 5182 52734 5234
rect 55570 5182 55582 5234
rect 55634 5182 55646 5234
rect 70130 5182 70142 5234
rect 70194 5182 70206 5234
rect 72258 5182 72270 5234
rect 72322 5182 72334 5234
rect 74386 5182 74398 5234
rect 74450 5182 74462 5234
rect 76514 5182 76526 5234
rect 76578 5182 76590 5234
rect 82226 5182 82238 5234
rect 82290 5182 82302 5234
rect 93202 5182 93214 5234
rect 93266 5182 93278 5234
rect 99586 5182 99598 5234
rect 99650 5182 99662 5234
rect 103282 5182 103294 5234
rect 103346 5182 103358 5234
rect 105410 5182 105422 5234
rect 105474 5182 105486 5234
rect 109106 5182 109118 5234
rect 109170 5182 109182 5234
rect 111234 5182 111246 5234
rect 111298 5182 111310 5234
rect 113362 5182 113374 5234
rect 113426 5182 113438 5234
rect 115490 5182 115502 5234
rect 115554 5182 115566 5234
rect 117842 5182 117854 5234
rect 117906 5182 117918 5234
rect 119970 5182 119982 5234
rect 120034 5182 120046 5234
rect 121314 5182 121326 5234
rect 121378 5182 121390 5234
rect 123442 5182 123454 5234
rect 123506 5182 123518 5234
rect 125010 5182 125022 5234
rect 125074 5182 125086 5234
rect 127138 5182 127150 5234
rect 127202 5182 127214 5234
rect 128482 5182 128494 5234
rect 128546 5182 128558 5234
rect 135874 5182 135886 5234
rect 135938 5182 135950 5234
rect 139346 5182 139358 5234
rect 139410 5182 139422 5234
rect 140914 5182 140926 5234
rect 140978 5182 140990 5234
rect 143042 5182 143054 5234
rect 143106 5182 143118 5234
rect 147298 5182 147310 5234
rect 147362 5182 147374 5234
rect 2034 5070 2046 5122
rect 2098 5070 2110 5122
rect 6514 5070 6526 5122
rect 6578 5070 6590 5122
rect 7298 5070 7310 5122
rect 7362 5070 7374 5122
rect 10098 5070 10110 5122
rect 10162 5070 10174 5122
rect 13906 5070 13918 5122
rect 13970 5070 13982 5122
rect 17938 5070 17950 5122
rect 18002 5070 18014 5122
rect 18722 5070 18734 5122
rect 18786 5070 18798 5122
rect 22530 5070 22542 5122
rect 22594 5070 22606 5122
rect 25890 5070 25902 5122
rect 25954 5070 25966 5122
rect 26674 5070 26686 5122
rect 26738 5070 26750 5122
rect 30370 5070 30382 5122
rect 30434 5070 30446 5122
rect 33954 5070 33966 5122
rect 34018 5070 34030 5122
rect 38322 5070 38334 5122
rect 38386 5070 38398 5122
rect 41794 5070 41806 5122
rect 41858 5070 41870 5122
rect 46386 5070 46398 5122
rect 46450 5070 46462 5122
rect 49858 5070 49870 5122
rect 49922 5070 49934 5122
rect 60386 5070 60398 5122
rect 60450 5070 60462 5122
rect 66658 5070 66670 5122
rect 66722 5070 66734 5122
rect 69458 5070 69470 5122
rect 69522 5070 69534 5122
rect 73714 5070 73726 5122
rect 73778 5070 73790 5122
rect 83906 5070 83918 5122
rect 83970 5070 83982 5122
rect 86706 5070 86718 5122
rect 86770 5070 86782 5122
rect 96114 5070 96126 5122
rect 96178 5070 96190 5122
rect 96674 5070 96686 5122
rect 96738 5070 96750 5122
rect 102610 5070 102622 5122
rect 102674 5070 102686 5122
rect 111906 5070 111918 5122
rect 111970 5070 111982 5122
rect 112690 5070 112702 5122
rect 112754 5070 112766 5122
rect 117058 5070 117070 5122
rect 117122 5070 117134 5122
rect 120642 5070 120654 5122
rect 120706 5070 120718 5122
rect 127922 5070 127934 5122
rect 127986 5070 127998 5122
rect 131282 5070 131294 5122
rect 131346 5070 131358 5122
rect 132962 5070 132974 5122
rect 133026 5070 133038 5122
rect 133746 5070 133758 5122
rect 133810 5070 133822 5122
rect 136434 5070 136446 5122
rect 136498 5070 136510 5122
rect 143826 5070 143838 5122
rect 143890 5070 143902 5122
rect 144498 5070 144510 5122
rect 144562 5070 144574 5122
rect 145170 5070 145182 5122
rect 145234 5070 145246 5122
rect 31154 4958 31166 5010
rect 31218 4958 31230 5010
rect 47058 4958 47070 5010
rect 47122 4958 47134 5010
rect 62178 4958 62190 5010
rect 62242 4958 62254 5010
rect 88946 4958 88958 5010
rect 89010 4958 89022 5010
rect 95330 4958 95342 5010
rect 95394 4958 95406 5010
rect 97458 4958 97470 5010
rect 97522 4958 97534 5010
rect 130610 4958 130622 5010
rect 130674 4958 130686 5010
rect 137218 4958 137230 5010
rect 137282 4958 137294 5010
rect 1344 4730 159092 4764
rect 1344 4678 40196 4730
rect 40248 4678 40320 4730
rect 40372 4678 40444 4730
rect 40496 4678 40568 4730
rect 40620 4678 40692 4730
rect 40744 4678 40816 4730
rect 40868 4678 40940 4730
rect 40992 4678 41064 4730
rect 41116 4678 79508 4730
rect 79560 4678 79632 4730
rect 79684 4678 79756 4730
rect 79808 4678 79880 4730
rect 79932 4678 80004 4730
rect 80056 4678 80128 4730
rect 80180 4678 80252 4730
rect 80304 4678 80376 4730
rect 80428 4678 118820 4730
rect 118872 4678 118944 4730
rect 118996 4678 119068 4730
rect 119120 4678 119192 4730
rect 119244 4678 119316 4730
rect 119368 4678 119440 4730
rect 119492 4678 119564 4730
rect 119616 4678 119688 4730
rect 119740 4678 158132 4730
rect 158184 4678 158256 4730
rect 158308 4678 158380 4730
rect 158432 4678 158504 4730
rect 158556 4678 158628 4730
rect 158680 4678 158752 4730
rect 158804 4678 158876 4730
rect 158928 4678 159000 4730
rect 159052 4678 159092 4730
rect 1344 4644 159092 4678
rect 6850 4398 6862 4450
rect 6914 4398 6926 4450
rect 13570 4398 13582 4450
rect 13634 4398 13646 4450
rect 30706 4398 30718 4450
rect 30770 4398 30782 4450
rect 37762 4398 37774 4450
rect 37826 4398 37838 4450
rect 43138 4398 43150 4450
rect 43202 4398 43214 4450
rect 46610 4398 46622 4450
rect 46674 4398 46686 4450
rect 63746 4398 63758 4450
rect 63810 4398 63822 4450
rect 65650 4398 65662 4450
rect 65714 4398 65726 4450
rect 105970 4398 105982 4450
rect 106034 4398 106046 4450
rect 109442 4398 109454 4450
rect 109506 4398 109518 4450
rect 115266 4398 115278 4450
rect 115330 4398 115342 4450
rect 118738 4398 118750 4450
rect 118802 4398 118814 4450
rect 121874 4398 121886 4450
rect 121938 4398 121950 4450
rect 131170 4398 131182 4450
rect 131234 4398 131246 4450
rect 134642 4398 134654 4450
rect 134706 4398 134718 4450
rect 5506 4286 5518 4338
rect 5570 4286 5582 4338
rect 6178 4286 6190 4338
rect 6242 4286 6254 4338
rect 12898 4286 12910 4338
rect 12962 4286 12974 4338
rect 22082 4286 22094 4338
rect 22146 4286 22158 4338
rect 29250 4286 29262 4338
rect 29314 4286 29326 4338
rect 29922 4286 29934 4338
rect 29986 4286 29998 4338
rect 37090 4286 37102 4338
rect 37154 4286 37166 4338
rect 42466 4286 42478 4338
rect 42530 4286 42542 4338
rect 45826 4286 45838 4338
rect 45890 4286 45902 4338
rect 53218 4286 53230 4338
rect 53282 4286 53294 4338
rect 53890 4286 53902 4338
rect 53954 4286 53966 4338
rect 60386 4286 60398 4338
rect 60450 4286 60462 4338
rect 70466 4286 70478 4338
rect 70530 4286 70542 4338
rect 73938 4286 73950 4338
rect 74002 4286 74014 4338
rect 83906 4286 83918 4338
rect 83970 4286 83982 4338
rect 89282 4286 89294 4338
rect 89346 4286 89358 4338
rect 100146 4286 100158 4338
rect 100210 4286 100222 4338
rect 105298 4286 105310 4338
rect 105362 4286 105374 4338
rect 108770 4286 108782 4338
rect 108834 4286 108846 4338
rect 116050 4286 116062 4338
rect 116114 4286 116126 4338
rect 119522 4286 119534 4338
rect 119586 4286 119598 4338
rect 121202 4286 121214 4338
rect 121266 4286 121278 4338
rect 124562 4286 124574 4338
rect 124626 4286 124638 4338
rect 131842 4286 131854 4338
rect 131906 4286 131918 4338
rect 135314 4286 135326 4338
rect 135378 4286 135390 4338
rect 139794 4286 139806 4338
rect 139858 4286 139870 4338
rect 143266 4286 143278 4338
rect 143330 4286 143342 4338
rect 2594 4174 2606 4226
rect 2658 4174 2670 4226
rect 4722 4174 4734 4226
rect 4786 4174 4798 4226
rect 8978 4174 8990 4226
rect 9042 4174 9054 4226
rect 15698 4174 15710 4226
rect 15762 4174 15774 4226
rect 22754 4174 22766 4226
rect 22818 4174 22830 4226
rect 24882 4174 24894 4226
rect 24946 4174 24958 4226
rect 26450 4174 26462 4226
rect 26514 4174 26526 4226
rect 28578 4174 28590 4226
rect 28642 4174 28654 4226
rect 32834 4174 32846 4226
rect 32898 4174 32910 4226
rect 39890 4174 39902 4226
rect 39954 4174 39966 4226
rect 45266 4174 45278 4226
rect 45330 4174 45342 4226
rect 48738 4174 48750 4226
rect 48802 4174 48814 4226
rect 50306 4174 50318 4226
rect 50370 4174 50382 4226
rect 52434 4174 52446 4226
rect 52498 4174 52510 4226
rect 54562 4174 54574 4226
rect 54626 4174 54638 4226
rect 56690 4174 56702 4226
rect 56754 4174 56766 4226
rect 78418 4174 78430 4226
rect 78482 4174 78494 4226
rect 88274 4174 88286 4226
rect 88338 4174 88350 4226
rect 93986 4174 93998 4226
rect 94050 4174 94062 4226
rect 97234 4174 97246 4226
rect 97298 4174 97310 4226
rect 99362 4174 99374 4226
rect 99426 4174 99438 4226
rect 108098 4174 108110 4226
rect 108162 4174 108174 4226
rect 111570 4174 111582 4226
rect 111634 4174 111646 4226
rect 113138 4174 113150 4226
rect 113202 4174 113214 4226
rect 116610 4174 116622 4226
rect 116674 4174 116686 4226
rect 124002 4174 124014 4226
rect 124066 4174 124078 4226
rect 125346 4174 125358 4226
rect 125410 4174 125422 4226
rect 127474 4174 127486 4226
rect 127538 4174 127550 4226
rect 129042 4174 129054 4226
rect 129106 4174 129118 4226
rect 132514 4174 132526 4226
rect 132578 4174 132590 4226
rect 136994 4174 137006 4226
rect 137058 4174 137070 4226
rect 139122 4174 139134 4226
rect 139186 4174 139198 4226
rect 140466 4174 140478 4226
rect 140530 4174 140542 4226
rect 142594 4174 142606 4226
rect 142658 4174 142670 4226
rect 1344 3946 158592 3980
rect 1344 3894 20540 3946
rect 20592 3894 20664 3946
rect 20716 3894 20788 3946
rect 20840 3894 20912 3946
rect 20964 3894 21036 3946
rect 21088 3894 21160 3946
rect 21212 3894 21284 3946
rect 21336 3894 21408 3946
rect 21460 3894 59852 3946
rect 59904 3894 59976 3946
rect 60028 3894 60100 3946
rect 60152 3894 60224 3946
rect 60276 3894 60348 3946
rect 60400 3894 60472 3946
rect 60524 3894 60596 3946
rect 60648 3894 60720 3946
rect 60772 3894 99164 3946
rect 99216 3894 99288 3946
rect 99340 3894 99412 3946
rect 99464 3894 99536 3946
rect 99588 3894 99660 3946
rect 99712 3894 99784 3946
rect 99836 3894 99908 3946
rect 99960 3894 100032 3946
rect 100084 3894 138476 3946
rect 138528 3894 138600 3946
rect 138652 3894 138724 3946
rect 138776 3894 138848 3946
rect 138900 3894 138972 3946
rect 139024 3894 139096 3946
rect 139148 3894 139220 3946
rect 139272 3894 139344 3946
rect 139396 3894 158592 3946
rect 1344 3860 158592 3894
rect 2034 3614 2046 3666
rect 2098 3614 2110 3666
rect 4162 3614 4174 3666
rect 4226 3614 4238 3666
rect 6626 3614 6638 3666
rect 6690 3614 6702 3666
rect 8754 3614 8766 3666
rect 8818 3614 8830 3666
rect 9650 3614 9662 3666
rect 9714 3614 9726 3666
rect 11778 3614 11790 3666
rect 11842 3614 11854 3666
rect 26338 3614 26350 3666
rect 26402 3614 26414 3666
rect 28466 3614 28478 3666
rect 28530 3614 28542 3666
rect 29474 3614 29486 3666
rect 29538 3614 29550 3666
rect 31602 3614 31614 3666
rect 31666 3614 31678 3666
rect 37874 3614 37886 3666
rect 37938 3614 37950 3666
rect 40002 3614 40014 3666
rect 40066 3614 40078 3666
rect 42018 3614 42030 3666
rect 42082 3614 42094 3666
rect 44146 3614 44158 3666
rect 44210 3614 44222 3666
rect 45938 3614 45950 3666
rect 46002 3614 46014 3666
rect 48066 3614 48078 3666
rect 48130 3614 48142 3666
rect 49858 3614 49870 3666
rect 49922 3614 49934 3666
rect 51986 3614 51998 3666
rect 52050 3614 52062 3666
rect 53778 3614 53790 3666
rect 53842 3614 53854 3666
rect 55906 3614 55918 3666
rect 55970 3614 55982 3666
rect 57698 3614 57710 3666
rect 57762 3614 57774 3666
rect 59826 3614 59838 3666
rect 59890 3614 59902 3666
rect 60834 3614 60846 3666
rect 60898 3614 60910 3666
rect 62962 3614 62974 3666
rect 63026 3614 63038 3666
rect 65538 3614 65550 3666
rect 65602 3614 65614 3666
rect 67666 3614 67678 3666
rect 67730 3614 67742 3666
rect 68450 3614 68462 3666
rect 68514 3614 68526 3666
rect 70578 3614 70590 3666
rect 70642 3614 70654 3666
rect 77298 3614 77310 3666
rect 77362 3614 77374 3666
rect 79426 3614 79438 3666
rect 79490 3614 79502 3666
rect 80994 3614 81006 3666
rect 81058 3614 81070 3666
rect 83122 3614 83134 3666
rect 83186 3614 83198 3666
rect 84914 3614 84926 3666
rect 84978 3614 84990 3666
rect 87042 3614 87054 3666
rect 87106 3614 87118 3666
rect 88834 3614 88846 3666
rect 88898 3614 88910 3666
rect 90962 3614 90974 3666
rect 91026 3614 91038 3666
rect 92754 3614 92766 3666
rect 92818 3614 92830 3666
rect 94882 3614 94894 3666
rect 94946 3614 94958 3666
rect 96674 3614 96686 3666
rect 96738 3614 96750 3666
rect 98802 3614 98814 3666
rect 98866 3614 98878 3666
rect 100594 3614 100606 3666
rect 100658 3614 100670 3666
rect 102722 3614 102734 3666
rect 102786 3614 102798 3666
rect 108434 3614 108446 3666
rect 108498 3614 108510 3666
rect 110562 3614 110574 3666
rect 110626 3614 110638 3666
rect 112354 3614 112366 3666
rect 112418 3614 112430 3666
rect 114482 3614 114494 3666
rect 114546 3614 114558 3666
rect 115490 3614 115502 3666
rect 115554 3614 115566 3666
rect 117618 3614 117630 3666
rect 117682 3614 117694 3666
rect 119410 3614 119422 3666
rect 119474 3614 119486 3666
rect 121538 3614 121550 3666
rect 121602 3614 121614 3666
rect 123330 3614 123342 3666
rect 123394 3614 123406 3666
rect 125458 3614 125470 3666
rect 125522 3614 125534 3666
rect 128034 3614 128046 3666
rect 128098 3614 128110 3666
rect 130162 3614 130174 3666
rect 130226 3614 130238 3666
rect 131954 3614 131966 3666
rect 132018 3614 132030 3666
rect 134082 3614 134094 3666
rect 134146 3614 134158 3666
rect 135874 3614 135886 3666
rect 135938 3614 135950 3666
rect 138002 3614 138014 3666
rect 138066 3614 138078 3666
rect 139794 3614 139806 3666
rect 139858 3614 139870 3666
rect 141922 3614 141934 3666
rect 141986 3614 141998 3666
rect 143714 3614 143726 3666
rect 143778 3614 143790 3666
rect 145842 3614 145854 3666
rect 145906 3614 145918 3666
rect 4834 3502 4846 3554
rect 4898 3502 4910 3554
rect 5842 3502 5854 3554
rect 5906 3502 5918 3554
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 25666 3502 25678 3554
rect 25730 3502 25742 3554
rect 32386 3502 32398 3554
rect 32450 3502 32462 3554
rect 37202 3502 37214 3554
rect 37266 3502 37278 3554
rect 41346 3502 41358 3554
rect 41410 3502 41422 3554
rect 45154 3502 45166 3554
rect 45218 3502 45230 3554
rect 49186 3502 49198 3554
rect 49250 3502 49262 3554
rect 53106 3502 53118 3554
rect 53170 3502 53182 3554
rect 57026 3502 57038 3554
rect 57090 3502 57102 3554
rect 63746 3502 63758 3554
rect 63810 3502 63822 3554
rect 64754 3502 64766 3554
rect 64818 3502 64830 3554
rect 71362 3502 71374 3554
rect 71426 3502 71438 3554
rect 76626 3502 76638 3554
rect 76690 3502 76702 3554
rect 80322 3502 80334 3554
rect 80386 3502 80398 3554
rect 84242 3502 84254 3554
rect 84306 3502 84318 3554
rect 88162 3502 88174 3554
rect 88226 3502 88238 3554
rect 92082 3502 92094 3554
rect 92146 3502 92158 3554
rect 95890 3502 95902 3554
rect 95954 3502 95966 3554
rect 99810 3502 99822 3554
rect 99874 3502 99886 3554
rect 107762 3502 107774 3554
rect 107826 3502 107838 3554
rect 111570 3502 111582 3554
rect 111634 3502 111646 3554
rect 118402 3502 118414 3554
rect 118466 3502 118478 3554
rect 122322 3502 122334 3554
rect 122386 3502 122398 3554
rect 126130 3502 126142 3554
rect 126194 3502 126206 3554
rect 127362 3502 127374 3554
rect 127426 3502 127438 3554
rect 131170 3502 131182 3554
rect 131234 3502 131246 3554
rect 135090 3502 135102 3554
rect 135154 3502 135166 3554
rect 139010 3502 139022 3554
rect 139074 3502 139086 3554
rect 142930 3502 142942 3554
rect 142994 3502 143006 3554
rect 1344 3162 159092 3196
rect 1344 3110 40196 3162
rect 40248 3110 40320 3162
rect 40372 3110 40444 3162
rect 40496 3110 40568 3162
rect 40620 3110 40692 3162
rect 40744 3110 40816 3162
rect 40868 3110 40940 3162
rect 40992 3110 41064 3162
rect 41116 3110 79508 3162
rect 79560 3110 79632 3162
rect 79684 3110 79756 3162
rect 79808 3110 79880 3162
rect 79932 3110 80004 3162
rect 80056 3110 80128 3162
rect 80180 3110 80252 3162
rect 80304 3110 80376 3162
rect 80428 3110 118820 3162
rect 118872 3110 118944 3162
rect 118996 3110 119068 3162
rect 119120 3110 119192 3162
rect 119244 3110 119316 3162
rect 119368 3110 119440 3162
rect 119492 3110 119564 3162
rect 119616 3110 119688 3162
rect 119740 3110 158132 3162
rect 158184 3110 158256 3162
rect 158308 3110 158380 3162
rect 158432 3110 158504 3162
rect 158556 3110 158628 3162
rect 158680 3110 158752 3162
rect 158804 3110 158876 3162
rect 158928 3110 159000 3162
rect 159052 3110 159092 3162
rect 1344 3076 159092 3110
<< via1 >>
rect 111582 6638 111634 6690
rect 112142 6638 112194 6690
rect 40196 6246 40248 6298
rect 40320 6246 40372 6298
rect 40444 6246 40496 6298
rect 40568 6246 40620 6298
rect 40692 6246 40744 6298
rect 40816 6246 40868 6298
rect 40940 6246 40992 6298
rect 41064 6246 41116 6298
rect 79508 6246 79560 6298
rect 79632 6246 79684 6298
rect 79756 6246 79808 6298
rect 79880 6246 79932 6298
rect 80004 6246 80056 6298
rect 80128 6246 80180 6298
rect 80252 6246 80304 6298
rect 80376 6246 80428 6298
rect 118820 6246 118872 6298
rect 118944 6246 118996 6298
rect 119068 6246 119120 6298
rect 119192 6246 119244 6298
rect 119316 6246 119368 6298
rect 119440 6246 119492 6298
rect 119564 6246 119616 6298
rect 119688 6246 119740 6298
rect 158132 6246 158184 6298
rect 158256 6246 158308 6298
rect 158380 6246 158432 6298
rect 158504 6246 158556 6298
rect 158628 6246 158680 6298
rect 158752 6246 158804 6298
rect 158876 6246 158928 6298
rect 159000 6246 159052 6298
rect 10670 5966 10722 6018
rect 2158 5854 2210 5906
rect 8878 5854 8930 5906
rect 9998 5854 10050 5906
rect 13918 5854 13970 5906
rect 17838 5854 17890 5906
rect 21646 5854 21698 5906
rect 25566 5854 25618 5906
rect 29486 5854 29538 5906
rect 33518 5854 33570 5906
rect 37326 5854 37378 5906
rect 41358 5854 41410 5906
rect 45278 5854 45330 5906
rect 49086 5854 49138 5906
rect 53006 5854 53058 5906
rect 57038 5854 57090 5906
rect 60846 5854 60898 5906
rect 64766 5854 64818 5906
rect 68686 5854 68738 5906
rect 72606 5854 72658 5906
rect 76638 5854 76690 5906
rect 80334 5854 80386 5906
rect 84142 5854 84194 5906
rect 90974 5854 91026 5906
rect 94894 5854 94946 5906
rect 98814 5854 98866 5906
rect 102734 5854 102786 5906
rect 103966 5854 104018 5906
rect 110574 5854 110626 5906
rect 114382 5854 114434 5906
rect 115614 5854 115666 5906
rect 119534 5854 119586 5906
rect 120206 5854 120258 5906
rect 123342 5854 123394 5906
rect 127262 5854 127314 5906
rect 131294 5854 131346 5906
rect 135102 5854 135154 5906
rect 139022 5854 139074 5906
rect 145742 5854 145794 5906
rect 2830 5742 2882 5794
rect 4958 5742 5010 5794
rect 5966 5742 6018 5794
rect 8094 5742 8146 5794
rect 12798 5742 12850 5794
rect 14590 5742 14642 5794
rect 16718 5742 16770 5794
rect 18510 5742 18562 5794
rect 20638 5742 20690 5794
rect 22430 5742 22482 5794
rect 24558 5742 24610 5794
rect 26350 5742 26402 5794
rect 28478 5742 28530 5794
rect 30270 5742 30322 5794
rect 32398 5742 32450 5794
rect 34190 5742 34242 5794
rect 36318 5742 36370 5794
rect 38110 5742 38162 5794
rect 40238 5742 40290 5794
rect 42030 5742 42082 5794
rect 44158 5742 44210 5794
rect 45950 5742 46002 5794
rect 48078 5742 48130 5794
rect 49870 5742 49922 5794
rect 51998 5742 52050 5794
rect 53790 5742 53842 5794
rect 55918 5742 55970 5794
rect 57710 5742 57762 5794
rect 59838 5742 59890 5794
rect 61630 5742 61682 5794
rect 63758 5742 63810 5794
rect 65550 5742 65602 5794
rect 67678 5742 67730 5794
rect 69470 5742 69522 5794
rect 71598 5742 71650 5794
rect 73390 5742 73442 5794
rect 75518 5742 75570 5794
rect 77310 5742 77362 5794
rect 79438 5742 79490 5794
rect 81006 5742 81058 5794
rect 83134 5742 83186 5794
rect 84926 5742 84978 5794
rect 87054 5742 87106 5794
rect 88062 5742 88114 5794
rect 90190 5742 90242 5794
rect 91982 5742 92034 5794
rect 94110 5742 94162 5794
rect 95902 5742 95954 5794
rect 98030 5742 98082 5794
rect 99822 5742 99874 5794
rect 101950 5742 102002 5794
rect 104750 5742 104802 5794
rect 106878 5742 106930 5794
rect 107662 5742 107714 5794
rect 109790 5742 109842 5794
rect 111582 5742 111634 5794
rect 113710 5742 113762 5794
rect 116286 5742 116338 5794
rect 118414 5742 118466 5794
rect 122334 5742 122386 5794
rect 124126 5742 124178 5794
rect 126254 5742 126306 5794
rect 128046 5742 128098 5794
rect 130174 5742 130226 5794
rect 131966 5742 132018 5794
rect 134094 5742 134146 5794
rect 135886 5742 135938 5794
rect 138014 5742 138066 5794
rect 139806 5742 139858 5794
rect 141934 5742 141986 5794
rect 142942 5742 142994 5794
rect 145070 5742 145122 5794
rect 20540 5462 20592 5514
rect 20664 5462 20716 5514
rect 20788 5462 20840 5514
rect 20912 5462 20964 5514
rect 21036 5462 21088 5514
rect 21160 5462 21212 5514
rect 21284 5462 21336 5514
rect 21408 5462 21460 5514
rect 59852 5462 59904 5514
rect 59976 5462 60028 5514
rect 60100 5462 60152 5514
rect 60224 5462 60276 5514
rect 60348 5462 60400 5514
rect 60472 5462 60524 5514
rect 60596 5462 60648 5514
rect 60720 5462 60772 5514
rect 99164 5462 99216 5514
rect 99288 5462 99340 5514
rect 99412 5462 99464 5514
rect 99536 5462 99588 5514
rect 99660 5462 99712 5514
rect 99784 5462 99836 5514
rect 99908 5462 99960 5514
rect 100032 5462 100084 5514
rect 138476 5462 138528 5514
rect 138600 5462 138652 5514
rect 138724 5462 138776 5514
rect 138848 5462 138900 5514
rect 138972 5462 139024 5514
rect 139096 5462 139148 5514
rect 139220 5462 139272 5514
rect 139344 5462 139396 5514
rect 2830 5182 2882 5234
rect 4958 5182 5010 5234
rect 9438 5182 9490 5234
rect 10782 5182 10834 5234
rect 12910 5182 12962 5234
rect 14702 5182 14754 5234
rect 16830 5182 16882 5234
rect 20862 5182 20914 5234
rect 23214 5182 23266 5234
rect 25342 5182 25394 5234
rect 28814 5182 28866 5234
rect 33294 5182 33346 5234
rect 34638 5182 34690 5234
rect 36766 5182 36818 5234
rect 39118 5182 39170 5234
rect 41246 5182 41298 5234
rect 42590 5182 42642 5234
rect 44718 5182 44770 5234
rect 49198 5182 49250 5234
rect 50542 5182 50594 5234
rect 52670 5182 52722 5234
rect 55582 5182 55634 5234
rect 70142 5182 70194 5234
rect 72270 5182 72322 5234
rect 74398 5182 74450 5234
rect 76526 5182 76578 5234
rect 82238 5182 82290 5234
rect 93214 5182 93266 5234
rect 99598 5182 99650 5234
rect 103294 5182 103346 5234
rect 105422 5182 105474 5234
rect 109118 5182 109170 5234
rect 111246 5182 111298 5234
rect 113374 5182 113426 5234
rect 115502 5182 115554 5234
rect 117854 5182 117906 5234
rect 119982 5182 120034 5234
rect 121326 5182 121378 5234
rect 123454 5182 123506 5234
rect 125022 5182 125074 5234
rect 127150 5182 127202 5234
rect 128494 5182 128546 5234
rect 135886 5182 135938 5234
rect 139358 5182 139410 5234
rect 140926 5182 140978 5234
rect 143054 5182 143106 5234
rect 147310 5182 147362 5234
rect 2046 5070 2098 5122
rect 6526 5070 6578 5122
rect 7310 5070 7362 5122
rect 10110 5070 10162 5122
rect 13918 5070 13970 5122
rect 17950 5070 18002 5122
rect 18734 5070 18786 5122
rect 22542 5070 22594 5122
rect 25902 5070 25954 5122
rect 26686 5070 26738 5122
rect 30382 5070 30434 5122
rect 33966 5070 34018 5122
rect 38334 5070 38386 5122
rect 41806 5070 41858 5122
rect 46398 5070 46450 5122
rect 49870 5070 49922 5122
rect 60398 5070 60450 5122
rect 66670 5070 66722 5122
rect 69470 5070 69522 5122
rect 73726 5070 73778 5122
rect 83918 5070 83970 5122
rect 86718 5070 86770 5122
rect 96126 5070 96178 5122
rect 96686 5070 96738 5122
rect 102622 5070 102674 5122
rect 111918 5070 111970 5122
rect 112702 5070 112754 5122
rect 117070 5070 117122 5122
rect 120654 5070 120706 5122
rect 127934 5070 127986 5122
rect 131294 5070 131346 5122
rect 132974 5070 133026 5122
rect 133758 5070 133810 5122
rect 136446 5070 136498 5122
rect 143838 5070 143890 5122
rect 144510 5070 144562 5122
rect 145182 5070 145234 5122
rect 31166 4958 31218 5010
rect 47070 4958 47122 5010
rect 62190 4958 62242 5010
rect 88958 4958 89010 5010
rect 95342 4958 95394 5010
rect 97470 4958 97522 5010
rect 130622 4958 130674 5010
rect 137230 4958 137282 5010
rect 40196 4678 40248 4730
rect 40320 4678 40372 4730
rect 40444 4678 40496 4730
rect 40568 4678 40620 4730
rect 40692 4678 40744 4730
rect 40816 4678 40868 4730
rect 40940 4678 40992 4730
rect 41064 4678 41116 4730
rect 79508 4678 79560 4730
rect 79632 4678 79684 4730
rect 79756 4678 79808 4730
rect 79880 4678 79932 4730
rect 80004 4678 80056 4730
rect 80128 4678 80180 4730
rect 80252 4678 80304 4730
rect 80376 4678 80428 4730
rect 118820 4678 118872 4730
rect 118944 4678 118996 4730
rect 119068 4678 119120 4730
rect 119192 4678 119244 4730
rect 119316 4678 119368 4730
rect 119440 4678 119492 4730
rect 119564 4678 119616 4730
rect 119688 4678 119740 4730
rect 158132 4678 158184 4730
rect 158256 4678 158308 4730
rect 158380 4678 158432 4730
rect 158504 4678 158556 4730
rect 158628 4678 158680 4730
rect 158752 4678 158804 4730
rect 158876 4678 158928 4730
rect 159000 4678 159052 4730
rect 6862 4398 6914 4450
rect 13582 4398 13634 4450
rect 30718 4398 30770 4450
rect 37774 4398 37826 4450
rect 43150 4398 43202 4450
rect 46622 4398 46674 4450
rect 63758 4398 63810 4450
rect 65662 4398 65714 4450
rect 105982 4398 106034 4450
rect 109454 4398 109506 4450
rect 115278 4398 115330 4450
rect 118750 4398 118802 4450
rect 121886 4398 121938 4450
rect 131182 4398 131234 4450
rect 134654 4398 134706 4450
rect 5518 4286 5570 4338
rect 6190 4286 6242 4338
rect 12910 4286 12962 4338
rect 22094 4286 22146 4338
rect 29262 4286 29314 4338
rect 29934 4286 29986 4338
rect 37102 4286 37154 4338
rect 42478 4286 42530 4338
rect 45838 4286 45890 4338
rect 53230 4286 53282 4338
rect 53902 4286 53954 4338
rect 60398 4286 60450 4338
rect 70478 4286 70530 4338
rect 73950 4286 74002 4338
rect 83918 4286 83970 4338
rect 89294 4286 89346 4338
rect 100158 4286 100210 4338
rect 105310 4286 105362 4338
rect 108782 4286 108834 4338
rect 116062 4286 116114 4338
rect 119534 4286 119586 4338
rect 121214 4286 121266 4338
rect 124574 4286 124626 4338
rect 131854 4286 131906 4338
rect 135326 4286 135378 4338
rect 139806 4286 139858 4338
rect 143278 4286 143330 4338
rect 2606 4174 2658 4226
rect 4734 4174 4786 4226
rect 8990 4174 9042 4226
rect 15710 4174 15762 4226
rect 22766 4174 22818 4226
rect 24894 4174 24946 4226
rect 26462 4174 26514 4226
rect 28590 4174 28642 4226
rect 32846 4174 32898 4226
rect 39902 4174 39954 4226
rect 45278 4174 45330 4226
rect 48750 4174 48802 4226
rect 50318 4174 50370 4226
rect 52446 4174 52498 4226
rect 54574 4174 54626 4226
rect 56702 4174 56754 4226
rect 78430 4174 78482 4226
rect 88286 4174 88338 4226
rect 93998 4174 94050 4226
rect 97246 4174 97298 4226
rect 99374 4174 99426 4226
rect 108110 4174 108162 4226
rect 111582 4174 111634 4226
rect 113150 4174 113202 4226
rect 116622 4174 116674 4226
rect 124014 4174 124066 4226
rect 125358 4174 125410 4226
rect 127486 4174 127538 4226
rect 129054 4174 129106 4226
rect 132526 4174 132578 4226
rect 137006 4174 137058 4226
rect 139134 4174 139186 4226
rect 140478 4174 140530 4226
rect 142606 4174 142658 4226
rect 20540 3894 20592 3946
rect 20664 3894 20716 3946
rect 20788 3894 20840 3946
rect 20912 3894 20964 3946
rect 21036 3894 21088 3946
rect 21160 3894 21212 3946
rect 21284 3894 21336 3946
rect 21408 3894 21460 3946
rect 59852 3894 59904 3946
rect 59976 3894 60028 3946
rect 60100 3894 60152 3946
rect 60224 3894 60276 3946
rect 60348 3894 60400 3946
rect 60472 3894 60524 3946
rect 60596 3894 60648 3946
rect 60720 3894 60772 3946
rect 99164 3894 99216 3946
rect 99288 3894 99340 3946
rect 99412 3894 99464 3946
rect 99536 3894 99588 3946
rect 99660 3894 99712 3946
rect 99784 3894 99836 3946
rect 99908 3894 99960 3946
rect 100032 3894 100084 3946
rect 138476 3894 138528 3946
rect 138600 3894 138652 3946
rect 138724 3894 138776 3946
rect 138848 3894 138900 3946
rect 138972 3894 139024 3946
rect 139096 3894 139148 3946
rect 139220 3894 139272 3946
rect 139344 3894 139396 3946
rect 2046 3614 2098 3666
rect 4174 3614 4226 3666
rect 6638 3614 6690 3666
rect 8766 3614 8818 3666
rect 9662 3614 9714 3666
rect 11790 3614 11842 3666
rect 26350 3614 26402 3666
rect 28478 3614 28530 3666
rect 29486 3614 29538 3666
rect 31614 3614 31666 3666
rect 37886 3614 37938 3666
rect 40014 3614 40066 3666
rect 42030 3614 42082 3666
rect 44158 3614 44210 3666
rect 45950 3614 46002 3666
rect 48078 3614 48130 3666
rect 49870 3614 49922 3666
rect 51998 3614 52050 3666
rect 53790 3614 53842 3666
rect 55918 3614 55970 3666
rect 57710 3614 57762 3666
rect 59838 3614 59890 3666
rect 60846 3614 60898 3666
rect 62974 3614 63026 3666
rect 65550 3614 65602 3666
rect 67678 3614 67730 3666
rect 68462 3614 68514 3666
rect 70590 3614 70642 3666
rect 77310 3614 77362 3666
rect 79438 3614 79490 3666
rect 81006 3614 81058 3666
rect 83134 3614 83186 3666
rect 84926 3614 84978 3666
rect 87054 3614 87106 3666
rect 88846 3614 88898 3666
rect 90974 3614 91026 3666
rect 92766 3614 92818 3666
rect 94894 3614 94946 3666
rect 96686 3614 96738 3666
rect 98814 3614 98866 3666
rect 100606 3614 100658 3666
rect 102734 3614 102786 3666
rect 108446 3614 108498 3666
rect 110574 3614 110626 3666
rect 112366 3614 112418 3666
rect 114494 3614 114546 3666
rect 115502 3614 115554 3666
rect 117630 3614 117682 3666
rect 119422 3614 119474 3666
rect 121550 3614 121602 3666
rect 123342 3614 123394 3666
rect 125470 3614 125522 3666
rect 128046 3614 128098 3666
rect 130174 3614 130226 3666
rect 131966 3614 132018 3666
rect 134094 3614 134146 3666
rect 135886 3614 135938 3666
rect 138014 3614 138066 3666
rect 139806 3614 139858 3666
rect 141934 3614 141986 3666
rect 143726 3614 143778 3666
rect 145854 3614 145906 3666
rect 4846 3502 4898 3554
rect 5854 3502 5906 3554
rect 12574 3502 12626 3554
rect 25678 3502 25730 3554
rect 32398 3502 32450 3554
rect 37214 3502 37266 3554
rect 41358 3502 41410 3554
rect 45166 3502 45218 3554
rect 49198 3502 49250 3554
rect 53118 3502 53170 3554
rect 57038 3502 57090 3554
rect 63758 3502 63810 3554
rect 64766 3502 64818 3554
rect 71374 3502 71426 3554
rect 76638 3502 76690 3554
rect 80334 3502 80386 3554
rect 84254 3502 84306 3554
rect 88174 3502 88226 3554
rect 92094 3502 92146 3554
rect 95902 3502 95954 3554
rect 99822 3502 99874 3554
rect 107774 3502 107826 3554
rect 111582 3502 111634 3554
rect 118414 3502 118466 3554
rect 122334 3502 122386 3554
rect 126142 3502 126194 3554
rect 127374 3502 127426 3554
rect 131182 3502 131234 3554
rect 135102 3502 135154 3554
rect 139022 3502 139074 3554
rect 142942 3502 142994 3554
rect 40196 3110 40248 3162
rect 40320 3110 40372 3162
rect 40444 3110 40496 3162
rect 40568 3110 40620 3162
rect 40692 3110 40744 3162
rect 40816 3110 40868 3162
rect 40940 3110 40992 3162
rect 41064 3110 41116 3162
rect 79508 3110 79560 3162
rect 79632 3110 79684 3162
rect 79756 3110 79808 3162
rect 79880 3110 79932 3162
rect 80004 3110 80056 3162
rect 80128 3110 80180 3162
rect 80252 3110 80304 3162
rect 80376 3110 80428 3162
rect 118820 3110 118872 3162
rect 118944 3110 118996 3162
rect 119068 3110 119120 3162
rect 119192 3110 119244 3162
rect 119316 3110 119368 3162
rect 119440 3110 119492 3162
rect 119564 3110 119616 3162
rect 119688 3110 119740 3162
rect 158132 3110 158184 3162
rect 158256 3110 158308 3162
rect 158380 3110 158432 3162
rect 158504 3110 158556 3162
rect 158628 3110 158680 3162
rect 158752 3110 158804 3162
rect 158876 3110 158928 3162
rect 159000 3110 159052 3162
<< metal2 >>
rect 1904 9200 2016 10000
rect 4592 9200 4704 10000
rect 7280 9200 7392 10000
rect 9968 9200 10080 10000
rect 12656 9200 12768 10000
rect 15344 9200 15456 10000
rect 18032 9200 18144 10000
rect 20720 9200 20832 10000
rect 23408 9200 23520 10000
rect 26096 9200 26208 10000
rect 28784 9200 28896 10000
rect 31472 9200 31584 10000
rect 34160 9200 34272 10000
rect 36848 9200 36960 10000
rect 39536 9200 39648 10000
rect 42224 9200 42336 10000
rect 44912 9200 45024 10000
rect 47600 9200 47712 10000
rect 50288 9200 50400 10000
rect 52976 9200 53088 10000
rect 55664 9200 55776 10000
rect 58352 9200 58464 10000
rect 61040 9200 61152 10000
rect 63728 9200 63840 10000
rect 66416 9200 66528 10000
rect 69104 9200 69216 10000
rect 71792 9200 71904 10000
rect 74480 9200 74592 10000
rect 77168 9200 77280 10000
rect 79856 9200 79968 10000
rect 82544 9200 82656 10000
rect 85232 9200 85344 10000
rect 87920 9200 88032 10000
rect 90608 9200 90720 10000
rect 93296 9200 93408 10000
rect 95984 9200 96096 10000
rect 98672 9200 98784 10000
rect 101360 9200 101472 10000
rect 104048 9200 104160 10000
rect 106736 9200 106848 10000
rect 109424 9200 109536 10000
rect 112112 9200 112224 10000
rect 114800 9200 114912 10000
rect 117488 9200 117600 10000
rect 120176 9200 120288 10000
rect 122864 9200 122976 10000
rect 125552 9200 125664 10000
rect 128240 9200 128352 10000
rect 130928 9200 131040 10000
rect 133616 9200 133728 10000
rect 136304 9200 136416 10000
rect 138992 9200 139104 10000
rect 141680 9200 141792 10000
rect 144368 9200 144480 10000
rect 147056 9200 147168 10000
rect 149744 9200 149856 10000
rect 152432 9200 152544 10000
rect 155120 9200 155232 10000
rect 157808 9200 157920 10000
rect 1932 3668 1988 9200
rect 2044 8260 2100 8270
rect 2044 5124 2100 8204
rect 4620 6468 4676 9200
rect 4620 6412 4900 6468
rect 2156 5906 2212 5918
rect 2156 5854 2158 5906
rect 2210 5854 2212 5906
rect 2156 5796 2212 5854
rect 2156 5730 2212 5740
rect 2828 5794 2884 5806
rect 2828 5742 2830 5794
rect 2882 5742 2884 5794
rect 2828 5236 2884 5742
rect 2044 4992 2100 5068
rect 2604 5234 2884 5236
rect 2604 5182 2830 5234
rect 2882 5182 2884 5234
rect 2604 5180 2884 5182
rect 4844 5236 4900 6412
rect 5964 6020 6020 6030
rect 4956 5794 5012 5806
rect 4956 5742 4958 5794
rect 5010 5742 5012 5794
rect 4956 5460 5012 5742
rect 5964 5794 6020 5964
rect 5964 5742 5966 5794
rect 6018 5742 6020 5794
rect 5964 5730 6020 5742
rect 4956 5404 5124 5460
rect 4956 5236 5012 5246
rect 4844 5234 5012 5236
rect 4844 5182 4958 5234
rect 5010 5182 5012 5234
rect 4844 5180 5012 5182
rect 2604 4226 2660 5180
rect 2828 5170 2884 5180
rect 4956 5170 5012 5180
rect 4732 5124 4788 5134
rect 4788 5068 4900 5124
rect 4732 5058 4788 5068
rect 2604 4174 2606 4226
rect 2658 4174 2660 4226
rect 2604 4162 2660 4174
rect 4172 4228 4228 4238
rect 2044 3668 2100 3678
rect 1932 3666 2100 3668
rect 1932 3614 2046 3666
rect 2098 3614 2100 3666
rect 1932 3612 2100 3614
rect 2044 3602 2100 3612
rect 4172 3666 4228 4172
rect 4732 4228 4788 4238
rect 4732 4134 4788 4172
rect 4172 3614 4174 3666
rect 4226 3614 4228 3666
rect 4172 3602 4228 3614
rect 4844 3556 4900 5068
rect 5068 4452 5124 5404
rect 7308 5348 7364 9200
rect 9996 7252 10052 9200
rect 9436 7196 10052 7252
rect 8876 5906 8932 5918
rect 8876 5854 8878 5906
rect 8930 5854 8932 5906
rect 8092 5794 8148 5806
rect 8092 5742 8094 5794
rect 8146 5742 8148 5794
rect 7308 5292 7476 5348
rect 6524 5124 6580 5134
rect 6524 5030 6580 5068
rect 7308 5124 7364 5134
rect 7308 5030 7364 5068
rect 5068 4386 5124 4396
rect 6636 4452 6692 4462
rect 5516 4340 5572 4350
rect 5516 4246 5572 4284
rect 6188 4340 6244 4350
rect 6188 4246 6244 4284
rect 6636 3666 6692 4396
rect 6860 4452 6916 4462
rect 6860 4358 6916 4396
rect 6636 3614 6638 3666
rect 6690 3614 6692 3666
rect 6636 3602 6692 3614
rect 7420 3668 7476 5292
rect 8092 5124 8148 5742
rect 8092 5058 8148 5068
rect 8876 5124 8932 5854
rect 8876 5058 8932 5068
rect 8988 5236 9044 5246
rect 8988 4226 9044 5180
rect 9436 5234 9492 7196
rect 12684 7028 12740 9200
rect 12684 6972 12964 7028
rect 10668 6020 10724 6030
rect 9996 5908 10052 5918
rect 9996 5814 10052 5852
rect 9436 5182 9438 5234
rect 9490 5182 9492 5234
rect 9436 5170 9492 5182
rect 10108 5684 10164 5694
rect 10108 5348 10164 5628
rect 10108 5122 10164 5292
rect 10668 5236 10724 5964
rect 12796 5796 12852 5806
rect 12796 5702 12852 5740
rect 10780 5236 10836 5246
rect 10668 5234 10836 5236
rect 10668 5182 10782 5234
rect 10834 5182 10836 5234
rect 10668 5180 10836 5182
rect 10780 5170 10836 5180
rect 12908 5234 12964 6972
rect 13916 5906 13972 5918
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 13580 5796 13636 5806
rect 12908 5182 12910 5234
rect 12962 5182 12964 5234
rect 12908 5170 12964 5182
rect 13020 5684 13076 5694
rect 10108 5070 10110 5122
rect 10162 5070 10164 5122
rect 10108 5058 10164 5070
rect 12572 4340 12628 4350
rect 8988 4174 8990 4226
rect 9042 4174 9044 4226
rect 8988 4162 9044 4174
rect 9660 4228 9716 4238
rect 7420 3602 7476 3612
rect 8764 3668 8820 3678
rect 8764 3574 8820 3612
rect 9660 3666 9716 4172
rect 9660 3614 9662 3666
rect 9714 3614 9716 3666
rect 9660 3602 9716 3614
rect 11788 4116 11844 4126
rect 11788 3666 11844 4060
rect 11788 3614 11790 3666
rect 11842 3614 11844 3666
rect 11788 3602 11844 3614
rect 5852 3556 5908 3566
rect 4844 3554 5908 3556
rect 4844 3502 4846 3554
rect 4898 3502 5854 3554
rect 5906 3502 5908 3554
rect 4844 3500 5908 3502
rect 4844 3490 4900 3500
rect 5852 3490 5908 3500
rect 12572 3556 12628 4284
rect 12908 4340 12964 4350
rect 13020 4340 13076 5628
rect 13580 5236 13636 5740
rect 13916 5684 13972 5854
rect 13916 5618 13972 5628
rect 14588 5794 14644 5806
rect 14588 5742 14590 5794
rect 14642 5742 14644 5794
rect 13580 4450 13636 5180
rect 13916 5124 13972 5134
rect 13916 5030 13972 5068
rect 14588 5012 14644 5742
rect 14700 5236 14756 5246
rect 14700 5142 14756 5180
rect 14588 4946 14644 4956
rect 13580 4398 13582 4450
rect 13634 4398 13636 4450
rect 13580 4386 13636 4398
rect 12908 4338 13076 4340
rect 12908 4286 12910 4338
rect 12962 4286 13076 4338
rect 12908 4284 13076 4286
rect 12908 4274 12964 4284
rect 15372 4228 15428 9200
rect 17836 5906 17892 5918
rect 17836 5854 17838 5906
rect 17890 5854 17892 5906
rect 16716 5796 16772 5806
rect 16716 5702 16772 5740
rect 17836 5684 17892 5854
rect 18060 5796 18116 9200
rect 18060 5730 18116 5740
rect 18508 5794 18564 5806
rect 18508 5742 18510 5794
rect 18562 5742 18564 5794
rect 17836 5618 17892 5628
rect 16828 5234 16884 5246
rect 16828 5182 16830 5234
rect 16882 5182 16884 5234
rect 16828 5012 16884 5182
rect 17948 5124 18004 5134
rect 17948 5030 18004 5068
rect 16828 4946 16884 4956
rect 18508 4788 18564 5742
rect 20636 5796 20692 5806
rect 20748 5796 20804 9200
rect 20636 5794 20804 5796
rect 20636 5742 20638 5794
rect 20690 5742 20804 5794
rect 20636 5740 20804 5742
rect 21644 5906 21700 5918
rect 21644 5854 21646 5906
rect 21698 5854 21700 5906
rect 21644 5796 21700 5854
rect 20636 5730 20692 5740
rect 20538 5516 21462 5526
rect 20538 5514 20556 5516
rect 20538 5462 20540 5514
rect 20538 5460 20556 5462
rect 20612 5460 20660 5516
rect 20716 5460 20764 5516
rect 20820 5514 20868 5516
rect 20924 5514 20972 5516
rect 20840 5462 20868 5514
rect 20964 5462 20972 5514
rect 20820 5460 20868 5462
rect 20924 5460 20972 5462
rect 21028 5514 21076 5516
rect 21132 5514 21180 5516
rect 21028 5462 21036 5514
rect 21132 5462 21160 5514
rect 21028 5460 21076 5462
rect 21132 5460 21180 5462
rect 21236 5460 21284 5516
rect 21340 5460 21388 5516
rect 21444 5514 21462 5516
rect 21460 5462 21462 5514
rect 21444 5460 21462 5462
rect 20538 5450 21462 5460
rect 20860 5234 20916 5246
rect 20860 5182 20862 5234
rect 20914 5182 20916 5234
rect 18732 5122 18788 5134
rect 18732 5070 18734 5122
rect 18786 5070 18788 5122
rect 18732 5012 18788 5070
rect 18732 4946 18788 4956
rect 18508 4722 18564 4732
rect 20860 4788 20916 5182
rect 21644 5124 21700 5740
rect 22428 5794 22484 5806
rect 22428 5742 22430 5794
rect 22482 5742 22484 5794
rect 21644 5058 21700 5068
rect 22092 5684 22148 5694
rect 20860 4722 20916 4732
rect 22092 4338 22148 5628
rect 22092 4286 22094 4338
rect 22146 4286 22148 4338
rect 22092 4274 22148 4286
rect 15708 4228 15764 4238
rect 15372 4226 15764 4228
rect 15372 4174 15710 4226
rect 15762 4174 15764 4226
rect 15372 4172 15764 4174
rect 22428 4228 22484 5742
rect 22540 5684 22596 5694
rect 22540 5124 22596 5628
rect 23212 5684 23268 5694
rect 23212 5234 23268 5628
rect 23212 5182 23214 5234
rect 23266 5182 23268 5234
rect 23212 5170 23268 5182
rect 22540 4992 22596 5068
rect 23436 4340 23492 9200
rect 25564 5906 25620 5918
rect 25564 5854 25566 5906
rect 25618 5854 25620 5906
rect 24556 5794 24612 5806
rect 24556 5742 24558 5794
rect 24610 5742 24612 5794
rect 24556 5684 24612 5742
rect 25564 5796 25620 5854
rect 25564 5730 25620 5740
rect 24556 5618 24612 5628
rect 25340 5234 25396 5246
rect 25340 5182 25342 5234
rect 25394 5182 25396 5234
rect 25340 4900 25396 5182
rect 25340 4834 25396 4844
rect 25900 5124 25956 5134
rect 25900 4452 25956 5068
rect 25900 4386 25956 4396
rect 23436 4274 23492 4284
rect 22764 4228 22820 4238
rect 22428 4226 22820 4228
rect 22428 4174 22766 4226
rect 22818 4174 22820 4226
rect 22428 4172 22820 4174
rect 15708 4162 15764 4172
rect 20538 3948 21462 3958
rect 20538 3946 20556 3948
rect 20538 3894 20540 3946
rect 20538 3892 20556 3894
rect 20612 3892 20660 3948
rect 20716 3892 20764 3948
rect 20820 3946 20868 3948
rect 20924 3946 20972 3948
rect 20840 3894 20868 3946
rect 20964 3894 20972 3946
rect 20820 3892 20868 3894
rect 20924 3892 20972 3894
rect 21028 3946 21076 3948
rect 21132 3946 21180 3948
rect 21028 3894 21036 3946
rect 21132 3894 21160 3946
rect 21028 3892 21076 3894
rect 21132 3892 21180 3894
rect 21236 3892 21284 3948
rect 21340 3892 21388 3948
rect 21444 3946 21462 3948
rect 21460 3894 21462 3946
rect 21444 3892 21462 3894
rect 20538 3882 21462 3892
rect 22764 3668 22820 4172
rect 24892 4228 24948 4238
rect 24892 4134 24948 4172
rect 26124 4228 26180 9200
rect 26348 5794 26404 5806
rect 26348 5742 26350 5794
rect 26402 5742 26404 5794
rect 26124 4162 26180 4172
rect 26236 5684 26292 5694
rect 26236 3668 26292 5628
rect 26348 5124 26404 5742
rect 28476 5794 28532 5806
rect 28476 5742 28478 5794
rect 28530 5742 28532 5794
rect 28476 5684 28532 5742
rect 28812 5684 28868 9200
rect 30380 6020 30436 6030
rect 29484 5906 29540 5918
rect 29484 5854 29486 5906
rect 29538 5854 29540 5906
rect 29484 5796 29540 5854
rect 29484 5730 29540 5740
rect 30268 5794 30324 5806
rect 30268 5742 30270 5794
rect 30322 5742 30324 5794
rect 28476 5618 28532 5628
rect 28700 5628 28868 5684
rect 30268 5684 30324 5742
rect 26348 5058 26404 5068
rect 26684 5124 26740 5134
rect 26684 5030 26740 5068
rect 28476 5124 28532 5134
rect 26460 4340 26516 4350
rect 26460 4226 26516 4284
rect 26460 4174 26462 4226
rect 26514 4174 26516 4226
rect 26460 4162 26516 4174
rect 26348 3668 26404 3678
rect 26236 3666 26404 3668
rect 26236 3614 26350 3666
rect 26402 3614 26404 3666
rect 26236 3612 26404 3614
rect 22764 3602 22820 3612
rect 26348 3602 26404 3612
rect 28476 3666 28532 5068
rect 28700 4900 28756 5628
rect 28812 5234 28868 5246
rect 28812 5182 28814 5234
rect 28866 5182 28868 5234
rect 28812 5012 28868 5182
rect 28812 4946 28868 4956
rect 28700 4834 28756 4844
rect 29260 4452 29316 4462
rect 29260 4338 29316 4396
rect 29260 4286 29262 4338
rect 29314 4286 29316 4338
rect 29260 4274 29316 4286
rect 29932 4452 29988 4462
rect 30268 4452 30324 5628
rect 30380 5796 30436 5964
rect 30380 5122 30436 5740
rect 30380 5070 30382 5122
rect 30434 5070 30436 5122
rect 30380 5058 30436 5070
rect 31164 5010 31220 5022
rect 31164 4958 31166 5010
rect 31218 4958 31220 5010
rect 31164 4788 31220 4958
rect 31500 5012 31556 9200
rect 34188 6020 34244 9200
rect 34076 5964 34244 6020
rect 33516 5908 33572 5918
rect 33516 5814 33572 5852
rect 32396 5794 32452 5806
rect 32396 5742 32398 5794
rect 32450 5742 32452 5794
rect 32396 5684 32452 5742
rect 32396 5618 32452 5628
rect 31500 4946 31556 4956
rect 33292 5234 33348 5246
rect 33292 5182 33294 5234
rect 33346 5182 33348 5234
rect 33292 4900 33348 5182
rect 33292 4834 33348 4844
rect 33964 5122 34020 5134
rect 33964 5070 33966 5122
rect 34018 5070 34020 5122
rect 33964 5012 34020 5070
rect 31164 4722 31220 4732
rect 30716 4452 30772 4462
rect 30268 4450 30772 4452
rect 30268 4398 30718 4450
rect 30770 4398 30772 4450
rect 30268 4396 30772 4398
rect 29932 4338 29988 4396
rect 30716 4386 30772 4396
rect 33964 4452 34020 4956
rect 33964 4386 34020 4396
rect 29932 4286 29934 4338
rect 29986 4286 29988 4338
rect 29932 4274 29988 4286
rect 32396 4340 32452 4350
rect 28588 4228 28644 4238
rect 28588 4134 28644 4172
rect 31612 4228 31668 4238
rect 28476 3614 28478 3666
rect 28530 3614 28532 3666
rect 28476 3602 28532 3614
rect 29484 3668 29540 3678
rect 29484 3574 29540 3612
rect 31612 3666 31668 4172
rect 31612 3614 31614 3666
rect 31666 3614 31668 3666
rect 12572 3462 12628 3500
rect 25676 3556 25732 3566
rect 25676 3462 25732 3500
rect 31612 3444 31668 3614
rect 32396 3556 32452 4284
rect 32844 4228 32900 4238
rect 32844 4134 32900 4172
rect 34076 4228 34132 5964
rect 34188 5794 34244 5806
rect 34188 5742 34190 5794
rect 34242 5742 34244 5794
rect 34188 5684 34244 5742
rect 36316 5794 36372 5806
rect 36316 5742 36318 5794
rect 36370 5742 36372 5794
rect 34188 5618 34244 5628
rect 34636 5684 34692 5694
rect 34636 5234 34692 5628
rect 34636 5182 34638 5234
rect 34690 5182 34692 5234
rect 34636 5170 34692 5182
rect 36316 5124 36372 5742
rect 36764 5236 36820 5246
rect 36876 5236 36932 9200
rect 37324 5908 37380 5918
rect 36764 5234 36932 5236
rect 36764 5182 36766 5234
rect 36818 5182 36932 5234
rect 36764 5180 36932 5182
rect 37212 5906 37380 5908
rect 37212 5854 37326 5906
rect 37378 5854 37380 5906
rect 37212 5852 37380 5854
rect 36764 5170 36820 5180
rect 36316 5058 36372 5068
rect 37212 5012 37268 5852
rect 37324 5842 37380 5852
rect 38108 5794 38164 5806
rect 38108 5742 38110 5794
rect 38162 5742 38164 5794
rect 38108 5236 38164 5742
rect 38108 5170 38164 5180
rect 38332 5796 38388 5806
rect 37100 4340 37156 4350
rect 37100 4246 37156 4284
rect 34076 4162 34132 4172
rect 32396 3424 32452 3500
rect 37212 3556 37268 4956
rect 37772 5124 37828 5134
rect 37772 4450 37828 5068
rect 38332 5122 38388 5740
rect 39116 5236 39172 5246
rect 39116 5142 39172 5180
rect 38332 5070 38334 5122
rect 38386 5070 38388 5122
rect 38332 5058 38388 5070
rect 37772 4398 37774 4450
rect 37826 4398 37828 4450
rect 37772 3668 37828 4398
rect 37884 3668 37940 3678
rect 37772 3666 37940 3668
rect 37772 3614 37886 3666
rect 37938 3614 37940 3666
rect 37772 3612 37940 3614
rect 37884 3602 37940 3612
rect 39564 3668 39620 9200
rect 40194 6300 41118 6310
rect 40194 6298 40212 6300
rect 40194 6246 40196 6298
rect 40194 6244 40212 6246
rect 40268 6244 40316 6300
rect 40372 6244 40420 6300
rect 40476 6298 40524 6300
rect 40580 6298 40628 6300
rect 40496 6246 40524 6298
rect 40620 6246 40628 6298
rect 40476 6244 40524 6246
rect 40580 6244 40628 6246
rect 40684 6298 40732 6300
rect 40788 6298 40836 6300
rect 40684 6246 40692 6298
rect 40788 6246 40816 6298
rect 40684 6244 40732 6246
rect 40788 6244 40836 6246
rect 40892 6244 40940 6300
rect 40996 6244 41044 6300
rect 41100 6298 41118 6300
rect 41116 6246 41118 6298
rect 41100 6244 41118 6246
rect 40194 6234 41118 6244
rect 41356 5908 41412 5918
rect 41356 5814 41412 5852
rect 40236 5794 40292 5806
rect 40236 5742 40238 5794
rect 40290 5742 40292 5794
rect 39900 5236 39956 5246
rect 39900 4226 39956 5180
rect 40236 5012 40292 5742
rect 42028 5794 42084 5806
rect 42028 5742 42030 5794
rect 42082 5742 42084 5794
rect 41244 5236 41300 5246
rect 41244 5142 41300 5180
rect 42028 5236 42084 5742
rect 42028 5170 42084 5180
rect 40236 4946 40292 4956
rect 41804 5122 41860 5134
rect 41804 5070 41806 5122
rect 41858 5070 41860 5122
rect 40194 4732 41118 4742
rect 40194 4730 40212 4732
rect 40194 4678 40196 4730
rect 40194 4676 40212 4678
rect 40268 4676 40316 4732
rect 40372 4676 40420 4732
rect 40476 4730 40524 4732
rect 40580 4730 40628 4732
rect 40496 4678 40524 4730
rect 40620 4678 40628 4730
rect 40476 4676 40524 4678
rect 40580 4676 40628 4678
rect 40684 4730 40732 4732
rect 40788 4730 40836 4732
rect 40684 4678 40692 4730
rect 40788 4678 40816 4730
rect 40684 4676 40732 4678
rect 40788 4676 40836 4678
rect 40892 4676 40940 4732
rect 40996 4676 41044 4732
rect 41100 4730 41118 4732
rect 41116 4678 41118 4730
rect 41100 4676 41118 4678
rect 40194 4666 41118 4676
rect 39900 4174 39902 4226
rect 39954 4174 39956 4226
rect 39900 4162 39956 4174
rect 39564 3602 39620 3612
rect 40012 3668 40068 3678
rect 40012 3574 40068 3612
rect 37212 3462 37268 3500
rect 41356 3556 41412 3566
rect 41356 3462 41412 3500
rect 41804 3556 41860 5070
rect 42140 5124 42196 5134
rect 42028 3668 42084 3678
rect 42140 3668 42196 5068
rect 42252 5012 42308 9200
rect 44940 7252 44996 9200
rect 44716 7196 44996 7252
rect 44156 5794 44212 5806
rect 44156 5742 44158 5794
rect 44210 5742 44212 5794
rect 42588 5236 42644 5246
rect 42588 5142 42644 5180
rect 42252 4946 42308 4956
rect 43148 5124 43204 5134
rect 43148 4450 43204 5068
rect 44156 5124 44212 5742
rect 44716 5234 44772 7196
rect 44716 5182 44718 5234
rect 44770 5182 44772 5234
rect 44716 5170 44772 5182
rect 45276 5906 45332 5918
rect 45276 5854 45278 5906
rect 45330 5854 45332 5906
rect 45276 5796 45332 5854
rect 44156 5058 44212 5068
rect 45276 5124 45332 5740
rect 45276 5058 45332 5068
rect 45948 5794 46004 5806
rect 45948 5742 45950 5794
rect 46002 5742 46004 5794
rect 43148 4398 43150 4450
rect 43202 4398 43204 4450
rect 43148 4386 43204 4398
rect 45948 4900 46004 5742
rect 46396 5124 46452 5134
rect 46396 5030 46452 5068
rect 47068 5012 47124 5022
rect 42476 4340 42532 4350
rect 42476 4246 42532 4284
rect 45836 4338 45892 4350
rect 45836 4286 45838 4338
rect 45890 4286 45892 4338
rect 45276 4228 45332 4238
rect 45276 4134 45332 4172
rect 45164 4116 45220 4126
rect 42028 3666 42196 3668
rect 42028 3614 42030 3666
rect 42082 3614 42196 3666
rect 42028 3612 42196 3614
rect 44156 3668 44212 3678
rect 42028 3602 42084 3612
rect 44156 3574 44212 3612
rect 41804 3490 41860 3500
rect 45164 3556 45220 4060
rect 45836 4116 45892 4286
rect 45836 4050 45892 4060
rect 45948 3666 46004 4844
rect 46620 5010 47124 5012
rect 46620 4958 47070 5010
rect 47122 4958 47124 5010
rect 46620 4956 47124 4958
rect 46620 4450 46676 4956
rect 47068 4946 47124 4956
rect 46620 4398 46622 4450
rect 46674 4398 46676 4450
rect 46620 4228 46676 4398
rect 46620 4162 46676 4172
rect 45948 3614 45950 3666
rect 46002 3614 46004 3666
rect 45948 3602 46004 3614
rect 47628 3668 47684 9200
rect 49084 5906 49140 5918
rect 49084 5854 49086 5906
rect 49138 5854 49140 5906
rect 48076 5796 48132 5806
rect 48076 5702 48132 5740
rect 48748 4452 48804 4462
rect 48748 4226 48804 4396
rect 48748 4174 48750 4226
rect 48802 4174 48804 4226
rect 48748 4162 48804 4174
rect 49084 4116 49140 5854
rect 49868 5796 49924 5806
rect 49868 5702 49924 5740
rect 49196 5348 49252 5358
rect 49196 5234 49252 5292
rect 49196 5182 49198 5234
rect 49250 5182 49252 5234
rect 49196 5170 49252 5182
rect 49756 5348 49812 5358
rect 47628 3602 47684 3612
rect 48076 4004 48132 4014
rect 48076 3666 48132 3948
rect 48076 3614 48078 3666
rect 48130 3614 48132 3666
rect 48076 3602 48132 3614
rect 49084 3556 49140 4060
rect 49756 3668 49812 5292
rect 49868 5124 49924 5134
rect 49868 5030 49924 5068
rect 50316 4452 50372 9200
rect 53004 6132 53060 9200
rect 52892 6076 53060 6132
rect 50540 5796 50596 5806
rect 50540 5234 50596 5740
rect 50540 5182 50542 5234
rect 50594 5182 50596 5234
rect 50540 5170 50596 5182
rect 51996 5794 52052 5806
rect 51996 5742 51998 5794
rect 52050 5742 52052 5794
rect 51996 5012 52052 5742
rect 51996 4946 52052 4956
rect 52668 5234 52724 5246
rect 52668 5182 52670 5234
rect 52722 5182 52724 5234
rect 50316 4386 50372 4396
rect 50316 4226 50372 4238
rect 50316 4174 50318 4226
rect 50370 4174 50372 4226
rect 49868 3668 49924 3678
rect 49756 3666 49924 3668
rect 49756 3614 49870 3666
rect 49922 3614 49924 3666
rect 49756 3612 49924 3614
rect 49868 3602 49924 3612
rect 49196 3556 49252 3566
rect 49084 3500 49196 3556
rect 45164 3424 45220 3500
rect 49196 3462 49252 3500
rect 50316 3444 50372 4174
rect 52444 4226 52500 4238
rect 52444 4174 52446 4226
rect 52498 4174 52500 4226
rect 52444 4116 52500 4174
rect 52444 4050 52500 4060
rect 51996 3780 52052 3790
rect 51996 3666 52052 3724
rect 51996 3614 51998 3666
rect 52050 3614 52052 3666
rect 51996 3602 52052 3614
rect 52668 3668 52724 5182
rect 52892 3780 52948 6076
rect 53004 5908 53060 5918
rect 53004 5236 53060 5852
rect 53788 5794 53844 5806
rect 53788 5742 53790 5794
rect 53842 5742 53844 5794
rect 53004 5170 53060 5180
rect 53116 5684 53172 5694
rect 52892 3714 52948 3724
rect 52668 3602 52724 3612
rect 31612 3378 31668 3388
rect 53116 3556 53172 5628
rect 53788 5348 53844 5742
rect 53788 5282 53844 5292
rect 55580 5236 55636 5246
rect 55580 5142 55636 5180
rect 53228 4338 53284 4350
rect 53228 4286 53230 4338
rect 53282 4286 53284 4338
rect 53228 4228 53284 4286
rect 53228 4162 53284 4172
rect 53900 4338 53956 4350
rect 53900 4286 53902 4338
rect 53954 4286 53956 4338
rect 53900 4228 53956 4286
rect 53788 3668 53844 3678
rect 53788 3574 53844 3612
rect 53116 3424 53172 3500
rect 53900 3556 53956 4172
rect 54572 4226 54628 4238
rect 54572 4174 54574 4226
rect 54626 4174 54628 4226
rect 54572 3668 54628 4174
rect 55692 4004 55748 9200
rect 57036 5906 57092 5918
rect 57036 5854 57038 5906
rect 57090 5854 57092 5906
rect 55916 5796 55972 5806
rect 55916 5702 55972 5740
rect 57036 5124 57092 5854
rect 57708 5796 57764 5806
rect 57708 5794 57876 5796
rect 57708 5742 57710 5794
rect 57762 5742 57876 5794
rect 57708 5740 57876 5742
rect 57708 5730 57764 5740
rect 56700 4676 56756 4686
rect 55692 3938 55748 3948
rect 55916 4228 55972 4238
rect 54572 3602 54628 3612
rect 55916 3666 55972 4172
rect 56700 4226 56756 4620
rect 57036 4564 57092 5068
rect 57036 4498 57092 4508
rect 57708 5012 57764 5022
rect 56700 4174 56702 4226
rect 56754 4174 56756 4226
rect 56700 4162 56756 4174
rect 55916 3614 55918 3666
rect 55970 3614 55972 3666
rect 55916 3602 55972 3614
rect 57708 3666 57764 4956
rect 57820 4676 57876 5740
rect 58380 4900 58436 9200
rect 60844 5906 60900 5918
rect 60844 5854 60846 5906
rect 60898 5854 60900 5906
rect 59836 5796 59892 5806
rect 59724 5794 59892 5796
rect 59724 5742 59838 5794
rect 59890 5742 59892 5794
rect 59724 5740 59892 5742
rect 59724 5012 59780 5740
rect 59836 5730 59892 5740
rect 60844 5684 60900 5854
rect 60844 5618 60900 5628
rect 59850 5516 60774 5526
rect 59850 5514 59868 5516
rect 59850 5462 59852 5514
rect 59850 5460 59868 5462
rect 59924 5460 59972 5516
rect 60028 5460 60076 5516
rect 60132 5514 60180 5516
rect 60236 5514 60284 5516
rect 60152 5462 60180 5514
rect 60276 5462 60284 5514
rect 60132 5460 60180 5462
rect 60236 5460 60284 5462
rect 60340 5514 60388 5516
rect 60444 5514 60492 5516
rect 60340 5462 60348 5514
rect 60444 5462 60472 5514
rect 60340 5460 60388 5462
rect 60444 5460 60492 5462
rect 60548 5460 60596 5516
rect 60652 5460 60700 5516
rect 60756 5514 60774 5516
rect 60772 5462 60774 5514
rect 60756 5460 60774 5462
rect 59850 5450 60774 5460
rect 59724 4946 59780 4956
rect 60396 5124 60452 5134
rect 58380 4834 58436 4844
rect 57820 4610 57876 4620
rect 60396 4338 60452 5068
rect 60396 4286 60398 4338
rect 60450 4286 60452 4338
rect 60396 4274 60452 4286
rect 61068 4228 61124 9200
rect 63756 6020 63812 9200
rect 63644 5964 63812 6020
rect 61628 5794 61684 5806
rect 61628 5742 61630 5794
rect 61682 5742 61684 5794
rect 61628 5012 61684 5742
rect 61628 4946 61684 4956
rect 62188 5010 62244 5022
rect 62188 4958 62190 5010
rect 62242 4958 62244 5010
rect 62188 4340 62244 4958
rect 63644 4900 63700 5964
rect 64764 5906 64820 5918
rect 64764 5854 64766 5906
rect 64818 5854 64820 5906
rect 63756 5794 63812 5806
rect 63756 5742 63758 5794
rect 63810 5742 63812 5794
rect 63756 5012 63812 5742
rect 63756 4946 63812 4956
rect 64764 5684 64820 5854
rect 63644 4834 63700 4844
rect 62188 4274 62244 4284
rect 63756 4452 63812 4462
rect 61068 4162 61124 4172
rect 59850 3948 60774 3958
rect 59850 3946 59868 3948
rect 59850 3894 59852 3946
rect 59850 3892 59868 3894
rect 59924 3892 59972 3948
rect 60028 3892 60076 3948
rect 60132 3946 60180 3948
rect 60236 3946 60284 3948
rect 60152 3894 60180 3946
rect 60276 3894 60284 3946
rect 60132 3892 60180 3894
rect 60236 3892 60284 3894
rect 60340 3946 60388 3948
rect 60444 3946 60492 3948
rect 60340 3894 60348 3946
rect 60444 3894 60472 3946
rect 60340 3892 60388 3894
rect 60444 3892 60492 3894
rect 60548 3892 60596 3948
rect 60652 3892 60700 3948
rect 60756 3946 60774 3948
rect 60772 3894 60774 3946
rect 60756 3892 60774 3894
rect 59850 3882 60774 3892
rect 60844 3892 60900 3902
rect 57708 3614 57710 3666
rect 57762 3614 57764 3666
rect 57708 3602 57764 3614
rect 59836 3668 59892 3678
rect 59836 3574 59892 3612
rect 60844 3666 60900 3836
rect 60844 3614 60846 3666
rect 60898 3614 60900 3666
rect 60844 3602 60900 3614
rect 62972 3668 63028 3678
rect 62972 3574 63028 3612
rect 53900 3490 53956 3500
rect 57036 3556 57092 3566
rect 57036 3462 57092 3500
rect 63756 3556 63812 4396
rect 63756 3424 63812 3500
rect 64764 3554 64820 5628
rect 65548 5794 65604 5806
rect 65548 5742 65550 5794
rect 65602 5742 65604 5794
rect 65548 3892 65604 5742
rect 66444 5012 66500 9200
rect 68684 5906 68740 5918
rect 68684 5854 68686 5906
rect 68738 5854 68740 5906
rect 67676 5794 67732 5806
rect 67676 5742 67678 5794
rect 67730 5742 67732 5794
rect 66444 4946 66500 4956
rect 66668 5124 66724 5134
rect 65660 4564 65716 4574
rect 65660 4450 65716 4508
rect 65660 4398 65662 4450
rect 65714 4398 65716 4450
rect 65660 4386 65716 4398
rect 66668 4340 66724 5068
rect 67676 5012 67732 5742
rect 67676 4946 67732 4956
rect 66668 4274 66724 4284
rect 68460 4900 68516 4910
rect 65548 3826 65604 3836
rect 65548 3668 65604 3678
rect 65548 3574 65604 3612
rect 67676 3668 67732 3678
rect 67676 3574 67732 3612
rect 68460 3666 68516 4844
rect 68684 4452 68740 5854
rect 68684 4386 68740 4396
rect 68460 3614 68462 3666
rect 68514 3614 68516 3666
rect 68460 3602 68516 3614
rect 69132 3668 69188 9200
rect 69468 5796 69524 5806
rect 69468 5702 69524 5740
rect 70140 5796 70196 5806
rect 69468 5572 69524 5582
rect 69468 5124 69524 5516
rect 70140 5234 70196 5740
rect 71596 5796 71652 5806
rect 71596 5702 71652 5740
rect 70140 5182 70142 5234
rect 70194 5182 70196 5234
rect 70140 5170 70196 5182
rect 69468 5030 69524 5068
rect 71820 5012 71876 9200
rect 72604 5908 72660 5918
rect 71820 4946 71876 4956
rect 72156 5906 72660 5908
rect 72156 5854 72606 5906
rect 72658 5854 72660 5906
rect 72156 5852 72660 5854
rect 72156 5124 72212 5852
rect 72604 5842 72660 5852
rect 73388 5796 73444 5806
rect 70588 4564 70644 4574
rect 70476 4340 70532 4350
rect 70476 4246 70532 4284
rect 69132 3602 69188 3612
rect 70588 3666 70644 4508
rect 70588 3614 70590 3666
rect 70642 3614 70644 3666
rect 70588 3602 70644 3614
rect 71372 3668 71428 3678
rect 64764 3502 64766 3554
rect 64818 3502 64820 3554
rect 64764 3490 64820 3502
rect 71372 3554 71428 3612
rect 72156 3668 72212 5068
rect 72268 5234 72324 5246
rect 72268 5182 72270 5234
rect 72322 5182 72324 5234
rect 72268 5012 72324 5182
rect 73388 5236 73444 5740
rect 73388 5170 73444 5180
rect 74396 5236 74452 5246
rect 74396 5142 74452 5180
rect 73724 5124 73780 5134
rect 73724 5030 73780 5068
rect 72268 4946 72324 4956
rect 74508 5012 74564 9200
rect 76636 5906 76692 5918
rect 76636 5854 76638 5906
rect 76690 5854 76692 5906
rect 75516 5796 75572 5806
rect 75516 5702 75572 5740
rect 74508 4946 74564 4956
rect 76524 5234 76580 5246
rect 76524 5182 76526 5234
rect 76578 5182 76580 5234
rect 76524 5012 76580 5182
rect 76636 5236 76692 5854
rect 77196 5796 77252 9200
rect 79884 6468 79940 9200
rect 79324 6412 79940 6468
rect 77196 5730 77252 5740
rect 77308 5794 77364 5806
rect 77308 5742 77310 5794
rect 77362 5742 77364 5794
rect 76636 5170 76692 5180
rect 76524 4946 76580 4956
rect 77308 5012 77364 5742
rect 72156 3602 72212 3612
rect 73948 4338 74004 4350
rect 73948 4286 73950 4338
rect 74002 4286 74004 4338
rect 71372 3502 71374 3554
rect 71426 3502 71428 3554
rect 71372 3490 71428 3502
rect 50316 3378 50372 3388
rect 40194 3164 41118 3174
rect 40194 3162 40212 3164
rect 40194 3110 40196 3162
rect 40194 3108 40212 3110
rect 40268 3108 40316 3164
rect 40372 3108 40420 3164
rect 40476 3162 40524 3164
rect 40580 3162 40628 3164
rect 40496 3110 40524 3162
rect 40620 3110 40628 3162
rect 40476 3108 40524 3110
rect 40580 3108 40628 3110
rect 40684 3162 40732 3164
rect 40788 3162 40836 3164
rect 40684 3110 40692 3162
rect 40788 3110 40816 3162
rect 40684 3108 40732 3110
rect 40788 3108 40836 3110
rect 40892 3108 40940 3164
rect 40996 3108 41044 3164
rect 41100 3162 41118 3164
rect 41116 3110 41118 3162
rect 41100 3108 41118 3110
rect 40194 3098 41118 3108
rect 73948 1764 74004 4286
rect 76636 3668 76692 3678
rect 76636 3554 76692 3612
rect 77308 3666 77364 4956
rect 78428 4340 78484 4350
rect 78428 4226 78484 4284
rect 78428 4174 78430 4226
rect 78482 4174 78484 4226
rect 78428 4162 78484 4174
rect 77308 3614 77310 3666
rect 77362 3614 77364 3666
rect 77308 3602 77364 3614
rect 79324 3668 79380 6412
rect 79506 6300 80430 6310
rect 79506 6298 79524 6300
rect 79506 6246 79508 6298
rect 79506 6244 79524 6246
rect 79580 6244 79628 6300
rect 79684 6244 79732 6300
rect 79788 6298 79836 6300
rect 79892 6298 79940 6300
rect 79808 6246 79836 6298
rect 79932 6246 79940 6298
rect 79788 6244 79836 6246
rect 79892 6244 79940 6246
rect 79996 6298 80044 6300
rect 80100 6298 80148 6300
rect 79996 6246 80004 6298
rect 80100 6246 80128 6298
rect 79996 6244 80044 6246
rect 80100 6244 80148 6246
rect 80204 6244 80252 6300
rect 80308 6244 80356 6300
rect 80412 6298 80430 6300
rect 80428 6246 80430 6298
rect 80412 6244 80430 6246
rect 79506 6234 80430 6244
rect 80332 5908 80388 5918
rect 79436 5796 79492 5806
rect 79436 5702 79492 5740
rect 80332 5124 80388 5852
rect 80332 5058 80388 5068
rect 81004 5796 81060 5806
rect 79506 4732 80430 4742
rect 79506 4730 79524 4732
rect 79506 4678 79508 4730
rect 79506 4676 79524 4678
rect 79580 4676 79628 4732
rect 79684 4676 79732 4732
rect 79788 4730 79836 4732
rect 79892 4730 79940 4732
rect 79808 4678 79836 4730
rect 79932 4678 79940 4730
rect 79788 4676 79836 4678
rect 79892 4676 79940 4678
rect 79996 4730 80044 4732
rect 80100 4730 80148 4732
rect 79996 4678 80004 4730
rect 80100 4678 80128 4730
rect 79996 4676 80044 4678
rect 80100 4676 80148 4678
rect 80204 4676 80252 4732
rect 80308 4676 80356 4732
rect 80412 4730 80430 4732
rect 80428 4678 80430 4730
rect 80412 4676 80430 4678
rect 79506 4666 80430 4676
rect 79436 3668 79492 3678
rect 79324 3666 79492 3668
rect 79324 3614 79438 3666
rect 79490 3614 79492 3666
rect 79324 3612 79492 3614
rect 79436 3602 79492 3612
rect 81004 3666 81060 5740
rect 82236 5234 82292 5246
rect 82236 5182 82238 5234
rect 82290 5182 82292 5234
rect 82236 5124 82292 5182
rect 82236 5058 82292 5068
rect 81004 3614 81006 3666
rect 81058 3614 81060 3666
rect 81004 3602 81060 3614
rect 82572 3668 82628 9200
rect 84140 5906 84196 5918
rect 84140 5854 84142 5906
rect 84194 5854 84196 5906
rect 83132 5796 83188 5806
rect 83132 5702 83188 5740
rect 84140 5684 84196 5854
rect 83916 5236 83972 5246
rect 83916 5122 83972 5180
rect 83916 5070 83918 5122
rect 83970 5070 83972 5122
rect 83916 4340 83972 5070
rect 83916 4208 83972 4284
rect 82572 3602 82628 3612
rect 83132 3668 83188 3678
rect 83132 3574 83188 3612
rect 76636 3502 76638 3554
rect 76690 3502 76692 3554
rect 76636 3490 76692 3502
rect 80332 3556 80388 3566
rect 80332 3462 80388 3500
rect 84140 3556 84196 5628
rect 84140 3490 84196 3500
rect 84252 5908 84308 5918
rect 84252 3668 84308 5852
rect 84252 3554 84308 3612
rect 84924 5796 84980 5806
rect 84924 3666 84980 5740
rect 85260 5796 85316 9200
rect 85260 5730 85316 5740
rect 87052 5796 87108 5806
rect 87948 5796 88004 9200
rect 88060 5796 88116 5806
rect 87948 5794 88116 5796
rect 87948 5742 88062 5794
rect 88114 5742 88116 5794
rect 87948 5740 88116 5742
rect 87052 5702 87108 5740
rect 88060 5730 88116 5740
rect 90188 5794 90244 5806
rect 90188 5742 90190 5794
rect 90242 5742 90244 5794
rect 86716 5236 86772 5246
rect 86716 5122 86772 5180
rect 86716 5070 86718 5122
rect 86770 5070 86772 5122
rect 86716 5058 86772 5070
rect 89292 5236 89348 5246
rect 88956 5010 89012 5022
rect 88956 4958 88958 5010
rect 89010 4958 89012 5010
rect 88284 4228 88340 4238
rect 88284 4134 88340 4172
rect 84924 3614 84926 3666
rect 84978 3614 84980 3666
rect 84924 3602 84980 3614
rect 87052 3780 87108 3790
rect 87052 3666 87108 3724
rect 88844 3780 88900 3790
rect 87052 3614 87054 3666
rect 87106 3614 87108 3666
rect 87052 3602 87108 3614
rect 88172 3668 88228 3678
rect 84252 3502 84254 3554
rect 84306 3502 84308 3554
rect 84252 3490 84308 3502
rect 88172 3554 88228 3612
rect 88844 3666 88900 3724
rect 88844 3614 88846 3666
rect 88898 3614 88900 3666
rect 88844 3602 88900 3614
rect 88172 3502 88174 3554
rect 88226 3502 88228 3554
rect 88172 3490 88228 3502
rect 88956 3556 89012 4958
rect 89292 4338 89348 5180
rect 89292 4286 89294 4338
rect 89346 4286 89348 4338
rect 89292 4274 89348 4286
rect 90188 3780 90244 5742
rect 90636 5796 90692 9200
rect 90636 5730 90692 5740
rect 90972 5908 91028 5918
rect 90972 5684 91028 5852
rect 91980 5796 92036 5806
rect 91980 5702 92036 5740
rect 90972 5618 91028 5628
rect 93212 5236 93268 5246
rect 93324 5236 93380 9200
rect 94892 5908 94948 5918
rect 94892 5814 94948 5852
rect 93212 5234 93380 5236
rect 93212 5182 93214 5234
rect 93266 5182 93380 5234
rect 93212 5180 93380 5182
rect 94108 5794 94164 5806
rect 94108 5742 94110 5794
rect 94162 5742 94164 5794
rect 93212 5170 93268 5180
rect 92092 4228 92148 4238
rect 90188 3714 90244 3724
rect 90972 3892 91028 3902
rect 90972 3666 91028 3836
rect 90972 3614 90974 3666
rect 91026 3614 91028 3666
rect 90972 3602 91028 3614
rect 92092 3780 92148 4172
rect 93996 4228 94052 4238
rect 88956 3490 89012 3500
rect 92092 3554 92148 3724
rect 92764 3892 92820 3902
rect 92764 3666 92820 3836
rect 92764 3614 92766 3666
rect 92818 3614 92820 3666
rect 92764 3602 92820 3614
rect 93996 3668 94052 4172
rect 94108 3892 94164 5742
rect 95900 5796 95956 5806
rect 96012 5796 96068 9200
rect 98700 6804 98756 9200
rect 98588 6748 98756 6804
rect 95900 5794 96068 5796
rect 95900 5742 95902 5794
rect 95954 5742 96068 5794
rect 95900 5740 96068 5742
rect 96124 5908 96180 5918
rect 95900 5730 95956 5740
rect 96124 5122 96180 5852
rect 98028 5794 98084 5806
rect 98028 5742 98030 5794
rect 98082 5742 98084 5794
rect 96124 5070 96126 5122
rect 96178 5070 96180 5122
rect 96124 5058 96180 5070
rect 96684 5124 96740 5134
rect 96684 5030 96740 5068
rect 94108 3826 94164 3836
rect 95340 5010 95396 5022
rect 95340 4958 95342 5010
rect 95394 4958 95396 5010
rect 93996 3602 94052 3612
rect 94892 3668 94948 3678
rect 94892 3574 94948 3612
rect 95340 3668 95396 4958
rect 97468 5010 97524 5022
rect 97468 4958 97470 5010
rect 97522 4958 97524 5010
rect 97244 4340 97300 4350
rect 97244 4226 97300 4284
rect 97244 4174 97246 4226
rect 97298 4174 97300 4226
rect 97244 4162 97300 4174
rect 95340 3602 95396 3612
rect 96684 3668 96740 3678
rect 97468 3668 97524 4958
rect 98028 3668 98084 5742
rect 98588 4340 98644 6748
rect 98812 5908 98868 5918
rect 98812 5814 98868 5852
rect 100156 5908 100212 5918
rect 99820 5796 99876 5806
rect 99820 5702 99876 5740
rect 99162 5516 100086 5526
rect 99162 5514 99180 5516
rect 99162 5462 99164 5514
rect 99162 5460 99180 5462
rect 99236 5460 99284 5516
rect 99340 5460 99388 5516
rect 99444 5514 99492 5516
rect 99548 5514 99596 5516
rect 99464 5462 99492 5514
rect 99588 5462 99596 5514
rect 99444 5460 99492 5462
rect 99548 5460 99596 5462
rect 99652 5514 99700 5516
rect 99756 5514 99804 5516
rect 99652 5462 99660 5514
rect 99756 5462 99784 5514
rect 99652 5460 99700 5462
rect 99756 5460 99804 5462
rect 99860 5460 99908 5516
rect 99964 5460 100012 5516
rect 100068 5514 100086 5516
rect 100084 5462 100086 5514
rect 100068 5460 100086 5462
rect 99162 5450 100086 5460
rect 98588 4274 98644 4284
rect 99596 5234 99652 5246
rect 99596 5182 99598 5234
rect 99650 5182 99652 5234
rect 99372 4226 99428 4238
rect 99372 4174 99374 4226
rect 99426 4174 99428 4226
rect 99372 4116 99428 4174
rect 99596 4116 99652 5182
rect 100156 4338 100212 5852
rect 101388 5796 101444 9200
rect 102732 5908 102788 5918
rect 102732 5814 102788 5852
rect 103964 5908 104020 5918
rect 103964 5814 104020 5852
rect 101388 5730 101444 5740
rect 101948 5794 102004 5806
rect 101948 5742 101950 5794
rect 102002 5742 102004 5794
rect 101948 5236 102004 5742
rect 104076 5796 104132 9200
rect 104076 5730 104132 5740
rect 104748 5794 104804 5806
rect 104748 5742 104750 5794
rect 104802 5742 104804 5794
rect 101948 5170 102004 5180
rect 102732 5236 102788 5246
rect 102620 5124 102676 5134
rect 102620 5030 102676 5068
rect 100156 4286 100158 4338
rect 100210 4286 100212 4338
rect 100156 4274 100212 4286
rect 99372 4060 100212 4116
rect 99162 3948 100086 3958
rect 99162 3946 99180 3948
rect 99162 3894 99164 3946
rect 99162 3892 99180 3894
rect 99236 3892 99284 3948
rect 99340 3892 99388 3948
rect 99444 3946 99492 3948
rect 99548 3946 99596 3948
rect 99464 3894 99492 3946
rect 99588 3894 99596 3946
rect 99444 3892 99492 3894
rect 99548 3892 99596 3894
rect 99652 3946 99700 3948
rect 99756 3946 99804 3948
rect 99652 3894 99660 3946
rect 99756 3894 99784 3946
rect 99652 3892 99700 3894
rect 99756 3892 99804 3894
rect 99860 3892 99908 3948
rect 99964 3892 100012 3948
rect 100068 3946 100086 3948
rect 100084 3894 100086 3946
rect 100068 3892 100086 3894
rect 99162 3882 100086 3892
rect 98812 3668 98868 3678
rect 97468 3666 98868 3668
rect 97468 3614 98814 3666
rect 98866 3614 98868 3666
rect 97468 3612 98868 3614
rect 100156 3668 100212 4060
rect 100604 3668 100660 3678
rect 100156 3666 100660 3668
rect 100156 3614 100606 3666
rect 100658 3614 100660 3666
rect 100156 3612 100660 3614
rect 96684 3574 96740 3612
rect 98812 3602 98868 3612
rect 100604 3602 100660 3612
rect 102732 3666 102788 5180
rect 103292 5236 103348 5246
rect 103292 5142 103348 5180
rect 104748 4452 104804 5742
rect 106764 5796 106820 9200
rect 107772 5908 107828 5918
rect 106876 5796 106932 5806
rect 106764 5794 106932 5796
rect 106764 5742 106878 5794
rect 106930 5742 106932 5794
rect 106764 5740 106932 5742
rect 106876 5730 106932 5740
rect 107660 5796 107716 5806
rect 107660 5702 107716 5740
rect 105420 5236 105476 5246
rect 105420 5142 105476 5180
rect 107772 5012 107828 5852
rect 104748 4386 104804 4396
rect 105980 4452 106036 4462
rect 105980 4358 106036 4396
rect 102732 3614 102734 3666
rect 102786 3614 102788 3666
rect 102732 3602 102788 3614
rect 105308 4340 105364 4350
rect 92092 3502 92094 3554
rect 92146 3502 92148 3554
rect 92092 3490 92148 3502
rect 95900 3556 95956 3566
rect 95900 3462 95956 3500
rect 99820 3556 99876 3566
rect 99820 3462 99876 3500
rect 105308 3444 105364 4284
rect 107772 3554 107828 4956
rect 109116 5234 109172 5246
rect 109116 5182 109118 5234
rect 109170 5182 109172 5234
rect 109116 4564 109172 5182
rect 109452 4676 109508 9200
rect 111580 6690 111636 6702
rect 111580 6638 111582 6690
rect 111634 6638 111636 6690
rect 110572 5906 110628 5918
rect 110572 5854 110574 5906
rect 110626 5854 110628 5906
rect 109788 5794 109844 5806
rect 109788 5742 109790 5794
rect 109842 5742 109844 5794
rect 109788 5572 109844 5742
rect 109788 5506 109844 5516
rect 110572 5012 110628 5854
rect 111580 5794 111636 6638
rect 112140 6690 112196 9200
rect 112140 6638 112142 6690
rect 112194 6638 112196 6690
rect 112140 6626 112196 6638
rect 114380 5906 114436 5918
rect 114380 5854 114382 5906
rect 114434 5854 114436 5906
rect 111580 5742 111582 5794
rect 111634 5742 111636 5794
rect 111580 5730 111636 5742
rect 111916 5796 111972 5806
rect 111244 5572 111300 5582
rect 111244 5234 111300 5516
rect 111244 5182 111246 5234
rect 111298 5182 111300 5234
rect 111244 5170 111300 5182
rect 111580 5348 111636 5358
rect 110572 4946 110628 4956
rect 109452 4610 109508 4620
rect 110572 4676 110628 4686
rect 109116 4498 109172 4508
rect 108108 4452 108164 4462
rect 108108 4226 108164 4396
rect 108108 4174 108110 4226
rect 108162 4174 108164 4226
rect 108108 4162 108164 4174
rect 108444 4452 108500 4462
rect 108444 3666 108500 4396
rect 109452 4452 109508 4462
rect 109452 4358 109508 4396
rect 108780 4340 108836 4350
rect 108780 4246 108836 4284
rect 108444 3614 108446 3666
rect 108498 3614 108500 3666
rect 108444 3602 108500 3614
rect 110572 3666 110628 4620
rect 111580 4226 111636 5292
rect 111580 4174 111582 4226
rect 111634 4174 111636 4226
rect 111580 4162 111636 4174
rect 111916 5122 111972 5740
rect 113708 5794 113764 5806
rect 113708 5742 113710 5794
rect 113762 5742 113764 5794
rect 111916 5070 111918 5122
rect 111970 5070 111972 5122
rect 111916 4228 111972 5070
rect 111916 4162 111972 4172
rect 112364 5348 112420 5358
rect 110572 3614 110574 3666
rect 110626 3614 110628 3666
rect 110572 3602 110628 3614
rect 111580 3780 111636 3790
rect 107772 3502 107774 3554
rect 107826 3502 107828 3554
rect 107772 3490 107828 3502
rect 111580 3556 111636 3724
rect 112364 3666 112420 5292
rect 113708 5348 113764 5742
rect 113708 5282 113764 5292
rect 113372 5236 113428 5246
rect 113372 5142 113428 5180
rect 112700 5124 112756 5134
rect 112700 5030 112756 5068
rect 114380 5012 114436 5854
rect 114380 4946 114436 4956
rect 114492 5236 114548 5246
rect 113148 4228 113204 4238
rect 113148 4134 113204 4172
rect 112364 3614 112366 3666
rect 112418 3614 112420 3666
rect 112364 3602 112420 3614
rect 114492 3666 114548 5180
rect 114828 4228 114884 9200
rect 115612 5906 115668 5918
rect 115612 5854 115614 5906
rect 115666 5854 115668 5906
rect 115612 5796 115668 5854
rect 115612 5730 115668 5740
rect 116284 5794 116340 5806
rect 116284 5742 116286 5794
rect 116338 5742 116340 5794
rect 115388 5572 115444 5582
rect 115276 5236 115332 5246
rect 115276 4450 115332 5180
rect 115276 4398 115278 4450
rect 115330 4398 115332 4450
rect 115276 4386 115332 4398
rect 114828 4162 114884 4172
rect 114492 3614 114494 3666
rect 114546 3614 114548 3666
rect 114492 3602 114548 3614
rect 115388 3668 115444 5516
rect 115500 5348 115556 5358
rect 115500 5234 115556 5292
rect 115500 5182 115502 5234
rect 115554 5182 115556 5234
rect 115500 5170 115556 5182
rect 116284 5236 116340 5742
rect 116284 5170 116340 5180
rect 117068 5124 117124 5134
rect 117068 5030 117124 5068
rect 116060 5012 116116 5022
rect 116060 4338 116116 4956
rect 116060 4286 116062 4338
rect 116114 4286 116116 4338
rect 116060 3892 116116 4286
rect 116620 4228 116676 4238
rect 116620 4134 116676 4172
rect 117516 4228 117572 9200
rect 120204 6468 120260 9200
rect 120092 6412 120260 6468
rect 118818 6300 119742 6310
rect 118818 6298 118836 6300
rect 118818 6246 118820 6298
rect 118818 6244 118836 6246
rect 118892 6244 118940 6300
rect 118996 6244 119044 6300
rect 119100 6298 119148 6300
rect 119204 6298 119252 6300
rect 119120 6246 119148 6298
rect 119244 6246 119252 6298
rect 119100 6244 119148 6246
rect 119204 6244 119252 6246
rect 119308 6298 119356 6300
rect 119412 6298 119460 6300
rect 119308 6246 119316 6298
rect 119412 6246 119440 6298
rect 119308 6244 119356 6246
rect 119412 6244 119460 6246
rect 119516 6244 119564 6300
rect 119620 6244 119668 6300
rect 119724 6298 119742 6300
rect 119740 6246 119742 6298
rect 119724 6244 119742 6246
rect 118818 6234 119742 6244
rect 118412 5908 118468 5918
rect 118412 5794 118468 5852
rect 118412 5742 118414 5794
rect 118466 5742 118468 5794
rect 118412 5730 118468 5742
rect 118636 5908 118692 5918
rect 117852 5236 117908 5246
rect 117852 5142 117908 5180
rect 117516 4162 117572 4172
rect 117628 4900 117684 4910
rect 116060 3826 116116 3836
rect 115500 3668 115556 3678
rect 115388 3666 115556 3668
rect 115388 3614 115502 3666
rect 115554 3614 115556 3666
rect 115388 3612 115556 3614
rect 115500 3602 115556 3612
rect 117628 3666 117684 4844
rect 118636 4452 118692 5852
rect 119532 5906 119588 5918
rect 119532 5854 119534 5906
rect 119586 5854 119588 5906
rect 119532 5796 119588 5854
rect 119532 5730 119588 5740
rect 119980 5234 120036 5246
rect 119980 5182 119982 5234
rect 120034 5182 120036 5234
rect 119980 5012 120036 5182
rect 119980 4946 120036 4956
rect 118818 4732 119742 4742
rect 118818 4730 118836 4732
rect 118818 4678 118820 4730
rect 118818 4676 118836 4678
rect 118892 4676 118940 4732
rect 118996 4676 119044 4732
rect 119100 4730 119148 4732
rect 119204 4730 119252 4732
rect 119120 4678 119148 4730
rect 119244 4678 119252 4730
rect 119100 4676 119148 4678
rect 119204 4676 119252 4678
rect 119308 4730 119356 4732
rect 119412 4730 119460 4732
rect 119308 4678 119316 4730
rect 119412 4678 119440 4730
rect 119308 4676 119356 4678
rect 119412 4676 119460 4678
rect 119516 4676 119564 4732
rect 119620 4676 119668 4732
rect 119724 4730 119742 4732
rect 119740 4678 119742 4730
rect 119724 4676 119742 4678
rect 118818 4666 119742 4676
rect 118748 4452 118804 4462
rect 118636 4450 118804 4452
rect 118636 4398 118750 4450
rect 118802 4398 118804 4450
rect 118636 4396 118804 4398
rect 118748 4386 118804 4396
rect 117628 3614 117630 3666
rect 117682 3614 117684 3666
rect 117628 3602 117684 3614
rect 118412 4340 118468 4350
rect 111580 3424 111636 3500
rect 118412 3554 118468 4284
rect 119532 4338 119588 4350
rect 119532 4286 119534 4338
rect 119586 4286 119588 4338
rect 119532 3892 119588 4286
rect 119532 3826 119588 3836
rect 119420 3668 119476 3678
rect 119420 3574 119476 3612
rect 120092 3668 120148 6412
rect 120204 5908 120260 5918
rect 120204 5814 120260 5852
rect 122332 5796 122388 5806
rect 121884 5794 122388 5796
rect 121884 5742 122334 5794
rect 122386 5742 122388 5794
rect 121884 5740 122388 5742
rect 121324 5460 121380 5470
rect 121324 5234 121380 5404
rect 121324 5182 121326 5234
rect 121378 5182 121380 5234
rect 121324 5170 121380 5182
rect 120652 5122 120708 5134
rect 120652 5070 120654 5122
rect 120706 5070 120708 5122
rect 120652 3892 120708 5070
rect 121884 4452 121940 5740
rect 122332 5730 122388 5740
rect 121548 4450 121940 4452
rect 121548 4398 121886 4450
rect 121938 4398 121940 4450
rect 121548 4396 121940 4398
rect 121212 4340 121268 4350
rect 121212 4246 121268 4284
rect 120652 3826 120708 3836
rect 120092 3602 120148 3612
rect 121548 3666 121604 4396
rect 121884 4386 121940 4396
rect 121548 3614 121550 3666
rect 121602 3614 121604 3666
rect 121548 3602 121604 3614
rect 122332 3892 122388 3902
rect 118412 3502 118414 3554
rect 118466 3502 118468 3554
rect 118412 3490 118468 3502
rect 122332 3554 122388 3836
rect 122892 3668 122948 9200
rect 123340 5908 123396 5918
rect 123340 5124 123396 5852
rect 124124 5794 124180 5806
rect 124124 5742 124126 5794
rect 124178 5742 124180 5794
rect 123340 5058 123396 5068
rect 123452 5234 123508 5246
rect 123452 5182 123454 5234
rect 123506 5182 123508 5234
rect 123452 4564 123508 5182
rect 123452 4498 123508 4508
rect 124124 5012 124180 5742
rect 124012 4228 124068 4238
rect 124012 4134 124068 4172
rect 124124 3780 124180 4956
rect 125020 5234 125076 5246
rect 125020 5182 125022 5234
rect 125074 5182 125076 5234
rect 125020 4900 125076 5182
rect 125580 5012 125636 9200
rect 127932 6020 127988 6030
rect 127260 5906 127316 5918
rect 127260 5854 127262 5906
rect 127314 5854 127316 5906
rect 126252 5794 126308 5806
rect 126252 5742 126254 5794
rect 126306 5742 126308 5794
rect 126252 5684 126308 5742
rect 126252 5618 126308 5628
rect 127148 5684 127204 5694
rect 127148 5234 127204 5628
rect 127148 5182 127150 5234
rect 127202 5182 127204 5234
rect 127148 5170 127204 5182
rect 125580 4946 125636 4956
rect 125020 4834 125076 4844
rect 124124 3714 124180 3724
rect 124572 4338 124628 4350
rect 124572 4286 124574 4338
rect 124626 4286 124628 4338
rect 122892 3602 122948 3612
rect 123340 3668 123396 3678
rect 123340 3574 123396 3612
rect 122332 3502 122334 3554
rect 122386 3502 122388 3554
rect 122332 3490 122388 3502
rect 124572 3556 124628 4286
rect 125356 4228 125412 4238
rect 125356 3668 125412 4172
rect 126140 3892 126196 3902
rect 125468 3668 125524 3678
rect 125356 3666 125524 3668
rect 125356 3614 125470 3666
rect 125522 3614 125524 3666
rect 125356 3612 125524 3614
rect 125468 3602 125524 3612
rect 124572 3490 124628 3500
rect 126140 3554 126196 3836
rect 127260 3892 127316 5854
rect 127932 5796 127988 5964
rect 127932 5122 127988 5740
rect 128044 5794 128100 5806
rect 128044 5742 128046 5794
rect 128098 5742 128100 5794
rect 128044 5236 128100 5742
rect 128044 5170 128100 5180
rect 127932 5070 127934 5122
rect 127986 5070 127988 5122
rect 127932 5058 127988 5070
rect 128268 4452 128324 9200
rect 130172 5794 130228 5806
rect 130172 5742 130174 5794
rect 130226 5742 130228 5794
rect 128492 5234 128548 5246
rect 128492 5182 128494 5234
rect 128546 5182 128548 5234
rect 128492 5012 128548 5182
rect 128492 4946 128548 4956
rect 130172 4788 130228 5742
rect 130172 4722 130228 4732
rect 130620 5010 130676 5022
rect 130620 4958 130622 5010
rect 130674 4958 130676 5010
rect 128268 4386 128324 4396
rect 129052 4452 129108 4462
rect 127484 4228 127540 4238
rect 127484 4134 127540 4172
rect 128044 4228 128100 4238
rect 127260 3826 127316 3836
rect 128044 3666 128100 4172
rect 129052 4226 129108 4396
rect 129052 4174 129054 4226
rect 129106 4174 129108 4226
rect 129052 4162 129108 4174
rect 130172 4452 130228 4462
rect 128044 3614 128046 3666
rect 128098 3614 128100 3666
rect 128044 3602 128100 3614
rect 130172 3666 130228 4396
rect 130620 4228 130676 4958
rect 130620 4162 130676 4172
rect 130956 4228 131012 9200
rect 131292 6020 131348 6030
rect 131292 5906 131348 5964
rect 131292 5854 131294 5906
rect 131346 5854 131348 5906
rect 131292 5842 131348 5854
rect 132972 5908 133028 5918
rect 131964 5794 132020 5806
rect 131964 5742 131966 5794
rect 132018 5742 132020 5794
rect 131292 5122 131348 5134
rect 131292 5070 131294 5122
rect 131346 5070 131348 5122
rect 131292 5012 131348 5070
rect 131180 4452 131236 4462
rect 131180 4358 131236 4396
rect 130956 4162 131012 4172
rect 130172 3614 130174 3666
rect 130226 3614 130228 3666
rect 130172 3602 130228 3614
rect 131180 3892 131236 3902
rect 131292 3892 131348 4956
rect 131964 4452 132020 5742
rect 132972 5122 133028 5852
rect 132972 5070 132974 5122
rect 133026 5070 133028 5122
rect 132972 5058 133028 5070
rect 131964 4386 132020 4396
rect 131236 3836 131348 3892
rect 131852 4338 131908 4350
rect 131852 4286 131854 4338
rect 131906 4286 131908 4338
rect 131852 3892 131908 4286
rect 132524 4228 132580 4238
rect 132524 4134 132580 4172
rect 133644 4228 133700 9200
rect 135100 5906 135156 5918
rect 135100 5854 135102 5906
rect 135154 5854 135156 5906
rect 134092 5794 134148 5806
rect 134092 5742 134094 5794
rect 134146 5742 134148 5794
rect 133756 5124 133812 5134
rect 133756 5030 133812 5068
rect 134092 5124 134148 5742
rect 134092 5058 134148 5068
rect 134652 5124 134708 5134
rect 134652 4450 134708 5068
rect 135100 5012 135156 5854
rect 135884 5794 135940 5806
rect 135884 5742 135886 5794
rect 135938 5742 135940 5794
rect 135884 5684 135940 5742
rect 135884 5618 135940 5628
rect 135884 5234 135940 5246
rect 135884 5182 135886 5234
rect 135938 5182 135940 5234
rect 135156 4956 135380 5012
rect 135100 4946 135156 4956
rect 134652 4398 134654 4450
rect 134706 4398 134708 4450
rect 134652 4386 134708 4398
rect 135324 4676 135380 4956
rect 135324 4338 135380 4620
rect 135324 4286 135326 4338
rect 135378 4286 135380 4338
rect 135324 4274 135380 4286
rect 133644 4162 133700 4172
rect 126140 3502 126142 3554
rect 126194 3502 126196 3554
rect 126140 3490 126196 3502
rect 127372 3556 127428 3566
rect 127372 3462 127428 3500
rect 131180 3554 131236 3836
rect 131852 3826 131908 3836
rect 135884 4116 135940 5182
rect 136332 5012 136388 9200
rect 139020 6132 139076 9200
rect 139020 6076 139188 6132
rect 139020 5908 139076 5918
rect 139020 5814 139076 5852
rect 138012 5796 138068 5806
rect 138012 5794 138180 5796
rect 138012 5742 138014 5794
rect 138066 5742 138180 5794
rect 138012 5740 138180 5742
rect 138012 5730 138068 5740
rect 138012 5348 138068 5358
rect 136332 4946 136388 4956
rect 136444 5122 136500 5134
rect 136444 5070 136446 5122
rect 136498 5070 136500 5122
rect 131964 3780 132020 3790
rect 131964 3666 132020 3724
rect 131964 3614 131966 3666
rect 132018 3614 132020 3666
rect 131964 3602 132020 3614
rect 134092 3780 134148 3790
rect 134092 3666 134148 3724
rect 134092 3614 134094 3666
rect 134146 3614 134148 3666
rect 134092 3602 134148 3614
rect 135884 3666 135940 4060
rect 136444 4676 136500 5070
rect 137228 5010 137284 5022
rect 137228 4958 137230 5010
rect 137282 4958 137284 5010
rect 137228 4900 137284 4958
rect 137228 4834 137284 4844
rect 136444 4004 136500 4620
rect 137004 4228 137060 4238
rect 137004 4134 137060 4172
rect 136444 3938 136500 3948
rect 135884 3614 135886 3666
rect 135938 3614 135940 3666
rect 135884 3602 135940 3614
rect 138012 3666 138068 5292
rect 138124 4676 138180 5740
rect 139132 5684 139188 6076
rect 139804 5794 139860 5806
rect 139804 5742 139806 5794
rect 139858 5742 139860 5794
rect 139132 5628 139524 5684
rect 138474 5516 139398 5526
rect 138474 5514 138492 5516
rect 138474 5462 138476 5514
rect 138474 5460 138492 5462
rect 138548 5460 138596 5516
rect 138652 5460 138700 5516
rect 138756 5514 138804 5516
rect 138860 5514 138908 5516
rect 138776 5462 138804 5514
rect 138900 5462 138908 5514
rect 138756 5460 138804 5462
rect 138860 5460 138908 5462
rect 138964 5514 139012 5516
rect 139068 5514 139116 5516
rect 138964 5462 138972 5514
rect 139068 5462 139096 5514
rect 138964 5460 139012 5462
rect 139068 5460 139116 5462
rect 139172 5460 139220 5516
rect 139276 5460 139324 5516
rect 139380 5514 139398 5516
rect 139396 5462 139398 5514
rect 139380 5460 139398 5462
rect 138474 5450 139398 5460
rect 139356 5234 139412 5246
rect 139356 5182 139358 5234
rect 139410 5182 139412 5234
rect 139356 4900 139412 5182
rect 139356 4834 139412 4844
rect 138124 4610 138180 4620
rect 138012 3614 138014 3666
rect 138066 3614 138068 3666
rect 138012 3602 138068 3614
rect 138348 4340 138404 4350
rect 131180 3502 131182 3554
rect 131234 3502 131236 3554
rect 131180 3490 131236 3502
rect 135100 3556 135156 3566
rect 135100 3462 135156 3500
rect 138348 3556 138404 4284
rect 139132 4228 139188 4238
rect 139132 4134 139188 4172
rect 139468 4228 139524 5628
rect 139804 5348 139860 5742
rect 141708 5796 141764 9200
rect 143836 5908 143892 5918
rect 141708 5730 141764 5740
rect 141932 5796 141988 5806
rect 142940 5796 142996 5806
rect 141932 5794 142100 5796
rect 141932 5742 141934 5794
rect 141986 5742 142100 5794
rect 141932 5740 142100 5742
rect 141932 5730 141988 5740
rect 139804 5282 139860 5292
rect 140924 5234 140980 5246
rect 140924 5182 140926 5234
rect 140978 5182 140980 5234
rect 140924 5012 140980 5182
rect 140924 4946 140980 4956
rect 141932 5124 141988 5134
rect 139468 4162 139524 4172
rect 139804 4338 139860 4350
rect 139804 4286 139806 4338
rect 139858 4286 139860 4338
rect 139804 4116 139860 4286
rect 140476 4228 140532 4238
rect 140476 4134 140532 4172
rect 139804 4050 139860 4060
rect 138474 3948 139398 3958
rect 138474 3946 138492 3948
rect 138474 3894 138476 3946
rect 138474 3892 138492 3894
rect 138548 3892 138596 3948
rect 138652 3892 138700 3948
rect 138756 3946 138804 3948
rect 138860 3946 138908 3948
rect 138776 3894 138804 3946
rect 138900 3894 138908 3946
rect 138756 3892 138804 3894
rect 138860 3892 138908 3894
rect 138964 3946 139012 3948
rect 139068 3946 139116 3948
rect 138964 3894 138972 3946
rect 139068 3894 139096 3946
rect 138964 3892 139012 3894
rect 139068 3892 139116 3894
rect 139172 3892 139220 3948
rect 139276 3892 139324 3948
rect 139380 3946 139398 3948
rect 139396 3894 139398 3946
rect 139380 3892 139398 3894
rect 138474 3882 139398 3892
rect 139804 3668 139860 3678
rect 139804 3574 139860 3612
rect 141932 3666 141988 5068
rect 141932 3614 141934 3666
rect 141986 3614 141988 3666
rect 141932 3602 141988 3614
rect 142044 3668 142100 5740
rect 142940 5702 142996 5740
rect 143052 5348 143108 5358
rect 143052 5234 143108 5292
rect 143052 5182 143054 5234
rect 143106 5182 143108 5234
rect 143052 5170 143108 5182
rect 143836 5122 143892 5852
rect 143836 5070 143838 5122
rect 143890 5070 143892 5122
rect 143724 4452 143780 4462
rect 143276 4338 143332 4350
rect 143276 4286 143278 4338
rect 143330 4286 143332 4338
rect 142044 3602 142100 3612
rect 142604 4226 142660 4238
rect 142604 4174 142606 4226
rect 142658 4174 142660 4226
rect 142604 3668 142660 4174
rect 142604 3602 142660 3612
rect 142940 4116 142996 4126
rect 138348 3490 138404 3500
rect 139020 3556 139076 3566
rect 139020 3462 139076 3500
rect 142940 3554 142996 4060
rect 143276 4116 143332 4286
rect 143276 4050 143332 4060
rect 143724 3666 143780 4396
rect 143836 4116 143892 5070
rect 143836 4050 143892 4060
rect 143724 3614 143726 3666
rect 143778 3614 143780 3666
rect 143724 3602 143780 3614
rect 144396 3668 144452 9200
rect 144508 6020 144564 6030
rect 144508 5122 144564 5964
rect 145740 5908 145796 5918
rect 145740 5814 145796 5852
rect 145068 5796 145124 5806
rect 145068 5794 145236 5796
rect 145068 5742 145070 5794
rect 145122 5742 145236 5794
rect 145068 5740 145236 5742
rect 145068 5730 145124 5740
rect 144508 5070 144510 5122
rect 144562 5070 144564 5122
rect 144508 5058 144564 5070
rect 145180 5124 145236 5740
rect 145180 5030 145236 5068
rect 147084 4564 147140 9200
rect 147084 4498 147140 4508
rect 147308 5234 147364 5246
rect 147308 5182 147310 5234
rect 147362 5182 147364 5234
rect 147308 5012 147364 5182
rect 147308 4452 147364 4956
rect 149772 4788 149828 9200
rect 149772 4722 149828 4732
rect 147308 4386 147364 4396
rect 152460 3780 152516 9200
rect 155148 4676 155204 9200
rect 157836 4900 157892 9200
rect 158130 6300 159054 6310
rect 158130 6298 158148 6300
rect 158130 6246 158132 6298
rect 158130 6244 158148 6246
rect 158204 6244 158252 6300
rect 158308 6244 158356 6300
rect 158412 6298 158460 6300
rect 158516 6298 158564 6300
rect 158432 6246 158460 6298
rect 158556 6246 158564 6298
rect 158412 6244 158460 6246
rect 158516 6244 158564 6246
rect 158620 6298 158668 6300
rect 158724 6298 158772 6300
rect 158620 6246 158628 6298
rect 158724 6246 158752 6298
rect 158620 6244 158668 6246
rect 158724 6244 158772 6246
rect 158828 6244 158876 6300
rect 158932 6244 158980 6300
rect 159036 6298 159054 6300
rect 159052 6246 159054 6298
rect 159036 6244 159054 6246
rect 158130 6234 159054 6244
rect 157836 4834 157892 4844
rect 158130 4732 159054 4742
rect 158130 4730 158148 4732
rect 158130 4678 158132 4730
rect 158130 4676 158148 4678
rect 158204 4676 158252 4732
rect 158308 4676 158356 4732
rect 158412 4730 158460 4732
rect 158516 4730 158564 4732
rect 158432 4678 158460 4730
rect 158556 4678 158564 4730
rect 158412 4676 158460 4678
rect 158516 4676 158564 4678
rect 158620 4730 158668 4732
rect 158724 4730 158772 4732
rect 158620 4678 158628 4730
rect 158724 4678 158752 4730
rect 158620 4676 158668 4678
rect 158724 4676 158772 4678
rect 158828 4676 158876 4732
rect 158932 4676 158980 4732
rect 159036 4730 159054 4732
rect 159052 4678 159054 4730
rect 159036 4676 159054 4678
rect 158130 4666 159054 4676
rect 155148 4610 155204 4620
rect 152460 3714 152516 3724
rect 144396 3602 144452 3612
rect 145852 3668 145908 3678
rect 145852 3574 145908 3612
rect 142940 3502 142942 3554
rect 142994 3502 142996 3554
rect 142940 3490 142996 3502
rect 105308 3378 105364 3388
rect 79506 3164 80430 3174
rect 79506 3162 79524 3164
rect 79506 3110 79508 3162
rect 79506 3108 79524 3110
rect 79580 3108 79628 3164
rect 79684 3108 79732 3164
rect 79788 3162 79836 3164
rect 79892 3162 79940 3164
rect 79808 3110 79836 3162
rect 79932 3110 79940 3162
rect 79788 3108 79836 3110
rect 79892 3108 79940 3110
rect 79996 3162 80044 3164
rect 80100 3162 80148 3164
rect 79996 3110 80004 3162
rect 80100 3110 80128 3162
rect 79996 3108 80044 3110
rect 80100 3108 80148 3110
rect 80204 3108 80252 3164
rect 80308 3108 80356 3164
rect 80412 3162 80430 3164
rect 80428 3110 80430 3162
rect 80412 3108 80430 3110
rect 79506 3098 80430 3108
rect 118818 3164 119742 3174
rect 118818 3162 118836 3164
rect 118818 3110 118820 3162
rect 118818 3108 118836 3110
rect 118892 3108 118940 3164
rect 118996 3108 119044 3164
rect 119100 3162 119148 3164
rect 119204 3162 119252 3164
rect 119120 3110 119148 3162
rect 119244 3110 119252 3162
rect 119100 3108 119148 3110
rect 119204 3108 119252 3110
rect 119308 3162 119356 3164
rect 119412 3162 119460 3164
rect 119308 3110 119316 3162
rect 119412 3110 119440 3162
rect 119308 3108 119356 3110
rect 119412 3108 119460 3110
rect 119516 3108 119564 3164
rect 119620 3108 119668 3164
rect 119724 3162 119742 3164
rect 119740 3110 119742 3162
rect 119724 3108 119742 3110
rect 118818 3098 119742 3108
rect 158130 3164 159054 3174
rect 158130 3162 158148 3164
rect 158130 3110 158132 3162
rect 158130 3108 158148 3110
rect 158204 3108 158252 3164
rect 158308 3108 158356 3164
rect 158412 3162 158460 3164
rect 158516 3162 158564 3164
rect 158432 3110 158460 3162
rect 158556 3110 158564 3162
rect 158412 3108 158460 3110
rect 158516 3108 158564 3110
rect 158620 3162 158668 3164
rect 158724 3162 158772 3164
rect 158620 3110 158628 3162
rect 158724 3110 158752 3162
rect 158620 3108 158668 3110
rect 158724 3108 158772 3110
rect 158828 3108 158876 3164
rect 158932 3108 158980 3164
rect 159036 3162 159054 3164
rect 159052 3110 159054 3162
rect 159036 3108 159054 3110
rect 158130 3098 159054 3108
rect 73948 1698 74004 1708
<< via2 >>
rect 2044 8204 2100 8260
rect 2156 5740 2212 5796
rect 2044 5122 2100 5124
rect 2044 5070 2046 5122
rect 2046 5070 2098 5122
rect 2098 5070 2100 5122
rect 2044 5068 2100 5070
rect 5964 5964 6020 6020
rect 4732 5068 4788 5124
rect 4172 4172 4228 4228
rect 4732 4226 4788 4228
rect 4732 4174 4734 4226
rect 4734 4174 4786 4226
rect 4786 4174 4788 4226
rect 4732 4172 4788 4174
rect 6524 5122 6580 5124
rect 6524 5070 6526 5122
rect 6526 5070 6578 5122
rect 6578 5070 6580 5122
rect 6524 5068 6580 5070
rect 7308 5122 7364 5124
rect 7308 5070 7310 5122
rect 7310 5070 7362 5122
rect 7362 5070 7364 5122
rect 7308 5068 7364 5070
rect 5068 4396 5124 4452
rect 6636 4396 6692 4452
rect 5516 4338 5572 4340
rect 5516 4286 5518 4338
rect 5518 4286 5570 4338
rect 5570 4286 5572 4338
rect 5516 4284 5572 4286
rect 6188 4338 6244 4340
rect 6188 4286 6190 4338
rect 6190 4286 6242 4338
rect 6242 4286 6244 4338
rect 6188 4284 6244 4286
rect 6860 4450 6916 4452
rect 6860 4398 6862 4450
rect 6862 4398 6914 4450
rect 6914 4398 6916 4450
rect 6860 4396 6916 4398
rect 8092 5068 8148 5124
rect 8876 5068 8932 5124
rect 8988 5180 9044 5236
rect 10668 6018 10724 6020
rect 10668 5966 10670 6018
rect 10670 5966 10722 6018
rect 10722 5966 10724 6018
rect 10668 5964 10724 5966
rect 9996 5906 10052 5908
rect 9996 5854 9998 5906
rect 9998 5854 10050 5906
rect 10050 5854 10052 5906
rect 9996 5852 10052 5854
rect 10108 5628 10164 5684
rect 10108 5292 10164 5348
rect 12796 5794 12852 5796
rect 12796 5742 12798 5794
rect 12798 5742 12850 5794
rect 12850 5742 12852 5794
rect 12796 5740 12852 5742
rect 13580 5740 13636 5796
rect 13020 5628 13076 5684
rect 12572 4284 12628 4340
rect 9660 4172 9716 4228
rect 7420 3612 7476 3668
rect 8764 3666 8820 3668
rect 8764 3614 8766 3666
rect 8766 3614 8818 3666
rect 8818 3614 8820 3666
rect 8764 3612 8820 3614
rect 11788 4060 11844 4116
rect 13916 5628 13972 5684
rect 13580 5180 13636 5236
rect 13916 5122 13972 5124
rect 13916 5070 13918 5122
rect 13918 5070 13970 5122
rect 13970 5070 13972 5122
rect 13916 5068 13972 5070
rect 14700 5234 14756 5236
rect 14700 5182 14702 5234
rect 14702 5182 14754 5234
rect 14754 5182 14756 5234
rect 14700 5180 14756 5182
rect 14588 4956 14644 5012
rect 16716 5794 16772 5796
rect 16716 5742 16718 5794
rect 16718 5742 16770 5794
rect 16770 5742 16772 5794
rect 16716 5740 16772 5742
rect 18060 5740 18116 5796
rect 17836 5628 17892 5684
rect 17948 5122 18004 5124
rect 17948 5070 17950 5122
rect 17950 5070 18002 5122
rect 18002 5070 18004 5122
rect 17948 5068 18004 5070
rect 16828 4956 16884 5012
rect 21644 5740 21700 5796
rect 20556 5514 20612 5516
rect 20556 5462 20592 5514
rect 20592 5462 20612 5514
rect 20556 5460 20612 5462
rect 20660 5514 20716 5516
rect 20660 5462 20664 5514
rect 20664 5462 20716 5514
rect 20660 5460 20716 5462
rect 20764 5514 20820 5516
rect 20868 5514 20924 5516
rect 20764 5462 20788 5514
rect 20788 5462 20820 5514
rect 20868 5462 20912 5514
rect 20912 5462 20924 5514
rect 20764 5460 20820 5462
rect 20868 5460 20924 5462
rect 20972 5460 21028 5516
rect 21076 5514 21132 5516
rect 21180 5514 21236 5516
rect 21076 5462 21088 5514
rect 21088 5462 21132 5514
rect 21180 5462 21212 5514
rect 21212 5462 21236 5514
rect 21076 5460 21132 5462
rect 21180 5460 21236 5462
rect 21284 5514 21340 5516
rect 21284 5462 21336 5514
rect 21336 5462 21340 5514
rect 21284 5460 21340 5462
rect 21388 5514 21444 5516
rect 21388 5462 21408 5514
rect 21408 5462 21444 5514
rect 21388 5460 21444 5462
rect 18732 4956 18788 5012
rect 18508 4732 18564 4788
rect 21644 5068 21700 5124
rect 22092 5628 22148 5684
rect 20860 4732 20916 4788
rect 22540 5628 22596 5684
rect 23212 5628 23268 5684
rect 22540 5122 22596 5124
rect 22540 5070 22542 5122
rect 22542 5070 22594 5122
rect 22594 5070 22596 5122
rect 22540 5068 22596 5070
rect 25564 5740 25620 5796
rect 24556 5628 24612 5684
rect 25340 4844 25396 4900
rect 25900 5122 25956 5124
rect 25900 5070 25902 5122
rect 25902 5070 25954 5122
rect 25954 5070 25956 5122
rect 25900 5068 25956 5070
rect 25900 4396 25956 4452
rect 23436 4284 23492 4340
rect 20556 3946 20612 3948
rect 20556 3894 20592 3946
rect 20592 3894 20612 3946
rect 20556 3892 20612 3894
rect 20660 3946 20716 3948
rect 20660 3894 20664 3946
rect 20664 3894 20716 3946
rect 20660 3892 20716 3894
rect 20764 3946 20820 3948
rect 20868 3946 20924 3948
rect 20764 3894 20788 3946
rect 20788 3894 20820 3946
rect 20868 3894 20912 3946
rect 20912 3894 20924 3946
rect 20764 3892 20820 3894
rect 20868 3892 20924 3894
rect 20972 3892 21028 3948
rect 21076 3946 21132 3948
rect 21180 3946 21236 3948
rect 21076 3894 21088 3946
rect 21088 3894 21132 3946
rect 21180 3894 21212 3946
rect 21212 3894 21236 3946
rect 21076 3892 21132 3894
rect 21180 3892 21236 3894
rect 21284 3946 21340 3948
rect 21284 3894 21336 3946
rect 21336 3894 21340 3946
rect 21284 3892 21340 3894
rect 21388 3946 21444 3948
rect 21388 3894 21408 3946
rect 21408 3894 21444 3946
rect 21388 3892 21444 3894
rect 24892 4226 24948 4228
rect 24892 4174 24894 4226
rect 24894 4174 24946 4226
rect 24946 4174 24948 4226
rect 24892 4172 24948 4174
rect 26124 4172 26180 4228
rect 26236 5628 26292 5684
rect 22764 3612 22820 3668
rect 30380 5964 30436 6020
rect 29484 5740 29540 5796
rect 28476 5628 28532 5684
rect 30268 5628 30324 5684
rect 26348 5068 26404 5124
rect 26684 5122 26740 5124
rect 26684 5070 26686 5122
rect 26686 5070 26738 5122
rect 26738 5070 26740 5122
rect 26684 5068 26740 5070
rect 28476 5068 28532 5124
rect 26460 4284 26516 4340
rect 28812 4956 28868 5012
rect 28700 4844 28756 4900
rect 29260 4396 29316 4452
rect 29932 4396 29988 4452
rect 30380 5740 30436 5796
rect 33516 5906 33572 5908
rect 33516 5854 33518 5906
rect 33518 5854 33570 5906
rect 33570 5854 33572 5906
rect 33516 5852 33572 5854
rect 32396 5628 32452 5684
rect 31500 4956 31556 5012
rect 33292 4844 33348 4900
rect 33964 4956 34020 5012
rect 31164 4732 31220 4788
rect 33964 4396 34020 4452
rect 32396 4284 32452 4340
rect 28588 4226 28644 4228
rect 28588 4174 28590 4226
rect 28590 4174 28642 4226
rect 28642 4174 28644 4226
rect 28588 4172 28644 4174
rect 31612 4172 31668 4228
rect 29484 3666 29540 3668
rect 29484 3614 29486 3666
rect 29486 3614 29538 3666
rect 29538 3614 29540 3666
rect 29484 3612 29540 3614
rect 12572 3554 12628 3556
rect 12572 3502 12574 3554
rect 12574 3502 12626 3554
rect 12626 3502 12628 3554
rect 12572 3500 12628 3502
rect 25676 3554 25732 3556
rect 25676 3502 25678 3554
rect 25678 3502 25730 3554
rect 25730 3502 25732 3554
rect 25676 3500 25732 3502
rect 31612 3388 31668 3444
rect 32844 4226 32900 4228
rect 32844 4174 32846 4226
rect 32846 4174 32898 4226
rect 32898 4174 32900 4226
rect 32844 4172 32900 4174
rect 34188 5628 34244 5684
rect 34636 5628 34692 5684
rect 36316 5068 36372 5124
rect 38108 5180 38164 5236
rect 38332 5740 38388 5796
rect 37212 4956 37268 5012
rect 37100 4338 37156 4340
rect 37100 4286 37102 4338
rect 37102 4286 37154 4338
rect 37154 4286 37156 4338
rect 37100 4284 37156 4286
rect 34076 4172 34132 4228
rect 32396 3554 32452 3556
rect 32396 3502 32398 3554
rect 32398 3502 32450 3554
rect 32450 3502 32452 3554
rect 32396 3500 32452 3502
rect 37772 5068 37828 5124
rect 39116 5234 39172 5236
rect 39116 5182 39118 5234
rect 39118 5182 39170 5234
rect 39170 5182 39172 5234
rect 39116 5180 39172 5182
rect 40212 6298 40268 6300
rect 40212 6246 40248 6298
rect 40248 6246 40268 6298
rect 40212 6244 40268 6246
rect 40316 6298 40372 6300
rect 40316 6246 40320 6298
rect 40320 6246 40372 6298
rect 40316 6244 40372 6246
rect 40420 6298 40476 6300
rect 40524 6298 40580 6300
rect 40420 6246 40444 6298
rect 40444 6246 40476 6298
rect 40524 6246 40568 6298
rect 40568 6246 40580 6298
rect 40420 6244 40476 6246
rect 40524 6244 40580 6246
rect 40628 6244 40684 6300
rect 40732 6298 40788 6300
rect 40836 6298 40892 6300
rect 40732 6246 40744 6298
rect 40744 6246 40788 6298
rect 40836 6246 40868 6298
rect 40868 6246 40892 6298
rect 40732 6244 40788 6246
rect 40836 6244 40892 6246
rect 40940 6298 40996 6300
rect 40940 6246 40992 6298
rect 40992 6246 40996 6298
rect 40940 6244 40996 6246
rect 41044 6298 41100 6300
rect 41044 6246 41064 6298
rect 41064 6246 41100 6298
rect 41044 6244 41100 6246
rect 41356 5906 41412 5908
rect 41356 5854 41358 5906
rect 41358 5854 41410 5906
rect 41410 5854 41412 5906
rect 41356 5852 41412 5854
rect 39900 5180 39956 5236
rect 41244 5234 41300 5236
rect 41244 5182 41246 5234
rect 41246 5182 41298 5234
rect 41298 5182 41300 5234
rect 41244 5180 41300 5182
rect 42028 5180 42084 5236
rect 40236 4956 40292 5012
rect 40212 4730 40268 4732
rect 40212 4678 40248 4730
rect 40248 4678 40268 4730
rect 40212 4676 40268 4678
rect 40316 4730 40372 4732
rect 40316 4678 40320 4730
rect 40320 4678 40372 4730
rect 40316 4676 40372 4678
rect 40420 4730 40476 4732
rect 40524 4730 40580 4732
rect 40420 4678 40444 4730
rect 40444 4678 40476 4730
rect 40524 4678 40568 4730
rect 40568 4678 40580 4730
rect 40420 4676 40476 4678
rect 40524 4676 40580 4678
rect 40628 4676 40684 4732
rect 40732 4730 40788 4732
rect 40836 4730 40892 4732
rect 40732 4678 40744 4730
rect 40744 4678 40788 4730
rect 40836 4678 40868 4730
rect 40868 4678 40892 4730
rect 40732 4676 40788 4678
rect 40836 4676 40892 4678
rect 40940 4730 40996 4732
rect 40940 4678 40992 4730
rect 40992 4678 40996 4730
rect 40940 4676 40996 4678
rect 41044 4730 41100 4732
rect 41044 4678 41064 4730
rect 41064 4678 41100 4730
rect 41044 4676 41100 4678
rect 39564 3612 39620 3668
rect 40012 3666 40068 3668
rect 40012 3614 40014 3666
rect 40014 3614 40066 3666
rect 40066 3614 40068 3666
rect 40012 3612 40068 3614
rect 37212 3554 37268 3556
rect 37212 3502 37214 3554
rect 37214 3502 37266 3554
rect 37266 3502 37268 3554
rect 37212 3500 37268 3502
rect 41356 3554 41412 3556
rect 41356 3502 41358 3554
rect 41358 3502 41410 3554
rect 41410 3502 41412 3554
rect 41356 3500 41412 3502
rect 42140 5068 42196 5124
rect 42588 5234 42644 5236
rect 42588 5182 42590 5234
rect 42590 5182 42642 5234
rect 42642 5182 42644 5234
rect 42588 5180 42644 5182
rect 42252 4956 42308 5012
rect 43148 5068 43204 5124
rect 45276 5740 45332 5796
rect 44156 5068 44212 5124
rect 45276 5068 45332 5124
rect 46396 5122 46452 5124
rect 46396 5070 46398 5122
rect 46398 5070 46450 5122
rect 46450 5070 46452 5122
rect 46396 5068 46452 5070
rect 45948 4844 46004 4900
rect 42476 4338 42532 4340
rect 42476 4286 42478 4338
rect 42478 4286 42530 4338
rect 42530 4286 42532 4338
rect 42476 4284 42532 4286
rect 45276 4226 45332 4228
rect 45276 4174 45278 4226
rect 45278 4174 45330 4226
rect 45330 4174 45332 4226
rect 45276 4172 45332 4174
rect 45164 4060 45220 4116
rect 44156 3666 44212 3668
rect 44156 3614 44158 3666
rect 44158 3614 44210 3666
rect 44210 3614 44212 3666
rect 44156 3612 44212 3614
rect 41804 3500 41860 3556
rect 45836 4060 45892 4116
rect 46620 4172 46676 4228
rect 48076 5794 48132 5796
rect 48076 5742 48078 5794
rect 48078 5742 48130 5794
rect 48130 5742 48132 5794
rect 48076 5740 48132 5742
rect 48748 4396 48804 4452
rect 49868 5794 49924 5796
rect 49868 5742 49870 5794
rect 49870 5742 49922 5794
rect 49922 5742 49924 5794
rect 49868 5740 49924 5742
rect 49196 5292 49252 5348
rect 49756 5292 49812 5348
rect 49084 4060 49140 4116
rect 47628 3612 47684 3668
rect 48076 3948 48132 4004
rect 45164 3554 45220 3556
rect 45164 3502 45166 3554
rect 45166 3502 45218 3554
rect 45218 3502 45220 3554
rect 45164 3500 45220 3502
rect 49868 5122 49924 5124
rect 49868 5070 49870 5122
rect 49870 5070 49922 5122
rect 49922 5070 49924 5122
rect 49868 5068 49924 5070
rect 50540 5740 50596 5796
rect 51996 4956 52052 5012
rect 50316 4396 50372 4452
rect 49196 3554 49252 3556
rect 49196 3502 49198 3554
rect 49198 3502 49250 3554
rect 49250 3502 49252 3554
rect 49196 3500 49252 3502
rect 52444 4060 52500 4116
rect 51996 3724 52052 3780
rect 53004 5906 53060 5908
rect 53004 5854 53006 5906
rect 53006 5854 53058 5906
rect 53058 5854 53060 5906
rect 53004 5852 53060 5854
rect 53004 5180 53060 5236
rect 53116 5628 53172 5684
rect 52892 3724 52948 3780
rect 52668 3612 52724 3668
rect 50316 3388 50372 3444
rect 53788 5292 53844 5348
rect 55580 5234 55636 5236
rect 55580 5182 55582 5234
rect 55582 5182 55634 5234
rect 55634 5182 55636 5234
rect 55580 5180 55636 5182
rect 53228 4172 53284 4228
rect 53900 4172 53956 4228
rect 53788 3666 53844 3668
rect 53788 3614 53790 3666
rect 53790 3614 53842 3666
rect 53842 3614 53844 3666
rect 53788 3612 53844 3614
rect 53116 3554 53172 3556
rect 53116 3502 53118 3554
rect 53118 3502 53170 3554
rect 53170 3502 53172 3554
rect 53116 3500 53172 3502
rect 55916 5794 55972 5796
rect 55916 5742 55918 5794
rect 55918 5742 55970 5794
rect 55970 5742 55972 5794
rect 55916 5740 55972 5742
rect 57036 5068 57092 5124
rect 56700 4620 56756 4676
rect 55692 3948 55748 4004
rect 55916 4172 55972 4228
rect 54572 3612 54628 3668
rect 57036 4508 57092 4564
rect 57708 4956 57764 5012
rect 60844 5628 60900 5684
rect 59868 5514 59924 5516
rect 59868 5462 59904 5514
rect 59904 5462 59924 5514
rect 59868 5460 59924 5462
rect 59972 5514 60028 5516
rect 59972 5462 59976 5514
rect 59976 5462 60028 5514
rect 59972 5460 60028 5462
rect 60076 5514 60132 5516
rect 60180 5514 60236 5516
rect 60076 5462 60100 5514
rect 60100 5462 60132 5514
rect 60180 5462 60224 5514
rect 60224 5462 60236 5514
rect 60076 5460 60132 5462
rect 60180 5460 60236 5462
rect 60284 5460 60340 5516
rect 60388 5514 60444 5516
rect 60492 5514 60548 5516
rect 60388 5462 60400 5514
rect 60400 5462 60444 5514
rect 60492 5462 60524 5514
rect 60524 5462 60548 5514
rect 60388 5460 60444 5462
rect 60492 5460 60548 5462
rect 60596 5514 60652 5516
rect 60596 5462 60648 5514
rect 60648 5462 60652 5514
rect 60596 5460 60652 5462
rect 60700 5514 60756 5516
rect 60700 5462 60720 5514
rect 60720 5462 60756 5514
rect 60700 5460 60756 5462
rect 59724 4956 59780 5012
rect 60396 5122 60452 5124
rect 60396 5070 60398 5122
rect 60398 5070 60450 5122
rect 60450 5070 60452 5122
rect 60396 5068 60452 5070
rect 58380 4844 58436 4900
rect 57820 4620 57876 4676
rect 61628 4956 61684 5012
rect 63756 4956 63812 5012
rect 64764 5628 64820 5684
rect 63644 4844 63700 4900
rect 62188 4284 62244 4340
rect 63756 4450 63812 4452
rect 63756 4398 63758 4450
rect 63758 4398 63810 4450
rect 63810 4398 63812 4450
rect 63756 4396 63812 4398
rect 61068 4172 61124 4228
rect 59868 3946 59924 3948
rect 59868 3894 59904 3946
rect 59904 3894 59924 3946
rect 59868 3892 59924 3894
rect 59972 3946 60028 3948
rect 59972 3894 59976 3946
rect 59976 3894 60028 3946
rect 59972 3892 60028 3894
rect 60076 3946 60132 3948
rect 60180 3946 60236 3948
rect 60076 3894 60100 3946
rect 60100 3894 60132 3946
rect 60180 3894 60224 3946
rect 60224 3894 60236 3946
rect 60076 3892 60132 3894
rect 60180 3892 60236 3894
rect 60284 3892 60340 3948
rect 60388 3946 60444 3948
rect 60492 3946 60548 3948
rect 60388 3894 60400 3946
rect 60400 3894 60444 3946
rect 60492 3894 60524 3946
rect 60524 3894 60548 3946
rect 60388 3892 60444 3894
rect 60492 3892 60548 3894
rect 60596 3946 60652 3948
rect 60596 3894 60648 3946
rect 60648 3894 60652 3946
rect 60596 3892 60652 3894
rect 60700 3946 60756 3948
rect 60700 3894 60720 3946
rect 60720 3894 60756 3946
rect 60700 3892 60756 3894
rect 60844 3836 60900 3892
rect 59836 3666 59892 3668
rect 59836 3614 59838 3666
rect 59838 3614 59890 3666
rect 59890 3614 59892 3666
rect 59836 3612 59892 3614
rect 62972 3666 63028 3668
rect 62972 3614 62974 3666
rect 62974 3614 63026 3666
rect 63026 3614 63028 3666
rect 62972 3612 63028 3614
rect 53900 3500 53956 3556
rect 57036 3554 57092 3556
rect 57036 3502 57038 3554
rect 57038 3502 57090 3554
rect 57090 3502 57092 3554
rect 57036 3500 57092 3502
rect 63756 3554 63812 3556
rect 63756 3502 63758 3554
rect 63758 3502 63810 3554
rect 63810 3502 63812 3554
rect 63756 3500 63812 3502
rect 66444 4956 66500 5012
rect 66668 5122 66724 5124
rect 66668 5070 66670 5122
rect 66670 5070 66722 5122
rect 66722 5070 66724 5122
rect 66668 5068 66724 5070
rect 65660 4508 65716 4564
rect 67676 4956 67732 5012
rect 66668 4284 66724 4340
rect 68460 4844 68516 4900
rect 65548 3836 65604 3892
rect 65548 3666 65604 3668
rect 65548 3614 65550 3666
rect 65550 3614 65602 3666
rect 65602 3614 65604 3666
rect 65548 3612 65604 3614
rect 67676 3666 67732 3668
rect 67676 3614 67678 3666
rect 67678 3614 67730 3666
rect 67730 3614 67732 3666
rect 67676 3612 67732 3614
rect 68684 4396 68740 4452
rect 69468 5794 69524 5796
rect 69468 5742 69470 5794
rect 69470 5742 69522 5794
rect 69522 5742 69524 5794
rect 69468 5740 69524 5742
rect 70140 5740 70196 5796
rect 69468 5516 69524 5572
rect 71596 5794 71652 5796
rect 71596 5742 71598 5794
rect 71598 5742 71650 5794
rect 71650 5742 71652 5794
rect 71596 5740 71652 5742
rect 69468 5122 69524 5124
rect 69468 5070 69470 5122
rect 69470 5070 69522 5122
rect 69522 5070 69524 5122
rect 69468 5068 69524 5070
rect 71820 4956 71876 5012
rect 73388 5794 73444 5796
rect 73388 5742 73390 5794
rect 73390 5742 73442 5794
rect 73442 5742 73444 5794
rect 73388 5740 73444 5742
rect 72156 5068 72212 5124
rect 70588 4508 70644 4564
rect 70476 4338 70532 4340
rect 70476 4286 70478 4338
rect 70478 4286 70530 4338
rect 70530 4286 70532 4338
rect 70476 4284 70532 4286
rect 69132 3612 69188 3668
rect 71372 3612 71428 3668
rect 73388 5180 73444 5236
rect 74396 5234 74452 5236
rect 74396 5182 74398 5234
rect 74398 5182 74450 5234
rect 74450 5182 74452 5234
rect 74396 5180 74452 5182
rect 73724 5122 73780 5124
rect 73724 5070 73726 5122
rect 73726 5070 73778 5122
rect 73778 5070 73780 5122
rect 73724 5068 73780 5070
rect 72268 4956 72324 5012
rect 75516 5794 75572 5796
rect 75516 5742 75518 5794
rect 75518 5742 75570 5794
rect 75570 5742 75572 5794
rect 75516 5740 75572 5742
rect 74508 4956 74564 5012
rect 77196 5740 77252 5796
rect 76636 5180 76692 5236
rect 76524 4956 76580 5012
rect 77308 4956 77364 5012
rect 72156 3612 72212 3668
rect 40212 3162 40268 3164
rect 40212 3110 40248 3162
rect 40248 3110 40268 3162
rect 40212 3108 40268 3110
rect 40316 3162 40372 3164
rect 40316 3110 40320 3162
rect 40320 3110 40372 3162
rect 40316 3108 40372 3110
rect 40420 3162 40476 3164
rect 40524 3162 40580 3164
rect 40420 3110 40444 3162
rect 40444 3110 40476 3162
rect 40524 3110 40568 3162
rect 40568 3110 40580 3162
rect 40420 3108 40476 3110
rect 40524 3108 40580 3110
rect 40628 3108 40684 3164
rect 40732 3162 40788 3164
rect 40836 3162 40892 3164
rect 40732 3110 40744 3162
rect 40744 3110 40788 3162
rect 40836 3110 40868 3162
rect 40868 3110 40892 3162
rect 40732 3108 40788 3110
rect 40836 3108 40892 3110
rect 40940 3162 40996 3164
rect 40940 3110 40992 3162
rect 40992 3110 40996 3162
rect 40940 3108 40996 3110
rect 41044 3162 41100 3164
rect 41044 3110 41064 3162
rect 41064 3110 41100 3162
rect 41044 3108 41100 3110
rect 76636 3612 76692 3668
rect 78428 4284 78484 4340
rect 79524 6298 79580 6300
rect 79524 6246 79560 6298
rect 79560 6246 79580 6298
rect 79524 6244 79580 6246
rect 79628 6298 79684 6300
rect 79628 6246 79632 6298
rect 79632 6246 79684 6298
rect 79628 6244 79684 6246
rect 79732 6298 79788 6300
rect 79836 6298 79892 6300
rect 79732 6246 79756 6298
rect 79756 6246 79788 6298
rect 79836 6246 79880 6298
rect 79880 6246 79892 6298
rect 79732 6244 79788 6246
rect 79836 6244 79892 6246
rect 79940 6244 79996 6300
rect 80044 6298 80100 6300
rect 80148 6298 80204 6300
rect 80044 6246 80056 6298
rect 80056 6246 80100 6298
rect 80148 6246 80180 6298
rect 80180 6246 80204 6298
rect 80044 6244 80100 6246
rect 80148 6244 80204 6246
rect 80252 6298 80308 6300
rect 80252 6246 80304 6298
rect 80304 6246 80308 6298
rect 80252 6244 80308 6246
rect 80356 6298 80412 6300
rect 80356 6246 80376 6298
rect 80376 6246 80412 6298
rect 80356 6244 80412 6246
rect 80332 5906 80388 5908
rect 80332 5854 80334 5906
rect 80334 5854 80386 5906
rect 80386 5854 80388 5906
rect 80332 5852 80388 5854
rect 79436 5794 79492 5796
rect 79436 5742 79438 5794
rect 79438 5742 79490 5794
rect 79490 5742 79492 5794
rect 79436 5740 79492 5742
rect 80332 5068 80388 5124
rect 81004 5794 81060 5796
rect 81004 5742 81006 5794
rect 81006 5742 81058 5794
rect 81058 5742 81060 5794
rect 81004 5740 81060 5742
rect 79524 4730 79580 4732
rect 79524 4678 79560 4730
rect 79560 4678 79580 4730
rect 79524 4676 79580 4678
rect 79628 4730 79684 4732
rect 79628 4678 79632 4730
rect 79632 4678 79684 4730
rect 79628 4676 79684 4678
rect 79732 4730 79788 4732
rect 79836 4730 79892 4732
rect 79732 4678 79756 4730
rect 79756 4678 79788 4730
rect 79836 4678 79880 4730
rect 79880 4678 79892 4730
rect 79732 4676 79788 4678
rect 79836 4676 79892 4678
rect 79940 4676 79996 4732
rect 80044 4730 80100 4732
rect 80148 4730 80204 4732
rect 80044 4678 80056 4730
rect 80056 4678 80100 4730
rect 80148 4678 80180 4730
rect 80180 4678 80204 4730
rect 80044 4676 80100 4678
rect 80148 4676 80204 4678
rect 80252 4730 80308 4732
rect 80252 4678 80304 4730
rect 80304 4678 80308 4730
rect 80252 4676 80308 4678
rect 80356 4730 80412 4732
rect 80356 4678 80376 4730
rect 80376 4678 80412 4730
rect 80356 4676 80412 4678
rect 82236 5068 82292 5124
rect 83132 5794 83188 5796
rect 83132 5742 83134 5794
rect 83134 5742 83186 5794
rect 83186 5742 83188 5794
rect 83132 5740 83188 5742
rect 84140 5628 84196 5684
rect 83916 5180 83972 5236
rect 83916 4338 83972 4340
rect 83916 4286 83918 4338
rect 83918 4286 83970 4338
rect 83970 4286 83972 4338
rect 83916 4284 83972 4286
rect 82572 3612 82628 3668
rect 83132 3666 83188 3668
rect 83132 3614 83134 3666
rect 83134 3614 83186 3666
rect 83186 3614 83188 3666
rect 83132 3612 83188 3614
rect 80332 3554 80388 3556
rect 80332 3502 80334 3554
rect 80334 3502 80386 3554
rect 80386 3502 80388 3554
rect 80332 3500 80388 3502
rect 84140 3500 84196 3556
rect 84252 5852 84308 5908
rect 84252 3612 84308 3668
rect 84924 5794 84980 5796
rect 84924 5742 84926 5794
rect 84926 5742 84978 5794
rect 84978 5742 84980 5794
rect 84924 5740 84980 5742
rect 85260 5740 85316 5796
rect 87052 5794 87108 5796
rect 87052 5742 87054 5794
rect 87054 5742 87106 5794
rect 87106 5742 87108 5794
rect 87052 5740 87108 5742
rect 86716 5180 86772 5236
rect 89292 5180 89348 5236
rect 88284 4226 88340 4228
rect 88284 4174 88286 4226
rect 88286 4174 88338 4226
rect 88338 4174 88340 4226
rect 88284 4172 88340 4174
rect 87052 3724 87108 3780
rect 88844 3724 88900 3780
rect 88172 3612 88228 3668
rect 90636 5740 90692 5796
rect 90972 5906 91028 5908
rect 90972 5854 90974 5906
rect 90974 5854 91026 5906
rect 91026 5854 91028 5906
rect 90972 5852 91028 5854
rect 91980 5794 92036 5796
rect 91980 5742 91982 5794
rect 91982 5742 92034 5794
rect 92034 5742 92036 5794
rect 91980 5740 92036 5742
rect 90972 5628 91028 5684
rect 94892 5906 94948 5908
rect 94892 5854 94894 5906
rect 94894 5854 94946 5906
rect 94946 5854 94948 5906
rect 94892 5852 94948 5854
rect 92092 4172 92148 4228
rect 90188 3724 90244 3780
rect 90972 3836 91028 3892
rect 93996 4226 94052 4228
rect 93996 4174 93998 4226
rect 93998 4174 94050 4226
rect 94050 4174 94052 4226
rect 93996 4172 94052 4174
rect 92092 3724 92148 3780
rect 88956 3500 89012 3556
rect 92764 3836 92820 3892
rect 96124 5852 96180 5908
rect 96684 5122 96740 5124
rect 96684 5070 96686 5122
rect 96686 5070 96738 5122
rect 96738 5070 96740 5122
rect 96684 5068 96740 5070
rect 94108 3836 94164 3892
rect 93996 3612 94052 3668
rect 94892 3666 94948 3668
rect 94892 3614 94894 3666
rect 94894 3614 94946 3666
rect 94946 3614 94948 3666
rect 94892 3612 94948 3614
rect 97244 4284 97300 4340
rect 95340 3612 95396 3668
rect 96684 3666 96740 3668
rect 96684 3614 96686 3666
rect 96686 3614 96738 3666
rect 96738 3614 96740 3666
rect 96684 3612 96740 3614
rect 98812 5906 98868 5908
rect 98812 5854 98814 5906
rect 98814 5854 98866 5906
rect 98866 5854 98868 5906
rect 98812 5852 98868 5854
rect 100156 5852 100212 5908
rect 99820 5794 99876 5796
rect 99820 5742 99822 5794
rect 99822 5742 99874 5794
rect 99874 5742 99876 5794
rect 99820 5740 99876 5742
rect 99180 5514 99236 5516
rect 99180 5462 99216 5514
rect 99216 5462 99236 5514
rect 99180 5460 99236 5462
rect 99284 5514 99340 5516
rect 99284 5462 99288 5514
rect 99288 5462 99340 5514
rect 99284 5460 99340 5462
rect 99388 5514 99444 5516
rect 99492 5514 99548 5516
rect 99388 5462 99412 5514
rect 99412 5462 99444 5514
rect 99492 5462 99536 5514
rect 99536 5462 99548 5514
rect 99388 5460 99444 5462
rect 99492 5460 99548 5462
rect 99596 5460 99652 5516
rect 99700 5514 99756 5516
rect 99804 5514 99860 5516
rect 99700 5462 99712 5514
rect 99712 5462 99756 5514
rect 99804 5462 99836 5514
rect 99836 5462 99860 5514
rect 99700 5460 99756 5462
rect 99804 5460 99860 5462
rect 99908 5514 99964 5516
rect 99908 5462 99960 5514
rect 99960 5462 99964 5514
rect 99908 5460 99964 5462
rect 100012 5514 100068 5516
rect 100012 5462 100032 5514
rect 100032 5462 100068 5514
rect 100012 5460 100068 5462
rect 98588 4284 98644 4340
rect 102732 5906 102788 5908
rect 102732 5854 102734 5906
rect 102734 5854 102786 5906
rect 102786 5854 102788 5906
rect 102732 5852 102788 5854
rect 103964 5906 104020 5908
rect 103964 5854 103966 5906
rect 103966 5854 104018 5906
rect 104018 5854 104020 5906
rect 103964 5852 104020 5854
rect 101388 5740 101444 5796
rect 104076 5740 104132 5796
rect 101948 5180 102004 5236
rect 102732 5180 102788 5236
rect 102620 5122 102676 5124
rect 102620 5070 102622 5122
rect 102622 5070 102674 5122
rect 102674 5070 102676 5122
rect 102620 5068 102676 5070
rect 99180 3946 99236 3948
rect 99180 3894 99216 3946
rect 99216 3894 99236 3946
rect 99180 3892 99236 3894
rect 99284 3946 99340 3948
rect 99284 3894 99288 3946
rect 99288 3894 99340 3946
rect 99284 3892 99340 3894
rect 99388 3946 99444 3948
rect 99492 3946 99548 3948
rect 99388 3894 99412 3946
rect 99412 3894 99444 3946
rect 99492 3894 99536 3946
rect 99536 3894 99548 3946
rect 99388 3892 99444 3894
rect 99492 3892 99548 3894
rect 99596 3892 99652 3948
rect 99700 3946 99756 3948
rect 99804 3946 99860 3948
rect 99700 3894 99712 3946
rect 99712 3894 99756 3946
rect 99804 3894 99836 3946
rect 99836 3894 99860 3946
rect 99700 3892 99756 3894
rect 99804 3892 99860 3894
rect 99908 3946 99964 3948
rect 99908 3894 99960 3946
rect 99960 3894 99964 3946
rect 99908 3892 99964 3894
rect 100012 3946 100068 3948
rect 100012 3894 100032 3946
rect 100032 3894 100068 3946
rect 100012 3892 100068 3894
rect 103292 5234 103348 5236
rect 103292 5182 103294 5234
rect 103294 5182 103346 5234
rect 103346 5182 103348 5234
rect 103292 5180 103348 5182
rect 107772 5852 107828 5908
rect 107660 5794 107716 5796
rect 107660 5742 107662 5794
rect 107662 5742 107714 5794
rect 107714 5742 107716 5794
rect 107660 5740 107716 5742
rect 105420 5234 105476 5236
rect 105420 5182 105422 5234
rect 105422 5182 105474 5234
rect 105474 5182 105476 5234
rect 105420 5180 105476 5182
rect 107772 4956 107828 5012
rect 104748 4396 104804 4452
rect 105980 4450 106036 4452
rect 105980 4398 105982 4450
rect 105982 4398 106034 4450
rect 106034 4398 106036 4450
rect 105980 4396 106036 4398
rect 105308 4338 105364 4340
rect 105308 4286 105310 4338
rect 105310 4286 105362 4338
rect 105362 4286 105364 4338
rect 105308 4284 105364 4286
rect 95900 3554 95956 3556
rect 95900 3502 95902 3554
rect 95902 3502 95954 3554
rect 95954 3502 95956 3554
rect 95900 3500 95956 3502
rect 99820 3554 99876 3556
rect 99820 3502 99822 3554
rect 99822 3502 99874 3554
rect 99874 3502 99876 3554
rect 99820 3500 99876 3502
rect 109788 5516 109844 5572
rect 111916 5740 111972 5796
rect 111244 5516 111300 5572
rect 111580 5292 111636 5348
rect 110572 4956 110628 5012
rect 109452 4620 109508 4676
rect 110572 4620 110628 4676
rect 109116 4508 109172 4564
rect 108108 4396 108164 4452
rect 108444 4396 108500 4452
rect 109452 4450 109508 4452
rect 109452 4398 109454 4450
rect 109454 4398 109506 4450
rect 109506 4398 109508 4450
rect 109452 4396 109508 4398
rect 108780 4338 108836 4340
rect 108780 4286 108782 4338
rect 108782 4286 108834 4338
rect 108834 4286 108836 4338
rect 108780 4284 108836 4286
rect 111916 4172 111972 4228
rect 112364 5292 112420 5348
rect 111580 3724 111636 3780
rect 113708 5292 113764 5348
rect 113372 5234 113428 5236
rect 113372 5182 113374 5234
rect 113374 5182 113426 5234
rect 113426 5182 113428 5234
rect 113372 5180 113428 5182
rect 112700 5122 112756 5124
rect 112700 5070 112702 5122
rect 112702 5070 112754 5122
rect 112754 5070 112756 5122
rect 112700 5068 112756 5070
rect 114380 4956 114436 5012
rect 114492 5180 114548 5236
rect 113148 4226 113204 4228
rect 113148 4174 113150 4226
rect 113150 4174 113202 4226
rect 113202 4174 113204 4226
rect 113148 4172 113204 4174
rect 115612 5740 115668 5796
rect 115388 5516 115444 5572
rect 115276 5180 115332 5236
rect 114828 4172 114884 4228
rect 115500 5292 115556 5348
rect 116284 5180 116340 5236
rect 117068 5122 117124 5124
rect 117068 5070 117070 5122
rect 117070 5070 117122 5122
rect 117122 5070 117124 5122
rect 117068 5068 117124 5070
rect 116060 4956 116116 5012
rect 116620 4226 116676 4228
rect 116620 4174 116622 4226
rect 116622 4174 116674 4226
rect 116674 4174 116676 4226
rect 116620 4172 116676 4174
rect 118836 6298 118892 6300
rect 118836 6246 118872 6298
rect 118872 6246 118892 6298
rect 118836 6244 118892 6246
rect 118940 6298 118996 6300
rect 118940 6246 118944 6298
rect 118944 6246 118996 6298
rect 118940 6244 118996 6246
rect 119044 6298 119100 6300
rect 119148 6298 119204 6300
rect 119044 6246 119068 6298
rect 119068 6246 119100 6298
rect 119148 6246 119192 6298
rect 119192 6246 119204 6298
rect 119044 6244 119100 6246
rect 119148 6244 119204 6246
rect 119252 6244 119308 6300
rect 119356 6298 119412 6300
rect 119460 6298 119516 6300
rect 119356 6246 119368 6298
rect 119368 6246 119412 6298
rect 119460 6246 119492 6298
rect 119492 6246 119516 6298
rect 119356 6244 119412 6246
rect 119460 6244 119516 6246
rect 119564 6298 119620 6300
rect 119564 6246 119616 6298
rect 119616 6246 119620 6298
rect 119564 6244 119620 6246
rect 119668 6298 119724 6300
rect 119668 6246 119688 6298
rect 119688 6246 119724 6298
rect 119668 6244 119724 6246
rect 118412 5852 118468 5908
rect 118636 5852 118692 5908
rect 117852 5234 117908 5236
rect 117852 5182 117854 5234
rect 117854 5182 117906 5234
rect 117906 5182 117908 5234
rect 117852 5180 117908 5182
rect 117516 4172 117572 4228
rect 117628 4844 117684 4900
rect 116060 3836 116116 3892
rect 119532 5740 119588 5796
rect 119980 4956 120036 5012
rect 118836 4730 118892 4732
rect 118836 4678 118872 4730
rect 118872 4678 118892 4730
rect 118836 4676 118892 4678
rect 118940 4730 118996 4732
rect 118940 4678 118944 4730
rect 118944 4678 118996 4730
rect 118940 4676 118996 4678
rect 119044 4730 119100 4732
rect 119148 4730 119204 4732
rect 119044 4678 119068 4730
rect 119068 4678 119100 4730
rect 119148 4678 119192 4730
rect 119192 4678 119204 4730
rect 119044 4676 119100 4678
rect 119148 4676 119204 4678
rect 119252 4676 119308 4732
rect 119356 4730 119412 4732
rect 119460 4730 119516 4732
rect 119356 4678 119368 4730
rect 119368 4678 119412 4730
rect 119460 4678 119492 4730
rect 119492 4678 119516 4730
rect 119356 4676 119412 4678
rect 119460 4676 119516 4678
rect 119564 4730 119620 4732
rect 119564 4678 119616 4730
rect 119616 4678 119620 4730
rect 119564 4676 119620 4678
rect 119668 4730 119724 4732
rect 119668 4678 119688 4730
rect 119688 4678 119724 4730
rect 119668 4676 119724 4678
rect 118412 4284 118468 4340
rect 111580 3554 111636 3556
rect 111580 3502 111582 3554
rect 111582 3502 111634 3554
rect 111634 3502 111636 3554
rect 111580 3500 111636 3502
rect 105308 3388 105364 3444
rect 119532 3836 119588 3892
rect 119420 3666 119476 3668
rect 119420 3614 119422 3666
rect 119422 3614 119474 3666
rect 119474 3614 119476 3666
rect 119420 3612 119476 3614
rect 120204 5906 120260 5908
rect 120204 5854 120206 5906
rect 120206 5854 120258 5906
rect 120258 5854 120260 5906
rect 120204 5852 120260 5854
rect 121324 5404 121380 5460
rect 121212 4338 121268 4340
rect 121212 4286 121214 4338
rect 121214 4286 121266 4338
rect 121266 4286 121268 4338
rect 121212 4284 121268 4286
rect 120652 3836 120708 3892
rect 120092 3612 120148 3668
rect 122332 3836 122388 3892
rect 123340 5906 123396 5908
rect 123340 5854 123342 5906
rect 123342 5854 123394 5906
rect 123394 5854 123396 5906
rect 123340 5852 123396 5854
rect 123340 5068 123396 5124
rect 123452 4508 123508 4564
rect 124124 4956 124180 5012
rect 124012 4226 124068 4228
rect 124012 4174 124014 4226
rect 124014 4174 124066 4226
rect 124066 4174 124068 4226
rect 124012 4172 124068 4174
rect 127932 5964 127988 6020
rect 126252 5628 126308 5684
rect 127148 5628 127204 5684
rect 125580 4956 125636 5012
rect 125020 4844 125076 4900
rect 124124 3724 124180 3780
rect 122892 3612 122948 3668
rect 123340 3666 123396 3668
rect 123340 3614 123342 3666
rect 123342 3614 123394 3666
rect 123394 3614 123396 3666
rect 123340 3612 123396 3614
rect 125356 4226 125412 4228
rect 125356 4174 125358 4226
rect 125358 4174 125410 4226
rect 125410 4174 125412 4226
rect 125356 4172 125412 4174
rect 126140 3836 126196 3892
rect 124572 3500 124628 3556
rect 127932 5740 127988 5796
rect 128044 5180 128100 5236
rect 128492 4956 128548 5012
rect 130172 4732 130228 4788
rect 128268 4396 128324 4452
rect 129052 4396 129108 4452
rect 127484 4226 127540 4228
rect 127484 4174 127486 4226
rect 127486 4174 127538 4226
rect 127538 4174 127540 4226
rect 127484 4172 127540 4174
rect 128044 4172 128100 4228
rect 127260 3836 127316 3892
rect 130172 4396 130228 4452
rect 130620 4172 130676 4228
rect 131292 5964 131348 6020
rect 132972 5852 133028 5908
rect 131292 4956 131348 5012
rect 131180 4450 131236 4452
rect 131180 4398 131182 4450
rect 131182 4398 131234 4450
rect 131234 4398 131236 4450
rect 131180 4396 131236 4398
rect 130956 4172 131012 4228
rect 131964 4396 132020 4452
rect 131180 3836 131236 3892
rect 132524 4226 132580 4228
rect 132524 4174 132526 4226
rect 132526 4174 132578 4226
rect 132578 4174 132580 4226
rect 132524 4172 132580 4174
rect 133756 5122 133812 5124
rect 133756 5070 133758 5122
rect 133758 5070 133810 5122
rect 133810 5070 133812 5122
rect 133756 5068 133812 5070
rect 134092 5068 134148 5124
rect 134652 5068 134708 5124
rect 135884 5628 135940 5684
rect 135100 4956 135156 5012
rect 135324 4620 135380 4676
rect 133644 4172 133700 4228
rect 131852 3836 131908 3892
rect 127372 3554 127428 3556
rect 127372 3502 127374 3554
rect 127374 3502 127426 3554
rect 127426 3502 127428 3554
rect 127372 3500 127428 3502
rect 139020 5906 139076 5908
rect 139020 5854 139022 5906
rect 139022 5854 139074 5906
rect 139074 5854 139076 5906
rect 139020 5852 139076 5854
rect 138012 5292 138068 5348
rect 136332 4956 136388 5012
rect 135884 4060 135940 4116
rect 131964 3724 132020 3780
rect 134092 3724 134148 3780
rect 137228 4844 137284 4900
rect 136444 4620 136500 4676
rect 137004 4226 137060 4228
rect 137004 4174 137006 4226
rect 137006 4174 137058 4226
rect 137058 4174 137060 4226
rect 137004 4172 137060 4174
rect 136444 3948 136500 4004
rect 138492 5514 138548 5516
rect 138492 5462 138528 5514
rect 138528 5462 138548 5514
rect 138492 5460 138548 5462
rect 138596 5514 138652 5516
rect 138596 5462 138600 5514
rect 138600 5462 138652 5514
rect 138596 5460 138652 5462
rect 138700 5514 138756 5516
rect 138804 5514 138860 5516
rect 138700 5462 138724 5514
rect 138724 5462 138756 5514
rect 138804 5462 138848 5514
rect 138848 5462 138860 5514
rect 138700 5460 138756 5462
rect 138804 5460 138860 5462
rect 138908 5460 138964 5516
rect 139012 5514 139068 5516
rect 139116 5514 139172 5516
rect 139012 5462 139024 5514
rect 139024 5462 139068 5514
rect 139116 5462 139148 5514
rect 139148 5462 139172 5514
rect 139012 5460 139068 5462
rect 139116 5460 139172 5462
rect 139220 5514 139276 5516
rect 139220 5462 139272 5514
rect 139272 5462 139276 5514
rect 139220 5460 139276 5462
rect 139324 5514 139380 5516
rect 139324 5462 139344 5514
rect 139344 5462 139380 5514
rect 139324 5460 139380 5462
rect 139356 4844 139412 4900
rect 138124 4620 138180 4676
rect 138348 4284 138404 4340
rect 135100 3554 135156 3556
rect 135100 3502 135102 3554
rect 135102 3502 135154 3554
rect 135154 3502 135156 3554
rect 135100 3500 135156 3502
rect 139132 4226 139188 4228
rect 139132 4174 139134 4226
rect 139134 4174 139186 4226
rect 139186 4174 139188 4226
rect 139132 4172 139188 4174
rect 143836 5852 143892 5908
rect 141708 5740 141764 5796
rect 139804 5292 139860 5348
rect 140924 4956 140980 5012
rect 141932 5068 141988 5124
rect 139468 4172 139524 4228
rect 140476 4226 140532 4228
rect 140476 4174 140478 4226
rect 140478 4174 140530 4226
rect 140530 4174 140532 4226
rect 140476 4172 140532 4174
rect 139804 4060 139860 4116
rect 138492 3946 138548 3948
rect 138492 3894 138528 3946
rect 138528 3894 138548 3946
rect 138492 3892 138548 3894
rect 138596 3946 138652 3948
rect 138596 3894 138600 3946
rect 138600 3894 138652 3946
rect 138596 3892 138652 3894
rect 138700 3946 138756 3948
rect 138804 3946 138860 3948
rect 138700 3894 138724 3946
rect 138724 3894 138756 3946
rect 138804 3894 138848 3946
rect 138848 3894 138860 3946
rect 138700 3892 138756 3894
rect 138804 3892 138860 3894
rect 138908 3892 138964 3948
rect 139012 3946 139068 3948
rect 139116 3946 139172 3948
rect 139012 3894 139024 3946
rect 139024 3894 139068 3946
rect 139116 3894 139148 3946
rect 139148 3894 139172 3946
rect 139012 3892 139068 3894
rect 139116 3892 139172 3894
rect 139220 3946 139276 3948
rect 139220 3894 139272 3946
rect 139272 3894 139276 3946
rect 139220 3892 139276 3894
rect 139324 3946 139380 3948
rect 139324 3894 139344 3946
rect 139344 3894 139380 3946
rect 139324 3892 139380 3894
rect 139804 3666 139860 3668
rect 139804 3614 139806 3666
rect 139806 3614 139858 3666
rect 139858 3614 139860 3666
rect 139804 3612 139860 3614
rect 142940 5794 142996 5796
rect 142940 5742 142942 5794
rect 142942 5742 142994 5794
rect 142994 5742 142996 5794
rect 142940 5740 142996 5742
rect 143052 5292 143108 5348
rect 143724 4396 143780 4452
rect 142044 3612 142100 3668
rect 142604 3612 142660 3668
rect 142940 4060 142996 4116
rect 138348 3500 138404 3556
rect 139020 3554 139076 3556
rect 139020 3502 139022 3554
rect 139022 3502 139074 3554
rect 139074 3502 139076 3554
rect 139020 3500 139076 3502
rect 143276 4060 143332 4116
rect 143836 4060 143892 4116
rect 144508 5964 144564 6020
rect 145740 5906 145796 5908
rect 145740 5854 145742 5906
rect 145742 5854 145794 5906
rect 145794 5854 145796 5906
rect 145740 5852 145796 5854
rect 145180 5122 145236 5124
rect 145180 5070 145182 5122
rect 145182 5070 145234 5122
rect 145234 5070 145236 5122
rect 145180 5068 145236 5070
rect 147084 4508 147140 4564
rect 147308 4956 147364 5012
rect 149772 4732 149828 4788
rect 147308 4396 147364 4452
rect 158148 6298 158204 6300
rect 158148 6246 158184 6298
rect 158184 6246 158204 6298
rect 158148 6244 158204 6246
rect 158252 6298 158308 6300
rect 158252 6246 158256 6298
rect 158256 6246 158308 6298
rect 158252 6244 158308 6246
rect 158356 6298 158412 6300
rect 158460 6298 158516 6300
rect 158356 6246 158380 6298
rect 158380 6246 158412 6298
rect 158460 6246 158504 6298
rect 158504 6246 158516 6298
rect 158356 6244 158412 6246
rect 158460 6244 158516 6246
rect 158564 6244 158620 6300
rect 158668 6298 158724 6300
rect 158772 6298 158828 6300
rect 158668 6246 158680 6298
rect 158680 6246 158724 6298
rect 158772 6246 158804 6298
rect 158804 6246 158828 6298
rect 158668 6244 158724 6246
rect 158772 6244 158828 6246
rect 158876 6298 158932 6300
rect 158876 6246 158928 6298
rect 158928 6246 158932 6298
rect 158876 6244 158932 6246
rect 158980 6298 159036 6300
rect 158980 6246 159000 6298
rect 159000 6246 159036 6298
rect 158980 6244 159036 6246
rect 157836 4844 157892 4900
rect 155148 4620 155204 4676
rect 158148 4730 158204 4732
rect 158148 4678 158184 4730
rect 158184 4678 158204 4730
rect 158148 4676 158204 4678
rect 158252 4730 158308 4732
rect 158252 4678 158256 4730
rect 158256 4678 158308 4730
rect 158252 4676 158308 4678
rect 158356 4730 158412 4732
rect 158460 4730 158516 4732
rect 158356 4678 158380 4730
rect 158380 4678 158412 4730
rect 158460 4678 158504 4730
rect 158504 4678 158516 4730
rect 158356 4676 158412 4678
rect 158460 4676 158516 4678
rect 158564 4676 158620 4732
rect 158668 4730 158724 4732
rect 158772 4730 158828 4732
rect 158668 4678 158680 4730
rect 158680 4678 158724 4730
rect 158772 4678 158804 4730
rect 158804 4678 158828 4730
rect 158668 4676 158724 4678
rect 158772 4676 158828 4678
rect 158876 4730 158932 4732
rect 158876 4678 158928 4730
rect 158928 4678 158932 4730
rect 158876 4676 158932 4678
rect 158980 4730 159036 4732
rect 158980 4678 159000 4730
rect 159000 4678 159036 4730
rect 158980 4676 159036 4678
rect 152460 3724 152516 3780
rect 144396 3612 144452 3668
rect 145852 3666 145908 3668
rect 145852 3614 145854 3666
rect 145854 3614 145906 3666
rect 145906 3614 145908 3666
rect 145852 3612 145908 3614
rect 79524 3162 79580 3164
rect 79524 3110 79560 3162
rect 79560 3110 79580 3162
rect 79524 3108 79580 3110
rect 79628 3162 79684 3164
rect 79628 3110 79632 3162
rect 79632 3110 79684 3162
rect 79628 3108 79684 3110
rect 79732 3162 79788 3164
rect 79836 3162 79892 3164
rect 79732 3110 79756 3162
rect 79756 3110 79788 3162
rect 79836 3110 79880 3162
rect 79880 3110 79892 3162
rect 79732 3108 79788 3110
rect 79836 3108 79892 3110
rect 79940 3108 79996 3164
rect 80044 3162 80100 3164
rect 80148 3162 80204 3164
rect 80044 3110 80056 3162
rect 80056 3110 80100 3162
rect 80148 3110 80180 3162
rect 80180 3110 80204 3162
rect 80044 3108 80100 3110
rect 80148 3108 80204 3110
rect 80252 3162 80308 3164
rect 80252 3110 80304 3162
rect 80304 3110 80308 3162
rect 80252 3108 80308 3110
rect 80356 3162 80412 3164
rect 80356 3110 80376 3162
rect 80376 3110 80412 3162
rect 80356 3108 80412 3110
rect 118836 3162 118892 3164
rect 118836 3110 118872 3162
rect 118872 3110 118892 3162
rect 118836 3108 118892 3110
rect 118940 3162 118996 3164
rect 118940 3110 118944 3162
rect 118944 3110 118996 3162
rect 118940 3108 118996 3110
rect 119044 3162 119100 3164
rect 119148 3162 119204 3164
rect 119044 3110 119068 3162
rect 119068 3110 119100 3162
rect 119148 3110 119192 3162
rect 119192 3110 119204 3162
rect 119044 3108 119100 3110
rect 119148 3108 119204 3110
rect 119252 3108 119308 3164
rect 119356 3162 119412 3164
rect 119460 3162 119516 3164
rect 119356 3110 119368 3162
rect 119368 3110 119412 3162
rect 119460 3110 119492 3162
rect 119492 3110 119516 3162
rect 119356 3108 119412 3110
rect 119460 3108 119516 3110
rect 119564 3162 119620 3164
rect 119564 3110 119616 3162
rect 119616 3110 119620 3162
rect 119564 3108 119620 3110
rect 119668 3162 119724 3164
rect 119668 3110 119688 3162
rect 119688 3110 119724 3162
rect 119668 3108 119724 3110
rect 158148 3162 158204 3164
rect 158148 3110 158184 3162
rect 158184 3110 158204 3162
rect 158148 3108 158204 3110
rect 158252 3162 158308 3164
rect 158252 3110 158256 3162
rect 158256 3110 158308 3162
rect 158252 3108 158308 3110
rect 158356 3162 158412 3164
rect 158460 3162 158516 3164
rect 158356 3110 158380 3162
rect 158380 3110 158412 3162
rect 158460 3110 158504 3162
rect 158504 3110 158516 3162
rect 158356 3108 158412 3110
rect 158460 3108 158516 3110
rect 158564 3108 158620 3164
rect 158668 3162 158724 3164
rect 158772 3162 158828 3164
rect 158668 3110 158680 3162
rect 158680 3110 158724 3162
rect 158772 3110 158804 3162
rect 158804 3110 158828 3162
rect 158668 3108 158724 3110
rect 158772 3108 158828 3110
rect 158876 3162 158932 3164
rect 158876 3110 158928 3162
rect 158928 3110 158932 3162
rect 158876 3108 158932 3110
rect 158980 3162 159036 3164
rect 158980 3110 159000 3162
rect 159000 3110 159036 3162
rect 158980 3108 159036 3110
rect 73948 1708 74004 1764
<< metal3 >>
rect 0 8260 800 8288
rect 0 8204 2044 8260
rect 2100 8204 2110 8260
rect 0 8176 800 8204
rect 40202 6244 40212 6300
rect 40268 6244 40316 6300
rect 40372 6244 40420 6300
rect 40476 6244 40524 6300
rect 40580 6244 40628 6300
rect 40684 6244 40732 6300
rect 40788 6244 40836 6300
rect 40892 6244 40940 6300
rect 40996 6244 41044 6300
rect 41100 6244 41110 6300
rect 79514 6244 79524 6300
rect 79580 6244 79628 6300
rect 79684 6244 79732 6300
rect 79788 6244 79836 6300
rect 79892 6244 79940 6300
rect 79996 6244 80044 6300
rect 80100 6244 80148 6300
rect 80204 6244 80252 6300
rect 80308 6244 80356 6300
rect 80412 6244 80422 6300
rect 118826 6244 118836 6300
rect 118892 6244 118940 6300
rect 118996 6244 119044 6300
rect 119100 6244 119148 6300
rect 119204 6244 119252 6300
rect 119308 6244 119356 6300
rect 119412 6244 119460 6300
rect 119516 6244 119564 6300
rect 119620 6244 119668 6300
rect 119724 6244 119734 6300
rect 158138 6244 158148 6300
rect 158204 6244 158252 6300
rect 158308 6244 158356 6300
rect 158412 6244 158460 6300
rect 158516 6244 158564 6300
rect 158620 6244 158668 6300
rect 158724 6244 158772 6300
rect 158828 6244 158876 6300
rect 158932 6244 158980 6300
rect 159036 6244 159046 6300
rect 5954 5964 5964 6020
rect 6020 5964 10668 6020
rect 10724 5964 10734 6020
rect 30370 5964 30380 6020
rect 30436 5964 33572 6020
rect 127922 5964 127932 6020
rect 127988 5964 131292 6020
rect 131348 5964 144508 6020
rect 144564 5964 144574 6020
rect 33516 5908 33572 5964
rect 8372 5852 9996 5908
rect 10052 5852 31948 5908
rect 33506 5852 33516 5908
rect 33572 5852 41356 5908
rect 41412 5852 53004 5908
rect 53060 5852 53070 5908
rect 80322 5852 80332 5908
rect 80388 5852 84252 5908
rect 84308 5852 84318 5908
rect 90962 5852 90972 5908
rect 91028 5852 94892 5908
rect 94948 5852 96124 5908
rect 96180 5852 98812 5908
rect 98868 5852 100156 5908
rect 100212 5852 102732 5908
rect 102788 5852 103964 5908
rect 104020 5852 107772 5908
rect 107828 5852 107838 5908
rect 118402 5852 118412 5908
rect 118468 5852 118636 5908
rect 118692 5852 120204 5908
rect 120260 5852 120270 5908
rect 123330 5852 123340 5908
rect 123396 5852 132972 5908
rect 133028 5852 139020 5908
rect 139076 5852 139086 5908
rect 143826 5852 143836 5908
rect 143892 5852 145740 5908
rect 145796 5852 145806 5908
rect 8372 5796 8428 5852
rect 31892 5796 31948 5852
rect 2146 5740 2156 5796
rect 2212 5740 8428 5796
rect 12786 5740 12796 5796
rect 12852 5740 13580 5796
rect 13636 5740 13646 5796
rect 16706 5740 16716 5796
rect 16772 5740 18060 5796
rect 18116 5740 18126 5796
rect 21634 5740 21644 5796
rect 21700 5740 25564 5796
rect 25620 5740 29484 5796
rect 29540 5740 30380 5796
rect 30436 5740 30446 5796
rect 31892 5740 38332 5796
rect 38388 5740 45276 5796
rect 45332 5740 45342 5796
rect 48066 5740 48076 5796
rect 48132 5740 49868 5796
rect 49924 5740 50540 5796
rect 50596 5740 50606 5796
rect 55906 5740 55916 5796
rect 55972 5740 69468 5796
rect 69524 5740 70140 5796
rect 70196 5740 70206 5796
rect 71586 5740 71596 5796
rect 71652 5740 73388 5796
rect 73444 5740 73454 5796
rect 75506 5740 75516 5796
rect 75572 5740 77196 5796
rect 77252 5740 77262 5796
rect 79426 5740 79436 5796
rect 79492 5740 81004 5796
rect 81060 5740 81070 5796
rect 83122 5740 83132 5796
rect 83188 5740 84924 5796
rect 84980 5740 84990 5796
rect 85250 5740 85260 5796
rect 85316 5740 87052 5796
rect 87108 5740 87118 5796
rect 90626 5740 90636 5796
rect 90692 5740 91980 5796
rect 92036 5740 92046 5796
rect 99810 5740 99820 5796
rect 99876 5740 101388 5796
rect 101444 5740 101454 5796
rect 104066 5740 104076 5796
rect 104132 5740 107660 5796
rect 107716 5740 107726 5796
rect 111906 5740 111916 5796
rect 111972 5740 115612 5796
rect 115668 5740 119532 5796
rect 119588 5740 127932 5796
rect 127988 5740 127998 5796
rect 141698 5740 141708 5796
rect 141764 5740 142940 5796
rect 142996 5740 143006 5796
rect 10098 5628 10108 5684
rect 10164 5628 13020 5684
rect 13076 5628 13916 5684
rect 13972 5628 17836 5684
rect 17892 5628 22092 5684
rect 22148 5628 22540 5684
rect 22596 5628 22606 5684
rect 23202 5628 23212 5684
rect 23268 5628 24556 5684
rect 24612 5628 26236 5684
rect 26292 5628 26302 5684
rect 28466 5628 28476 5684
rect 28532 5628 30268 5684
rect 30324 5628 30334 5684
rect 32386 5628 32396 5684
rect 32452 5628 34188 5684
rect 34244 5628 34636 5684
rect 34692 5628 34702 5684
rect 53106 5628 53116 5684
rect 53172 5628 60844 5684
rect 60900 5628 64764 5684
rect 64820 5628 64830 5684
rect 84130 5628 84140 5684
rect 84196 5628 90972 5684
rect 91028 5628 91038 5684
rect 126242 5628 126252 5684
rect 126308 5628 127148 5684
rect 127204 5628 135884 5684
rect 135940 5628 135950 5684
rect 64764 5572 64820 5628
rect 64764 5516 69468 5572
rect 69524 5516 69534 5572
rect 109778 5516 109788 5572
rect 109844 5516 111244 5572
rect 111300 5516 115388 5572
rect 115444 5516 115454 5572
rect 20546 5460 20556 5516
rect 20612 5460 20660 5516
rect 20716 5460 20764 5516
rect 20820 5460 20868 5516
rect 20924 5460 20972 5516
rect 21028 5460 21076 5516
rect 21132 5460 21180 5516
rect 21236 5460 21284 5516
rect 21340 5460 21388 5516
rect 21444 5460 21454 5516
rect 59858 5460 59868 5516
rect 59924 5460 59972 5516
rect 60028 5460 60076 5516
rect 60132 5460 60180 5516
rect 60236 5460 60284 5516
rect 60340 5460 60388 5516
rect 60444 5460 60492 5516
rect 60548 5460 60596 5516
rect 60652 5460 60700 5516
rect 60756 5460 60766 5516
rect 99170 5460 99180 5516
rect 99236 5460 99284 5516
rect 99340 5460 99388 5516
rect 99444 5460 99492 5516
rect 99548 5460 99596 5516
rect 99652 5460 99700 5516
rect 99756 5460 99804 5516
rect 99860 5460 99908 5516
rect 99964 5460 100012 5516
rect 100068 5460 100078 5516
rect 138482 5460 138492 5516
rect 138548 5460 138596 5516
rect 138652 5460 138700 5516
rect 138756 5460 138804 5516
rect 138860 5460 138908 5516
rect 138964 5460 139012 5516
rect 139068 5460 139116 5516
rect 139172 5460 139220 5516
rect 139276 5460 139324 5516
rect 139380 5460 139390 5516
rect 114212 5404 121324 5460
rect 121380 5404 121390 5460
rect 8372 5292 10108 5348
rect 10164 5292 10174 5348
rect 49186 5292 49196 5348
rect 49252 5292 49756 5348
rect 49812 5292 53788 5348
rect 53844 5292 53854 5348
rect 111570 5292 111580 5348
rect 111636 5292 112364 5348
rect 112420 5292 113708 5348
rect 113764 5292 113774 5348
rect 8372 5236 8428 5292
rect 114212 5236 114268 5404
rect 115490 5292 115500 5348
rect 115556 5292 117908 5348
rect 138002 5292 138012 5348
rect 138068 5292 139804 5348
rect 139860 5292 143052 5348
rect 143108 5292 143118 5348
rect 117852 5236 117908 5292
rect 6524 5180 8428 5236
rect 8652 5180 8988 5236
rect 9044 5180 9054 5236
rect 13570 5180 13580 5236
rect 13636 5180 14700 5236
rect 14756 5180 14766 5236
rect 38098 5180 38108 5236
rect 38164 5180 39116 5236
rect 39172 5180 39900 5236
rect 39956 5180 39966 5236
rect 41234 5180 41244 5236
rect 41300 5180 42028 5236
rect 42084 5180 42588 5236
rect 42644 5180 42654 5236
rect 52994 5180 53004 5236
rect 53060 5180 55580 5236
rect 55636 5180 55646 5236
rect 73378 5180 73388 5236
rect 73444 5180 74396 5236
rect 74452 5180 74462 5236
rect 76626 5180 76636 5236
rect 76692 5180 82292 5236
rect 83906 5180 83916 5236
rect 83972 5180 86716 5236
rect 86772 5180 89292 5236
rect 89348 5180 89358 5236
rect 101938 5180 101948 5236
rect 102004 5180 102732 5236
rect 102788 5180 103292 5236
rect 103348 5180 103358 5236
rect 105410 5180 105420 5236
rect 105476 5180 113372 5236
rect 113428 5180 114268 5236
rect 114482 5180 114492 5236
rect 114548 5180 115276 5236
rect 115332 5180 116284 5236
rect 116340 5180 116350 5236
rect 117842 5180 117852 5236
rect 117908 5180 128044 5236
rect 128100 5180 128110 5236
rect 6524 5124 6580 5180
rect 8652 5124 8708 5180
rect 82236 5124 82292 5180
rect 2034 5068 2044 5124
rect 2100 5068 4732 5124
rect 4788 5068 6524 5124
rect 6580 5068 6590 5124
rect 7298 5068 7308 5124
rect 7364 5068 8092 5124
rect 8148 5068 8708 5124
rect 8866 5068 8876 5124
rect 8932 5068 13916 5124
rect 13972 5068 17948 5124
rect 18004 5068 21644 5124
rect 21700 5068 21710 5124
rect 22530 5068 22540 5124
rect 22596 5068 25900 5124
rect 25956 5068 25966 5124
rect 26338 5068 26348 5124
rect 26404 5068 26684 5124
rect 26740 5068 28476 5124
rect 28532 5068 28542 5124
rect 36306 5068 36316 5124
rect 36372 5068 37772 5124
rect 37828 5068 37838 5124
rect 42130 5068 42140 5124
rect 42196 5068 43148 5124
rect 43204 5068 44156 5124
rect 44212 5068 44222 5124
rect 45266 5068 45276 5124
rect 45332 5068 46396 5124
rect 46452 5068 49868 5124
rect 49924 5068 57036 5124
rect 57092 5068 57102 5124
rect 60386 5068 60396 5124
rect 60452 5068 66668 5124
rect 66724 5068 66734 5124
rect 69458 5068 69468 5124
rect 69524 5068 72156 5124
rect 72212 5068 72222 5124
rect 73714 5068 73724 5124
rect 73780 5068 80332 5124
rect 80388 5068 80398 5124
rect 82226 5068 82236 5124
rect 82292 5068 96684 5124
rect 96740 5068 102620 5124
rect 102676 5068 112700 5124
rect 112756 5068 117068 5124
rect 117124 5068 123340 5124
rect 123396 5068 123406 5124
rect 133746 5068 133756 5124
rect 133812 5068 134092 5124
rect 134148 5068 134652 5124
rect 134708 5068 134718 5124
rect 141922 5068 141932 5124
rect 141988 5068 145180 5124
rect 145236 5068 145246 5124
rect 0 5012 800 5040
rect 159200 5012 160000 5040
rect 0 4956 980 5012
rect 14578 4956 14588 5012
rect 14644 4956 16828 5012
rect 16884 4956 18732 5012
rect 18788 4956 18798 5012
rect 28802 4956 28812 5012
rect 28868 4956 31500 5012
rect 31556 4956 31566 5012
rect 33954 4956 33964 5012
rect 34020 4956 37212 5012
rect 37268 4956 37278 5012
rect 40226 4956 40236 5012
rect 40292 4956 42252 5012
rect 42308 4956 42318 5012
rect 51986 4956 51996 5012
rect 52052 4956 55468 5012
rect 57698 4956 57708 5012
rect 57764 4956 59724 5012
rect 59780 4956 61628 5012
rect 61684 4956 61694 5012
rect 63746 4956 63756 5012
rect 63812 4956 66444 5012
rect 66500 4956 66510 5012
rect 67666 4956 67676 5012
rect 67732 4956 71820 5012
rect 71876 4956 71886 5012
rect 72258 4956 72268 5012
rect 72324 4956 74508 5012
rect 74564 4956 74574 5012
rect 76514 4956 76524 5012
rect 76580 4956 77308 5012
rect 77364 4956 77374 5012
rect 107762 4956 107772 5012
rect 107828 4956 110572 5012
rect 110628 4956 114380 5012
rect 114436 4956 116060 5012
rect 116116 4956 116126 5012
rect 119970 4956 119980 5012
rect 120036 4956 124124 5012
rect 124180 4956 124190 5012
rect 125570 4956 125580 5012
rect 125636 4956 128492 5012
rect 128548 4956 128558 5012
rect 131282 4956 131292 5012
rect 131348 4956 135100 5012
rect 135156 4956 135166 5012
rect 136322 4956 136332 5012
rect 136388 4956 140924 5012
rect 140980 4956 140990 5012
rect 147298 4956 147308 5012
rect 147364 4956 160000 5012
rect 0 4928 800 4956
rect 924 4676 980 4956
rect 55412 4900 55468 4956
rect 159200 4928 160000 4956
rect 25330 4844 25340 4900
rect 25396 4844 28700 4900
rect 28756 4844 28766 4900
rect 33282 4844 33292 4900
rect 33348 4844 45948 4900
rect 46004 4844 46014 4900
rect 55412 4844 58380 4900
rect 58436 4844 58446 4900
rect 63634 4844 63644 4900
rect 63700 4844 68460 4900
rect 68516 4844 68526 4900
rect 117618 4844 117628 4900
rect 117684 4844 125020 4900
rect 125076 4844 137228 4900
rect 137284 4844 137294 4900
rect 139346 4844 139356 4900
rect 139412 4844 157836 4900
rect 157892 4844 157902 4900
rect 18498 4732 18508 4788
rect 18564 4732 20860 4788
rect 20916 4732 31164 4788
rect 31220 4732 31230 4788
rect 130162 4732 130172 4788
rect 130228 4732 149772 4788
rect 149828 4732 149838 4788
rect 40202 4676 40212 4732
rect 40268 4676 40316 4732
rect 40372 4676 40420 4732
rect 40476 4676 40524 4732
rect 40580 4676 40628 4732
rect 40684 4676 40732 4732
rect 40788 4676 40836 4732
rect 40892 4676 40940 4732
rect 40996 4676 41044 4732
rect 41100 4676 41110 4732
rect 79514 4676 79524 4732
rect 79580 4676 79628 4732
rect 79684 4676 79732 4732
rect 79788 4676 79836 4732
rect 79892 4676 79940 4732
rect 79996 4676 80044 4732
rect 80100 4676 80148 4732
rect 80204 4676 80252 4732
rect 80308 4676 80356 4732
rect 80412 4676 80422 4732
rect 118826 4676 118836 4732
rect 118892 4676 118940 4732
rect 118996 4676 119044 4732
rect 119100 4676 119148 4732
rect 119204 4676 119252 4732
rect 119308 4676 119356 4732
rect 119412 4676 119460 4732
rect 119516 4676 119564 4732
rect 119620 4676 119668 4732
rect 119724 4676 119734 4732
rect 158138 4676 158148 4732
rect 158204 4676 158252 4732
rect 158308 4676 158356 4732
rect 158412 4676 158460 4732
rect 158516 4676 158564 4732
rect 158620 4676 158668 4732
rect 158724 4676 158772 4732
rect 158828 4676 158876 4732
rect 158932 4676 158980 4732
rect 159036 4676 159046 4732
rect 700 4620 980 4676
rect 56690 4620 56700 4676
rect 56756 4620 57820 4676
rect 57876 4620 67228 4676
rect 109442 4620 109452 4676
rect 109508 4620 110572 4676
rect 110628 4620 110638 4676
rect 135314 4620 135324 4676
rect 135380 4620 136444 4676
rect 136500 4620 136510 4676
rect 138114 4620 138124 4676
rect 138180 4620 155148 4676
rect 155204 4620 155214 4676
rect 700 4228 756 4620
rect 67172 4564 67228 4620
rect 57026 4508 57036 4564
rect 57092 4508 65660 4564
rect 65716 4508 65726 4564
rect 67172 4508 70588 4564
rect 70644 4508 70654 4564
rect 105980 4508 109116 4564
rect 109172 4508 109182 4564
rect 123442 4508 123452 4564
rect 123508 4508 147084 4564
rect 147140 4508 147150 4564
rect 105980 4452 106036 4508
rect 5058 4396 5068 4452
rect 5124 4396 6636 4452
rect 6692 4396 6860 4452
rect 6916 4396 6926 4452
rect 25890 4396 25900 4452
rect 25956 4396 29260 4452
rect 29316 4396 29932 4452
rect 29988 4396 33964 4452
rect 34020 4396 34030 4452
rect 48738 4396 48748 4452
rect 48804 4396 50316 4452
rect 50372 4396 50382 4452
rect 63746 4396 63756 4452
rect 63812 4396 68684 4452
rect 68740 4396 68750 4452
rect 104738 4396 104748 4452
rect 104804 4396 105980 4452
rect 106036 4396 106046 4452
rect 108098 4396 108108 4452
rect 108164 4396 108444 4452
rect 108500 4396 109452 4452
rect 109508 4396 109518 4452
rect 128258 4396 128268 4452
rect 128324 4396 129052 4452
rect 129108 4396 129118 4452
rect 130162 4396 130172 4452
rect 130228 4396 131180 4452
rect 131236 4396 131964 4452
rect 132020 4396 132030 4452
rect 143714 4396 143724 4452
rect 143780 4396 147308 4452
rect 147364 4396 147374 4452
rect 5506 4284 5516 4340
rect 5572 4284 6188 4340
rect 6244 4284 12572 4340
rect 12628 4284 12638 4340
rect 23426 4284 23436 4340
rect 23492 4284 26460 4340
rect 26516 4284 26526 4340
rect 32386 4284 32396 4340
rect 32452 4284 37100 4340
rect 37156 4284 42476 4340
rect 42532 4284 62188 4340
rect 62244 4284 62254 4340
rect 66658 4284 66668 4340
rect 66724 4284 70476 4340
rect 70532 4284 78428 4340
rect 78484 4284 83916 4340
rect 83972 4284 83982 4340
rect 97234 4284 97244 4340
rect 97300 4284 98588 4340
rect 98644 4284 98654 4340
rect 105298 4284 105308 4340
rect 105364 4284 108780 4340
rect 108836 4284 118412 4340
rect 118468 4284 121212 4340
rect 121268 4284 138348 4340
rect 138404 4284 138414 4340
rect 700 4172 868 4228
rect 4162 4172 4172 4228
rect 4228 4172 4732 4228
rect 4788 4172 9660 4228
rect 9716 4172 9726 4228
rect 24882 4172 24892 4228
rect 24948 4172 26124 4228
rect 26180 4172 26190 4228
rect 28578 4172 28588 4228
rect 28644 4172 31612 4228
rect 31668 4172 31678 4228
rect 32834 4172 32844 4228
rect 32900 4172 34076 4228
rect 34132 4172 34142 4228
rect 45266 4172 45276 4228
rect 45332 4172 46620 4228
rect 46676 4172 46686 4228
rect 53218 4172 53228 4228
rect 53284 4172 53900 4228
rect 53956 4172 53966 4228
rect 55906 4172 55916 4228
rect 55972 4172 61068 4228
rect 61124 4172 61134 4228
rect 88274 4172 88284 4228
rect 88340 4172 92092 4228
rect 92148 4172 92158 4228
rect 93986 4172 93996 4228
rect 94052 4172 111916 4228
rect 111972 4172 111982 4228
rect 113138 4172 113148 4228
rect 113204 4172 114828 4228
rect 114884 4172 114894 4228
rect 116610 4172 116620 4228
rect 116676 4172 117516 4228
rect 117572 4172 117582 4228
rect 124002 4172 124012 4228
rect 124068 4172 125356 4228
rect 125412 4172 125422 4228
rect 127474 4172 127484 4228
rect 127540 4172 128044 4228
rect 128100 4172 130620 4228
rect 130676 4172 130686 4228
rect 130946 4172 130956 4228
rect 131012 4172 132524 4228
rect 132580 4172 132590 4228
rect 133634 4172 133644 4228
rect 133700 4172 137004 4228
rect 137060 4172 137070 4228
rect 137228 4172 139132 4228
rect 139188 4172 139198 4228
rect 139458 4172 139468 4228
rect 139524 4172 140476 4228
rect 140532 4172 140542 4228
rect 812 4116 868 4172
rect 137228 4116 137284 4172
rect 812 4060 11788 4116
rect 11844 4060 11854 4116
rect 45154 4060 45164 4116
rect 45220 4060 45836 4116
rect 45892 4060 49084 4116
rect 49140 4060 49150 4116
rect 52434 4060 52444 4116
rect 52500 4060 60900 4116
rect 135874 4060 135884 4116
rect 135940 4060 137284 4116
rect 137732 4060 139804 4116
rect 139860 4060 142940 4116
rect 142996 4060 143276 4116
rect 143332 4060 143836 4116
rect 143892 4060 143902 4116
rect 48066 3948 48076 4004
rect 48132 3948 55692 4004
rect 55748 3948 55758 4004
rect 20546 3892 20556 3948
rect 20612 3892 20660 3948
rect 20716 3892 20764 3948
rect 20820 3892 20868 3948
rect 20924 3892 20972 3948
rect 21028 3892 21076 3948
rect 21132 3892 21180 3948
rect 21236 3892 21284 3948
rect 21340 3892 21388 3948
rect 21444 3892 21454 3948
rect 59858 3892 59868 3948
rect 59924 3892 59972 3948
rect 60028 3892 60076 3948
rect 60132 3892 60180 3948
rect 60236 3892 60284 3948
rect 60340 3892 60388 3948
rect 60444 3892 60492 3948
rect 60548 3892 60596 3948
rect 60652 3892 60700 3948
rect 60756 3892 60766 3948
rect 60844 3892 60900 4060
rect 137732 4004 137788 4060
rect 136434 3948 136444 4004
rect 136500 3948 137788 4004
rect 99170 3892 99180 3948
rect 99236 3892 99284 3948
rect 99340 3892 99388 3948
rect 99444 3892 99492 3948
rect 99548 3892 99596 3948
rect 99652 3892 99700 3948
rect 99756 3892 99804 3948
rect 99860 3892 99908 3948
rect 99964 3892 100012 3948
rect 100068 3892 100078 3948
rect 138482 3892 138492 3948
rect 138548 3892 138596 3948
rect 138652 3892 138700 3948
rect 138756 3892 138804 3948
rect 138860 3892 138908 3948
rect 138964 3892 139012 3948
rect 139068 3892 139116 3948
rect 139172 3892 139220 3948
rect 139276 3892 139324 3948
rect 139380 3892 139390 3948
rect 60834 3836 60844 3892
rect 60900 3836 65548 3892
rect 65604 3836 65614 3892
rect 90962 3836 90972 3892
rect 91028 3836 92764 3892
rect 92820 3836 94108 3892
rect 94164 3836 94174 3892
rect 116050 3836 116060 3892
rect 116116 3836 119532 3892
rect 119588 3836 120652 3892
rect 120708 3836 122332 3892
rect 122388 3836 126140 3892
rect 126196 3836 127260 3892
rect 127316 3836 131180 3892
rect 131236 3836 131852 3892
rect 131908 3836 131918 3892
rect 51986 3724 51996 3780
rect 52052 3724 52892 3780
rect 52948 3724 52958 3780
rect 87042 3724 87052 3780
rect 87108 3724 88844 3780
rect 88900 3724 90188 3780
rect 90244 3724 90254 3780
rect 92082 3724 92092 3780
rect 92148 3724 111580 3780
rect 111636 3724 111646 3780
rect 124114 3724 124124 3780
rect 124180 3724 131964 3780
rect 132020 3724 132030 3780
rect 134082 3724 134092 3780
rect 134148 3724 152460 3780
rect 152516 3724 152526 3780
rect 7410 3612 7420 3668
rect 7476 3612 8764 3668
rect 8820 3612 8830 3668
rect 22754 3612 22764 3668
rect 22820 3612 29484 3668
rect 29540 3612 29550 3668
rect 39554 3612 39564 3668
rect 39620 3612 40012 3668
rect 40068 3612 40078 3668
rect 44146 3612 44156 3668
rect 44212 3612 47628 3668
rect 47684 3612 47694 3668
rect 52658 3612 52668 3668
rect 52724 3612 53788 3668
rect 53844 3612 54572 3668
rect 54628 3612 54638 3668
rect 59826 3612 59836 3668
rect 59892 3612 62972 3668
rect 63028 3612 65548 3668
rect 65604 3612 65614 3668
rect 67666 3612 67676 3668
rect 67732 3612 69132 3668
rect 69188 3612 69198 3668
rect 71362 3612 71372 3668
rect 71428 3612 72156 3668
rect 72212 3612 76636 3668
rect 76692 3612 80388 3668
rect 82562 3612 82572 3668
rect 82628 3612 83132 3668
rect 83188 3612 83198 3668
rect 84242 3612 84252 3668
rect 84308 3612 88172 3668
rect 88228 3612 93996 3668
rect 94052 3612 94062 3668
rect 94882 3612 94892 3668
rect 94948 3612 95340 3668
rect 95396 3612 96684 3668
rect 96740 3612 96750 3668
rect 119410 3612 119420 3668
rect 119476 3612 120092 3668
rect 120148 3612 120158 3668
rect 122882 3612 122892 3668
rect 122948 3612 123340 3668
rect 123396 3612 123406 3668
rect 139794 3612 139804 3668
rect 139860 3612 142044 3668
rect 142100 3612 142604 3668
rect 142660 3612 142670 3668
rect 144386 3612 144396 3668
rect 144452 3612 145852 3668
rect 145908 3612 145918 3668
rect 80332 3556 80388 3612
rect 12562 3500 12572 3556
rect 12628 3500 25676 3556
rect 25732 3500 32396 3556
rect 32452 3500 32462 3556
rect 37202 3500 37212 3556
rect 37268 3500 41356 3556
rect 41412 3500 41804 3556
rect 41860 3500 45164 3556
rect 45220 3500 45230 3556
rect 49186 3500 49196 3556
rect 49252 3500 53116 3556
rect 53172 3500 53182 3556
rect 53890 3500 53900 3556
rect 53956 3500 57036 3556
rect 57092 3500 63756 3556
rect 63812 3500 63822 3556
rect 80322 3500 80332 3556
rect 80388 3500 84140 3556
rect 84196 3500 84206 3556
rect 88946 3500 88956 3556
rect 89012 3500 95900 3556
rect 95956 3500 99820 3556
rect 99876 3500 99886 3556
rect 111570 3500 111580 3556
rect 111636 3500 124572 3556
rect 124628 3500 127372 3556
rect 127428 3500 135100 3556
rect 135156 3500 135166 3556
rect 138338 3500 138348 3556
rect 138404 3500 139020 3556
rect 139076 3500 139086 3556
rect 99820 3444 99876 3500
rect 31602 3388 31612 3444
rect 31668 3388 50316 3444
rect 50372 3388 50382 3444
rect 99820 3388 105308 3444
rect 105364 3388 105374 3444
rect 40202 3108 40212 3164
rect 40268 3108 40316 3164
rect 40372 3108 40420 3164
rect 40476 3108 40524 3164
rect 40580 3108 40628 3164
rect 40684 3108 40732 3164
rect 40788 3108 40836 3164
rect 40892 3108 40940 3164
rect 40996 3108 41044 3164
rect 41100 3108 41110 3164
rect 79514 3108 79524 3164
rect 79580 3108 79628 3164
rect 79684 3108 79732 3164
rect 79788 3108 79836 3164
rect 79892 3108 79940 3164
rect 79996 3108 80044 3164
rect 80100 3108 80148 3164
rect 80204 3108 80252 3164
rect 80308 3108 80356 3164
rect 80412 3108 80422 3164
rect 118826 3108 118836 3164
rect 118892 3108 118940 3164
rect 118996 3108 119044 3164
rect 119100 3108 119148 3164
rect 119204 3108 119252 3164
rect 119308 3108 119356 3164
rect 119412 3108 119460 3164
rect 119516 3108 119564 3164
rect 119620 3108 119668 3164
rect 119724 3108 119734 3164
rect 158138 3108 158148 3164
rect 158204 3108 158252 3164
rect 158308 3108 158356 3164
rect 158412 3108 158460 3164
rect 158516 3108 158564 3164
rect 158620 3108 158668 3164
rect 158724 3108 158772 3164
rect 158828 3108 158876 3164
rect 158932 3108 158980 3164
rect 159036 3108 159046 3164
rect 0 1764 800 1792
rect 0 1708 73948 1764
rect 74004 1708 74014 1764
rect 0 1680 800 1708
<< via3 >>
rect 40212 6244 40268 6300
rect 40316 6244 40372 6300
rect 40420 6244 40476 6300
rect 40524 6244 40580 6300
rect 40628 6244 40684 6300
rect 40732 6244 40788 6300
rect 40836 6244 40892 6300
rect 40940 6244 40996 6300
rect 41044 6244 41100 6300
rect 79524 6244 79580 6300
rect 79628 6244 79684 6300
rect 79732 6244 79788 6300
rect 79836 6244 79892 6300
rect 79940 6244 79996 6300
rect 80044 6244 80100 6300
rect 80148 6244 80204 6300
rect 80252 6244 80308 6300
rect 80356 6244 80412 6300
rect 118836 6244 118892 6300
rect 118940 6244 118996 6300
rect 119044 6244 119100 6300
rect 119148 6244 119204 6300
rect 119252 6244 119308 6300
rect 119356 6244 119412 6300
rect 119460 6244 119516 6300
rect 119564 6244 119620 6300
rect 119668 6244 119724 6300
rect 158148 6244 158204 6300
rect 158252 6244 158308 6300
rect 158356 6244 158412 6300
rect 158460 6244 158516 6300
rect 158564 6244 158620 6300
rect 158668 6244 158724 6300
rect 158772 6244 158828 6300
rect 158876 6244 158932 6300
rect 158980 6244 159036 6300
rect 20556 5460 20612 5516
rect 20660 5460 20716 5516
rect 20764 5460 20820 5516
rect 20868 5460 20924 5516
rect 20972 5460 21028 5516
rect 21076 5460 21132 5516
rect 21180 5460 21236 5516
rect 21284 5460 21340 5516
rect 21388 5460 21444 5516
rect 59868 5460 59924 5516
rect 59972 5460 60028 5516
rect 60076 5460 60132 5516
rect 60180 5460 60236 5516
rect 60284 5460 60340 5516
rect 60388 5460 60444 5516
rect 60492 5460 60548 5516
rect 60596 5460 60652 5516
rect 60700 5460 60756 5516
rect 99180 5460 99236 5516
rect 99284 5460 99340 5516
rect 99388 5460 99444 5516
rect 99492 5460 99548 5516
rect 99596 5460 99652 5516
rect 99700 5460 99756 5516
rect 99804 5460 99860 5516
rect 99908 5460 99964 5516
rect 100012 5460 100068 5516
rect 138492 5460 138548 5516
rect 138596 5460 138652 5516
rect 138700 5460 138756 5516
rect 138804 5460 138860 5516
rect 138908 5460 138964 5516
rect 139012 5460 139068 5516
rect 139116 5460 139172 5516
rect 139220 5460 139276 5516
rect 139324 5460 139380 5516
rect 40212 4676 40268 4732
rect 40316 4676 40372 4732
rect 40420 4676 40476 4732
rect 40524 4676 40580 4732
rect 40628 4676 40684 4732
rect 40732 4676 40788 4732
rect 40836 4676 40892 4732
rect 40940 4676 40996 4732
rect 41044 4676 41100 4732
rect 79524 4676 79580 4732
rect 79628 4676 79684 4732
rect 79732 4676 79788 4732
rect 79836 4676 79892 4732
rect 79940 4676 79996 4732
rect 80044 4676 80100 4732
rect 80148 4676 80204 4732
rect 80252 4676 80308 4732
rect 80356 4676 80412 4732
rect 118836 4676 118892 4732
rect 118940 4676 118996 4732
rect 119044 4676 119100 4732
rect 119148 4676 119204 4732
rect 119252 4676 119308 4732
rect 119356 4676 119412 4732
rect 119460 4676 119516 4732
rect 119564 4676 119620 4732
rect 119668 4676 119724 4732
rect 158148 4676 158204 4732
rect 158252 4676 158308 4732
rect 158356 4676 158412 4732
rect 158460 4676 158516 4732
rect 158564 4676 158620 4732
rect 158668 4676 158724 4732
rect 158772 4676 158828 4732
rect 158876 4676 158932 4732
rect 158980 4676 159036 4732
rect 20556 3892 20612 3948
rect 20660 3892 20716 3948
rect 20764 3892 20820 3948
rect 20868 3892 20924 3948
rect 20972 3892 21028 3948
rect 21076 3892 21132 3948
rect 21180 3892 21236 3948
rect 21284 3892 21340 3948
rect 21388 3892 21444 3948
rect 59868 3892 59924 3948
rect 59972 3892 60028 3948
rect 60076 3892 60132 3948
rect 60180 3892 60236 3948
rect 60284 3892 60340 3948
rect 60388 3892 60444 3948
rect 60492 3892 60548 3948
rect 60596 3892 60652 3948
rect 60700 3892 60756 3948
rect 99180 3892 99236 3948
rect 99284 3892 99340 3948
rect 99388 3892 99444 3948
rect 99492 3892 99548 3948
rect 99596 3892 99652 3948
rect 99700 3892 99756 3948
rect 99804 3892 99860 3948
rect 99908 3892 99964 3948
rect 100012 3892 100068 3948
rect 138492 3892 138548 3948
rect 138596 3892 138652 3948
rect 138700 3892 138756 3948
rect 138804 3892 138860 3948
rect 138908 3892 138964 3948
rect 139012 3892 139068 3948
rect 139116 3892 139172 3948
rect 139220 3892 139276 3948
rect 139324 3892 139380 3948
rect 40212 3108 40268 3164
rect 40316 3108 40372 3164
rect 40420 3108 40476 3164
rect 40524 3108 40580 3164
rect 40628 3108 40684 3164
rect 40732 3108 40788 3164
rect 40836 3108 40892 3164
rect 40940 3108 40996 3164
rect 41044 3108 41100 3164
rect 79524 3108 79580 3164
rect 79628 3108 79684 3164
rect 79732 3108 79788 3164
rect 79836 3108 79892 3164
rect 79940 3108 79996 3164
rect 80044 3108 80100 3164
rect 80148 3108 80204 3164
rect 80252 3108 80308 3164
rect 80356 3108 80412 3164
rect 118836 3108 118892 3164
rect 118940 3108 118996 3164
rect 119044 3108 119100 3164
rect 119148 3108 119204 3164
rect 119252 3108 119308 3164
rect 119356 3108 119412 3164
rect 119460 3108 119516 3164
rect 119564 3108 119620 3164
rect 119668 3108 119724 3164
rect 158148 3108 158204 3164
rect 158252 3108 158308 3164
rect 158356 3108 158412 3164
rect 158460 3108 158516 3164
rect 158564 3108 158620 3164
rect 158668 3108 158724 3164
rect 158772 3108 158828 3164
rect 158876 3108 158932 3164
rect 158980 3108 159036 3164
<< metal4 >>
rect 20500 5516 21500 6332
rect 20500 5460 20556 5516
rect 20612 5460 20660 5516
rect 20716 5460 20764 5516
rect 20820 5460 20868 5516
rect 20924 5460 20972 5516
rect 21028 5460 21076 5516
rect 21132 5460 21180 5516
rect 21236 5460 21284 5516
rect 21340 5460 21388 5516
rect 21444 5460 21500 5516
rect 20500 3948 21500 5460
rect 20500 3892 20556 3948
rect 20612 3892 20660 3948
rect 20716 3892 20764 3948
rect 20820 3892 20868 3948
rect 20924 3892 20972 3948
rect 21028 3892 21076 3948
rect 21132 3892 21180 3948
rect 21236 3892 21284 3948
rect 21340 3892 21388 3948
rect 21444 3892 21500 3948
rect 20500 3076 21500 3892
rect 40156 6300 41156 6332
rect 40156 6244 40212 6300
rect 40268 6244 40316 6300
rect 40372 6244 40420 6300
rect 40476 6244 40524 6300
rect 40580 6244 40628 6300
rect 40684 6244 40732 6300
rect 40788 6244 40836 6300
rect 40892 6244 40940 6300
rect 40996 6244 41044 6300
rect 41100 6244 41156 6300
rect 40156 4732 41156 6244
rect 40156 4676 40212 4732
rect 40268 4676 40316 4732
rect 40372 4676 40420 4732
rect 40476 4676 40524 4732
rect 40580 4676 40628 4732
rect 40684 4676 40732 4732
rect 40788 4676 40836 4732
rect 40892 4676 40940 4732
rect 40996 4676 41044 4732
rect 41100 4676 41156 4732
rect 40156 3164 41156 4676
rect 40156 3108 40212 3164
rect 40268 3108 40316 3164
rect 40372 3108 40420 3164
rect 40476 3108 40524 3164
rect 40580 3108 40628 3164
rect 40684 3108 40732 3164
rect 40788 3108 40836 3164
rect 40892 3108 40940 3164
rect 40996 3108 41044 3164
rect 41100 3108 41156 3164
rect 40156 3076 41156 3108
rect 59812 5516 60812 6332
rect 59812 5460 59868 5516
rect 59924 5460 59972 5516
rect 60028 5460 60076 5516
rect 60132 5460 60180 5516
rect 60236 5460 60284 5516
rect 60340 5460 60388 5516
rect 60444 5460 60492 5516
rect 60548 5460 60596 5516
rect 60652 5460 60700 5516
rect 60756 5460 60812 5516
rect 59812 3948 60812 5460
rect 59812 3892 59868 3948
rect 59924 3892 59972 3948
rect 60028 3892 60076 3948
rect 60132 3892 60180 3948
rect 60236 3892 60284 3948
rect 60340 3892 60388 3948
rect 60444 3892 60492 3948
rect 60548 3892 60596 3948
rect 60652 3892 60700 3948
rect 60756 3892 60812 3948
rect 59812 3076 60812 3892
rect 79468 6300 80468 6332
rect 79468 6244 79524 6300
rect 79580 6244 79628 6300
rect 79684 6244 79732 6300
rect 79788 6244 79836 6300
rect 79892 6244 79940 6300
rect 79996 6244 80044 6300
rect 80100 6244 80148 6300
rect 80204 6244 80252 6300
rect 80308 6244 80356 6300
rect 80412 6244 80468 6300
rect 79468 4732 80468 6244
rect 79468 4676 79524 4732
rect 79580 4676 79628 4732
rect 79684 4676 79732 4732
rect 79788 4676 79836 4732
rect 79892 4676 79940 4732
rect 79996 4676 80044 4732
rect 80100 4676 80148 4732
rect 80204 4676 80252 4732
rect 80308 4676 80356 4732
rect 80412 4676 80468 4732
rect 79468 3164 80468 4676
rect 79468 3108 79524 3164
rect 79580 3108 79628 3164
rect 79684 3108 79732 3164
rect 79788 3108 79836 3164
rect 79892 3108 79940 3164
rect 79996 3108 80044 3164
rect 80100 3108 80148 3164
rect 80204 3108 80252 3164
rect 80308 3108 80356 3164
rect 80412 3108 80468 3164
rect 79468 3076 80468 3108
rect 99124 5516 100124 6332
rect 99124 5460 99180 5516
rect 99236 5460 99284 5516
rect 99340 5460 99388 5516
rect 99444 5460 99492 5516
rect 99548 5460 99596 5516
rect 99652 5460 99700 5516
rect 99756 5460 99804 5516
rect 99860 5460 99908 5516
rect 99964 5460 100012 5516
rect 100068 5460 100124 5516
rect 99124 3948 100124 5460
rect 99124 3892 99180 3948
rect 99236 3892 99284 3948
rect 99340 3892 99388 3948
rect 99444 3892 99492 3948
rect 99548 3892 99596 3948
rect 99652 3892 99700 3948
rect 99756 3892 99804 3948
rect 99860 3892 99908 3948
rect 99964 3892 100012 3948
rect 100068 3892 100124 3948
rect 99124 3076 100124 3892
rect 118780 6300 119780 6332
rect 118780 6244 118836 6300
rect 118892 6244 118940 6300
rect 118996 6244 119044 6300
rect 119100 6244 119148 6300
rect 119204 6244 119252 6300
rect 119308 6244 119356 6300
rect 119412 6244 119460 6300
rect 119516 6244 119564 6300
rect 119620 6244 119668 6300
rect 119724 6244 119780 6300
rect 118780 4732 119780 6244
rect 118780 4676 118836 4732
rect 118892 4676 118940 4732
rect 118996 4676 119044 4732
rect 119100 4676 119148 4732
rect 119204 4676 119252 4732
rect 119308 4676 119356 4732
rect 119412 4676 119460 4732
rect 119516 4676 119564 4732
rect 119620 4676 119668 4732
rect 119724 4676 119780 4732
rect 118780 3164 119780 4676
rect 118780 3108 118836 3164
rect 118892 3108 118940 3164
rect 118996 3108 119044 3164
rect 119100 3108 119148 3164
rect 119204 3108 119252 3164
rect 119308 3108 119356 3164
rect 119412 3108 119460 3164
rect 119516 3108 119564 3164
rect 119620 3108 119668 3164
rect 119724 3108 119780 3164
rect 118780 3076 119780 3108
rect 138436 5516 139436 6332
rect 138436 5460 138492 5516
rect 138548 5460 138596 5516
rect 138652 5460 138700 5516
rect 138756 5460 138804 5516
rect 138860 5460 138908 5516
rect 138964 5460 139012 5516
rect 139068 5460 139116 5516
rect 139172 5460 139220 5516
rect 139276 5460 139324 5516
rect 139380 5460 139436 5516
rect 138436 3948 139436 5460
rect 138436 3892 138492 3948
rect 138548 3892 138596 3948
rect 138652 3892 138700 3948
rect 138756 3892 138804 3948
rect 138860 3892 138908 3948
rect 138964 3892 139012 3948
rect 139068 3892 139116 3948
rect 139172 3892 139220 3948
rect 139276 3892 139324 3948
rect 139380 3892 139436 3948
rect 138436 3076 139436 3892
rect 158092 6300 159092 6332
rect 158092 6244 158148 6300
rect 158204 6244 158252 6300
rect 158308 6244 158356 6300
rect 158412 6244 158460 6300
rect 158516 6244 158564 6300
rect 158620 6244 158668 6300
rect 158724 6244 158772 6300
rect 158828 6244 158876 6300
rect 158932 6244 158980 6300
rect 159036 6244 159092 6300
rect 158092 4732 159092 6244
rect 158092 4676 158148 4732
rect 158204 4676 158252 4732
rect 158308 4676 158356 4732
rect 158412 4676 158460 4732
rect 158516 4676 158564 4732
rect 158620 4676 158668 4732
rect 158724 4676 158772 4732
rect 158828 4676 158876 4732
rect 158932 4676 158980 4732
rect 159036 4676 159092 4732
rect 158092 3164 159092 4676
rect 158092 3108 158148 3164
rect 158204 3108 158252 3164
rect 158308 3108 158356 3164
rect 158412 3108 158460 3164
rect 158516 3108 158564 3164
rect 158620 3108 158668 3164
rect 158724 3108 158772 3164
rect 158828 3108 158876 3164
rect 158932 3108 158980 3164
rect 159036 3108 159092 3164
rect 158092 3076 159092 3108
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1667941163
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1667941163
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1667941163
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102
timestamp 1667941163
transform 1 0 12768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 13328 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142
timestamp 1667941163
transform 1 0 17248 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_177
timestamp 1667941163
transform 1 0 21168 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1667941163
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_212
timestamp 1667941163
transform 1 0 25088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_214
timestamp 1667941163
transform 1 0 25312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1667941163
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_247
timestamp 1667941163
transform 1 0 29008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_249
timestamp 1667941163
transform 1 0 29232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1667941163
transform 1 0 32928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1667941163
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1667941163
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1667941163
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1667941163
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_352
timestamp 1667941163
transform 1 0 40768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_354
timestamp 1667941163
transform 1 0 40992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1667941163
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_387
timestamp 1667941163
transform 1 0 44688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_389
timestamp 1667941163
transform 1 0 44912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1667941163
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_422
timestamp 1667941163
transform 1 0 48608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_424
timestamp 1667941163
transform 1 0 48832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1667941163
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_457
timestamp 1667941163
transform 1 0 52528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_459
timestamp 1667941163
transform 1 0 52752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1667941163
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_492
timestamp 1667941163
transform 1 0 56448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_494
timestamp 1667941163
transform 1 0 56672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1667941163
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_527
timestamp 1667941163
transform 1 0 60368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_529
timestamp 1667941163
transform 1 0 60592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1667941163
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_562
timestamp 1667941163
transform 1 0 64288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_564
timestamp 1667941163
transform 1 0 64512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1667941163
transform 1 0 67872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1667941163
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_627
timestamp 1667941163
transform 1 0 71568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1667941163
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_632
timestamp 1667941163
transform 1 0 72128 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1667941163
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_667
timestamp 1667941163
transform 1 0 76048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_669
timestamp 1667941163
transform 1 0 76272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_699
timestamp 1667941163
transform 1 0 79632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1667941163
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_732
timestamp 1667941163
transform 1 0 83328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_734
timestamp 1667941163
transform 1 0 83552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_737
timestamp 1667941163
transform 1 0 83888 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_767
timestamp 1667941163
transform 1 0 87248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_769
timestamp 1667941163
transform 1 0 87472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1667941163
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_802
timestamp 1667941163
transform 1 0 91168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_804
timestamp 1667941163
transform 1 0 91392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1667941163
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_837
timestamp 1667941163
transform 1 0 95088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1667941163
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_842
timestamp 1667941163
transform 1 0 95648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_872
timestamp 1667941163
transform 1 0 99008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1667941163
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1667941163
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_907
timestamp 1667941163
transform 1 0 102928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_909
timestamp 1667941163
transform 1 0 103152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_912
timestamp 1667941163
transform 1 0 103488 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_944
timestamp 1667941163
transform 1 0 107072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_947
timestamp 1667941163
transform 1 0 107408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_977
timestamp 1667941163
transform 1 0 110768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1667941163
transform 1 0 110992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1667941163
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1012
timestamp 1667941163
transform 1 0 114688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1667941163
transform 1 0 114912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1667941163
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1047
timestamp 1667941163
transform 1 0 118608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1049
timestamp 1667941163
transform 1 0 118832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1052
timestamp 1667941163
transform 1 0 119168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1082
timestamp 1667941163
transform 1 0 122528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1667941163
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1667941163
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1117
timestamp 1667941163
transform 1 0 126448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1119
timestamp 1667941163
transform 1 0 126672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1667941163
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1152
timestamp 1667941163
transform 1 0 130368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1667941163
transform 1 0 130592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1667941163
transform 1 0 130928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1187
timestamp 1667941163
transform 1 0 134288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1189
timestamp 1667941163
transform 1 0 134512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1192
timestamp 1667941163
transform 1 0 134848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1222
timestamp 1667941163
transform 1 0 138208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1224
timestamp 1667941163
transform 1 0 138432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1667941163
transform 1 0 138768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1257
timestamp 1667941163
transform 1 0 142128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1259
timestamp 1667941163
transform 1 0 142352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1262
timestamp 1667941163
transform 1 0 142688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1292
timestamp 1667941163
transform 1 0 146048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1294
timestamp 1667941163
transform 1 0 146272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1297
timestamp 1667941163
transform 1 0 146608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1329
timestamp 1667941163
transform 1 0 150192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1332
timestamp 1667941163
transform 1 0 150528 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1364
timestamp 1667941163
transform 1 0 154112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1367
timestamp 1667941163
transform 1 0 154448 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1399
timestamp 1667941163
transform 1 0 158032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_39
timestamp 1667941163
transform 1 0 5712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_73 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 9520 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_89
timestamp 1667941163
transform 1 0 11312 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_97 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 12208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_130
timestamp 1667941163
transform 1 0 15904 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_138
timestamp 1667941163
transform 1 0 16800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_144
timestamp 1667941163
transform 1 0 17472 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_176
timestamp 1667941163
transform 1 0 21056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_180
timestamp 1667941163
transform 1 0 21504 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_182
timestamp 1667941163
transform 1 0 21728 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_215
timestamp 1667941163
transform 1 0 25424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_252
timestamp 1667941163
transform 1 0 29568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1667941163
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_286
timestamp 1667941163
transform 1 0 33376 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_302
timestamp 1667941163
transform 1 0 35168 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_310
timestamp 1667941163
transform 1 0 36064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_314
timestamp 1667941163
transform 1 0 36512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_316
timestamp 1667941163
transform 1 0 36736 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_346
timestamp 1667941163
transform 1 0 40096 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1667941163
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_357
timestamp 1667941163
transform 1 0 41328 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_394
timestamp 1667941163
transform 1 0 45472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1667941163
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_428
timestamp 1667941163
transform 1 0 49280 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_465
timestamp 1667941163
transform 1 0 53424 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1667941163
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_499
timestamp 1667941163
transform 1 0 57232 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_515
timestamp 1667941163
transform 1 0 59024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1667941163
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1667941163
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_621
timestamp 1667941163
transform 1 0 70896 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_637
timestamp 1667941163
transform 1 0 72688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1667941163
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_692
timestamp 1667941163
transform 1 0 78848 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_708
timestamp 1667941163
transform 1 0 80640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_712
timestamp 1667941163
transform 1 0 81088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_728
timestamp 1667941163
transform 1 0 82880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1667941163
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_783
timestamp 1667941163
transform 1 0 89040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_834
timestamp 1667941163
transform 1 0 94752 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_850
timestamp 1667941163
transform 1 0 96544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_854
timestamp 1667941163
transform 1 0 96992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_884
timestamp 1667941163
transform 1 0 100352 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_916
timestamp 1667941163
transform 1 0 103936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_920
timestamp 1667941163
transform 1 0 104384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_922
timestamp 1667941163
transform 1 0 104608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_925
timestamp 1667941163
transform 1 0 104944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_955
timestamp 1667941163
transform 1 0 108304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_986
timestamp 1667941163
transform 1 0 111776 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1667941163
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1026
timestamp 1667941163
transform 1 0 116256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1057
timestamp 1667941163
transform 1 0 119728 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1067
timestamp 1667941163
transform 1 0 120848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1097
timestamp 1667941163
transform 1 0 124208 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1128
timestamp 1667941163
transform 1 0 127680 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1667941163
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1168
timestamp 1667941163
transform 1 0 132160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1199
timestamp 1667941163
transform 1 0 135632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1209
timestamp 1667941163
transform 1 0 136752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1239
timestamp 1667941163
transform 1 0 140112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1270
timestamp 1667941163
transform 1 0 143584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1280 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 144704 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1344
timestamp 1667941163
transform 1 0 151872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1348
timestamp 1667941163
transform 1 0 152320 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_1351
timestamp 1667941163
transform 1 0 152656 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1383
timestamp 1667941163
transform 1 0 156240 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1399
timestamp 1667941163
transform 1 0 158032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1401
timestamp 1667941163
transform 1 0 158256 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_2
timestamp 1667941163
transform 1 0 1568 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_4
timestamp 1667941163
transform 1 0 1792 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_37
timestamp 1667941163
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_74
timestamp 1667941163
transform 1 0 9632 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_108
timestamp 1667941163
transform 1 0 13440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_110
timestamp 1667941163
transform 1 0 13664 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_140
timestamp 1667941163
transform 1 0 17024 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_144
timestamp 1667941163
transform 1 0 17472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_146
timestamp 1667941163
transform 1 0 17696 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_179
timestamp 1667941163
transform 1 0 21392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_216
timestamp 1667941163
transform 1 0 25536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1667941163
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_250
timestamp 1667941163
transform 1 0 29344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_287
timestamp 1667941163
transform 1 0 33488 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1667941163
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_321
timestamp 1667941163
transform 1 0 37296 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_358
timestamp 1667941163
transform 1 0 41440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1667941163
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_392
timestamp 1667941163
transform 1 0 45248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_429
timestamp 1667941163
transform 1 0 49392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1667941163
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_463
timestamp 1667941163
transform 1 0 53200 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_479
timestamp 1667941163
transform 1 0 54992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1667941163
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1667941163
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_585
timestamp 1667941163
transform 1 0 66864 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_601
timestamp 1667941163
transform 1 0 68656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1667941163
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_635
timestamp 1667941163
transform 1 0 72464 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_643
timestamp 1667941163
transform 1 0 73360 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1667941163
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_676
timestamp 1667941163
transform 1 0 77056 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_692
timestamp 1667941163
transform 1 0 78848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1667941163
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_747
timestamp 1667941163
transform 1 0 85008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_798
timestamp 1667941163
transform 1 0 90720 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_814
timestamp 1667941163
transform 1 0 92512 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_818
timestamp 1667941163
transform 1 0 92960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_848
timestamp 1667941163
transform 1 0 96320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_879
timestamp 1667941163
transform 1 0 99792 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_889
timestamp 1667941163
transform 1 0 100912 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_897
timestamp 1667941163
transform 1 0 101808 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_901
timestamp 1667941163
transform 1 0 102256 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_931
timestamp 1667941163
transform 1 0 105616 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_947
timestamp 1667941163
transform 1 0 107408 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_955
timestamp 1667941163
transform 1 0 108304 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1667941163
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_960
timestamp 1667941163
transform 1 0 108864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_990
timestamp 1667941163
transform 1 0 112224 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1021
timestamp 1667941163
transform 1 0 115696 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1667941163
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1061
timestamp 1667941163
transform 1 0 120176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1092
timestamp 1667941163
transform 1 0 123648 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1102
timestamp 1667941163
transform 1 0 124768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1132
timestamp 1667941163
transform 1 0 128128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1163
timestamp 1667941163
transform 1 0 131600 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1173
timestamp 1667941163
transform 1 0 132720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1203
timestamp 1667941163
transform 1 0 136080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1234
timestamp 1667941163
transform 1 0 139552 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1244
timestamp 1667941163
transform 1 0 140672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1274
timestamp 1667941163
transform 1 0 144032 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1305
timestamp 1667941163
transform 1 0 147504 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1315
timestamp 1667941163
transform 1 0 148624 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1379
timestamp 1667941163
transform 1 0 155792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1383
timestamp 1667941163
transform 1 0 156240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1386
timestamp 1667941163
transform 1 0 156576 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_2
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_4
timestamp 1667941163
transform 1 0 1792 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_34
timestamp 1667941163
transform 1 0 5152 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_37
timestamp 1667941163
transform 1 0 5488 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_39
timestamp 1667941163
transform 1 0 5712 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_69
timestamp 1667941163
transform 1 0 9072 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_72
timestamp 1667941163
transform 1 0 9408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_74
timestamp 1667941163
transform 1 0 9632 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_104
timestamp 1667941163
transform 1 0 12992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_107
timestamp 1667941163
transform 1 0 13328 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_109
timestamp 1667941163
transform 1 0 13552 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_139
timestamp 1667941163
transform 1 0 16912 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_142
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1667941163
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_174
timestamp 1667941163
transform 1 0 20832 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_177
timestamp 1667941163
transform 1 0 21168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_179
timestamp 1667941163
transform 1 0 21392 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1667941163
transform 1 0 24752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_212
timestamp 1667941163
transform 1 0 25088 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_214
timestamp 1667941163
transform 1 0 25312 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_244
timestamp 1667941163
transform 1 0 28672 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_247
timestamp 1667941163
transform 1 0 29008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_249
timestamp 1667941163
transform 1 0 29232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 32592 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1667941163
transform 1 0 32928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_284
timestamp 1667941163
transform 1 0 33152 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_314
timestamp 1667941163
transform 1 0 36512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_317
timestamp 1667941163
transform 1 0 36848 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_319
timestamp 1667941163
transform 1 0 37072 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1667941163
transform 1 0 40432 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_352
timestamp 1667941163
transform 1 0 40768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1667941163
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_384
timestamp 1667941163
transform 1 0 44352 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_387
timestamp 1667941163
transform 1 0 44688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_389
timestamp 1667941163
transform 1 0 44912 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1667941163
transform 1 0 48272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_422
timestamp 1667941163
transform 1 0 48608 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_424
timestamp 1667941163
transform 1 0 48832 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_454
timestamp 1667941163
transform 1 0 52192 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_457
timestamp 1667941163
transform 1 0 52528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_459
timestamp 1667941163
transform 1 0 52752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_489
timestamp 1667941163
transform 1 0 56112 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_492
timestamp 1667941163
transform 1 0 56448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_494
timestamp 1667941163
transform 1 0 56672 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_524
timestamp 1667941163
transform 1 0 60032 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_527
timestamp 1667941163
transform 1 0 60368 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_529
timestamp 1667941163
transform 1 0 60592 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_559
timestamp 1667941163
transform 1 0 63952 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_562
timestamp 1667941163
transform 1 0 64288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_564
timestamp 1667941163
transform 1 0 64512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_594
timestamp 1667941163
transform 1 0 67872 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_597
timestamp 1667941163
transform 1 0 68208 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_599
timestamp 1667941163
transform 1 0 68432 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_629
timestamp 1667941163
transform 1 0 71792 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_632
timestamp 1667941163
transform 1 0 72128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_634
timestamp 1667941163
transform 1 0 72352 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_664
timestamp 1667941163
transform 1 0 75712 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_667
timestamp 1667941163
transform 1 0 76048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_669
timestamp 1667941163
transform 1 0 76272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_699
timestamp 1667941163
transform 1 0 79632 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_702
timestamp 1667941163
transform 1 0 79968 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_732
timestamp 1667941163
transform 1 0 83328 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_734
timestamp 1667941163
transform 1 0 83552 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_737
timestamp 1667941163
transform 1 0 83888 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_767
timestamp 1667941163
transform 1 0 87248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_769
timestamp 1667941163
transform 1 0 87472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_772
timestamp 1667941163
transform 1 0 87808 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_802
timestamp 1667941163
transform 1 0 91168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_804
timestamp 1667941163
transform 1 0 91392 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_807
timestamp 1667941163
transform 1 0 91728 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_837
timestamp 1667941163
transform 1 0 95088 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_839
timestamp 1667941163
transform 1 0 95312 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_842
timestamp 1667941163
transform 1 0 95648 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_872
timestamp 1667941163
transform 1 0 99008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_874
timestamp 1667941163
transform 1 0 99232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_877
timestamp 1667941163
transform 1 0 99568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_907
timestamp 1667941163
transform 1 0 102928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_909
timestamp 1667941163
transform 1 0 103152 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_912
timestamp 1667941163
transform 1 0 103488 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_914
timestamp 1667941163
transform 1 0 103712 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_944
timestamp 1667941163
transform 1 0 107072 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_947
timestamp 1667941163
transform 1 0 107408 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_977
timestamp 1667941163
transform 1 0 110768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_979
timestamp 1667941163
transform 1 0 110992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_982
timestamp 1667941163
transform 1 0 111328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1012
timestamp 1667941163
transform 1 0 114688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1014
timestamp 1667941163
transform 1 0 114912 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1017
timestamp 1667941163
transform 1 0 115248 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1047
timestamp 1667941163
transform 1 0 118608 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1049
timestamp 1667941163
transform 1 0 118832 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1052
timestamp 1667941163
transform 1 0 119168 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1082
timestamp 1667941163
transform 1 0 122528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1084
timestamp 1667941163
transform 1 0 122752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1087
timestamp 1667941163
transform 1 0 123088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1117
timestamp 1667941163
transform 1 0 126448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1119
timestamp 1667941163
transform 1 0 126672 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1122
timestamp 1667941163
transform 1 0 127008 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1152
timestamp 1667941163
transform 1 0 130368 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1154
timestamp 1667941163
transform 1 0 130592 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1157
timestamp 1667941163
transform 1 0 130928 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1187
timestamp 1667941163
transform 1 0 134288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1189
timestamp 1667941163
transform 1 0 134512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1192
timestamp 1667941163
transform 1 0 134848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1222
timestamp 1667941163
transform 1 0 138208 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1224
timestamp 1667941163
transform 1 0 138432 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1227
timestamp 1667941163
transform 1 0 138768 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1257
timestamp 1667941163
transform 1 0 142128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1259
timestamp 1667941163
transform 1 0 142352 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1262
timestamp 1667941163
transform 1 0 142688 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1292
timestamp 1667941163
transform 1 0 146048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1294
timestamp 1667941163
transform 1 0 146272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1297
timestamp 1667941163
transform 1 0 146608 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1329
timestamp 1667941163
transform 1 0 150192 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1332
timestamp 1667941163
transform 1 0 150528 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1364
timestamp 1667941163
transform 1 0 154112 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1367
timestamp 1667941163
transform 1 0 154448 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1399
timestamp 1667941163
transform 1 0 158032 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 158592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 158592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 158592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 158592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_8 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_9
timestamp 1667941163
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_10
timestamp 1667941163
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_11
timestamp 1667941163
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_12
timestamp 1667941163
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_13
timestamp 1667941163
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_14
timestamp 1667941163
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_15
timestamp 1667941163
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_16
timestamp 1667941163
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_17
timestamp 1667941163
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18
timestamp 1667941163
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1667941163
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1667941163
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1667941163
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1667941163
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_23
timestamp 1667941163
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24
timestamp 1667941163
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1667941163
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1667941163
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1667941163
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1667941163
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1667941163
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1667941163
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1667941163
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1667941163
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1667941163
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1667941163
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1667941163
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1667941163
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1667941163
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1667941163
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1667941163
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1667941163
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1667941163
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1667941163
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1667941163
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1667941163
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1667941163
transform 1 0 150304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1667941163
transform 1 0 154224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1667941163
transform 1 0 158144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1667941163
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1667941163
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1667941163
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1667941163
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1667941163
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1667941163
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1667941163
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1667941163
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1667941163
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1667941163
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1667941163
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1667941163
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1667941163
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1667941163
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1667941163
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1667941163
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1667941163
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1667941163
transform 1 0 152432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1667941163
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1667941163
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1667941163
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1667941163
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1667941163
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1667941163
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1667941163
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1667941163
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1667941163
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1667941163
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1667941163
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1667941163
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1667941163
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1667941163
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_81
timestamp 1667941163
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_82
timestamp 1667941163
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_83
timestamp 1667941163
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1667941163
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1667941163
transform 1 0 148400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1667941163
transform 1 0 156352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1667941163
transform 1 0 5264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1667941163
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1667941163
transform 1 0 13104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1667941163
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1667941163
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1667941163
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1667941163
transform 1 0 28784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1667941163
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1667941163
transform 1 0 36624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1667941163
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1667941163
transform 1 0 44464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1667941163
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1667941163
transform 1 0 52304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1667941163
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1667941163
transform 1 0 60144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1667941163
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1667941163
transform 1 0 67984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1667941163
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1667941163
transform 1 0 75824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1667941163
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1667941163
transform 1 0 83664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1667941163
transform 1 0 87584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1667941163
transform 1 0 91504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1667941163
transform 1 0 95424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1667941163
transform 1 0 99344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1667941163
transform 1 0 103264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1667941163
transform 1 0 107184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1667941163
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1667941163
transform 1 0 115024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1667941163
transform 1 0 118944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1667941163
transform 1 0 122864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1667941163
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1667941163
transform 1 0 130704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1667941163
transform 1 0 134624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1667941163
transform 1 0 138544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1667941163
transform 1 0 142464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1667941163
transform 1 0 146384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1667941163
transform 1 0 150304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1667941163
transform 1 0 154224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1667941163
transform 1 0 158144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _000_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 25760 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _001_
timestamp 1667941163
transform 1 0 29792 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _002_
timestamp 1667941163
transform 1 0 33712 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _003_
timestamp 1667941163
transform 1 0 36960 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _004_
timestamp 1667941163
transform 1 0 37184 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _005_
timestamp 1667941163
transform 1 0 41664 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _006_
timestamp 1667941163
transform 1 0 41104 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _007_
timestamp 1667941163
transform 1 0 45696 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _008_
timestamp 1667941163
transform 1 0 48944 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _009_
timestamp 1667941163
transform 1 0 69216 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _010_
timestamp 1667941163
transform 1 0 72464 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _011_
timestamp 1667941163
transform 1 0 76384 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _012_
timestamp 1667941163
transform 1 0 80080 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _013_
timestamp 1667941163
transform 1 0 84000 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _014_
timestamp 1667941163
transform -1 0 91168 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _015_
timestamp 1667941163
transform -1 0 95088 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _016_
timestamp 1667941163
transform -1 0 96320 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _017_
timestamp 1667941163
transform -1 0 99008 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _018_
timestamp 1667941163
transform -1 0 100352 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _019_
timestamp 1667941163
transform -1 0 102928 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _020_
timestamp 1667941163
transform 1 0 120400 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _021_
timestamp 1667941163
transform 1 0 127120 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _022_
timestamp 1667941163
transform 1 0 131040 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _023_
timestamp 1667941163
transform 1 0 134960 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _024_
timestamp 1667941163
transform 1 0 136304 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _025_
timestamp 1667941163
transform -1 0 110768 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _026_
timestamp 1667941163
transform 1 0 103824 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _027_
timestamp 1667941163
transform 1 0 107520 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _028_
timestamp 1667941163
transform -1 0 114688 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _029_
timestamp 1667941163
transform -1 0 116256 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _030_
timestamp 1667941163
transform -1 0 119728 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _031_
timestamp 1667941163
transform -1 0 122528 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _032_
timestamp 1667941163
transform -1 0 126448 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _033_
timestamp 1667941163
transform -1 0 131600 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _034_
timestamp 1667941163
transform -1 0 132160 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _035_
timestamp 1667941163
transform -1 0 135632 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _036_
timestamp 1667941163
transform -1 0 140112 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _037_
timestamp 1667941163
transform -1 0 144032 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _038_
timestamp 1667941163
transform -1 0 143584 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _039_
timestamp 1667941163
transform -1 0 146048 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _040_
timestamp 1667941163
transform 1 0 142800 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _041_
timestamp 1667941163
transform -1 0 12768 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _042_
timestamp 1667941163
transform -1 0 5712 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _043_
timestamp 1667941163
transform 1 0 1904 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _044_
timestamp 1667941163
transform 1 0 5936 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _045_
timestamp 1667941163
transform -1 0 9072 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _046_
timestamp 1667941163
transform 1 0 9744 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _047_
timestamp 1667941163
transform 1 0 13776 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _048_
timestamp 1667941163
transform 1 0 17808 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _049_
timestamp 1667941163
transform 1 0 30240 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _050_
timestamp 1667941163
transform 1 0 45024 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _051_
timestamp 1667941163
transform 1 0 49616 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _052_
timestamp 1667941163
transform 1 0 53648 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _053_
timestamp 1667941163
transform 1 0 56784 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _054_
timestamp 1667941163
transform 1 0 56784 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _055_
timestamp 1667941163
transform -1 0 63952 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _056_
timestamp 1667941163
transform -1 0 53424 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _057_
timestamp 1667941163
transform -1 0 32592 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _058_
timestamp 1667941163
transform 1 0 21504 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _059_
timestamp 1667941163
transform 1 0 25424 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _060_
timestamp 1667941163
transform 1 0 25424 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _061_
timestamp 1667941163
transform 1 0 29344 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _062_
timestamp 1667941163
transform 1 0 33264 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _063_
timestamp 1667941163
transform 1 0 36848 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _064_
timestamp 1667941163
transform 1 0 38192 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _065_
timestamp 1667941163
transform 1 0 41104 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _066_
timestamp 1667941163
transform 1 0 42224 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _067_
timestamp 1667941163
transform 1 0 46144 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _068_
timestamp 1667941163
transform 1 0 52864 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _069_
timestamp 1667941163
transform 1 0 68544 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _070_
timestamp 1667941163
transform 1 0 73472 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _071_
timestamp 1667941163
transform 1 0 76384 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _072_
timestamp 1667941163
transform 1 0 80080 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _073_
timestamp 1667941163
transform 1 0 84000 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _074_
timestamp 1667941163
transform 1 0 87920 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _075_
timestamp 1667941163
transform 1 0 91840 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _076_
timestamp 1667941163
transform 1 0 95760 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _077_
timestamp 1667941163
transform 1 0 96544 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _078_
timestamp 1667941163
transform 1 0 99680 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _079_
timestamp 1667941163
transform 1 0 102368 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _080_
timestamp 1667941163
transform 1 0 112448 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _081_
timestamp 1667941163
transform 1 0 116928 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _082_
timestamp 1667941163
transform 1 0 123200 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _083_
timestamp 1667941163
transform -1 0 128128 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _084_
timestamp 1667941163
transform -1 0 118608 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _085_
timestamp 1667941163
transform -1 0 112224 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _086_
timestamp 1667941163
transform 1 0 105056 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _087_
timestamp 1667941163
transform 1 0 108528 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _088_
timestamp 1667941163
transform 1 0 111440 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _089_
timestamp 1667941163
transform 1 0 115360 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _090_
timestamp 1667941163
transform 1 0 119280 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _091_
timestamp 1667941163
transform 1 0 120960 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _092_
timestamp 1667941163
transform 1 0 124432 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _093_
timestamp 1667941163
transform 1 0 127120 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _094_
timestamp 1667941163
transform 1 0 131040 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _095_
timestamp 1667941163
transform 1 0 132832 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _096_
timestamp 1667941163
transform 1 0 134960 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _097_
timestamp 1667941163
transform 1 0 138880 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _098_
timestamp 1667941163
transform 1 0 138880 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _099_
timestamp 1667941163
transform 1 0 144256 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _100_
timestamp 1667941163
transform -1 0 5152 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _101_
timestamp 1667941163
transform 1 0 1904 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _102_
timestamp 1667941163
transform 1 0 5712 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _103_
timestamp 1667941163
transform 1 0 6384 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _104_
timestamp 1667941163
transform 1 0 9856 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _105_
timestamp 1667941163
transform 1 0 12656 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _106_
timestamp 1667941163
transform 1 0 13664 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _107_
timestamp 1667941163
transform 1 0 17584 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _108_
timestamp 1667941163
transform 1 0 45024 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _109_
timestamp 1667941163
transform 1 0 48944 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _110_
timestamp 1667941163
transform 1 0 52864 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _111_
timestamp 1667941163
transform -1 0 71568 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _112_
timestamp 1667941163
transform 1 0 60704 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _113_
timestamp 1667941163
transform 1 0 64624 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _114_
timestamp 1667941163
transform 1 0 64624 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _115_
timestamp 1667941163
transform -1 0 29568 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _116_
timestamp 1667941163
transform 1 0 21840 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _117_
timestamp 1667941163
transform 1 0 22288 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_sclk pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 73248 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_sclk
timestamp 1667941163
transform -1 0 66864 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_sclk
timestamp 1667941163
transform 1 0 59248 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_sclk
timestamp 1667941163
transform -1 0 70896 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_sclk
timestamp 1667941163
transform -1 0 60816 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_sclk
timestamp 1667941163
transform 1 0 83104 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_sclk
timestamp 1667941163
transform 1 0 85120 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_sclk
timestamp 1667941163
transform -1 0 84672 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_sclk
timestamp 1667941163
transform 1 0 89152 0 -1 4704
box -86 -86 5686 870
<< labels >>
flabel metal3 s 0 8176 800 8288 0 FreeSans 448 0 0 0 latch
port 0 nsew signal input
flabel metal3 s 0 1680 800 1792 0 FreeSans 448 0 0 0 sclk
port 1 nsew signal input
flabel metal3 s 0 4928 800 5040 0 FreeSans 448 0 0 0 sdin
port 2 nsew signal input
flabel metal3 s 159200 4928 160000 5040 0 FreeSans 448 0 0 0 sr_out
port 3 nsew signal tristate
flabel metal2 s 23408 9200 23520 10000 0 FreeSans 448 90 0 0 tune_s1_series_gy[0]
port 4 nsew signal tristate
flabel metal2 s 26096 9200 26208 10000 0 FreeSans 448 90 0 0 tune_s1_series_gy[1]
port 5 nsew signal tristate
flabel metal2 s 28784 9200 28896 10000 0 FreeSans 448 90 0 0 tune_s1_series_gy[2]
port 6 nsew signal tristate
flabel metal2 s 31472 9200 31584 10000 0 FreeSans 448 90 0 0 tune_s1_series_gy[3]
port 7 nsew signal tristate
flabel metal2 s 34160 9200 34272 10000 0 FreeSans 448 90 0 0 tune_s1_series_gy[4]
port 8 nsew signal tristate
flabel metal2 s 36848 9200 36960 10000 0 FreeSans 448 90 0 0 tune_s1_series_gy[5]
port 9 nsew signal tristate
flabel metal2 s 39536 9200 39648 10000 0 FreeSans 448 90 0 0 tune_s1_series_gygy[0]
port 10 nsew signal tristate
flabel metal2 s 42224 9200 42336 10000 0 FreeSans 448 90 0 0 tune_s1_series_gygy[1]
port 11 nsew signal tristate
flabel metal2 s 44912 9200 45024 10000 0 FreeSans 448 90 0 0 tune_s1_series_gygy[2]
port 12 nsew signal tristate
flabel metal2 s 47600 9200 47712 10000 0 FreeSans 448 90 0 0 tune_s1_series_gygy[3]
port 13 nsew signal tristate
flabel metal2 s 50288 9200 50400 10000 0 FreeSans 448 90 0 0 tune_s1_series_gygy[4]
port 14 nsew signal tristate
flabel metal2 s 52976 9200 53088 10000 0 FreeSans 448 90 0 0 tune_s1_series_gygy[5]
port 15 nsew signal tristate
flabel metal2 s 1904 9200 2016 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[0]
port 16 nsew signal tristate
flabel metal2 s 4592 9200 4704 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[1]
port 17 nsew signal tristate
flabel metal2 s 7280 9200 7392 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[2]
port 18 nsew signal tristate
flabel metal2 s 9968 9200 10080 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[3]
port 19 nsew signal tristate
flabel metal2 s 12656 9200 12768 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[4]
port 20 nsew signal tristate
flabel metal2 s 15344 9200 15456 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[5]
port 21 nsew signal tristate
flabel metal2 s 18032 9200 18144 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[6]
port 22 nsew signal tristate
flabel metal2 s 20720 9200 20832 10000 0 FreeSans 448 90 0 0 tune_s1_shunt[7]
port 23 nsew signal tristate
flabel metal2 s 55664 9200 55776 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[0]
port 24 nsew signal tristate
flabel metal2 s 58352 9200 58464 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[1]
port 25 nsew signal tristate
flabel metal2 s 61040 9200 61152 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[2]
port 26 nsew signal tristate
flabel metal2 s 63728 9200 63840 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[3]
port 27 nsew signal tristate
flabel metal2 s 66416 9200 66528 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[4]
port 28 nsew signal tristate
flabel metal2 s 69104 9200 69216 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[5]
port 29 nsew signal tristate
flabel metal2 s 71792 9200 71904 10000 0 FreeSans 448 90 0 0 tune_s1_shunt_gy[6]
port 30 nsew signal tristate
flabel metal2 s 104048 9200 104160 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[0]
port 31 nsew signal tristate
flabel metal2 s 106736 9200 106848 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[1]
port 32 nsew signal tristate
flabel metal2 s 109424 9200 109536 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[2]
port 33 nsew signal tristate
flabel metal2 s 112112 9200 112224 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[3]
port 34 nsew signal tristate
flabel metal2 s 114800 9200 114912 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[4]
port 35 nsew signal tristate
flabel metal2 s 117488 9200 117600 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[5]
port 36 nsew signal tristate
flabel metal2 s 120176 9200 120288 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[6]
port 37 nsew signal tristate
flabel metal2 s 122864 9200 122976 10000 0 FreeSans 448 90 0 0 tune_s2_series_gy[7]
port 38 nsew signal tristate
flabel metal2 s 125552 9200 125664 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[0]
port 39 nsew signal tristate
flabel metal2 s 128240 9200 128352 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[1]
port 40 nsew signal tristate
flabel metal2 s 130928 9200 131040 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[2]
port 41 nsew signal tristate
flabel metal2 s 133616 9200 133728 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[3]
port 42 nsew signal tristate
flabel metal2 s 136304 9200 136416 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[4]
port 43 nsew signal tristate
flabel metal2 s 138992 9200 139104 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[5]
port 44 nsew signal tristate
flabel metal2 s 141680 9200 141792 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[6]
port 45 nsew signal tristate
flabel metal2 s 144368 9200 144480 10000 0 FreeSans 448 90 0 0 tune_s2_series_gygy[7]
port 46 nsew signal tristate
flabel metal2 s 74480 9200 74592 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[0]
port 47 nsew signal tristate
flabel metal2 s 101360 9200 101472 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[10]
port 48 nsew signal tristate
flabel metal2 s 77168 9200 77280 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[1]
port 49 nsew signal tristate
flabel metal2 s 79856 9200 79968 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[2]
port 50 nsew signal tristate
flabel metal2 s 82544 9200 82656 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[3]
port 51 nsew signal tristate
flabel metal2 s 85232 9200 85344 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[4]
port 52 nsew signal tristate
flabel metal2 s 87920 9200 88032 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[5]
port 53 nsew signal tristate
flabel metal2 s 90608 9200 90720 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[6]
port 54 nsew signal tristate
flabel metal2 s 93296 9200 93408 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[7]
port 55 nsew signal tristate
flabel metal2 s 95984 9200 96096 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[8]
port 56 nsew signal tristate
flabel metal2 s 98672 9200 98784 10000 0 FreeSans 448 90 0 0 tune_s2_shunt[9]
port 57 nsew signal tristate
flabel metal2 s 147056 9200 147168 10000 0 FreeSans 448 90 0 0 tune_s2_shunt_gy[0]
port 58 nsew signal tristate
flabel metal2 s 149744 9200 149856 10000 0 FreeSans 448 90 0 0 tune_s2_shunt_gy[1]
port 59 nsew signal tristate
flabel metal2 s 152432 9200 152544 10000 0 FreeSans 448 90 0 0 tune_s2_shunt_gy[2]
port 60 nsew signal tristate
flabel metal2 s 155120 9200 155232 10000 0 FreeSans 448 90 0 0 tune_s2_shunt_gy[3]
port 61 nsew signal tristate
flabel metal2 s 157808 9200 157920 10000 0 FreeSans 448 90 0 0 tune_s2_shunt_gy[4]
port 62 nsew signal tristate
flabel metal4 s 20500 3076 21500 6332 0 FreeSans 5120 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 59812 3076 60812 6332 0 FreeSans 5120 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 99124 3076 100124 6332 0 FreeSans 5120 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 138436 3076 139436 6332 0 FreeSans 5120 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 40156 3076 41156 6332 0 FreeSans 5120 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 79468 3076 80468 6332 0 FreeSans 5120 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 118780 3076 119780 6332 0 FreeSans 5120 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 158092 3076 159092 6332 0 FreeSans 5120 90 0 0 vss
port 64 nsew ground bidirectional
rlabel metal1 79968 5488 79968 5488 0 vdd
rlabel metal1 80218 6272 80218 6272 0 vss
rlabel metal2 78456 4256 78456 4256 0 clknet_0_sclk
rlabel metal3 5880 4312 5880 4312 0 clknet_3_0__leaf_sclk
rlabel metal2 53928 3920 53928 3920 0 clknet_3_1__leaf_sclk
rlabel metal2 2184 5824 2184 5824 0 clknet_3_2__leaf_sclk
rlabel metal2 21672 5488 21672 5488 0 clknet_3_3__leaf_sclk
rlabel metal2 92120 3640 92120 3640 0 clknet_3_4__leaf_sclk
rlabel metal3 97888 3528 97888 3528 0 clknet_3_5__leaf_sclk
rlabel metal2 76664 5544 76664 5544 0 clknet_3_6__leaf_sclk
rlabel metal2 94024 3920 94024 3920 0 clknet_3_7__leaf_sclk
rlabel metal2 2072 6664 2072 6664 0 latch
rlabel metal2 73976 3024 73976 3024 0 sclk
rlabel metal3 854 4984 854 4984 0 sdin
rlabel metal2 4200 3920 4200 3920 0 sr\[0\]
rlabel metal3 53256 3640 53256 3640 0 sr\[10\]
rlabel metal2 70616 4088 70616 4088 0 sr\[11\]
rlabel metal2 59808 5768 59808 5768 0 sr\[12\]
rlabel metal3 61432 3640 61432 3640 0 sr\[13\]
rlabel metal2 52472 4144 52472 4144 0 sr\[14\]
rlabel metal2 31640 3920 31640 3920 0 sr\[15\]
rlabel metal2 22792 3920 22792 3920 0 sr\[16\]
rlabel metal2 24584 5712 24584 5712 0 sr\[17\]
rlabel metal3 27608 5096 27608 5096 0 sr\[18\]
rlabel metal2 30296 5096 30296 5096 0 sr\[19\]
rlabel metal2 2856 5488 2856 5488 0 sr\[1\]
rlabel metal2 34216 5712 34216 5712 0 sr\[20\]
rlabel metal2 37800 4760 37800 4760 0 sr\[21\]
rlabel metal3 38640 5208 38640 5208 0 sr\[22\]
rlabel metal2 42056 5488 42056 5488 0 sr\[23\]
rlabel metal2 44184 5432 44184 5432 0 sr\[24\]
rlabel metal2 46648 4704 46648 4704 0 sr\[25\]
rlabel metal2 49224 5264 49224 5264 0 sr\[26\]
rlabel metal2 70168 5488 70168 5488 0 sr\[27\]
rlabel metal2 73416 5488 73416 5488 0 sr\[28\]
rlabel metal2 77336 4704 77336 4704 0 sr\[29\]
rlabel metal3 5992 4424 5992 4424 0 sr\[2\]
rlabel metal2 81032 4704 81032 4704 0 sr\[30\]
rlabel metal2 84952 4704 84952 4704 0 sr\[31\]
rlabel metal2 88872 3696 88872 3696 0 sr\[32\]
rlabel metal2 92792 3752 92792 3752 0 sr\[33\]
rlabel metal3 95816 3640 95816 3640 0 sr\[34\]
rlabel metal2 97496 4312 97496 4312 0 sr\[35\]
rlabel metal2 99400 4144 99400 4144 0 sr\[36\]
rlabel metal2 101976 5488 101976 5488 0 sr\[37\]
rlabel metal2 121352 5320 121352 5320 0 sr\[38\]
rlabel metal2 115528 5264 115528 5264 0 sr\[39\]
rlabel metal2 8120 5432 8120 5432 0 sr\[3\]
rlabel metal2 124152 4760 124152 4760 0 sr\[40\]
rlabel metal2 127176 5432 127176 5432 0 sr\[41\]
rlabel metal2 125048 5040 125048 5040 0 sr\[42\]
rlabel metal2 115472 3640 115472 3640 0 sr\[43\]
rlabel metal3 105392 4424 105392 4424 0 sr\[44\]
rlabel metal2 108136 4312 108136 4312 0 sr\[45\]
rlabel metal2 112392 4480 112392 4480 0 sr\[46\]
rlabel metal2 115304 4816 115304 4816 0 sr\[47\]
rlabel metal2 118440 5824 118440 5824 0 sr\[48\]
rlabel metal2 121912 5096 121912 5096 0 sr\[49\]
rlabel metal2 5992 5880 5992 5880 0 sr\[4\]
rlabel metal3 124712 4200 124712 4200 0 sr\[50\]
rlabel metal3 129080 4200 129080 4200 0 sr\[51\]
rlabel metal3 131600 4424 131600 4424 0 sr\[52\]
rlabel metal3 134232 5096 134232 5096 0 sr\[53\]
rlabel metal2 135912 3864 135912 3864 0 sr\[54\]
rlabel metal2 139832 5544 139832 5544 0 sr\[55\]
rlabel metal2 142632 3920 142632 3920 0 sr\[56\]
rlabel metal3 143584 5096 143584 5096 0 sr\[57\]
rlabel metal2 13608 5096 13608 5096 0 sr\[5\]
rlabel metal2 16856 5096 16856 5096 0 sr\[6\]
rlabel metal2 20888 4984 20888 4984 0 sr\[7\]
rlabel metal2 45976 4704 45976 4704 0 sr\[8\]
rlabel metal3 49000 5768 49000 5768 0 sr\[9\]
rlabel metal2 147336 4816 147336 4816 0 sr_out
rlabel metal2 26488 4256 26488 4256 0 tune_s1_series_gy[0]
rlabel metal3 25536 4200 25536 4200 0 tune_s1_series_gy[1]
rlabel metal2 25368 5040 25368 5040 0 tune_s1_series_gy[2]
rlabel metal2 28840 5096 28840 5096 0 tune_s1_series_gy[3]
rlabel metal3 33488 4200 33488 4200 0 tune_s1_series_gy[4]
rlabel metal2 36848 5208 36848 5208 0 tune_s1_series_gy[5]
rlabel metal3 39816 3640 39816 3640 0 tune_s1_series_gygy[0]
rlabel metal2 40264 5376 40264 5376 0 tune_s1_series_gygy[1]
rlabel metal2 44744 6216 44744 6216 0 tune_s1_series_gygy[2]
rlabel metal3 45920 3640 45920 3640 0 tune_s1_series_gygy[3]
rlabel metal2 48776 4312 48776 4312 0 tune_s1_series_gygy[4]
rlabel metal2 52024 3696 52024 3696 0 tune_s1_series_gygy[5]
rlabel metal2 2016 3640 2016 3640 0 tune_s1_shunt[0]
rlabel metal2 4928 5208 4928 5208 0 tune_s1_shunt[1]
rlabel metal2 7448 4480 7448 4480 0 tune_s1_shunt[2]
rlabel metal2 9464 6216 9464 6216 0 tune_s1_shunt[3]
rlabel metal2 12936 6104 12936 6104 0 tune_s1_shunt[4]
rlabel metal2 15568 4200 15568 4200 0 tune_s1_shunt[5]
rlabel metal3 17416 5768 17416 5768 0 tune_s1_shunt[6]
rlabel metal2 20720 5768 20720 5768 0 tune_s1_shunt[7]
rlabel metal2 48104 3808 48104 3808 0 tune_s1_shunt_gy[0]
rlabel metal2 52024 5376 52024 5376 0 tune_s1_shunt_gy[1]
rlabel metal2 55944 3920 55944 3920 0 tune_s1_shunt_gy[2]
rlabel metal2 68488 4256 68488 4256 0 tune_s1_shunt_gy[3]
rlabel metal2 63784 5376 63784 5376 0 tune_s1_shunt_gy[4]
rlabel metal3 68432 3640 68432 3640 0 tune_s1_shunt_gy[5]
rlabel metal2 67704 5376 67704 5376 0 tune_s1_shunt_gy[6]
rlabel metal3 105896 5768 105896 5768 0 tune_s2_series_gy[0]
rlabel metal2 106848 5768 106848 5768 0 tune_s2_series_gy[1]
rlabel metal2 110600 4144 110600 4144 0 tune_s2_series_gy[2]
rlabel metal2 111608 6216 111608 6216 0 tune_s2_series_gy[3]
rlabel metal2 114856 6706 114856 6706 0 tune_s2_series_gy[4]
rlabel metal3 117096 4200 117096 4200 0 tune_s2_series_gy[5]
rlabel metal3 119784 3640 119784 3640 0 tune_s2_series_gy[6]
rlabel metal3 123144 3640 123144 3640 0 tune_s2_series_gy[7]
rlabel metal2 125608 7098 125608 7098 0 tune_s2_series_gygy[0]
rlabel metal2 129080 4312 129080 4312 0 tune_s2_series_gygy[1]
rlabel metal3 131768 4200 131768 4200 0 tune_s2_series_gygy[2]
rlabel metal3 135352 4200 135352 4200 0 tune_s2_series_gygy[3]
rlabel metal2 140952 5096 140952 5096 0 tune_s2_series_gygy[4]
rlabel metal3 140000 4200 140000 4200 0 tune_s2_series_gygy[5]
rlabel metal3 142352 5768 142352 5768 0 tune_s2_series_gygy[6]
rlabel metal3 145152 3640 145152 3640 0 tune_s2_series_gygy[7]
rlabel metal2 72296 5096 72296 5096 0 tune_s2_shunt[0]
rlabel metal3 100632 5768 100632 5768 0 tune_s2_shunt[10]
rlabel metal3 76384 5768 76384 5768 0 tune_s2_shunt[1]
rlabel metal2 79408 3640 79408 3640 0 tune_s2_shunt[2]
rlabel metal3 82880 3640 82880 3640 0 tune_s2_shunt[3]
rlabel metal3 86184 5768 86184 5768 0 tune_s2_shunt[4]
rlabel metal2 88032 5768 88032 5768 0 tune_s2_shunt[5]
rlabel metal2 90664 7490 90664 7490 0 tune_s2_shunt[6]
rlabel metal2 93296 5208 93296 5208 0 tune_s2_shunt[7]
rlabel metal2 95984 5768 95984 5768 0 tune_s2_shunt[8]
rlabel metal2 97272 4256 97272 4256 0 tune_s2_shunt[9]
rlabel metal2 123480 4872 123480 4872 0 tune_s2_shunt_gy[0]
rlabel metal2 130200 5264 130200 5264 0 tune_s2_shunt_gy[1]
rlabel metal2 134120 3696 134120 3696 0 tune_s2_shunt_gy[2]
rlabel metal2 138096 5768 138096 5768 0 tune_s2_shunt_gy[3]
rlabel metal2 139384 5040 139384 5040 0 tune_s2_shunt_gy[4]
<< properties >>
string FIXED_BBOX 0 0 160000 10000
<< end >>
