** sch_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/chebyshev_test_l1_pex_1.sch
**.subckt chebyshev_test_l1_pex_1
C1 vip GND 41.67p m=1
C2 vin GND 41.67p m=1
C3 net12 GND 10.32p m=1
C4 net2 GND 10.32p m=1
C5 net1 GND 1p m=1
C6 net13 GND 1p m=1
C7 net3 GND 3.8p m=1
C8 net14 GND 3.8p m=1
V1 vdd GND 1.8
C10 net4 GND 30p m=1
C12 net7 GND 12.16p m=1
C13 net5 GND 0.8p m=1
C14 net15 GND 0.8p m=1
C15 net8 GND 2p m=1
C16 net16 GND 2p m=1
C9 net6 GND 30p m=1
C11 net17 GND 12.16p m=1
x6 vdd GND vip vin net1 net13 net6 net4 net12 net2 net14 net3 filterstage_pex
x1 vdd GND net6 net4 net5 net15 net11 net10 net17 net7 net16 net8 filterstage_pex
V2 net9 GND PULSE(0 1.8 0 1n 1n {tau/2} {tau})
x2 vip vdd GND vin vdd net9 GND GND GND GND GND GND GND GND injector_pex
x3 vdd GND vop_buf net10 net11 von_buf vop voxor von active_load_pex
**** begin user architecture code


* .ac dec 1000 1e6 1e9
.param tau=100n
.tran 5ns {10*tau}
.save all
.control
run
display
* let vod = vop-von
* plot vdb(vod)
plot vop von
plot vop_buf von_buf voxor
.endc



.include /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends

* expanding   symbol:  filterstage_pex.sym # of pins=12
** sym_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/filterstage_pex.sym
** sch_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/filterstage_pex.sch
.subckt filterstage_pex vdd vss nbusin_nshunt pbusin_pshunt nshunt_gy pshunt_gy nbusout pbusout
+ pseries_gy nseries_gy pseries_gygy nseries_gygy
*.iopin vdd
*.iopin vss
*.iopin nbusin_nshunt
*.iopin pbusin_pshunt
*.iopin nbusout
*.iopin pbusout
*.iopin pseries_gy
*.iopin nseries_gy
*.iopin pseries_gygy
*.iopin nseries_gygy
*.iopin nshunt_gy
*.iopin pshunt_gy
**** begin user architecture code

.subckt filterstage_flat nbusin_nshunt nbusout nseries_gy nseries_gygy nshunt_gy pbusin_pshunt
+  pbusout pseries_gy pseries_gygy pshunt_gy vss vdd
X0 a_3932_14487# a_3844_14584# vss vss nfet_06v0 w=0.82u l=1u
X1 pbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X2 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X3 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X4 a_3932_11351# a_3844_11448# vss vss nfet_06v0 w=0.82u l=1u
X5 vss nbusin_nshunt pbusin_pshunt vss nfet_06v0 w=0.82u l=0.6u
X6 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X7 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X8 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X9 nshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X10 vdd a_8412_13352# a_8324_13396# vdd pfet_06v0 w=1.22u l=1u
X11 a_13564_14487# a_13476_14584# vss vss nfet_06v0 w=0.82u l=1u
X12 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X13 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X14 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X15 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X16 vdd a_17372_16055# a_17284_16152# vdd pfet_06v0 w=1.22u l=1u
X17 a_10988_14920# a_10900_14964# vss vss nfet_06v0 w=0.82u l=1u
X18 vdd a_1692_14487# a_1604_14584# vdd pfet_06v0 w=1.22u l=1u
X19 vdd a_1692_11351# a_1604_11448# vdd pfet_06v0 w=1.22u l=1u
X20 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X21 vdd a_14348_16055# a_14260_16152# vdd pfet_06v0 w=1.22u l=1u
X22 vdd a_16812_14920# a_16724_14964# vdd pfet_06v0 w=1.22u l=1u
X23 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X24 vss pbusin_pshunt nshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X25 a_21292_3511# a_21204_3608# vss vss nfet_06v0 w=0.82u l=1u
X26 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X27 pshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X28 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X29 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X30 a_10876_16055# a_10788_16152# vss vss nfet_06v0 w=0.82u l=1u
X31 vss pshunt_gy pshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X32 pseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X33 vss nseries_gy nbusin_nshunt vss nfet_06v0 w=0.82u l=0.6u
X34 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X35 vdd a_20844_11784# a_20756_11828# vdd pfet_06v0 w=1.22u l=1u
X36 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X37 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X38 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X39 vdd a_21516_14487# a_21428_14584# vdd pfet_06v0 w=1.22u l=1u
X40 vdd a_8860_13352# a_8772_13396# vdd pfet_06v0 w=1.22u l=1u
X41 vdd a_21516_11351# a_21428_11448# vdd pfet_06v0 w=1.22u l=1u
X42 vdd pshunt_gy nshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X43 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X44 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X45 vdd a_12220_16055# a_12132_16152# vdd pfet_06v0 w=1.22u l=1u
X46 a_18268_16055# a_18180_16152# vss vss nfet_06v0 w=0.82u l=1u
X47 a_6620_14920# a_6532_14964# vss vss nfet_06v0 w=0.82u l=1u
X48 a_10988_14487# a_10900_14584# vss vss nfet_06v0 w=0.82u l=1u
X49 a_10988_11351# a_10900_11448# vss vss nfet_06v0 w=0.82u l=1u
X50 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X51 vdd a_11660_8215# a_11572_8312# vdd pfet_06v0 w=1.22u l=1u
X52 a_8748_14487# a_8660_14584# vss vss nfet_06v0 w=0.82u l=1u
X53 vdd a_14796_16055# a_14708_16152# vdd pfet_06v0 w=1.22u l=1u
X54 vdd a_17932_14487# a_17844_14584# vdd pfet_06v0 w=1.22u l=1u
X55 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X56 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X57 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X58 vdd a_14908_14487# a_14820_14584# vdd pfet_06v0 w=1.22u l=1u
X59 vdd a_15468_13352# a_15380_13396# vdd pfet_06v0 w=1.22u l=1u
X60 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X61 nseries_gygy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X62 vdd a_1692_13352# a_1604_13396# vdd pfet_06v0 w=1.22u l=1u
X63 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X64 a_13228_14920# a_13140_14964# vss vss nfet_06v0 w=0.82u l=1u
X65 a_10540_11784# a_10452_11828# vss vss nfet_06v0 w=0.82u l=1u
X66 a_21740_11784# a_21652_11828# vss vss nfet_06v0 w=0.82u l=1u
X67 a_16812_3944# a_16724_3988# vss vss nfet_06v0 w=0.82u l=1u
X68 vdd a_11548_3944# a_11460_3988# vdd pfet_06v0 w=1.22u l=1u
X69 vdd a_10876_5079# a_10788_5176# vdd pfet_06v0 w=1.22u l=1u
X70 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X71 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X72 a_16140_16055# a_16052_16152# vss vss nfet_06v0 w=0.82u l=1u
X73 vdd a_21964_14487# a_21876_14584# vdd pfet_06v0 w=1.22u l=1u
X74 nbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X75 vdd a_21964_11351# a_21876_11448# vdd pfet_06v0 w=1.22u l=1u
X76 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X77 vdd a_4828_14920# a_4740_14964# vdd pfet_06v0 w=1.22u l=1u
X78 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X79 pbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X80 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X81 a_9644_8648# a_9556_8692# vss vss nfet_06v0 w=0.82u l=1u
X82 a_20284_14920# a_20196_14964# vss vss nfet_06v0 w=0.82u l=1u
X83 vdd a_20844_12919# a_20756_13016# vdd pfet_06v0 w=1.22u l=1u
X84 vdd a_4828_11784# a_4740_11828# vdd pfet_06v0 w=1.22u l=1u
X85 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X86 vdd a_21516_13352# a_21428_13396# vdd pfet_06v0 w=1.22u l=1u
X87 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X88 vdd a_7404_16055# a_7316_16152# vdd pfet_06v0 w=1.22u l=1u
X89 vdd a_7404_12919# a_7316_13016# vdd pfet_06v0 w=1.22u l=1u
X90 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X91 a_16252_14487# a_16164_14584# vss vss nfet_06v0 w=0.82u l=1u
X92 pseries_gygy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X93 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X94 a_3932_16055# a_3844_16152# vss vss nfet_06v0 w=0.82u l=1u
X95 a_13676_14920# a_13588_14964# vss vss nfet_06v0 w=0.82u l=1u
X96 vdd a_4380_14487# a_4292_14584# vdd pfet_06v0 w=1.22u l=1u
X97 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X98 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X99 vdd a_4380_11351# a_4292_11448# vdd pfet_06v0 w=1.22u l=1u
X100 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X101 a_5724_11784# a_5636_11828# vss vss nfet_06v0 w=0.82u l=1u
X102 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X103 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X104 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X105 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X106 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X107 vdd nseries_gy pbusout vdd pfet_06v0 w=1.22u l=0.5u
X108 vdd a_21964_13352# a_21876_13396# vdd pfet_06v0 w=1.22u l=1u
X109 a_5612_12919# a_5524_13016# vss vss nfet_06v0 w=0.82u l=1u
X110 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X111 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X112 vdd a_4828_16055# a_4740_16152# vdd pfet_06v0 w=1.22u l=1u
X113 vdd a_7852_16055# a_7764_16152# vdd pfet_06v0 w=1.22u l=1u
X114 vdd a_12332_14920# a_12244_14964# vdd pfet_06v0 w=1.22u l=1u
X115 vdd a_7852_12919# a_7764_13016# vdd pfet_06v0 w=1.22u l=1u
X116 vdd a_12332_11784# a_12244_11828# vdd pfet_06v0 w=1.22u l=1u
X117 vdd a_4828_12919# a_4740_13016# vdd pfet_06v0 w=1.22u l=1u
X118 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X119 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X120 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X121 a_7068_13352# a_6980_13396# vss vss nfet_06v0 w=0.82u l=1u
X122 vdd a_4380_13352# a_4292_13396# vdd pfet_06v0 w=1.22u l=1u
X123 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X124 a_8748_16055# a_8660_16152# vss vss nfet_06v0 w=0.82u l=1u
X125 a_2140_14920# a_2052_14964# vss vss nfet_06v0 w=0.82u l=1u
X126 vss nseries_gygy pseries_gygy vss nfet_06v0 w=0.82u l=0.6u
X127 vdd a_9196_14487# a_9108_14584# vdd pfet_06v0 w=1.22u l=1u
X128 vdd a_12780_14920# a_12692_14964# vdd pfet_06v0 w=1.22u l=1u
X129 vdd a_12780_11784# a_12692_11828# vdd pfet_06v0 w=1.22u l=1u
X130 vss nseries_gy nbusin_nshunt vss nfet_06v0 w=0.82u l=0.6u
X131 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X132 vdd a_20508_16055# a_20420_16152# vdd pfet_06v0 w=1.22u l=1u
X133 vdd a_7516_14920# a_7428_14964# vdd pfet_06v0 w=1.22u l=1u
X134 vdd a_7516_11784# a_7428_11828# vdd pfet_06v0 w=1.22u l=1u
X135 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X136 vdd a_12332_12919# a_12244_13016# vdd pfet_06v0 w=1.22u l=1u
X137 vdd a_3036_10216# a_2948_10260# vdd pfet_06v0 w=1.22u l=1u
X138 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X139 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X140 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X141 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X142 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X143 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X144 a_16364_14920# a_16276_14964# vss vss nfet_06v0 w=0.82u l=1u
X145 a_2140_14487# a_2052_14584# vss vss nfet_06v0 w=0.82u l=1u
X146 a_2140_11351# a_2052_11448# vss vss nfet_06v0 w=0.82u l=1u
X147 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X148 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X149 a_13564_5079# a_13476_5176# vss vss nfet_06v0 w=0.82u l=1u
X150 a_8412_11784# a_8324_11828# vss vss nfet_06v0 w=0.82u l=1u
X151 a_10540_12919# a_10452_13016# vss vss nfet_06v0 w=0.82u l=1u
X152 vdd a_7964_14920# a_7876_14964# vdd pfet_06v0 w=1.22u l=1u
X153 vdd a_7964_11784# a_7876_11828# vdd pfet_06v0 w=1.22u l=1u
X154 vdd a_12780_12919# a_12692_13016# vdd pfet_06v0 w=1.22u l=1u
X155 a_8300_12919# a_8212_13016# vss vss nfet_06v0 w=0.82u l=1u
X156 vdd a_8636_11351# a_8548_11448# vdd pfet_06v0 w=1.22u l=1u
X157 vdd a_3484_10216# a_3396_10260# vdd pfet_06v0 w=1.22u l=1u
X158 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X159 vdd a_15020_14920# a_14932_14964# vdd pfet_06v0 w=1.22u l=1u
X160 vdd a_17596_14920# a_17508_14964# vdd pfet_06v0 w=1.22u l=1u
X161 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X162 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X163 a_8860_11784# a_8772_11828# vss vss nfet_06v0 w=0.82u l=1u
X164 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X165 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X166 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X167 vdd a_22076_9783# a_21988_9880# vdd pfet_06v0 w=1.22u l=1u
X168 vdd a_22076_6647# a_21988_6744# vdd pfet_06v0 w=1.22u l=1u
X169 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X170 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X171 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X172 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X173 a_1692_11784# a_1604_11828# vss vss nfet_06v0 w=0.82u l=1u
X174 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X175 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X176 vdd pshunt_gy nshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X177 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X178 a_16812_8648# a_16724_8692# vss vss nfet_06v0 w=0.82u l=1u
X179 a_15804_14487# a_15716_14584# vss vss nfet_06v0 w=0.82u l=1u
X180 nbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X181 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X182 vdd a_20172_14487# a_20084_14584# vdd pfet_06v0 w=1.22u l=1u
X183 a_11436_13352# a_11348_13396# vss vss nfet_06v0 w=0.82u l=1u
X184 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X185 vdd a_19612_16055# a_19524_16152# vdd pfet_06v0 w=1.22u l=1u
X186 vdd a_3036_14920# a_2948_14964# vdd pfet_06v0 w=1.22u l=1u
X187 vdd a_3932_14487# a_3844_14584# vdd pfet_06v0 w=1.22u l=1u
X188 vdd a_3932_11351# a_3844_11448# vdd pfet_06v0 w=1.22u l=1u
X189 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X190 a_19948_12919# a_19860_13016# vss vss nfet_06v0 w=0.82u l=1u
X191 vdd a_3036_11784# a_2948_11828# vdd pfet_06v0 w=1.22u l=1u
X192 vdd nbusin_nshunt pbusin_pshunt vdd pfet_06v0 w=1.22u l=0.5u
X193 pbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X194 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X195 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X196 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X197 vdd a_13564_14487# a_13476_14584# vdd pfet_06v0 w=1.22u l=1u
X198 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X199 pbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X200 a_2140_16055# a_2052_16152# vss vss nfet_06v0 w=0.82u l=1u
X201 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X202 a_1692_6647# a_1604_6744# vss vss nfet_06v0 w=0.82u l=1u
X203 pbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X204 pseries_gygy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X205 vdd pbusin_pshunt nshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X206 a_1692_3511# a_1604_3608# vss vss nfet_06v0 w=0.82u l=1u
X207 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X208 vdd a_21292_3511# a_21204_3608# vdd pfet_06v0 w=1.22u l=1u
X209 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X210 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X211 vdd pshunt_gy pshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X212 a_11884_13352# a_11796_13396# vss vss nfet_06v0 w=0.82u l=1u
X213 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X214 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X215 vdd a_3484_14920# a_3396_14964# vdd pfet_06v0 w=1.22u l=1u
X216 a_9644_13352# a_9556_13396# vss vss nfet_06v0 w=0.82u l=1u
X217 vdd a_3484_11784# a_3396_11828# vdd pfet_06v0 w=1.22u l=1u
X218 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X219 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X220 vdd a_20172_13352# a_20084_13396# vdd pfet_06v0 w=1.22u l=1u
X221 vdd a_3036_16055# a_2948_16152# vdd pfet_06v0 w=1.22u l=1u
X222 vdd a_6060_16055# a_5972_16152# vdd pfet_06v0 w=1.22u l=1u
X223 vdd a_3932_13352# a_3844_13396# vdd pfet_06v0 w=1.22u l=1u
X224 vdd a_6060_12919# a_5972_13016# vdd pfet_06v0 w=1.22u l=1u
X225 nshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X226 vdd a_3036_12919# a_2948_13016# vdd pfet_06v0 w=1.22u l=1u
X227 vdd a_10988_14487# a_10900_14584# vdd pfet_06v0 w=1.22u l=1u
X228 a_19276_13352# a_19188_13396# vss vss nfet_06v0 w=0.82u l=1u
X229 vdd a_10988_11351# a_10900_11448# vdd pfet_06v0 w=1.22u l=1u
X230 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X231 vdd a_8748_14487# a_8660_14584# vdd pfet_06v0 w=1.22u l=1u
X232 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X233 a_7068_14920# a_6980_14964# vss vss nfet_06v0 w=0.82u l=1u
X234 a_4380_11784# a_4292_11828# vss vss nfet_06v0 w=0.82u l=1u
X235 vdd a_20844_8215# a_20756_8312# vdd pfet_06v0 w=1.22u l=1u
X236 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X237 vdd nbusout nseries_gy vdd pfet_06v0 w=1.22u l=0.5u
X238 vdd a_21292_8648# a_21204_8692# vdd pfet_06v0 w=1.22u l=1u
X239 nshunt_gy pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X240 pbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X241 vdd a_3484_16055# a_3396_16152# vdd pfet_06v0 w=1.22u l=1u
X242 a_18940_14920# a_18852_14964# vss vss nfet_06v0 w=0.82u l=1u
X243 a_14124_13352# a_14036_13396# vss vss nfet_06v0 w=0.82u l=1u
X244 nseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X245 nseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X246 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X247 a_15916_14920# a_15828_14964# vss vss nfet_06v0 w=0.82u l=1u
X248 vdd a_3484_12919# a_3396_13016# vdd pfet_06v0 w=1.22u l=1u
X249 pseries_gygy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X250 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X251 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X252 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X253 vdd a_10988_13352# a_10900_13396# vdd pfet_06v0 w=1.22u l=1u
X254 vdd a_16252_14487# a_16164_14584# vdd pfet_06v0 w=1.22u l=1u
X255 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X256 vdd a_21516_8215# a_21428_8312# vdd pfet_06v0 w=1.22u l=1u
X257 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X258 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X259 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X260 a_1692_12919# a_1604_13016# vss vss nfet_06v0 w=0.82u l=1u
X261 a_14572_13352# a_14484_13396# vss vss nfet_06v0 w=0.82u l=1u
X262 pbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X263 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X264 a_1692_8215# a_1604_8312# vss vss nfet_06v0 w=0.82u l=1u
X265 vdd a_6172_14920# a_6084_14964# vdd pfet_06v0 w=1.22u l=1u
X266 vdd a_6172_11784# a_6084_11828# vdd pfet_06v0 w=1.22u l=1u
X267 vdd a_8860_3944# a_8772_3988# vdd pfet_06v0 w=1.22u l=1u
X268 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X269 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X270 vdd a_6620_13352# a_6532_13396# vdd pfet_06v0 w=1.22u l=1u
X271 a_21516_12919# a_21428_13016# vss vss nfet_06v0 w=0.82u l=1u
X272 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X273 a_6508_14487# a_6420_14584# vss vss nfet_06v0 w=0.82u l=1u
X274 vdd a_2588_9783# a_2500_9880# vdd pfet_06v0 w=1.22u l=1u
X275 a_20620_13352# a_20532_13396# vss vss nfet_06v0 w=0.82u l=1u
X276 vdd a_13228_13352# a_13140_13396# vdd pfet_06v0 w=1.22u l=1u
X277 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X278 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X279 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X280 vdd a_21516_7080# a_21428_7124# vdd pfet_06v0 w=1.22u l=1u
X281 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X282 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X283 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X284 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X285 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X286 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X287 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X288 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X289 a_21964_12919# a_21876_13016# vss vss nfet_06v0 w=0.82u l=1u
X290 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X291 a_6956_14487# a_6868_14584# vss vss nfet_06v0 w=0.82u l=1u
X292 vss nseries_gygy nseries_gygy vss nfet_06v0 w=0.82u l=0.6u
X293 a_2588_13352# a_2500_13396# vss vss nfet_06v0 w=0.82u l=1u
X294 vdd a_13676_13352# a_13588_13396# vdd pfet_06v0 w=1.22u l=1u
X295 a_14012_14487# a_13924_14584# vss vss nfet_06v0 w=0.82u l=1u
X296 a_2588_10216# a_2500_10260# vss vss nfet_06v0 w=0.82u l=1u
X297 vdd a_2588_8648# a_2500_8692# vdd pfet_06v0 w=1.22u l=1u
X298 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X299 vdd a_21964_8215# a_21876_8312# vdd pfet_06v0 w=1.22u l=1u
X300 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X301 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X302 pshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X303 nshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X304 a_11436_14920# a_11348_14964# vss vss nfet_06v0 w=0.82u l=1u
X305 vdd a_2140_14487# a_2052_14584# vdd pfet_06v0 w=1.22u l=1u
X306 vdd a_2140_11351# a_2052_11448# vdd pfet_06v0 w=1.22u l=1u
X307 a_20844_8648# a_20756_8692# vss vss nfet_06v0 w=0.82u l=1u
X308 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X309 pbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X310 a_4380_12919# a_4292_13016# vss vss nfet_06v0 w=0.82u l=1u
X311 a_11324_16055# a_11236_16152# vss vss nfet_06v0 w=0.82u l=1u
X312 vdd a_19836_14920# a_19748_14964# vdd pfet_06v0 w=1.22u l=1u
X313 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X314 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X315 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X316 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X317 nbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X318 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X319 vdd a_5612_16055# a_5524_16152# vdd pfet_06v0 w=1.22u l=1u
X320 vdd a_5612_12919# a_5524_13016# vdd pfet_06v0 w=1.22u l=1u
X321 a_14460_14487# a_14372_14584# vss vss nfet_06v0 w=0.82u l=1u
X322 a_18828_13352# a_18740_13396# vss vss nfet_06v0 w=0.82u l=1u
X323 a_11436_14487# a_11348_14584# vss vss nfet_06v0 w=0.82u l=1u
X324 a_10092_13352# a_10004_13396# vss vss nfet_06v0 w=0.82u l=1u
X325 a_11436_11351# a_11348_11448# vss vss nfet_06v0 w=0.82u l=1u
X326 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X327 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X328 a_11884_14920# a_11796_14964# vss vss nfet_06v0 w=0.82u l=1u
X329 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X330 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X331 vdd a_15244_16055# a_15156_16152# vdd pfet_06v0 w=1.22u l=1u
X332 a_9644_14920# a_9556_14964# vss vss nfet_06v0 w=0.82u l=1u
X333 nbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X334 nshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X335 vdd a_21964_7080# a_21876_7124# vdd pfet_06v0 w=1.22u l=1u
X336 a_3932_11784# a_3844_11828# vss vss nfet_06v0 w=0.82u l=1u
X337 nseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X338 a_11772_16055# a_11684_16152# vss vss nfet_06v0 w=0.82u l=1u
X339 vdd a_2140_13352# a_2052_13396# vdd pfet_06v0 w=1.22u l=1u
X340 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X341 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X342 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X343 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X344 a_6508_16055# a_6420_16152# vss vss nfet_06v0 w=0.82u l=1u
X345 a_9532_16055# a_9444_16152# vss vss nfet_06v0 w=0.82u l=1u
X346 vdd a_10540_14920# a_10452_14964# vdd pfet_06v0 w=1.22u l=1u
X347 vdd a_21740_11784# a_21652_11828# vdd pfet_06v0 w=1.22u l=1u
X348 vdd a_16812_3944# a_16724_3988# vdd pfet_06v0 w=1.22u l=1u
X349 vdd a_10540_11784# a_10452_11828# vdd pfet_06v0 w=1.22u l=1u
X350 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X351 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X352 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X353 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X354 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X355 a_19164_16055# a_19076_16152# vss vss nfet_06v0 w=0.82u l=1u
X356 a_11884_14487# a_11796_14584# vss vss nfet_06v0 w=0.82u l=1u
X357 a_9196_12919# a_9108_13016# vss vss nfet_06v0 w=0.82u l=1u
X358 a_2140_3511# a_2052_3608# vss vss nfet_06v0 w=0.82u l=1u
X359 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X360 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X361 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X362 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X363 a_9644_14487# a_9556_14584# vss vss nfet_06v0 w=0.82u l=1u
X364 vdd a_12668_16055# a_12580_16152# vdd pfet_06v0 w=1.22u l=1u
X365 vdd a_15692_16055# a_15604_16152# vdd pfet_06v0 w=1.22u l=1u
X366 a_5276_13352# a_5188_13396# vss vss nfet_06v0 w=0.82u l=1u
X367 vdd a_15804_14487# a_15716_14584# vdd pfet_06v0 w=1.22u l=1u
X368 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X369 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X370 vss nseries_gy pseries_gygy vss nfet_06v0 w=0.82u l=0.6u
X371 pbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X372 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X373 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X374 a_14124_14920# a_14036_14964# vss vss nfet_06v0 w=0.82u l=1u
X375 a_19276_14487# a_19188_14584# vss vss nfet_06v0 w=0.82u l=1u
X376 a_6956_16055# a_6868_16152# vss vss nfet_06v0 w=0.82u l=1u
X377 a_9980_16055# a_9892_16152# vss vss nfet_06v0 w=0.82u l=1u
X378 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X379 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X380 vdd a_13564_5079# a_13476_5176# vdd pfet_06v0 w=1.22u l=1u
X381 a_10988_11784# a_10900_11828# vss vss nfet_06v0 w=0.82u l=1u
X382 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X383 vdd a_5724_14920# a_5636_14964# vdd pfet_06v0 w=1.22u l=1u
X384 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X385 vdd a_21740_16055# a_21652_16152# vdd pfet_06v0 w=1.22u l=1u
X386 a_16588_16055# a_16500_16152# vss vss nfet_06v0 w=0.82u l=1u
X387 a_21180_14920# a_21092_14964# vss vss nfet_06v0 w=0.82u l=1u
X388 vdd a_5724_11784# a_5636_11828# vdd pfet_06v0 w=1.22u l=1u
X389 vdd a_1692_9783# a_1604_9880# vdd pfet_06v0 w=1.22u l=1u
X390 vdd a_1692_3511# a_1604_3608# vdd pfet_06v0 w=1.22u l=1u
X391 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X392 vdd a_1692_6647# a_1604_6744# vdd pfet_06v0 w=1.22u l=1u
X393 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X394 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X395 vdd a_10540_12919# a_10452_13016# vdd pfet_06v0 w=1.22u l=1u
X396 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X397 vdd a_8300_16055# a_8212_16152# vdd pfet_06v0 w=1.22u l=1u
X398 vdd a_8300_12919# a_8212_13016# vdd pfet_06v0 w=1.22u l=1u
X399 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X400 a_14124_11351# a_14036_11448# vss vss nfet_06v0 w=0.82u l=1u
X401 a_14572_14920# a_14484_14964# vss vss nfet_06v0 w=0.82u l=1u
X402 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X403 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X404 a_6620_11784# a_6532_11828# vss vss nfet_06v0 w=0.82u l=1u
X405 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X406 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X407 a_20844_9783# a_20756_9880# vss vss nfet_06v0 w=0.82u l=1u
X408 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X409 vdd a_1692_10216# a_1604_10260# vdd pfet_06v0 w=1.22u l=1u
X410 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X411 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X412 a_13228_11784# a_13140_11828# vss vss nfet_06v0 w=0.82u l=1u
X413 vdd a_1692_8648# a_1604_8692# vdd pfet_06v0 w=1.22u l=1u
X414 nseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X415 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X416 vdd nseries_gygy pseries_gygy vdd pfet_06v0 w=1.22u l=0.5u
X417 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X418 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X419 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X420 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X421 vdd a_10988_9783# a_10900_9880# vdd pfet_06v0 w=1.22u l=1u
X422 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X423 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X424 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X425 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X426 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X427 a_12108_3511# a_12020_3608# vss vss nfet_06v0 w=0.82u l=1u
X428 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X429 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X430 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X431 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X432 a_2140_8215# a_2052_8312# vss vss nfet_06v0 w=0.82u l=1u
X433 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X434 a_13900_16055# a_13812_16152# vss vss nfet_06v0 w=0.82u l=1u
X435 a_19388_14920# a_19300_14964# vss vss nfet_06v0 w=0.82u l=1u
X436 vdd a_19948_12919# a_19860_13016# vdd pfet_06v0 w=1.22u l=1u
X437 a_3932_12919# a_3844_13016# vss vss nfet_06v0 w=0.82u l=1u
X438 a_20620_14487# a_20532_14584# vss vss nfet_06v0 w=0.82u l=1u
X439 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X440 a_13676_11784# a_13588_11828# vss vss nfet_06v0 w=0.82u l=1u
X441 a_20620_11351# a_20532_11448# vss vss nfet_06v0 w=0.82u l=1u
X442 a_2588_14920# a_2500_14964# vss vss nfet_06v0 w=0.82u l=1u
X443 vdd a_8412_14920# a_8324_14964# vdd pfet_06v0 w=1.22u l=1u
X444 nseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X445 pseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X446 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X447 vdd a_8412_11784# a_8324_11828# vdd pfet_06v0 w=1.22u l=1u
X448 vdd a_3036_9783# a_2948_9880# vdd pfet_06v0 w=1.22u l=1u
X449 pshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X450 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X451 a_13564_12919# a_13476_13016# vss vss nfet_06v0 w=0.82u l=1u
X452 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X453 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X454 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X455 pshunt_gy pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X456 vdd a_18044_14920# a_17956_14964# vdd pfet_06v0 w=1.22u l=1u
X457 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X458 pseries_gygy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X459 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X460 vdd a_17820_16055# a_17732_16152# vdd pfet_06v0 w=1.22u l=1u
X461 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X462 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X463 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X464 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X465 a_2588_14487# a_2500_14584# vss vss nfet_06v0 w=0.82u l=1u
X466 a_2588_11351# a_2500_11448# vss vss nfet_06v0 w=0.82u l=1u
X467 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X468 vdd a_8860_14920# a_8772_14964# vdd pfet_06v0 w=1.22u l=1u
X469 vdd a_22076_14920# a_21988_14964# vdd pfet_06v0 w=1.22u l=1u
X470 vdd a_7068_13352# a_6980_13396# vdd pfet_06v0 w=1.22u l=1u
X471 vdd a_8860_11784# a_8772_11828# vdd pfet_06v0 w=1.22u l=1u
X472 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X473 a_10092_14920# a_10004_14964# vss vss nfet_06v0 w=0.82u l=1u
X474 vdd a_6508_14487# a_6420_14584# vdd pfet_06v0 w=1.22u l=1u
X475 vdd a_4380_10216# a_4292_10260# vdd pfet_06v0 w=1.22u l=1u
X476 nseries_gygy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X477 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X478 a_10988_12919# a_10900_13016# vss vss nfet_06v0 w=0.82u l=1u
X479 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X480 pshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X481 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X482 a_8748_12919# a_8660_13016# vss vss nfet_06v0 w=0.82u l=1u
X483 a_2140_11784# a_2052_11828# vss vss nfet_06v0 w=0.82u l=1u
X484 a_18716_16055# a_18628_16152# vss vss nfet_06v0 w=0.82u l=1u
X485 vdd a_15468_14920# a_15380_14964# vdd pfet_06v0 w=1.22u l=1u
X486 vdd a_18492_14920# a_18404_14964# vdd pfet_06v0 w=1.22u l=1u
X487 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X488 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X489 vdd a_1692_14920# a_1604_14964# vdd pfet_06v0 w=1.22u l=1u
X490 a_21068_13352# a_20980_13396# vss vss nfet_06v0 w=0.82u l=1u
X491 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X492 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X493 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X494 a_12556_3511# a_12468_3608# vss vss nfet_06v0 w=0.82u l=1u
X495 a_4828_13352# a_4740_13396# vss vss nfet_06v0 w=0.82u l=1u
X496 vdd a_1692_11784# a_1604_11828# vdd pfet_06v0 w=1.22u l=1u
X497 a_4828_10216# a_4740_10260# vss vss nfet_06v0 w=0.82u l=1u
X498 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X499 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X500 a_18828_14487# a_18740_14584# vss vss nfet_06v0 w=0.82u l=1u
X501 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X502 a_10092_14487# a_10004_14584# vss vss nfet_06v0 w=0.82u l=1u
X503 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X504 vdd a_6956_14487# a_6868_14584# vdd pfet_06v0 w=1.22u l=1u
X505 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X506 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X507 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X508 vdd a_3484_9783# a_3396_9880# vdd pfet_06v0 w=1.22u l=1u
X509 a_5276_14920# a_5188_14964# vss vss nfet_06v0 w=0.82u l=1u
X510 a_20732_14920# a_20644_14964# vss vss nfet_06v0 w=0.82u l=1u
X511 vdd a_14012_14487# a_13924_14584# vdd pfet_06v0 w=1.22u l=1u
X512 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X513 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X514 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X515 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X516 pbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X517 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X518 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X519 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X520 vdd a_1692_16055# a_1604_16152# vdd pfet_06v0 w=1.22u l=1u
X521 a_12332_13352# a_12244_13396# vss vss nfet_06v0 w=0.82u l=1u
X522 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X523 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X524 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X525 vdd a_1692_12919# a_1604_13016# vdd pfet_06v0 w=1.22u l=1u
X526 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X527 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X528 vdd a_11436_14487# a_11348_14584# vdd pfet_06v0 w=1.22u l=1u
X529 vdd a_14460_14487# a_14372_14584# vdd pfet_06v0 w=1.22u l=1u
X530 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X531 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X532 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X533 vdd a_11436_11351# a_11348_11448# vdd pfet_06v0 w=1.22u l=1u
X534 vss pshunt_gy nshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X535 vdd a_21516_12919# a_21428_13016# vdd pfet_06v0 w=1.22u l=1u
X536 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X537 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X538 a_2588_16055# a_2500_16152# vss vss nfet_06v0 w=0.82u l=1u
X539 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X540 a_21740_8648# a_21652_8692# vss vss nfet_06v0 w=0.82u l=1u
X541 a_12780_13352# a_12692_13396# vss vss nfet_06v0 w=0.82u l=1u
X542 vdd a_4380_14920# a_4292_14964# vdd pfet_06v0 w=1.22u l=1u
X543 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X544 a_7516_13352# a_7428_13396# vss vss nfet_06v0 w=0.82u l=1u
X545 vdd a_4380_11784# a_4292_11828# vdd pfet_06v0 w=1.22u l=1u
X546 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X547 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X548 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X549 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X550 vdd a_11884_14487# a_11796_14584# vdd pfet_06v0 w=1.22u l=1u
X551 vdd a_2140_9783# a_2052_9880# vdd pfet_06v0 w=1.22u l=1u
X552 vdd a_2140_3511# a_2052_3608# vdd pfet_06v0 w=1.22u l=1u
X553 vdd a_9644_14487# a_9556_14584# vdd pfet_06v0 w=1.22u l=1u
X554 vdd a_21964_12919# a_21876_13016# vdd pfet_06v0 w=1.22u l=1u
X555 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X556 a_8860_3511# a_8772_3608# vss vss nfet_06v0 w=0.82u l=1u
X557 vdd a_11436_13352# a_11348_13396# vdd pfet_06v0 w=1.22u l=1u
X558 pbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X559 vdd nseries_gy pseries_gygy vdd pfet_06v0 w=1.22u l=0.5u
X560 a_21292_16055# a_21204_16152# vss vss nfet_06v0 w=0.82u l=1u
X561 vdd a_19276_14487# a_19188_14584# vdd pfet_06v0 w=1.22u l=1u
X562 a_7964_13352# a_7876_13396# vss vss nfet_06v0 w=0.82u l=1u
X563 a_2140_12919# a_2052_13016# vss vss nfet_06v0 w=0.82u l=1u
X564 vdd a_4380_16055# a_4292_16152# vdd pfet_06v0 w=1.22u l=1u
X565 a_15020_13352# a_14932_13396# vss vss nfet_06v0 w=0.82u l=1u
X566 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X567 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X568 a_16812_14920# a_16724_14964# vss vss nfet_06v0 w=0.82u l=1u
X569 vdd a_4380_12919# a_4292_13016# vdd pfet_06v0 w=1.22u l=1u
X570 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X571 pbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X572 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X573 nbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X574 vdd a_11884_13352# a_11796_13396# vdd pfet_06v0 w=1.22u l=1u
X575 vdd a_2140_8648# a_2052_8692# vdd pfet_06v0 w=1.22u l=1u
X576 vdd a_21628_14920# a_21540_14964# vdd pfet_06v0 w=1.22u l=1u
X577 vdd a_9644_13352# a_9556_13396# vdd pfet_06v0 w=1.22u l=1u
X578 vdd a_14124_11351# a_14036_11448# vdd pfet_06v0 w=1.22u l=1u
X579 vdd a_3932_10216# a_3844_10260# vdd pfet_06v0 w=1.22u l=1u
X580 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X581 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X582 vdd a_19276_13352# a_19188_13396# vdd pfet_06v0 w=1.22u l=1u
X583 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X584 nbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X585 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X586 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X587 nseries_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X588 vdd a_20060_16055# a_19972_16152# vdd pfet_06v0 w=1.22u l=1u
X589 a_7068_11784# a_6980_11828# vss vss nfet_06v0 w=0.82u l=1u
X590 a_12892_6647# a_12804_6744# vss vss nfet_06v0 w=0.82u l=1u
X591 a_20396_12919# a_20308_13016# vss vss nfet_06v0 w=0.82u l=1u
X592 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X593 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X594 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X595 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X596 vss nbusin_nshunt pshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X597 pshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X598 vdd a_13452_16055# a_13364_16152# vdd pfet_06v0 w=1.22u l=1u
X599 a_7404_14487# a_7316_14584# vss vss nfet_06v0 w=0.82u l=1u
X600 vdd a_9196_12919# a_9108_13016# vdd pfet_06v0 w=1.22u l=1u
X601 vdd a_10428_16055# a_10340_16152# vdd pfet_06v0 w=1.22u l=1u
X602 a_3036_13352# a_2948_13396# vss vss nfet_06v0 w=0.82u l=1u
X603 vdd a_14124_13352# a_14036_13396# vdd pfet_06v0 w=1.22u l=1u
X604 a_3036_10216# a_2948_10260# vss vss nfet_06v0 w=0.82u l=1u
X605 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X606 vdd a_12108_3511# a_12020_3608# vdd pfet_06v0 w=1.22u l=1u
X607 a_4828_14920# a_4740_14964# vss vss nfet_06v0 w=0.82u l=1u
X608 nseries_gygy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X609 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X610 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X611 pseries_gygy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X612 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X613 vdd a_20620_14487# a_20532_14584# vdd pfet_06v0 w=1.22u l=1u
X614 vdd a_20620_11351# a_20532_11448# vdd pfet_06v0 w=1.22u l=1u
X615 pseries_gygy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X616 a_13564_6647# a_13476_6744# vss vss nfet_06v0 w=0.82u l=1u
X617 a_14348_16055# a_14260_16152# vss vss nfet_06v0 w=0.82u l=1u
X618 a_17372_16055# a_17284_16152# vss vss nfet_06v0 w=0.82u l=1u
X619 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X620 a_7852_14487# a_7764_14584# vss vss nfet_06v0 w=0.82u l=1u
X621 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X622 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X623 vdd a_10876_16055# a_10788_16152# vdd pfet_06v0 w=1.22u l=1u
X624 a_4828_14487# a_4740_14584# vss vss nfet_06v0 w=0.82u l=1u
X625 a_3484_13352# a_3396_13396# vss vss nfet_06v0 w=0.82u l=1u
X626 vdd a_14572_13352# a_14484_13396# vdd pfet_06v0 w=1.22u l=1u
X627 a_4828_11351# a_4740_11448# vss vss nfet_06v0 w=0.82u l=1u
X628 a_3484_10216# a_3396_10260# vss vss nfet_06v0 w=0.82u l=1u
X629 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X630 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X631 pbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X632 pseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X633 a_12332_14920# a_12244_14964# vss vss nfet_06v0 w=0.82u l=1u
X634 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X635 nbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X636 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X637 vdd a_2588_14487# a_2500_14584# vdd pfet_06v0 w=1.22u l=1u
X638 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X639 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X640 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X641 vdd a_18268_16055# a_18180_16152# vdd pfet_06v0 w=1.22u l=1u
X642 a_12220_16055# a_12132_16152# vss vss nfet_06v0 w=0.82u l=1u
X643 vdd a_2588_11351# a_2500_11448# vdd pfet_06v0 w=1.22u l=1u
X644 nbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X645 pbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X646 a_11660_8215# a_11572_8312# vss vss nfet_06v0 w=0.82u l=1u
X647 vdd a_3932_14920# a_3844_14964# vdd pfet_06v0 w=1.22u l=1u
X648 a_14796_16055# a_14708_16152# vss vss nfet_06v0 w=0.82u l=1u
X649 vdd a_20620_13352# a_20532_13396# vdd pfet_06v0 w=1.22u l=1u
X650 vdd a_3932_11784# a_3844_11828# vdd pfet_06v0 w=1.22u l=1u
X651 nshunt_gy pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X652 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X653 vss nseries_gy pbusout vss nfet_06v0 w=0.82u l=0.6u
X654 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X655 a_19724_13352# a_19636_13396# vss vss nfet_06v0 w=0.82u l=1u
X656 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X657 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X658 a_12332_14487# a_12244_14584# vss vss nfet_06v0 w=0.82u l=1u
X659 nbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X660 a_12780_14920# a_12692_14964# vss vss nfet_06v0 w=0.82u l=1u
X661 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X662 vdd a_12556_3511# a_12468_3608# vdd pfet_06v0 w=1.22u l=1u
X663 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X664 vdd a_16140_16055# a_16052_16152# vdd pfet_06v0 w=1.22u l=1u
X665 pseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X666 a_7516_14920# a_7428_14964# vss vss nfet_06v0 w=0.82u l=1u
X667 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X668 vdd a_10092_14487# a_10004_14584# vdd pfet_06v0 w=1.22u l=1u
X669 vdd a_18828_14487# a_18740_14584# vdd pfet_06v0 w=1.22u l=1u
X670 a_7404_16055# a_7316_16152# vss vss nfet_06v0 w=0.82u l=1u
X671 vdd a_2588_13352# a_2500_13396# vdd pfet_06v0 w=1.22u l=1u
X672 nbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X673 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X674 vdd a_3932_16055# a_3844_16152# vdd pfet_06v0 w=1.22u l=1u
X675 vdd a_3932_12919# a_3844_13016# vdd pfet_06v0 w=1.22u l=1u
X676 a_11436_11784# a_11348_11828# vss vss nfet_06v0 w=0.82u l=1u
X677 pshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X678 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X679 nbusin_nshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X680 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X681 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X682 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X683 vdd a_10988_14920# a_10900_14964# vdd pfet_06v0 w=1.22u l=1u
X684 a_12780_14487# a_12692_14584# vss vss nfet_06v0 w=0.82u l=1u
X685 vdd a_10988_11784# a_10900_11828# vdd pfet_06v0 w=1.22u l=1u
X686 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X687 a_6172_13352# a_6084_13396# vss vss nfet_06v0 w=0.82u l=1u
X688 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X689 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X690 a_7964_14920# a_7876_14964# vss vss nfet_06v0 w=0.82u l=1u
X691 vdd a_13564_12919# a_13476_13016# vdd pfet_06v0 w=1.22u l=1u
X692 a_13452_3511# a_13364_3608# vss vss nfet_06v0 w=0.82u l=1u
X693 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X694 a_15020_14920# a_14932_14964# vss vss nfet_06v0 w=0.82u l=1u
X695 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X696 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X697 a_7852_16055# a_7764_16152# vss vss nfet_06v0 w=0.82u l=1u
X698 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X699 a_4828_16055# a_4740_16152# vss vss nfet_06v0 w=0.82u l=1u
X700 a_17596_14920# a_17508_14964# vss vss nfet_06v0 w=0.82u l=1u
X701 nshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X702 vdd a_10092_13352# a_10004_13396# vdd pfet_06v0 w=1.22u l=1u
X703 vdd a_18828_13352# a_18740_13396# vdd pfet_06v0 w=1.22u l=1u
X704 a_11884_11784# a_11796_11828# vss vss nfet_06v0 w=0.82u l=1u
X705 vdd a_6620_14920# a_6532_14964# vdd pfet_06v0 w=1.22u l=1u
X706 a_9644_11784# a_9556_11828# vss vss nfet_06v0 w=0.82u l=1u
X707 vss pshunt_gy pbusin_pshunt vss nfet_06v0 w=0.82u l=0.6u
X708 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X709 vdd a_6620_11784# a_6532_11828# vdd pfet_06v0 w=1.22u l=1u
X710 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X711 a_22076_5079# a_21988_5176# vss vss nfet_06v0 w=0.82u l=1u
X712 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X713 vdd a_2140_10216# a_2052_10260# vdd pfet_06v0 w=1.22u l=1u
X714 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X715 vdd a_10988_12919# a_10900_13016# vdd pfet_06v0 w=1.22u l=1u
X716 a_6508_12919# a_6420_13016# vss vss nfet_06v0 w=0.82u l=1u
X717 vdd a_8748_16055# a_8660_16152# vdd pfet_06v0 w=1.22u l=1u
X718 vdd a_13228_14920# a_13140_14964# vdd pfet_06v0 w=1.22u l=1u
X719 vdd a_13228_11784# a_13140_11828# vdd pfet_06v0 w=1.22u l=1u
X720 vdd a_8748_12919# a_8660_13016# vdd pfet_06v0 w=1.22u l=1u
X721 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X722 vdd nseries_gy nbusin_nshunt vdd pfet_06v0 w=1.22u l=0.5u
X723 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X724 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X725 vdd a_9644_8648# a_9556_8692# vdd pfet_06v0 w=1.22u l=1u
X726 pseries_gygy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X727 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X728 a_20508_16055# a_20420_16152# vss vss nfet_06v0 w=0.82u l=1u
X729 vdd a_20284_14920# a_20196_14964# vdd pfet_06v0 w=1.22u l=1u
X730 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X731 vdd a_5276_13352# a_5188_13396# vdd pfet_06v0 w=1.22u l=1u
X732 pbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X733 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X734 vdd a_8860_3511# a_8772_3608# vdd pfet_06v0 w=1.22u l=1u
X735 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X736 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X737 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X738 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X739 a_3036_14920# a_2948_14964# vss vss nfet_06v0 w=0.82u l=1u
X740 a_6956_12919# a_6868_13016# vss vss nfet_06v0 w=0.82u l=1u
X741 vdd a_13676_14920# a_13588_14964# vdd pfet_06v0 w=1.22u l=1u
X742 vdd a_13676_11784# a_13588_11828# vdd pfet_06v0 w=1.22u l=1u
X743 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X744 a_14012_12919# a_13924_13016# vss vss nfet_06v0 w=0.82u l=1u
X745 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X746 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X747 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X748 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X749 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X750 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X751 vdd nseries_gy nbusin_nshunt vdd pfet_06v0 w=1.22u l=0.5u
X752 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X753 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X754 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X755 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X756 a_6060_14487# a_5972_14584# vss vss nfet_06v0 w=0.82u l=1u
X757 vss nbusin_nshunt pbusin_pshunt vss nfet_06v0 w=0.82u l=0.6u
X758 a_3036_14487# a_2948_14584# vss vss nfet_06v0 w=0.82u l=1u
X759 a_3036_11351# a_2948_11448# vss vss nfet_06v0 w=0.82u l=1u
X760 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X761 a_3484_14920# a_3396_14964# vss vss nfet_06v0 w=0.82u l=1u
X762 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X763 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X764 a_11436_12919# a_11348_13016# vss vss nfet_06v0 w=0.82u l=1u
X765 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X766 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X767 a_10540_13352# a_10452_13396# vss vss nfet_06v0 w=0.82u l=1u
X768 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X769 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X770 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X771 vdd a_2140_14920# a_2052_14964# vdd pfet_06v0 w=1.22u l=1u
X772 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X773 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X774 a_21516_7080# a_21428_7124# vss vss nfet_06v0 w=0.82u l=1u
X775 vdd a_2140_11784# a_2052_11828# vdd pfet_06v0 w=1.22u l=1u
X776 vdd a_12892_6647# a_12804_6744# vdd pfet_06v0 w=1.22u l=1u
X777 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X778 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X779 a_21292_8648# a_21204_8692# vss vss nfet_06v0 w=0.82u l=1u
X780 a_3484_14487# a_3396_14584# vss vss nfet_06v0 w=0.82u l=1u
X781 a_3484_11351# a_3396_11448# vss vss nfet_06v0 w=0.82u l=1u
X782 vss pshunt_gy nshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X783 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X784 vdd nbusin_nshunt pshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X785 vdd a_7404_14487# a_7316_14584# vdd pfet_06v0 w=1.22u l=1u
X786 a_11884_12919# a_11796_13016# vss vss nfet_06v0 w=0.82u l=1u
X787 a_19612_16055# a_19524_16152# vss vss nfet_06v0 w=0.82u l=1u
X788 a_9644_12919# a_9556_13016# vss vss nfet_06v0 w=0.82u l=1u
X789 nbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X790 vdd a_16364_14920# a_16276_14964# vdd pfet_06v0 w=1.22u l=1u
X791 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X792 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X793 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X794 a_5724_13352# a_5636_13396# vss vss nfet_06v0 w=0.82u l=1u
X795 a_2588_11784# a_2500_11828# vss vss nfet_06v0 w=0.82u l=1u
X796 nshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X797 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X798 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X799 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X800 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X801 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X802 vdd a_2140_16055# a_2052_16152# vdd pfet_06v0 w=1.22u l=1u
X803 vdd a_2140_12919# a_2052_13016# vdd pfet_06v0 w=1.22u l=1u
X804 vdd a_13564_6647# a_13476_6744# vdd pfet_06v0 w=1.22u l=1u
X805 a_19724_14487# a_19636_14584# vss vss nfet_06v0 w=0.82u l=1u
X806 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X807 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X808 pbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X809 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X810 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X811 vdd a_4828_14487# a_4740_14584# vdd pfet_06v0 w=1.22u l=1u
X812 vdd a_7852_14487# a_7764_14584# vdd pfet_06v0 w=1.22u l=1u
X813 nbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X814 pshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X815 vdd a_4828_11351# a_4740_11448# vdd pfet_06v0 w=1.22u l=1u
X816 a_6172_14920# a_6084_14964# vss vss nfet_06v0 w=0.82u l=1u
X817 pseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X818 pseries_gy pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X819 a_6060_16055# a_5972_16152# vss vss nfet_06v0 w=0.82u l=1u
X820 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X821 a_3036_16055# a_2948_16152# vss vss nfet_06v0 w=0.82u l=1u
X822 a_21292_11784# a_21204_11828# vss vss nfet_06v0 w=0.82u l=1u
X823 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X824 a_10092_11784# a_10004_11828# vss vss nfet_06v0 w=0.82u l=1u
X825 nseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X826 a_21964_7080# a_21876_7124# vss vss nfet_06v0 w=0.82u l=1u
X827 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X828 vss nseries_gygy nseries_gygy vss nfet_06v0 w=0.82u l=0.6u
X829 a_1692_3944# a_1604_3988# vss vss nfet_06v0 w=0.82u l=1u
X830 a_22076_9783# a_21988_9880# vss vss nfet_06v0 w=0.82u l=1u
X831 a_20844_8215# a_20756_8312# vss vss nfet_06v0 w=0.82u l=1u
X832 vdd nseries_gy pbusout vdd pfet_06v0 w=1.22u l=0.5u
X833 nbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X834 vdd a_12332_14487# a_12244_14584# vdd pfet_06v0 w=1.22u l=1u
X835 vdd a_21068_13352# a_20980_13396# vdd pfet_06v0 w=1.22u l=1u
X836 vdd a_20396_12919# a_20308_13016# vdd pfet_06v0 w=1.22u l=1u
X837 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X838 vdd a_4828_13352# a_4740_13396# vdd pfet_06v0 w=1.22u l=1u
X839 pseries_gy pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X840 vdd a_16812_8648# a_16724_8692# vdd pfet_06v0 w=1.22u l=1u
X841 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X842 a_3484_16055# a_3396_16152# vss vss nfet_06v0 w=0.82u l=1u
X843 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X844 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X845 a_8412_13352# a_8324_13396# vss vss nfet_06v0 w=0.82u l=1u
X846 a_5276_11784# a_5188_11828# vss vss nfet_06v0 w=0.82u l=1u
X847 a_2588_8648# a_2500_8692# vss vss nfet_06v0 w=0.82u l=1u
X848 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X849 pshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X850 vdd a_12780_14487# a_12692_14584# vdd pfet_06v0 w=1.22u l=1u
X851 nbusout pbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X852 a_21516_8215# a_21428_8312# vss vss nfet_06v0 w=0.82u l=1u
X853 a_19836_14920# a_19748_14964# vss vss nfet_06v0 w=0.82u l=1u
X854 a_5612_14487# a_5524_14584# vss vss nfet_06v0 w=0.82u l=1u
X855 a_5612_11351# a_5524_11448# vss vss nfet_06v0 w=0.82u l=1u
X856 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X857 vdd a_12332_13352# a_12244_13396# vdd pfet_06v0 w=1.22u l=1u
X858 vdd a_13452_3511# a_13364_3608# vdd pfet_06v0 w=1.22u l=1u
X859 vdd a_1692_8215# a_1604_8312# vdd pfet_06v0 w=1.22u l=1u
X860 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X861 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X862 a_8860_13352# a_8772_13396# vss vss nfet_06v0 w=0.82u l=1u
X863 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X864 vdd pshunt_gy pbusin_pshunt vdd pfet_06v0 w=1.22u l=0.5u
X865 a_2588_12919# a_2500_13016# vss vss nfet_06v0 w=0.82u l=1u
X866 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X867 pshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X868 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X869 a_15468_13352# a_15380_13396# vss vss nfet_06v0 w=0.82u l=1u
X870 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X871 vdd a_7068_14920# a_6980_14964# vdd pfet_06v0 w=1.22u l=1u
X872 a_1692_13352# a_1604_13396# vss vss nfet_06v0 w=0.82u l=1u
X873 vdd a_12780_13352# a_12692_13396# vdd pfet_06v0 w=1.22u l=1u
X874 vdd a_7068_11784# a_6980_11828# vdd pfet_06v0 w=1.22u l=1u
X875 a_1692_10216# a_1604_10260# vss vss nfet_06v0 w=0.82u l=1u
X876 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X877 a_20620_6647# a_20532_6744# vss vss nfet_06v0 w=0.82u l=1u
X878 a_10540_14920# a_10452_14964# vss vss nfet_06v0 w=0.82u l=1u
X879 vdd a_7516_13352# a_7428_13396# vdd pfet_06v0 w=1.22u l=1u
X880 vss nbusout nseries_gy vss nfet_06v0 w=0.82u l=0.6u
X881 a_20620_3511# a_20532_3608# vss vss nfet_06v0 w=0.82u l=1u
X882 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X883 vdd a_18940_14920# a_18852_14964# vdd pfet_06v0 w=1.22u l=1u
X884 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X885 vdd a_15916_14920# a_15828_14964# vdd pfet_06v0 w=1.22u l=1u
X886 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X887 a_21516_13352# a_21428_13396# vss vss nfet_06v0 w=0.82u l=1u
X888 pseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X889 vdd nseries_gygy nseries_gygy vdd pfet_06v0 w=1.22u l=0.5u
X890 nbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X891 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X892 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X893 a_10092_12919# a_10004_13016# vss vss nfet_06v0 w=0.82u l=1u
X894 a_21964_8215# a_21876_8312# vss vss nfet_06v0 w=0.82u l=1u
X895 a_10540_14487# a_10452_14584# vss vss nfet_06v0 w=0.82u l=1u
X896 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X897 a_1692_5079# a_1604_5176# vss vss nfet_06v0 w=0.82u l=1u
X898 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X899 vdd a_7964_13352# a_7876_13396# vdd pfet_06v0 w=1.22u l=1u
X900 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X901 a_8300_14487# a_8212_14584# vss vss nfet_06v0 w=0.82u l=1u
X902 nseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X903 vdd a_11324_16055# a_11236_16152# vdd pfet_06v0 w=1.22u l=1u
X904 a_5724_14920# a_5636_14964# vss vss nfet_06v0 w=0.82u l=1u
X905 vdd a_15020_13352# a_14932_13396# vdd pfet_06v0 w=1.22u l=1u
X906 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X907 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X908 a_21964_13352# a_21876_13396# vss vss nfet_06v0 w=0.82u l=1u
X909 vss nbusin_nshunt pshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X910 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X911 a_5612_16055# a_5524_16152# vss vss nfet_06v0 w=0.82u l=1u
X912 vdd nbusin_nshunt pbusin_pshunt vdd pfet_06v0 w=1.22u l=0.5u
X913 vdd a_3036_14487# a_2948_14584# vdd pfet_06v0 w=1.22u l=1u
X914 vdd a_6060_14487# a_5972_14584# vdd pfet_06v0 w=1.22u l=1u
X915 a_20844_11784# a_20756_11828# vss vss nfet_06v0 w=0.82u l=1u
X916 vdd a_3036_11351# a_2948_11448# vdd pfet_06v0 w=1.22u l=1u
X917 vss pbusin_pshunt nshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X918 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X919 a_15244_16055# a_15156_16152# vss vss nfet_06v0 w=0.82u l=1u
X920 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X921 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X922 a_2588_9783# a_2500_9880# vss vss nfet_06v0 w=0.82u l=1u
X923 vdd a_20844_9783# a_20756_9880# vdd pfet_06v0 w=1.22u l=1u
X924 vdd a_22076_5079# a_21988_5176# vdd pfet_06v0 w=1.22u l=1u
X925 nseries_gy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X926 vdd a_11772_16055# a_11684_16152# vdd pfet_06v0 w=1.22u l=1u
X927 a_4380_13352# a_4292_13396# vss vss nfet_06v0 w=0.82u l=1u
X928 a_4380_10216# a_4292_10260# vss vss nfet_06v0 w=0.82u l=1u
X929 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X930 vdd a_9532_16055# a_9444_16152# vdd pfet_06v0 w=1.22u l=1u
X931 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X932 nseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X933 vdd a_6508_16055# a_6420_16152# vdd pfet_06v0 w=1.22u l=1u
X934 vdd a_6508_12919# a_6420_13016# vdd pfet_06v0 w=1.22u l=1u
X935 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X936 a_18380_14487# a_18292_14584# vss vss nfet_06v0 w=0.82u l=1u
X937 a_1692_8648# a_1604_8692# vss vss nfet_06v0 w=0.82u l=1u
X938 a_11548_3944# a_11460_3988# vss vss nfet_06v0 w=0.82u l=1u
X939 a_15356_14487# a_15268_14584# vss vss nfet_06v0 w=0.82u l=1u
X940 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X941 vdd a_3484_14487# a_3396_14584# vdd pfet_06v0 w=1.22u l=1u
X942 vss pbusin_pshunt nshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X943 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X944 vdd a_19164_16055# a_19076_16152# vdd pfet_06v0 w=1.22u l=1u
X945 vdd a_3484_11351# a_3396_11448# vdd pfet_06v0 w=1.22u l=1u
X946 a_4828_11784# a_4740_11828# vss vss nfet_06v0 w=0.82u l=1u
X947 pbusin_pshunt pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X948 a_15692_16055# a_15604_16152# vss vss nfet_06v0 w=0.82u l=1u
X949 vdd a_3036_13352# a_2948_13396# vdd pfet_06v0 w=1.22u l=1u
X950 nseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X951 a_12668_16055# a_12580_16152# vss vss nfet_06v0 w=0.82u l=1u
X952 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X953 vdd a_9980_16055# a_9892_16152# vdd pfet_06v0 w=1.22u l=1u
X954 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X955 vdd a_6956_16055# a_6868_16152# vdd pfet_06v0 w=1.22u l=1u
X956 vdd a_11436_14920# a_11348_14964# vdd pfet_06v0 w=1.22u l=1u
X957 vdd a_6956_12919# a_6868_13016# vdd pfet_06v0 w=1.22u l=1u
X958 vdd a_11436_11784# a_11348_11828# vdd pfet_06v0 w=1.22u l=1u
X959 vdd a_20844_8648# a_20756_8692# vdd pfet_06v0 w=1.22u l=1u
X960 a_21740_3511# a_21652_3608# vss vss nfet_06v0 w=0.82u l=1u
X961 nshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X962 a_8412_14920# a_8324_14964# vss vss nfet_06v0 w=0.82u l=1u
X963 vdd a_14012_12919# a_13924_13016# vdd pfet_06v0 w=1.22u l=1u
X964 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X965 vdd a_16588_16055# a_16500_16152# vdd pfet_06v0 w=1.22u l=1u
X966 a_21740_16055# a_21652_16152# vss vss nfet_06v0 w=0.82u l=1u
X967 vdd a_19724_14487# a_19636_14584# vdd pfet_06v0 w=1.22u l=1u
X968 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X969 pseries_gygy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X970 pseries_gy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X971 a_8300_16055# a_8212_16152# vss vss nfet_06v0 w=0.82u l=1u
X972 vdd a_3484_13352# a_3396_13396# vdd pfet_06v0 w=1.22u l=1u
X973 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X974 pshunt_gy pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X975 a_18044_14920# a_17956_14964# vss vss nfet_06v0 w=0.82u l=1u
X976 a_12332_11784# a_12244_11828# vss vss nfet_06v0 w=0.82u l=1u
X977 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X978 pseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X979 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X980 vdd a_11884_14920# a_11796_14964# vdd pfet_06v0 w=1.22u l=1u
X981 vdd a_11884_11784# a_11796_11828# vdd pfet_06v0 w=1.22u l=1u
X982 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X983 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X984 vdd a_9644_14920# a_9556_14964# vdd pfet_06v0 w=1.22u l=1u
X985 a_8860_14920# a_8772_14964# vss vss nfet_06v0 w=0.82u l=1u
X986 a_22076_14920# a_21988_14964# vss vss nfet_06v0 w=0.82u l=1u
X987 vdd a_9644_11784# a_9556_11828# vdd pfet_06v0 w=1.22u l=1u
X988 pshunt_gy pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X989 vss pshunt_gy nshunt_gy vss nfet_06v0 w=0.82u l=0.6u
X990 vdd a_11436_12919# a_11348_13016# vdd pfet_06v0 w=1.22u l=1u
X991 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X992 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X993 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X994 nshunt_gy nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X995 nshunt_gy pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X996 nseries_gy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X997 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X998 nbusout nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X999 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1000 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1001 pbusin_pshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1002 a_15468_14920# a_15380_14964# vss vss nfet_06v0 w=0.82u l=1u
X1003 a_18492_14920# a_18404_14964# vss vss nfet_06v0 w=0.82u l=1u
X1004 vdd a_19724_13352# a_19636_13396# vdd pfet_06v0 w=1.22u l=1u
X1005 a_10876_5079# a_10788_5176# vss vss nfet_06v0 w=0.82u l=1u
X1006 a_1692_14920# a_1604_14964# vss vss nfet_06v0 w=0.82u l=1u
X1007 a_12780_11784# a_12692_11828# vss vss nfet_06v0 w=0.82u l=1u
X1008 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1009 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1010 a_7516_11784# a_7428_11828# vss vss nfet_06v0 w=0.82u l=1u
X1011 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X1012 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1013 a_20844_12919# a_20756_13016# vss vss nfet_06v0 w=0.82u l=1u
X1014 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1015 vdd a_2140_8215# a_2052_8312# vdd pfet_06v0 w=1.22u l=1u
X1016 nseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1017 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1018 vdd a_11884_12919# a_11796_13016# vdd pfet_06v0 w=1.22u l=1u
X1019 a_7404_12919# a_7316_13016# vss vss nfet_06v0 w=0.82u l=1u
X1020 vdd a_2588_10216# a_2500_10260# vdd pfet_06v0 w=1.22u l=1u
X1021 vdd a_14124_14920# a_14036_14964# vdd pfet_06v0 w=1.22u l=1u
X1022 vdd a_9644_12919# a_9556_13016# vdd pfet_06v0 w=1.22u l=1u
X1023 vdd a_13900_16055# a_13812_16152# vdd pfet_06v0 w=1.22u l=1u
X1024 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1025 a_1692_14487# a_1604_14584# vss vss nfet_06v0 w=0.82u l=1u
X1026 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1027 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1028 a_1692_11351# a_1604_11448# vss vss nfet_06v0 w=0.82u l=1u
X1029 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1030 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1031 vdd a_21180_14920# a_21092_14964# vdd pfet_06v0 w=1.22u l=1u
X1032 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1033 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1034 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1035 a_1692_9783# a_1604_9880# vss vss nfet_06v0 w=0.82u l=1u
X1036 vdd a_5612_14487# a_5524_14584# vdd pfet_06v0 w=1.22u l=1u
X1037 vdd a_6172_13352# a_6084_13396# vdd pfet_06v0 w=1.22u l=1u
X1038 a_7964_11784# a_7876_11828# vss vss nfet_06v0 w=0.82u l=1u
X1039 vdd a_5612_11351# a_5524_11448# vdd pfet_06v0 w=1.22u l=1u
X1040 a_17820_16055# a_17732_16152# vss vss nfet_06v0 w=0.82u l=1u
X1041 a_4828_12919# a_4740_13016# vss vss nfet_06v0 w=0.82u l=1u
X1042 a_7852_12919# a_7764_13016# vss vss nfet_06v0 w=0.82u l=1u
X1043 vdd a_14572_14920# a_14484_14964# vdd pfet_06v0 w=1.22u l=1u
X1044 a_21516_14487# a_21428_14584# vss vss nfet_06v0 w=0.82u l=1u
X1045 nbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1046 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1047 a_20172_13352# a_20084_13396# vss vss nfet_06v0 w=0.82u l=1u
X1048 a_21516_11351# a_21428_11448# vss vss nfet_06v0 w=0.82u l=1u
X1049 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1050 pseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1051 a_3932_13352# a_3844_13396# vss vss nfet_06v0 w=0.82u l=1u
X1052 a_3932_10216# a_3844_10260# vss vss nfet_06v0 w=0.82u l=1u
X1053 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1054 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1055 nbusin_nshunt nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1056 a_14908_14487# a_14820_14584# vss vss nfet_06v0 w=0.82u l=1u
X1057 a_17932_14487# a_17844_14584# vss vss nfet_06v0 w=0.82u l=1u
X1058 nseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1059 pbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1060 pshunt_gy pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1061 vdd a_18716_16055# a_18628_16152# vdd pfet_06v0 w=1.22u l=1u
X1062 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1063 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1064 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1065 pshunt_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1066 a_4380_14920# a_4292_14964# vss vss nfet_06v0 w=0.82u l=1u
X1067 nseries_gy nseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1068 vdd a_20620_3511# a_20532_3608# vdd pfet_06v0 w=1.22u l=1u
X1069 pshunt_gy nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1070 vdd a_20620_6647# a_20532_6744# vdd pfet_06v0 w=1.22u l=1u
X1071 a_21964_14487# a_21876_14584# vss vss nfet_06v0 w=0.82u l=1u
X1072 a_10988_9783# a_10900_9880# vss vss nfet_06v0 w=0.82u l=1u
X1073 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1074 a_21964_11351# a_21876_11448# vss vss nfet_06v0 w=0.82u l=1u
X1075 a_12332_12919# a_12244_13016# vss vss nfet_06v0 w=0.82u l=1u
X1076 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1077 pseries_gy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1078 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1079 a_3036_11784# a_2948_11828# vss vss nfet_06v0 w=0.82u l=1u
X1080 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1081 vdd a_19388_14920# a_19300_14964# vdd pfet_06v0 w=1.22u l=1u
X1082 a_10988_13352# a_10900_13396# vss vss nfet_06v0 w=0.82u l=1u
X1083 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1084 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1085 a_4380_14487# a_4292_14584# vss vss nfet_06v0 w=0.82u l=1u
X1086 nseries_gy nbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1087 vdd a_2588_14920# a_2500_14964# vdd pfet_06v0 w=1.22u l=1u
X1088 vdd a_2588_11784# a_2500_11828# vdd pfet_06v0 w=1.22u l=1u
X1089 a_4380_11351# a_4292_11448# vss vss nfet_06v0 w=0.82u l=1u
X1090 vdd a_10540_14487# a_10452_14584# vdd pfet_06v0 w=1.22u l=1u
X1091 pbusin_pshunt pshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1092 nshunt_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1093 vdd a_8300_14487# a_8212_14584# vdd pfet_06v0 w=1.22u l=1u
X1094 a_3036_9783# a_2948_9880# vss vss nfet_06v0 w=0.82u l=1u
X1095 nbusin_nshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1096 pseries_gygy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1097 a_1692_16055# a_1604_16152# vss vss nfet_06v0 w=0.82u l=1u
X1098 a_12780_12919# a_12692_13016# vss vss nfet_06v0 w=0.82u l=1u
X1099 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1100 vss nseries_gy pbusout vss nfet_06v0 w=0.82u l=0.6u
X1101 pseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X1102 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1103 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1104 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1105 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1106 a_3484_11784# a_3396_11828# vss vss nfet_06v0 w=0.82u l=1u
X1107 a_2140_8648# a_2052_8692# vss vss nfet_06v0 w=0.82u l=1u
X1108 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1109 vdd nbusin_nshunt pshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X1110 a_21628_14920# a_21540_14964# vss vss nfet_06v0 w=0.82u l=1u
X1111 a_6620_13352# a_6532_13396# vss vss nfet_06v0 w=0.82u l=1u
X1112 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1113 vdd pbusin_pshunt nshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X1114 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1115 nbusout pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1116 vdd a_2588_16055# a_2500_16152# vdd pfet_06v0 w=1.22u l=1u
X1117 vdd a_10092_14920# a_10004_14964# vdd pfet_06v0 w=1.22u l=1u
X1118 a_13228_13352# a_13140_13396# vss vss nfet_06v0 w=0.82u l=1u
X1119 vdd a_10092_11784# a_10004_11828# vdd pfet_06v0 w=1.22u l=1u
X1120 vdd a_21292_11784# a_21204_11828# vdd pfet_06v0 w=1.22u l=1u
X1121 vdd a_2588_12919# a_2500_13016# vdd pfet_06v0 w=1.22u l=1u
X1122 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X1123 vdd nseries_gygy nseries_gygy vdd pfet_06v0 w=1.22u l=0.5u
X1124 vdd a_10540_13352# a_10452_13396# vdd pfet_06v0 w=1.22u l=1u
X1125 pshunt_gy pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1126 nbusin_nshunt nshunt_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1127 vdd a_1692_3944# a_1604_3988# vdd pfet_06v0 w=1.22u l=1u
X1128 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1129 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1130 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1131 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1132 a_9196_14487# a_9108_14584# vss vss nfet_06v0 w=0.82u l=1u
X1133 pseries_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1134 vdd a_15356_14487# a_15268_14584# vdd pfet_06v0 w=1.22u l=1u
X1135 vdd a_18380_14487# a_18292_14584# vdd pfet_06v0 w=1.22u l=1u
X1136 pseries_gygy pseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X1137 pseries_gy nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1138 nbusin_nshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1139 nseries_gy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1140 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1141 nshunt_gy pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1142 nbusout pbusout vss vss nfet_06v0 w=0.82u l=0.6u
X1143 vdd pbusin_pshunt nshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X1144 nseries_gygy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X1145 pbusout nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1146 pbusout nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1147 a_13676_13352# a_13588_13396# vss vss nfet_06v0 w=0.82u l=1u
X1148 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1149 vdd a_21292_16055# a_21204_16152# vdd pfet_06v0 w=1.22u l=1u
X1150 vdd a_5276_14920# a_5188_14964# vdd pfet_06v0 w=1.22u l=1u
X1151 vdd a_20732_14920# a_20644_14964# vdd pfet_06v0 w=1.22u l=1u
X1152 vdd a_5276_11784# a_5188_11828# vdd pfet_06v0 w=1.22u l=1u
X1153 a_3484_9783# a_3396_9880# vss vss nfet_06v0 w=0.82u l=1u
X1154 nseries_gy nseries_gygy vss vss nfet_06v0 w=0.82u l=0.6u
X1155 vdd a_10092_12919# a_10004_13016# vdd pfet_06v0 w=1.22u l=1u
X1156 vdd a_5724_13352# a_5636_13396# vdd pfet_06v0 w=1.22u l=1u
X1157 nbusin_nshunt nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1158 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1159 vdd a_21740_3511# a_21652_3608# vdd pfet_06v0 w=1.22u l=1u
X1160 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1161 vdd a_1692_5079# a_1604_5176# vdd pfet_06v0 w=1.22u l=1u
X1162 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1163 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1164 pbusin_pshunt nbusin_nshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1165 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1166 nbusin_nshunt nshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1167 a_4380_16055# a_4292_16152# vss vss nfet_06v0 w=0.82u l=1u
X1168 a_8636_11351# a_8548_11448# vss vss nfet_06v0 w=0.82u l=1u
X1169 pbusin_pshunt pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1170 pseries_gygy nseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1171 a_6172_11784# a_6084_11828# vss vss nfet_06v0 w=0.82u l=1u
X1172 a_8860_3944# a_8772_3988# vss vss nfet_06v0 w=0.82u l=1u
X1173 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1174 nseries_gygy pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1175 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1176 nseries_gygy pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1177 pbusout nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X1178 a_6060_12919# a_5972_13016# vss vss nfet_06v0 w=0.82u l=1u
X1179 pbusin_pshunt pbusin_pshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1180 a_3036_12919# a_2948_13016# vss vss nfet_06v0 w=0.82u l=1u
X1181 pseries_gygy nseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1182 pshunt_gy nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1183 pshunt_gy pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1184 nshunt_gy pshunt_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1185 vdd pshunt_gy nshunt_gy vdd pfet_06v0 w=1.22u l=0.5u
X1186 a_3932_14920# a_3844_14964# vss vss nfet_06v0 w=0.82u l=1u
X1187 a_2140_13352# a_2052_13396# vss vss nfet_06v0 w=0.82u l=1u
X1188 a_2140_10216# a_2052_10260# vss vss nfet_06v0 w=0.82u l=1u
X1189 vdd a_21740_8648# a_21652_8692# vdd pfet_06v0 w=1.22u l=1u
X1190 pbusin_pshunt pseries_gy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1191 a_22076_6647# a_21988_6744# vss vss nfet_06v0 w=0.82u l=1u
X1192 nseries_gy nbusout vdd vdd pfet_06v0 w=1.22u l=0.5u
X1193 a_20060_16055# a_19972_16152# vss vss nfet_06v0 w=0.82u l=1u
X1194 nbusout pseries_gy vss vss nfet_06v0 w=0.82u l=0.6u
X1195 nbusin_nshunt pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1196 pbusin_pshunt nbusin_nshunt vss vss nfet_06v0 w=0.82u l=0.6u
X1197 vdd a_4828_10216# a_4740_10260# vdd pfet_06v0 w=1.22u l=1u
X1198 pseries_gy pseries_gygy vdd vdd pfet_06v0 w=1.22u l=0.5u
X1199 a_2140_9783# a_2052_9880# vss vss nfet_06v0 w=0.82u l=1u
X1200 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
X1201 a_10428_16055# a_10340_16152# vss vss nfet_06v0 w=0.82u l=1u
X1202 a_13452_16055# a_13364_16152# vss vss nfet_06v0 w=0.82u l=1u
X1203 a_20172_14487# a_20084_14584# vss vss nfet_06v0 w=0.82u l=1u
X1204 a_3484_12919# a_3396_13016# vss vss nfet_06v0 w=0.82u l=1u
X1205 nseries_gy pbusin_pshunt vdd vdd pfet_06v0 w=1.22u l=0.5u
C0 pseries_gy nseries_gygy 2.99fF
C1 pseries_gy pbusin_pshunt 3.33fF
C2 pbusin_pshunt nshunt_gy 4.12fF
C3 pseries_gy nbusin_nshunt 3.34fF
C4 nbusin_nshunt nshunt_gy 3.27fF
C5 nbusin_nshunt pbusin_pshunt 10.19fF
C6 vdd nseries_gy 13.55fF
C7 nseries_gy pbusout 4.01fF
C8 vdd nbusout 4.58fF
C9 nseries_gy pseries_gy 12.91fF
C10 vdd pshunt_gy 4.38fF
C11 pbusout nbusout 3.32fF
C12 vdd pseries_gygy 4.25fF
C13 nseries_gy nseries_gygy 4.21fF
C14 nseries_gy pbusin_pshunt 2.92fF
C15 nseries_gy nbusin_nshunt 4.30fF
C16 nbusout pseries_gy 3.12fF
C17 pshunt_gy nshunt_gy 6.42fF
C18 pseries_gy pseries_gygy 2.70fF
C19 nseries_gygy pseries_gygy 3.04fF
C20 pshunt_gy pbusin_pshunt 3.45fF
C21 pshunt_gy nbusin_nshunt 2.94fF
C22 vdd pbusout 4.55fF
C23 nseries_gy nbusout 3.77fF
C24 vdd pseries_gy 13.09fF
C25 vdd nshunt_gy 4.16fF
C26 vdd nseries_gygy 4.40fF
C27 vdd pbusin_pshunt 8.62fF
C28 pbusout pseries_gy 3.40fF
C29 vdd nbusin_nshunt 9.39fF
C30 nseries_gy pseries_gygy 4.58fF
C31 pseries_gygy vss 13.48fF
C32 nshunt_gy vss 12.95fF
C33 nseries_gygy vss 13.27fF
C34 pbusin_pshunt vss 25.10fF
C35 nbusin_nshunt vss 25.81fF
C36 pshunt_gy vss 13.24fF
C37 pseries_gy vss 37.10fF
C38 nbusout vss 12.47fF
C39 pbusout vss 13.01fF
C40 nseries_gy vss 38.25fF
C41 vdd vss 523.92fF
.ends

XDUT nbusin_nshunt nbusout nseries_gy nseries_gygy nshunt_gy pbusin_pshunt  pbusout pseries_gy
+ pseries_gygy pshunt_gy vss vdd filterstage_flat


**** end user architecture code
.ends


* expanding   symbol:  injector_pex.sym # of pins=14
** sym_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/injector_pex.sym
** sch_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/injector_pex.sch
.subckt injector_pex outp vdd vss outn enable signal trim_n[0] trim_n[1] trim_n[2] trim_n[3]
+ trim_p[0] trim_p[1] trim_p[2] trim_p[3]
*.ipin enable
*.ipin signal
*.ipin trim_n[0]
*.ipin trim_n[1]
*.ipin trim_n[2]
*.ipin trim_n[3]
*.ipin trim_p[0]
*.ipin trim_p[1]
*.ipin trim_p[2]
*.ipin trim_p[3]
*.iopin vss
*.iopin vdd
*.iopin outp
*.iopin outn
**** begin user architecture code

* NGSPICE file created from injector_flat.ext - technology: gf180mcuC

.subckt injector_flat enable outn outp signal trim_n[0] trim_n[1] trim_n[2] trim_n[3]  trim_p[0]
+ trim_p[1] trim_p[2] trim_p[3] vss vdd
X0 _13_ a_8301_4728# vdd vdd pfet_06v0 w=1.22u l=0.5u
X1 vdd a_9644_7080# a_9556_7124# vdd pfet_06v0 w=1.22u l=1u
X2 a_3055_3728# a_2612_3229# vdd vdd pfet_06v0 w=0.62u l=0.5u
X3 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X4 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X5 vdd trim_p[0] a_2388_7933# vdd pfet_06v0 w=0.62u l=0.5u
X6 _09_ a_6285_4728# vdd vdd pfet_06v0 w=1.22u l=0.5u
X7 vdd a_3036_5079# a_2948_5176# vdd pfet_06v0 w=1.22u l=1u
X8 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X9 a_5948_7080# a_5860_7124# vss vss nfet_06v0 w=0.82u l=1u
X10 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X11 vdd _20_ outp vdd pfet_06v0 w=1.22u l=0.5u
X12 vss trim_p[1] a_7204_7933# vss nfet_06v0 w=0.36u l=0.6u
X13 a_15496_8308# trim_p[3] vdd vdd pfet_06v0 w=0.62u l=0.5u
X14 outp _18_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X15 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X16 a_3820_5512# a_3732_5556# vss vss nfet_06v0 w=0.82u l=1u
X17 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X18 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X19 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X20 vdd a_5052_7080# a_4964_7124# vdd pfet_06v0 w=1.22u l=1u
X21 a_8573_7889# _00_ vss vss nfet_06v0 w=0.36u l=0.6u
X22 a_14703_8432# a_15496_8308# a_14723_7933# vdd pfet_06v0 w=0.62u l=0.5u
X23 a_3932_6647# a_3844_6744# vss vss nfet_06v0 w=0.82u l=1u
X24 a_7636_7675# a_7204_7156# vss vss nfet_06v0 w=0.36u l=0.6u
X25 _06_ a_14237_3944# vdd vdd pfet_06v0 w=1.22u l=0.5u
X26 vdd a_3484_5079# a_3396_5176# vdd pfet_06v0 w=1.22u l=1u
X27 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X28 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X29 vdd _15_ outn vdd pfet_06v0 w=1.22u l=0.5u
X30 a_9869_3160# a_9869_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X31 a_16280_3604# trim_n[3] vss vss nfet_06v0 w=0.36u l=0.6u
X32 a_6621_3160# a_6621_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X33 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X34 vdd _26_ a_11124_3229# vdd pfet_06v0 w=0.62u l=0.5u
X35 vdd a_2140_3944# a_2052_3988# vdd pfet_06v0 w=1.22u l=1u
X36 vdd a_3981_4417# a_3004_4020# vdd pfet_06v0 w=0.62u l=0.5u
X37 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X38 vss signal_n a_2161_6296# vss nfet_06v0 w=0.36u l=0.6u
X39 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X40 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X41 outp a_14703_8432# vdd vdd pfet_06v0 w=1.095u l=0.5u
X42 a_16280_3604# trim_n[3] vdd vdd pfet_06v0 w=0.62u l=0.5u
X43 outn a_7555_4539# vss vss nfet_06v0 w=0.82u l=0.6u
X44 a_16700_3944# a_16612_3988# vss vss nfet_06v0 w=0.82u l=1u
X45 vdd a_2140_5079# a_2052_5176# vdd pfet_06v0 w=1.22u l=1u
X46 vss a_3757_7889# a_2820_7933# vss nfet_06v0 w=0.36u l=0.6u
X47 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X48 vdd a_8573_7553# a_7596_7156# vdd pfet_06v0 w=0.62u l=0.5u
X49 a_16851_4797# a_16388_4797# vss vss nfet_06v0 w=0.36u l=0.6u
X50 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X51 a_15487_3728# a_16280_3604# a_15507_3229# vdd pfet_06v0 w=0.62u l=0.5u
X52 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X53 vdd a_3004_4020# outn vdd pfet_06v0 w=1.095u l=0.5u
X54 a_12463_3988# a_12020_4539# vdd vdd pfet_06v0 w=0.62u l=0.5u
X55 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X56 vdd a_4828_6647# a_4740_6744# vdd pfet_06v0 w=1.22u l=1u
X57 vss _22_ a_2612_3229# vss nfet_06v0 w=0.36u l=0.6u
X58 vss signal a_1924_6040# vss nfet_06v0 w=0.365u l=0.6u
X59 vss _07_ outn vss nfet_06v0 w=0.82u l=0.6u
X60 a_12360_8308# trim_p[2] vss vss nfet_06v0 w=0.36u l=0.6u
X61 _10_ a_10093_3944# vdd vdd pfet_06v0 w=1.22u l=0.5u
X62 vdd a_6060_8215# a_5972_8312# vdd pfet_06v0 w=1.22u l=1u
X63 _03_ a_1716_6040# vdd vdd pfet_06v0 w=1.215u l=0.5u
X64 a_12780_5079# a_12692_5176# vss vss nfet_06v0 w=0.82u l=1u
X65 vdd a_17932_8215# a_17844_8312# vdd pfet_06v0 w=1.22u l=1u
X66 _03_ a_1716_6040# vss vss nfet_06v0 w=0.815u l=0.6u
X67 vdd a_8573_7889# a_7596_8400# vdd pfet_06v0 w=0.62u l=0.5u
X68 a_7667_3229# trim_n[1] a_7647_3728# vss nfet_06v0 w=0.36u l=0.6u
X69 a_10541_3160# a_10541_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X70 a_4268_5512# a_4180_5556# vss vss nfet_06v0 w=0.82u l=1u
X71 outn _09_ vss vss nfet_06v0 w=0.82u l=0.6u
X72 a_12483_4539# a_12020_4539# vss vss nfet_06v0 w=0.36u l=0.6u
X73 a_7667_3229# a_7204_3229# vss vss nfet_06v0 w=0.36u l=0.6u
X74 vss _25_ a_12020_4539# vss nfet_06v0 w=0.36u l=0.6u
X75 a_3004_4020# trim_n[0] vdd vdd pfet_06v0 w=0.62u l=0.5u
X76 a_1692_6647# a_1604_6744# vss vss nfet_06v0 w=0.82u l=1u
X77 vss trim_p[2] a_12020_7156# vss nfet_06v0 w=0.36u l=0.6u
X78 vss a_16280_3604# a_15507_3229# vss nfet_06v0 w=0.36u l=0.6u
X79 a_3055_3728# a_3848_3604# a_3075_3229# vdd pfet_06v0 w=0.62u l=0.5u
X80 _28_ a_5501_5512# vdd vdd pfet_06v0 w=1.22u l=0.5u
X81 vss _00_ outn vss nfet_06v0 w=0.82u l=0.6u
X82 a_8189_5512# a_8189_5512# vss vss nfet_06v0 w=0.82u l=0.6u
X83 a_3757_7889# _00_ vss vss nfet_06v0 w=0.36u l=0.6u
X84 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X85 a_8573_7553# _00_ vdd vdd pfet_06v0 w=0.62u l=0.5u
X86 a_2161_6296# _00_ vss vss nfet_06v0 w=0.36u l=0.6u
X87 outn a_14835_7675# vss vss nfet_06v0 w=0.82u l=0.6u
X88 a_6844_7080# a_6756_7124# vss vss nfet_06v0 w=0.82u l=1u
X89 vdd a_9644_3944# a_9556_3988# vdd pfet_06v0 w=1.22u l=1u
X90 vdd a_4716_5512# a_4628_5556# vdd pfet_06v0 w=1.22u l=1u
X91 a_5612_6647# a_5524_6744# vss vss nfet_06v0 w=0.82u l=1u
X92 a_14815_7124# a_15608_7112# a_14835_7675# vdd pfet_06v0 w=0.62u l=0.5u
X93 a_7596_7156# trim_p[1] a_7636_7675# vss nfet_06v0 w=0.36u l=0.6u
X94 vss _00_ outn vss nfet_06v0 w=0.82u l=0.6u
X95 vdd a_3932_6647# a_3844_6744# vdd pfet_06v0 w=1.22u l=1u
X96 vss a_2820_7675# outp vss nfet_06v0 w=0.82u l=0.6u
X97 vdd trim_n[1] a_7535_3988# vdd pfet_06v0 w=0.62u l=0.5u
X98 vdd signal a_1716_6040# vdd pfet_06v0 w=0.6u l=0.5u
X99 a_12412_7156# trim_p[2] a_12452_7675# vss nfet_06v0 w=0.36u l=0.6u
X100 _05_ a_9869_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X101 _25_ a_6621_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X102 a_16831_5296# a_17624_5172# a_16851_4797# vdd pfet_06v0 w=0.62u l=0.5u
X103 vdd a_7596_7156# outn vdd pfet_06v0 w=1.095u l=0.5u
X104 vss a_17699_6040# a_17699_6040# vss nfet_06v0 w=0.82u l=0.6u
X105 vdd trim_n[1] a_7647_3728# vdd pfet_06v0 w=0.62u l=0.5u
X106 a_2780_7156# trim_p[0] vdd vdd pfet_06v0 w=0.62u l=0.5u
X107 vdd _00_ outp vdd pfet_06v0 w=1.22u l=0.5u
X108 vdd a_14012_7080# a_13924_7124# vdd pfet_06v0 w=1.22u l=1u
X109 a_5500_7080# a_5412_7124# vss vss nfet_06v0 w=0.82u l=1u
X110 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X111 a_8573_7889# _00_ vdd vdd pfet_06v0 w=0.62u l=0.5u
X112 vdd a_3296_6296# _02_ vdd pfet_06v0 w=1.22u l=0.5u
X113 a_3372_5512# a_3284_5556# vss vss nfet_06v0 w=0.82u l=1u
X114 vss a_12360_8308# a_11587_7933# vss nfet_06v0 w=0.36u l=0.6u
X115 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X116 a_2820_7933# a_2388_7933# a_2780_8400# vdd pfet_06v0 w=0.62u l=0.5u
X117 a_5612_8215# a_5524_8312# vss vss nfet_06v0 w=0.82u l=1u
X118 a_2161_6296# signal_n a_2553_6875# vdd pfet_06v0 w=0.565u l=0.5u
X119 a_11587_3229# a_11124_3229# vss vss nfet_06v0 w=0.36u l=0.6u
X120 vdd trim_n[0] a_3055_3728# vdd pfet_06v0 w=0.62u l=0.5u
X121 vdd signal signal_n vdd pfet_06v0 w=1.22u l=0.5u
X122 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X123 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X124 a_15507_3229# trim_n[3] a_15487_3728# vss nfet_06v0 w=0.36u l=0.6u
X125 vss a_2820_7933# outn vss nfet_06v0 w=0.82u l=0.6u
X126 outp _10_ vss vss nfet_06v0 w=0.82u l=0.6u
X127 vdd a_3820_5512# a_3732_5556# vdd pfet_06v0 w=1.22u l=1u
X128 outp _06_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X129 vdd a_7596_8400# outp vdd pfet_06v0 w=1.095u l=0.5u
X130 a_14237_3160# a_14237_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X131 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X132 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X133 a_3296_6296# _03_ vss vss nfet_06v0 w=0.36u l=0.6u
X134 a_16831_5296# a_16388_4797# vdd vdd pfet_06v0 w=0.62u l=0.5u
X135 outn _05_ vss vss nfet_06v0 w=0.82u l=0.6u
X136 vdd a_6947_4772# _11_ vdd pfet_06v0 w=1.22u l=0.5u
X137 outp _12_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X138 outn a_12483_4539# vss vss nfet_06v0 w=0.82u l=0.6u
X139 _16_ a_10541_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X140 a_4829_4728# a_4829_4728# vss vss nfet_06v0 w=0.82u l=0.6u
X141 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X142 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X143 a_7647_3728# a_7204_3229# vdd vdd pfet_06v0 w=0.62u l=0.5u
X144 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X145 a_12452_7675# a_12020_7156# vss vss nfet_06v0 w=0.36u l=0.6u
X146 vdd trim_n[2] a_11567_3728# vdd pfet_06v0 w=0.62u l=0.5u
X147 vdd a_1692_6647# a_1604_6744# vdd pfet_06v0 w=1.22u l=1u
X148 vdd _00_ outp vdd pfet_06v0 w=1.22u l=0.5u
X149 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X150 a_3757_7553# _00_ vdd vdd pfet_06v0 w=0.62u l=0.5u
X151 vdd _07_ outn vdd pfet_06v0 w=1.22u l=0.5u
X152 a_12668_6647# a_12580_6744# vss vss nfet_06v0 w=0.82u l=1u
X153 vdd a_12780_5079# a_12692_5176# vdd pfet_06v0 w=1.22u l=1u
X154 vdd _27_ a_15044_3229# vdd pfet_06v0 w=0.62u l=0.5u
X155 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X156 vdd a_16700_3944# a_16612_3988# vdd pfet_06v0 w=1.22u l=1u
X157 vdd a_5612_6647# a_5524_6744# vdd pfet_06v0 w=1.22u l=1u
X158 a_11587_7933# trim_p[2] a_11567_8432# vss nfet_06v0 w=0.36u l=0.6u
X159 a_9644_5512# a_9556_5556# vss vss nfet_06v0 w=0.82u l=1u
X160 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X161 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X162 a_5837_3944# a_5837_3944# vss vss nfet_06v0 w=0.82u l=0.6u
X163 vss _28_ a_16388_4797# vss nfet_06v0 w=0.36u l=0.6u
X164 a_2780_8400# trim_p[0] a_2820_7933# vss nfet_06v0 w=0.36u l=0.6u
X165 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X166 vdd a_6835_6340# _15_ vdd pfet_06v0 w=1.22u l=0.5u
X167 a_6509_3944# a_6509_3944# vss vss nfet_06v0 w=0.82u l=0.6u
X168 a_3757_7889# _00_ vdd vdd pfet_06v0 w=0.62u l=0.5u
X169 a_1716_6040# enable vdd vdd pfet_06v0 w=0.6u l=0.5u
X170 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X171 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X172 outp _08_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X173 a_16365_5512# a_16365_5512# vss vss nfet_06v0 w=0.82u l=0.6u
X174 a_14723_7933# trim_p[3] a_14703_8432# vss nfet_06v0 w=0.36u l=0.6u
X175 a_6396_7080# a_6308_7124# vss vss nfet_06v0 w=0.82u l=1u
X176 a_11567_3728# a_11124_3229# vdd vdd pfet_06v0 w=0.62u l=0.5u
X177 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X178 a_4640_7864# _04_ vss vss nfet_06v0 w=0.36u l=0.6u
X179 vdd a_4268_5512# a_4180_5556# vdd pfet_06v0 w=1.22u l=1u
X180 a_9644_7080# a_9556_7124# vss vss nfet_06v0 w=0.82u l=1u
X181 vss a_17475_3204# a_17475_3204# vss nfet_06v0 w=0.82u l=0.6u
X182 vss trim_p[1] a_7204_7156# vss nfet_06v0 w=0.36u l=0.6u
X183 a_3981_4417# _21_ vdd vdd pfet_06v0 w=0.62u l=0.5u
X184 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X185 vss a_7636_7675# outn vss nfet_06v0 w=0.82u l=0.6u
X186 vdd trim_n[2] a_12463_3988# vdd pfet_06v0 w=0.62u l=0.5u
X187 outn _17_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X188 outn _17_ vss vss nfet_06v0 w=0.82u l=0.6u
X189 a_8573_7553# _00_ vss vss nfet_06v0 w=0.36u l=0.6u
X190 a_7596_7156# trim_p[1] vdd vdd pfet_06v0 w=0.62u l=0.5u
X191 vdd _00_ outp vdd pfet_06v0 w=1.22u l=0.5u
X192 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X193 vdd _00_ outn vdd pfet_06v0 w=1.22u l=0.5u
X194 _08_ a_8189_5512# vdd vdd pfet_06v0 w=1.22u l=0.5u
X195 a_4380_6647# a_4292_6744# vss vss nfet_06v0 w=0.82u l=1u
X196 _18_ a_14237_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X197 outp _16_ vss vss nfet_06v0 w=0.82u l=0.6u
X198 a_12412_7156# trim_p[2] vdd vdd pfet_06v0 w=0.62u l=0.5u
X199 a_5052_7080# a_4964_7124# vss vss nfet_06v0 w=0.82u l=1u
X200 a_15496_8308# trim_p[3] vss vss nfet_06v0 w=0.36u l=0.6u
X201 vss a_2161_6296# _04_ vss nfet_06v0 w=0.82u l=0.6u
X202 a_16812_5512# a_16724_5556# vss vss nfet_06v0 w=0.82u l=1u
X203 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X204 a_13389_7553# _00_ vdd vdd pfet_06v0 w=0.62u l=0.5u
X205 vdd _00_ outn vdd pfet_06v0 w=1.22u l=0.5u
X206 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X207 a_3981_4417# _21_ vss vss nfet_06v0 w=0.36u l=0.6u
X208 a_7636_7933# a_7204_7933# a_7596_8400# vdd pfet_06v0 w=0.62u l=0.5u
X209 a_7535_3988# a_8328_3976# a_7555_4539# vdd pfet_06v0 w=0.62u l=0.5u
X210 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X211 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X212 vss _23_ a_7092_4539# vss nfet_06v0 w=0.36u l=0.6u
X213 vdd trim_p[1] a_7204_7933# vdd pfet_06v0 w=0.62u l=0.5u
X214 vdd _00_ a_11124_7933# vdd pfet_06v0 w=0.62u l=0.5u
X215 a_8328_3976# trim_n[1] vss vss nfet_06v0 w=0.36u l=0.6u
X216 vss a_3757_7553# a_2820_7675# vss nfet_06v0 w=0.36u l=0.6u
X217 a_2820_7933# a_2388_7933# vss vss nfet_06v0 w=0.36u l=0.6u
X218 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X219 vdd trim_p[0] a_2388_7156# vdd pfet_06v0 w=0.62u l=0.5u
X220 vdd trim_p[2] a_11567_8432# vdd pfet_06v0 w=0.62u l=0.5u
X221 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X222 vss a_7636_7933# outp vss nfet_06v0 w=0.82u l=0.6u
X223 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X224 vdd a_3372_5512# a_3284_5556# vdd pfet_06v0 w=1.22u l=1u
X225 outp a_7647_3728# vdd vdd pfet_06v0 w=1.095u l=0.5u
X226 vss _11_ outn vss nfet_06v0 w=0.82u l=0.6u
X227 vdd a_12668_6647# a_12580_6744# vdd pfet_06v0 w=1.22u l=1u
X228 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X229 vss _00_ a_14372_7675# vss nfet_06v0 w=0.36u l=0.6u
X230 _17_ a_4829_4728# vdd vdd pfet_06v0 w=1.22u l=0.5u
X231 _00_ enable vdd vdd pfet_06v0 w=1.22u l=0.5u
X232 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X233 vdd a_15683_4772# _14_ vdd pfet_06v0 w=1.22u l=0.5u
X234 vss _26_ a_11124_3229# vss nfet_06v0 w=0.36u l=0.6u
X235 outp a_7667_3229# vss vss nfet_06v0 w=0.82u l=0.6u
X236 vdd _00_ a_14260_7933# vdd pfet_06v0 w=0.62u l=0.5u
X237 vdd _25_ a_12020_4539# vdd pfet_06v0 w=0.62u l=0.5u
X238 outp a_3055_3728# vdd vdd pfet_06v0 w=1.095u l=0.5u
X239 a_15507_3229# a_15044_3229# vss vss nfet_06v0 w=0.36u l=0.6u
X240 vdd trim_p[3] a_14703_8432# vdd pfet_06v0 w=0.62u l=0.5u
X241 vss a_15496_8308# a_14723_7933# vss nfet_06v0 w=0.36u l=0.6u
X242 outp a_3075_3229# vss vss nfet_06v0 w=0.82u l=0.6u
X243 vss a_8573_7889# a_7636_7933# vss nfet_06v0 w=0.36u l=0.6u
X244 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X245 a_3757_7553# _00_ vss vss nfet_06v0 w=0.36u l=0.6u
X246 vdd _23_ a_7092_4539# vdd pfet_06v0 w=0.62u l=0.5u
X247 outp a_16831_5296# vdd vdd pfet_06v0 w=1.095u l=0.5u
X248 vss trim_p[0] a_2388_7933# vss nfet_06v0 w=0.36u l=0.6u
X249 a_6060_6647# a_5972_6744# vss vss nfet_06v0 w=0.82u l=1u
X250 outp a_11567_3728# vdd vdd pfet_06v0 w=1.095u l=0.5u
X251 a_14684_3511# a_14596_3608# vss vss nfet_06v0 w=0.82u l=1u
X252 vdd a_4380_6647# a_4292_6744# vdd pfet_06v0 w=1.22u l=1u
X253 a_3075_3229# trim_n[0] a_3055_3728# vss nfet_06v0 w=0.36u l=0.6u
X254 a_17932_3511# a_17844_3608# vss vss nfet_06v0 w=0.82u l=1u
X255 a_4604_3944# a_4516_3988# vss vss nfet_06v0 w=0.82u l=1u
X256 vdd trim_n[3] a_15487_3728# vdd pfet_06v0 w=0.62u l=0.5u
X257 outn _13_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X258 vdd a_9644_5512# a_9556_5556# vdd pfet_06v0 w=1.22u l=1u
X259 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X260 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X261 _23_ a_5837_3944# vdd vdd pfet_06v0 w=1.22u l=0.5u
X262 a_11587_7933# a_11124_7933# vss vss nfet_06v0 w=0.36u l=0.6u
X263 outn _19_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X264 outp a_11587_3229# vss vss nfet_06v0 w=0.82u l=0.6u
X265 outn a_15487_3728# vdd vdd pfet_06v0 w=1.095u l=0.5u
X266 vdd a_5948_7080# a_5860_7124# vdd pfet_06v0 w=1.22u l=1u
X267 a_4157_4728# a_4157_4728# vss vss nfet_06v0 w=0.82u l=0.6u
X268 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X269 vss a_3981_4417# a_3044_4539# vss nfet_06v0 w=0.36u l=0.6u
X270 vdd a_17699_6040# _20_ vdd pfet_06v0 w=1.22u l=0.5u
X271 _19_ a_6509_3944# vdd vdd pfet_06v0 w=1.22u l=0.5u
X272 outp _18_ vss vss nfet_06v0 w=0.82u l=0.6u
X273 a_14012_7080# a_13924_7124# vss vss nfet_06v0 w=0.82u l=1u
X274 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X275 a_6060_8215# a_5972_8312# vss vss nfet_06v0 w=0.82u l=1u
X276 vdd a_3757_7553# a_2780_7156# vdd pfet_06v0 w=0.62u l=0.5u
X277 vss a_3044_4539# outn vss nfet_06v0 w=0.82u l=0.6u
X278 a_17932_8215# a_17844_8312# vss vss nfet_06v0 w=0.82u l=1u
X279 _12_ a_16365_5512# vdd vdd pfet_06v0 w=1.22u l=0.5u
X280 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X281 vss signal signal_n vss nfet_06v0 w=0.82u l=0.6u
X282 outn a_11587_7933# vss vss nfet_06v0 w=0.82u l=0.6u
X283 a_14723_7933# a_14260_7933# vss vss nfet_06v0 w=0.36u l=0.6u
X284 a_12463_3988# a_13256_3976# a_12483_4539# vdd pfet_06v0 w=0.62u l=0.5u
X285 vdd _22_ a_2612_3229# vdd pfet_06v0 w=0.62u l=0.5u
X286 a_5165_3944# a_5165_3944# vss vss nfet_06v0 w=0.82u l=0.6u
X287 a_7636_7933# a_7204_7933# vss vss nfet_06v0 w=0.36u l=0.6u
X288 vdd _00_ a_14372_7675# vdd pfet_06v0 w=0.62u l=0.5u
X289 vdd trim_n[0] a_2612_4020# vdd pfet_06v0 w=0.62u l=0.5u
X290 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X291 vss a_12452_7675# outp vss nfet_06v0 w=0.82u l=0.6u
X292 vss _24_ a_7204_3229# vss nfet_06v0 w=0.36u l=0.6u
X293 a_2588_5079# a_2500_5176# vss vss nfet_06v0 w=0.82u l=1u
X294 outp _10_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X295 a_7555_4539# trim_n[1] a_7535_3988# vss nfet_06v0 w=0.36u l=0.6u
X296 a_15487_3728# a_15044_3229# vdd vdd pfet_06v0 w=0.62u l=0.5u
X297 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X298 a_13389_7553# _00_ vss vss nfet_06v0 w=0.36u l=0.6u
X299 outn a_11567_8432# vdd vdd pfet_06v0 w=1.095u l=0.5u
X300 a_13256_3976# trim_n[2] vss vss nfet_06v0 w=0.36u l=0.6u
X301 a_8440_3604# trim_n[1] vss vss nfet_06v0 w=0.36u l=0.6u
X302 a_1692_3944# a_1604_3988# vss vss nfet_06v0 w=0.82u l=1u
X303 vdd trim_p[2] a_12020_7156# vdd pfet_06v0 w=0.62u l=0.5u
X304 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X305 vdd a_3757_7889# a_2780_8400# vdd pfet_06v0 w=0.62u l=0.5u
X306 a_8328_3976# trim_n[1] vdd vdd pfet_06v0 w=0.62u l=0.5u
X307 vdd a_16812_5512# a_16724_5556# vdd pfet_06v0 w=1.22u l=1u
X308 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X309 vss a_6947_4772# a_6947_4772# vss nfet_06v0 w=0.82u l=0.6u
X310 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X311 a_4829_3160# a_4829_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X312 vdd trim_n[3] a_16831_5296# vdd pfet_06v0 w=0.62u l=0.5u
X313 a_8440_3604# trim_n[1] vdd vdd pfet_06v0 w=0.62u l=0.5u
X314 a_2820_7675# a_2388_7156# a_2780_7156# vdd pfet_06v0 w=0.62u l=0.5u
X315 vss _14_ outp vss nfet_06v0 w=0.82u l=0.6u
X316 a_3848_3604# trim_n[0] vss vss nfet_06v0 w=0.36u l=0.6u
X317 vss a_17624_5172# a_16851_4797# vss nfet_06v0 w=0.36u l=0.6u
X318 a_14835_7675# trim_p[3] a_14815_7124# vss nfet_06v0 w=0.36u l=0.6u
X319 outp _06_ vss vss nfet_06v0 w=0.82u l=0.6u
X320 vss _00_ outp vss nfet_06v0 w=0.82u l=0.6u
X321 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X322 vdd a_6060_6647# a_5972_6744# vdd pfet_06v0 w=1.22u l=1u
X323 vdd a_14684_3511# a_14596_3608# vdd pfet_06v0 w=1.22u l=1u
X324 a_7647_3728# a_8440_3604# a_7667_3229# vdd pfet_06v0 w=0.62u l=0.5u
X325 vdd a_17932_3511# a_17844_3608# vdd pfet_06v0 w=1.22u l=1u
X326 vdd _11_ outn vdd pfet_06v0 w=1.22u l=0.5u
X327 outp _08_ vss vss nfet_06v0 w=0.82u l=0.6u
X328 a_3044_4539# a_2612_4020# vss vss nfet_06v0 w=0.36u l=0.6u
X329 a_2780_7156# trim_p[0] a_2820_7675# vss nfet_06v0 w=0.36u l=0.6u
X330 vdd a_5612_8215# a_5524_8312# vdd pfet_06v0 w=1.22u l=1u
X331 a_3848_3604# trim_n[0] vdd vdd pfet_06v0 w=0.62u l=0.5u
X332 outp _12_ vss vss nfet_06v0 w=0.82u l=0.6u
X333 a_14815_7124# a_14372_7675# vdd vdd pfet_06v0 w=0.62u l=0.5u
X334 a_2780_8400# trim_p[0] vdd vdd pfet_06v0 w=0.62u l=0.5u
X335 a_1692_5079# a_1604_5176# vss vss nfet_06v0 w=0.82u l=1u
X336 a_2553_6875# _00_ vdd vdd pfet_06v0 w=0.565u l=0.5u
X337 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X338 a_15608_7112# trim_p[3] vss vss nfet_06v0 w=0.36u l=0.6u
X339 vdd a_2780_7156# outp vdd pfet_06v0 w=1.095u l=0.5u
X340 a_5949_3160# a_5949_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X341 a_12360_3604# trim_n[2] vss vss nfet_06v0 w=0.36u l=0.6u
X342 outn a_7535_3988# vdd vdd pfet_06v0 w=1.095u l=0.5u
X343 a_15608_7112# trim_p[3] vdd vdd pfet_06v0 w=0.62u l=0.5u
X344 outp a_16851_4797# vss vss nfet_06v0 w=0.82u l=0.6u
X345 a_1924_6040# enable a_1716_6040# vss nfet_06v0 w=0.365u l=0.6u
X346 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X347 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X348 a_5612_5079# a_5524_5176# vss vss nfet_06v0 w=0.82u l=1u
X349 vdd a_6844_7080# a_6756_7124# vdd pfet_06v0 w=1.22u l=1u
X350 vss a_13256_3976# a_12483_4539# vss nfet_06v0 w=0.36u l=0.6u
X351 vss a_8440_3604# a_7667_3229# vss nfet_06v0 w=0.36u l=0.6u
X352 vss _27_ a_15044_3229# vss nfet_06v0 w=0.36u l=0.6u
X353 a_17624_5172# trim_n[3] vdd vdd pfet_06v0 w=0.62u l=0.5u
X354 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X355 a_8301_4728# a_8301_4728# vss vss nfet_06v0 w=0.82u l=0.6u
X356 a_14237_3944# a_14237_3944# vss vss nfet_06v0 w=0.82u l=0.6u
X357 a_11567_8432# a_11124_7933# vdd vdd pfet_06v0 w=0.62u l=0.5u
X358 vss _15_ outn vss nfet_06v0 w=0.82u l=0.6u
X359 a_12360_3604# trim_n[2] vdd vdd pfet_06v0 w=0.62u l=0.5u
X360 a_6285_4728# a_6285_4728# vss vss nfet_06v0 w=0.82u l=0.6u
X361 a_3036_5079# a_2948_5176# vss vss nfet_06v0 w=0.82u l=1u
X362 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X363 outn _09_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X364 outp _01_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X365 a_2140_3944# a_2052_3988# vss vss nfet_06v0 w=0.82u l=1u
X366 vss _00_ outp vss nfet_06v0 w=0.82u l=0.6u
X367 vss a_6835_6340# a_6835_6340# vss nfet_06v0 w=0.82u l=0.6u
X368 a_7596_8400# trim_p[1] a_7636_7933# vss nfet_06v0 w=0.36u l=0.6u
X369 _21_ a_4157_4728# vdd vdd pfet_06v0 w=1.22u l=0.5u
X370 vdd a_2780_8400# outn vdd pfet_06v0 w=1.095u l=0.5u
X371 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X372 a_11567_3728# a_12360_3604# a_11587_3229# vdd pfet_06v0 w=0.62u l=0.5u
X373 vss a_3848_3604# a_3075_3229# vss nfet_06v0 w=0.36u l=0.6u
X374 a_16851_4797# trim_n[3] a_16831_5296# vss nfet_06v0 w=0.36u l=0.6u
X375 vss a_8328_3976# a_7555_4539# vss nfet_06v0 w=0.36u l=0.6u
X376 vdd a_5500_7080# a_5412_7124# vdd pfet_06v0 w=1.22u l=1u
X377 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X378 a_2029_3160# a_2029_3160# vss vss nfet_06v0 w=0.82u l=0.6u
X379 outn _02_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X380 outn _02_ vss vss nfet_06v0 w=0.82u l=0.6u
X381 vdd a_4604_3944# a_4516_3988# vdd pfet_06v0 w=1.22u l=1u
X382 outp _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X383 vss trim_n[0] a_2612_4020# vss nfet_06v0 w=0.36u l=0.6u
X384 outn _00_ vss vss nfet_06v0 w=0.82u l=0.6u
X385 a_3484_5079# a_3396_5176# vss vss nfet_06v0 w=0.82u l=1u
X386 a_2820_7675# a_2388_7156# vss vss nfet_06v0 w=0.36u l=0.6u
X387 _00_ enable vss vss nfet_06v0 w=0.82u l=0.6u
X388 vdd a_13389_7553# a_12412_7156# vdd pfet_06v0 w=0.62u l=0.5u
X389 vdd a_4640_7864# _01_ vdd pfet_06v0 w=1.22u l=0.5u
X390 outp _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X391 a_3075_3229# a_2612_3229# vss vss nfet_06v0 w=0.36u l=0.6u
X392 _24_ a_4829_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X393 a_14703_8432# a_14260_7933# vdd vdd pfet_06v0 w=0.62u l=0.5u
X394 outn _00_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X395 vss _20_ outp vss nfet_06v0 w=0.82u l=0.6u
X396 vss _00_ a_11124_7933# vss nfet_06v0 w=0.36u l=0.6u
X397 a_3296_6296# _03_ vdd vdd pfet_06v0 w=0.565u l=0.5u
X398 vss a_15608_7112# a_14835_7675# vss nfet_06v0 w=0.36u l=0.6u
X399 vdd a_2588_5079# a_2500_5176# vdd pfet_06v0 w=1.22u l=1u
X400 a_10093_3944# a_10093_3944# vss vss nfet_06v0 w=0.82u l=0.6u
X401 vss a_12360_3604# a_11587_3229# vss nfet_06v0 w=0.36u l=0.6u
X402 outn a_15507_3229# vss vss nfet_06v0 w=0.82u l=0.6u
X403 vdd a_12412_7156# outp vdd pfet_06v0 w=1.095u l=0.5u
X404 a_12483_4539# trim_n[2] a_12463_3988# vss nfet_06v0 w=0.36u l=0.6u
X405 a_2140_5079# a_2052_5176# vss vss nfet_06v0 w=0.82u l=1u
X406 a_7535_3988# a_7092_4539# vdd vdd pfet_06v0 w=0.62u l=0.5u
X407 a_13256_3976# trim_n[2] vdd vdd pfet_06v0 w=0.62u l=0.5u
X408 vss a_15683_4772# a_15683_4772# vss nfet_06v0 w=0.82u l=0.6u
X409 outp _01_ vss vss nfet_06v0 w=0.82u l=0.6u
X410 _27_ a_5165_3944# vdd vdd pfet_06v0 w=1.22u l=0.5u
X411 vdd _14_ outp vdd pfet_06v0 w=1.22u l=0.5u
X412 a_5501_5512# a_5501_5512# vss vss nfet_06v0 w=0.82u l=0.6u
X413 a_7636_7675# a_7204_7156# a_7596_7156# vdd pfet_06v0 w=0.62u l=0.5u
X414 vss _00_ a_14260_7933# vss nfet_06v0 w=0.36u l=0.6u
X415 vss _00_ outp vss nfet_06v0 w=0.82u l=0.6u
X416 a_12452_7675# a_12020_7156# a_12412_7156# vdd pfet_06v0 w=0.62u l=0.5u
X417 _26_ a_5949_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X418 vdd trim_p[1] a_7204_7156# vdd pfet_06v0 w=0.62u l=0.5u
X419 vss a_8573_7553# a_7636_7675# vss nfet_06v0 w=0.36u l=0.6u
X420 vss a_3296_6296# _02_ vss nfet_06v0 w=0.82u l=0.6u
X421 vdd a_1692_3944# a_1604_3988# vdd pfet_06v0 w=1.22u l=1u
X422 vss a_13389_7553# a_12452_7675# vss nfet_06v0 w=0.36u l=0.6u
X423 a_9644_3944# a_9556_3988# vss vss nfet_06v0 w=0.82u l=1u
X424 a_4716_5512# a_4628_5556# vss vss nfet_06v0 w=0.82u l=1u
X425 a_7555_4539# a_7092_4539# vss vss nfet_06v0 w=0.36u l=0.6u
X426 vdd _28_ a_16388_4797# vdd pfet_06v0 w=0.62u l=0.5u
X427 vdd trim_p[3] a_14815_7124# vdd pfet_06v0 w=0.62u l=0.5u
X428 vss trim_p[0] a_2388_7156# vss nfet_06v0 w=0.36u l=0.6u
X429 outn _05_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X430 a_7596_8400# trim_p[1] vdd vdd pfet_06v0 w=0.62u l=0.5u
X431 vss a_4640_7864# _01_ vss nfet_06v0 w=0.82u l=0.6u
X432 outn _19_ vss vss nfet_06v0 w=0.82u l=0.6u
X433 vdd a_17475_3204# _07_ vdd pfet_06v0 w=1.22u l=0.5u
X434 a_17624_5172# trim_n[3] vss vss nfet_06v0 w=0.36u l=0.6u
X435 vdd a_1692_5079# a_1604_5176# vdd pfet_06v0 w=1.22u l=1u
X436 a_4828_6647# a_4740_6744# vss vss nfet_06v0 w=0.82u l=1u
X437 a_12360_8308# trim_p[2] vdd vdd pfet_06v0 w=0.62u l=0.5u
X438 outn a_14815_7124# vdd vdd pfet_06v0 w=1.095u l=0.5u
X439 vdd _24_ a_7204_3229# vdd pfet_06v0 w=0.62u l=0.5u
X440 outp a_14723_7933# vss vss nfet_06v0 w=0.82u l=0.6u
X441 a_3004_4020# trim_n[0] a_3044_4539# vss nfet_06v0 w=0.36u l=0.6u
X442 a_4640_7864# _04_ vdd vdd pfet_06v0 w=0.565u l=0.5u
X443 a_11567_8432# a_12360_8308# a_11587_7933# vdd pfet_06v0 w=0.62u l=0.5u
X444 _22_ a_2029_3160# vdd vdd pfet_06v0 w=1.22u l=0.5u
X445 outp _16_ vdd vdd pfet_06v0 w=1.22u l=0.5u
X446 outn a_12463_3988# vdd vdd pfet_06v0 w=1.095u l=0.5u
X447 outn _13_ vss vss nfet_06v0 w=0.82u l=0.6u
X448 vdd a_5612_5079# a_5524_5176# vdd pfet_06v0 w=1.22u l=1u
X449 a_14835_7675# a_14372_7675# vss vss nfet_06v0 w=0.36u l=0.6u
X450 a_11587_3229# trim_n[2] a_11567_3728# vss nfet_06v0 w=0.36u l=0.6u
X451 a_3044_4539# a_2612_4020# a_3004_4020# vdd pfet_06v0 w=0.62u l=0.5u
X452 vdd a_2161_6296# _04_ vdd pfet_06v0 w=1.22u l=0.5u
X453 vdd a_6396_7080# a_6308_7124# vdd pfet_06v0 w=1.22u l=1u
C0 _27_ _07_ 2.90fF
C1 outp vdd 5.81fF
C2 _10_ _19_ 3.02fF
C3 outn vdd 5.93fF
C4 _00_ vdd 3.45fF
C5 _00_ _17_ 2.81fF
C6 _08_ outn 3.45fF
C7 outp outn 5.06fF
C8 _00_ outp 6.12fF
C9 _28_ outn 2.17fF
C10 _00_ _28_ 2.35fF
C11 _16_ _00_ 2.42fF
C12 _00_ outn 6.24fF
C13 trim_n[2] vss 2.73fF
C14 trim_n[1] vss 2.75fF
C15 trim_n[0] vss 2.69fF
C16 trim_n[3] vss 2.90fF
C17 trim_p[3] vss 2.63fF
C18 trim_p[2] vss 2.71fF
C19 trim_p[1] vss 2.58fF
C20 outn vss 7.10fF
C21 trim_p[0] vss 2.57fF
C22 outp vss 7.76fF
C23 vdd vss 178.33fF
C24 _00_ vss 22.42fF $ **FLOATING
.ends



XDUT enable outn outp signal trim_n[0] trim_n[1] trim_n[2] trim_n[3]  trim_p[0] trim_p[1] trim_p[2]
+ trim_p[3] vss vdd injector_flat


**** end user architecture code
.ends


* expanding   symbol:  active_load_pex.sym # of pins=9
** sym_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/active_load_pex.sym
** sch_path: /home/andylithia/openmpw/Project-Futo-Chip1/xschem/active_load_pex.sch
.subckt active_load_pex vdd vss outpn pbus nbus outnn outp outxor outn
*.iopin vdd
*.iopin vss
*.iopin pbus
*.iopin nbus
*.iopin outp
*.iopin outn
*.opin outpn
*.opin outnn
*.opin outxor
**** begin user architecture code

* NGSPICE file created from active_load_flat.ext - technology: gf180mcuC

.subckt active_load_flat nbus outn outnn outp outpn outxor pbus vdd vss
X0 vss outn outp vss nfet_06v0 w=0.82u l=0.6u
X1 pbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X2 outp nbus vss vss nfet_06v0 w=0.82u l=0.6u
X3 vdd a_8300_8215# a_8212_8312# vdd pfet_06v0 w=1.22u l=1u
X4 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X5 vdd a_7068_7080# a_6980_7124# vdd pfet_06v0 w=1.22u l=1u
X6 vdd a_9532_8215# a_9444_8312# vdd pfet_06v0 w=1.22u l=1u
X7 pbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X8 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X9 vdd a_8860_7080# a_8772_7124# vdd pfet_06v0 w=1.22u l=1u
X10 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X11 outxor a_9016_6876# vss vss nfet_06v0 w=0.82u l=0.6u
X12 outn outn vss vss nfet_06v0 w=0.82u l=0.6u
X13 vdd a_8748_5079# a_8660_5176# vdd pfet_06v0 w=1.22u l=1u
X14 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X15 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X16 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X17 outp nbus vss vss nfet_06v0 w=0.82u l=0.6u
X18 vdd a_9980_8215# a_9892_8312# vdd pfet_06v0 w=1.22u l=1u
X19 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X20 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X21 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X22 pbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X23 a_6956_5512# a_6868_5556# vss vss nfet_06v0 w=0.82u l=1u
X24 nbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X25 vdd outn outn vdd pfet_06v0 w=1.22u l=0.5u
X26 a_6172_5079# a_6084_5176# vss vss nfet_06v0 w=0.82u l=1u
X27 vdd a_6060_8215# a_5972_8312# vdd pfet_06v0 w=1.22u l=1u
X28 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X29 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X30 a_1692_7080# a_1604_7124# vss vss nfet_06v0 w=0.82u l=1u
X31 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X32 a_6508_8215# a_6420_8312# vss vss nfet_06v0 w=0.82u l=1u
X33 nbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X34 a_9912_6340# outpn outxor vss nfet_06v0 w=0.82u l=0.6u
X35 pbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X36 vdd outn outnn vdd pfet_06v0 w=1.22u l=0.5u
X37 a_6956_8215# a_6868_8312# vss vss nfet_06v0 w=0.82u l=1u
X38 a_7516_7080# a_7428_7124# vss vss nfet_06v0 w=0.82u l=1u
X39 a_1692_8215# a_1604_8312# vss vss nfet_06v0 w=0.82u l=1u
X40 vdd a_8860_3944# a_8772_3988# vdd pfet_06v0 w=1.22u l=1u
X41 pbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X42 a_7516_6647# a_7428_6744# vss vss nfet_06v0 w=0.82u l=1u
X43 vdd a_5052_3944# a_4964_3988# vdd pfet_06v0 w=1.22u l=1u
X44 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X45 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X46 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X47 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X48 a_5612_8215# a_5524_8312# vss vss nfet_06v0 w=0.82u l=1u
X49 a_7964_7080# a_7876_7124# vss vss nfet_06v0 w=0.82u l=1u
X50 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X51 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X52 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X53 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X54 a_7964_6647# a_7876_6744# vss vss nfet_06v0 w=0.82u l=1u
X55 vss outnn a_9912_6340# vss nfet_06v0 w=0.82u l=0.6u
X56 a_8748_8215# a_8660_8312# vss vss nfet_06v0 w=0.82u l=1u
X57 a_6620_7080# a_6532_7124# vss vss nfet_06v0 w=0.82u l=1u
X58 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X59 outn pbus vss vss nfet_06v0 w=0.82u l=0.6u
X60 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X61 outp nbus vss vss nfet_06v0 w=0.82u l=0.6u
X62 outp outp vss vss nfet_06v0 w=0.82u l=0.6u
X63 outn pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X64 vdd a_6172_5079# a_6084_5176# vdd pfet_06v0 w=1.22u l=1u
X65 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X66 nbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X67 vdd a_6956_5512# a_6868_5556# vdd pfet_06v0 w=1.22u l=1u
X68 outp nbus vss vss nfet_06v0 w=0.82u l=0.6u
X69 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X70 a_7404_8215# a_7316_8312# vss vss nfet_06v0 w=0.82u l=1u
X71 outp outp vdd vdd pfet_06v0 w=1.22u l=0.5u
X72 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X73 outxor outpn a_9688_6744# vdd pfet_06v0 w=1.22u l=0.5u
X74 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X75 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X76 outp outp vdd vdd pfet_06v0 w=1.22u l=0.5u
X77 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X78 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X79 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X80 outp outn vdd vdd pfet_06v0 w=1.22u l=0.5u
X81 a_8860_5512# a_8772_5556# vss vss nfet_06v0 w=0.82u l=1u
X82 a_7852_8215# a_7764_8312# vss vss nfet_06v0 w=0.82u l=1u
X83 a_8412_7080# a_8324_7124# vss vss nfet_06v0 w=0.82u l=1u
X84 vdd a_7516_6647# a_7428_6744# vdd pfet_06v0 w=1.22u l=1u
X85 nbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X86 outn outn vss vss nfet_06v0 w=0.82u l=0.6u
X87 vss outpn a_9016_6876# vss nfet_06v0 w=0.36u l=0.6u
X88 vss nbus pbus vss nfet_06v0 w=0.82u l=0.6u
X89 a_7068_7080# a_6980_7124# vss vss nfet_06v0 w=0.82u l=1u
X90 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X91 vdd a_7964_6647# a_7876_6744# vdd pfet_06v0 w=1.22u l=1u
X92 a_8860_7080# a_8772_7124# vss vss nfet_06v0 w=0.82u l=1u
X93 vdd pbus pbus vdd pfet_06v0 w=1.22u l=0.5u
X94 a_9204_6876# outnn a_9016_6876# vdd pfet_06v0 w=0.56u l=0.5u
X95 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X96 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X97 vdd pbus pbus vdd pfet_06v0 w=1.22u l=0.5u
X98 a_9532_3511# a_9444_3608# vss vss nfet_06v0 w=0.82u l=1u
X99 nbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X100 nbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X101 a_8300_8215# a_8212_8312# vss vss nfet_06v0 w=0.82u l=1u
X102 outn outp vss vss nfet_06v0 w=0.82u l=0.6u
X103 a_6172_3511# a_6084_3608# vss vss nfet_06v0 w=0.82u l=1u
X104 outn outn vdd vdd pfet_06v0 w=1.22u l=0.5u
X105 a_9532_8215# a_9444_8312# vss vss nfet_06v0 w=0.82u l=1u
X106 nbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X107 outn pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X108 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X109 vdd nbus pbus vdd pfet_06v0 w=1.22u l=0.5u
X110 pbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X111 a_9980_8215# a_9892_8312# vss vss nfet_06v0 w=0.82u l=1u
X112 nbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X113 outn pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X114 outn outp vss vss nfet_06v0 w=0.82u l=0.6u
X115 outn outn vdd vdd pfet_06v0 w=1.22u l=0.5u
X116 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X117 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X118 a_9688_6744# a_9016_6876# vdd vdd pfet_06v0 w=1.22u l=0.5u
X119 pbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X120 vdd outn outp vdd pfet_06v0 w=1.22u l=0.5u
X121 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X122 outp outp vdd vdd pfet_06v0 w=1.22u l=0.5u
X123 vss outp outpn vss nfet_06v0 w=0.82u l=0.6u
X124 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X125 vdd a_9532_3511# a_9444_3608# vdd pfet_06v0 w=1.22u l=1u
X126 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X127 vdd a_8860_5512# a_8772_5556# vdd pfet_06v0 w=1.22u l=1u
X128 a_6060_8215# a_5972_8312# vss vss nfet_06v0 w=0.82u l=1u
X129 outn pbus vss vss nfet_06v0 w=0.82u l=0.6u
X130 outp nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X131 outp nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X132 vdd a_6508_8215# a_6420_8312# vdd pfet_06v0 w=1.22u l=1u
X133 vdd a_6172_3511# a_6084_3608# vdd pfet_06v0 w=1.22u l=1u
X134 pbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X135 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X136 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X137 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X138 vdd a_6956_8215# a_6868_8312# vdd pfet_06v0 w=1.22u l=1u
X139 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X140 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X141 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X142 vdd a_1692_8215# a_1604_8312# vdd pfet_06v0 w=1.22u l=1u
X143 pbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X144 pbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X145 vdd a_5612_8215# a_5524_8312# vdd pfet_06v0 w=1.22u l=1u
X146 vdd a_1692_7080# a_1604_7124# vdd pfet_06v0 w=1.22u l=1u
X147 outp outp vss vss nfet_06v0 w=0.82u l=0.6u
X148 a_9016_6876# outnn vss vss nfet_06v0 w=0.36u l=0.6u
X149 a_1692_5079# a_1604_5176# vss vss nfet_06v0 w=0.82u l=1u
X150 outp outn vss vss nfet_06v0 w=0.82u l=0.6u
X151 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X152 vdd a_8748_8215# a_8660_8312# vdd pfet_06v0 w=1.22u l=1u
X153 vdd a_7516_7080# a_7428_7124# vdd pfet_06v0 w=1.22u l=1u
X154 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X155 vdd outp outpn vdd pfet_06v0 w=1.22u l=0.5u
X156 a_9688_6744# outnn outxor vdd pfet_06v0 w=1.22u l=0.5u
X157 vdd a_7404_8215# a_7316_8312# vdd pfet_06v0 w=1.22u l=1u
X158 vss pbus pbus vss nfet_06v0 w=0.82u l=0.6u
X159 a_8748_5079# a_8660_5176# vss vss nfet_06v0 w=0.82u l=1u
X160 pbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X161 vdd a_7964_7080# a_7876_7124# vdd pfet_06v0 w=1.22u l=1u
X162 outn pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X163 vss pbus pbus vss nfet_06v0 w=0.82u l=0.6u
X164 outp outp vdd vdd pfet_06v0 w=1.22u l=0.5u
X165 nbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X166 vdd a_7852_8215# a_7764_8312# vdd pfet_06v0 w=1.22u l=1u
X167 nbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X168 vdd a_6620_7080# a_6532_7124# vdd pfet_06v0 w=1.22u l=1u
X169 outn outp vdd vdd pfet_06v0 w=1.22u l=0.5u
X170 nbus pbus vss vss nfet_06v0 w=0.82u l=0.6u
X171 outn pbus vss vss nfet_06v0 w=0.82u l=0.6u
X172 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X173 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X174 outn outn vss vss nfet_06v0 w=0.82u l=0.6u
X175 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X176 vdd outpn a_9204_6876# vdd pfet_06v0 w=0.56u l=0.5u
X177 outn pbus vss vss nfet_06v0 w=0.82u l=0.6u
X178 outp outp vss vss nfet_06v0 w=0.82u l=0.6u
X179 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X180 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X181 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X182 vss outn outnn vss nfet_06v0 w=0.82u l=0.6u
X183 outn outn vdd vdd pfet_06v0 w=1.22u l=0.5u
X184 outp outp vss vss nfet_06v0 w=0.82u l=0.6u
X185 vdd a_1692_5079# a_1604_5176# vdd pfet_06v0 w=1.22u l=1u
X186 outp nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X187 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X188 nbus nbus vss vss nfet_06v0 w=0.82u l=0.6u
X189 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X190 vss outn outn vss nfet_06v0 w=0.82u l=0.6u
X191 outn outp vdd vdd pfet_06v0 w=1.22u l=0.5u
X192 a_8860_3944# a_8772_3988# vss vss nfet_06v0 w=0.82u l=1u
X193 a_5052_3944# a_4964_3988# vss vss nfet_06v0 w=0.82u l=1u
X194 nbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X195 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X196 nbus nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X197 vdd a_8412_7080# a_8324_7124# vdd pfet_06v0 w=1.22u l=1u
X198 pbus pbus vdd vdd pfet_06v0 w=1.22u l=0.5u
X199 outp nbus vdd vdd pfet_06v0 w=1.22u l=0.5u
C0 pbus vdd 5.47fF
C1 vdd outn 2.39fF
C2 vdd nbus 5.46fF
C3 vdd outp 2.79fF
C4 pbus nbus 4.17fF
C5 outp outn 2.09fF
C6 outp vss 6.09fF
C7 outn vss 5.91fF
C8 pbus vss 16.82fF
C9 nbus vss 16.68fF
C10 vdd vss 101.68fF
.ends



XDUT nbus outn outnn outp outpn outxor pbus vdd vss active_load_flat


**** end user architecture code
.ends

.GLOBAL GND
.end
