magic
tech gf180mcuC
magscale 1 2
timestamp 1669947198
<< metal4 >>
rect 13000 47062 25160 47702
rect 41160 47382 53000 47702
rect 40840 47062 53000 47382
rect 13000 46742 25480 47062
rect 40520 46742 53000 47062
rect 13000 46102 25800 46742
rect 40200 46102 53000 46742
rect 13000 45782 26120 46102
rect 39880 45782 53000 46102
rect 13000 45462 26440 45782
rect 39560 45462 53000 45782
rect 13000 44822 26760 45462
rect 39240 44822 53000 45462
rect 13000 44502 27080 44822
rect 38920 44502 53000 44822
rect 13000 43862 27400 44502
rect 38600 43862 53000 44502
rect 13000 43542 27720 43862
rect 38280 43542 53000 43862
rect 13000 43222 28040 43542
rect 37960 43222 53000 43542
rect 13000 42582 28360 43222
rect 37640 42582 53000 43222
rect 13000 42262 28680 42582
rect 37320 42262 53000 42582
rect 13000 41942 29000 42262
rect 37000 41942 53000 42262
rect 13000 41302 29320 41942
rect 36680 41302 53000 41942
rect 13000 40982 29640 41302
rect 36360 40982 53000 41302
rect 13000 40342 29960 40982
rect 36040 40342 53000 40982
rect 13000 40022 30280 40342
rect 35720 40022 53000 40342
rect 13000 39702 30600 40022
rect 35400 39702 53000 40022
rect 15880 39382 30920 39702
rect 16200 39062 30920 39382
rect 35080 39382 50120 39702
rect 35080 39062 49800 39382
rect 16200 38742 31240 39062
rect 34760 38742 49800 39062
rect 16200 38422 31560 38742
rect 34440 38422 49800 38742
rect 16200 37782 31880 38422
rect 34120 37782 49800 38422
rect 16200 37462 32200 37782
rect 33800 37462 49800 37782
rect 16200 36822 32520 37462
rect 33480 36822 49800 37462
rect 16200 36502 32840 36822
rect 33160 36502 49800 36822
rect 16200 34902 49800 36502
rect 16200 27542 24840 34902
rect 25160 34582 40840 34902
rect 25480 34262 40520 34582
rect 25800 33622 40200 34262
rect 26120 33302 39880 33622
rect 26440 32982 39560 33302
rect 26760 32342 39240 32982
rect 27080 32022 38920 32342
rect 27400 31702 38600 32022
rect 27720 31062 38280 31702
rect 28040 30742 37960 31062
rect 28360 30422 37640 30742
rect 28680 29782 37320 30422
rect 29000 29462 37000 29782
rect 29320 28822 36680 29462
rect 29640 28502 36360 28822
rect 29960 28182 36040 28502
rect 30280 27542 35720 28182
rect 41160 27542 49800 34902
rect 15880 27222 24840 27542
rect 30600 27222 35400 27542
rect 41160 27222 50120 27542
rect 13000 19222 28040 27222
rect 30920 26902 35080 27222
rect 31240 26262 34760 26902
rect 31560 25942 34440 26262
rect 31880 25622 34120 25942
rect 32200 24982 33800 25622
rect 32520 24662 33480 24982
rect 32840 24342 33160 24662
rect 37960 19222 53000 27222
tri 5920 12215 7440 13735 se
rect 7440 12215 8428 13735
rect 9492 12215 10480 13735
tri 10480 12215 12000 13735 sw
rect 31000 12215 35560 13735
tri 36320 12215 37840 13735 se
rect 37840 12215 40130 13735
tri 40130 12215 41650 13735 sw
tri 42400 12975 43160 13735 se
rect 43160 12975 47720 13735
tri 47720 12975 48480 13735 sw
rect 42400 12215 48480 12975
tri 49240 12215 50760 13735 se
rect 50760 12215 51748 13735
rect 52812 12215 53800 13735
tri 53800 12215 55320 13735 sw
rect 5920 7655 7440 12215
tri 7440 11455 8200 12215 nw
tri 9720 11455 10480 12215 ne
tri 7440 7655 8200 8415 sw
tri 9720 7655 10480 8415 se
rect 10480 7655 12000 12215
tri 18840 11455 19600 12215 se
rect 19600 11455 23400 12215
tri 23400 11455 24160 12215 sw
rect 12760 9935 16560 11455
tri 16560 9935 18080 11455 sw
rect 12760 9175 14280 9935
tri 15800 9175 16560 9935 ne
tri 5920 6135 7440 7655 ne
rect 7440 6135 10480 7655
tri 10480 6135 12000 7655 nw
rect 12760 7655 14280 8415
tri 15800 7655 16560 8415 se
rect 16560 7655 18080 9935
rect 12760 6135 16560 7655
tri 16560 6135 18080 7655 nw
rect 18840 10695 24160 11455
rect 18840 7655 20360 10695
rect 22640 9935 24160 10695
rect 21424 9175 24160 9935
rect 21424 8415 23400 9175
tri 23400 8415 24160 9175 nw
rect 24760 11035 26280 11455
tri 26620 11035 27040 11455 se
rect 27040 11035 28560 11455
tri 28560 11035 28980 11455 sw
rect 24760 9935 28980 11035
tri 28980 9935 30080 11035 sw
rect 18840 6895 24160 7655
tri 18840 6135 19600 6895 ne
rect 19600 6135 23400 6895
tri 23400 6135 24160 6895 nw
rect 24760 6135 26280 9935
tri 26280 9175 27040 9935 nw
tri 27800 9175 28560 9935 ne
rect 28560 6135 30080 9935
rect 31000 10695 32520 12215
rect 31000 9175 34040 10695
rect 36320 9175 37840 12215
tri 37840 11455 38600 12215 nw
tri 39370 11455 40130 12215 ne
rect 40130 9175 41640 12215
rect 42400 10695 43920 12215
rect 42400 9935 47720 10695
tri 47720 9935 48480 10695 sw
tri 42400 9175 43160 9935 ne
rect 43160 9175 48480 9935
rect 31000 6135 32520 9175
rect 36320 7655 38600 9175
rect 39360 7655 41640 9175
rect 46960 7655 48480 9175
rect 36320 6135 37840 7655
rect 40130 6135 41640 7655
rect 42400 6895 48480 7655
tri 42400 6135 43160 6895 ne
rect 43160 6135 47720 6895
tri 47720 6135 48480 6895 nw
rect 49240 7655 50760 12215
tri 50760 11455 51520 12215 nw
tri 53040 11455 53800 12215 ne
tri 50760 7655 51520 8415 sw
tri 53040 7655 53800 8415 se
rect 53800 7655 55320 12215
tri 49240 6135 50760 7655 ne
rect 50760 6135 53800 7655
tri 53800 6135 55320 7655 nw
tri 56080 12215 57600 13735 se
rect 57600 12215 59880 13735
tri 59880 12215 61400 13735 sw
rect 56080 7655 57600 12215
tri 57600 11455 58360 12215 nw
tri 59120 11455 59880 12215 ne
rect 59880 10695 61400 12215
tri 57600 7655 58360 8415 sw
tri 59120 7655 59880 8415 se
rect 59880 7655 61400 9175
tri 56080 6135 57600 7655 ne
rect 57600 6135 59880 7655
tri 59880 6135 61400 7655 nw
rect 12760 3855 14280 6135
<< fillblock >>
rect 0 0 66000 50000
<< end >>
