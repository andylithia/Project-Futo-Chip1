magic
tech gf180mcuC
magscale 1 10
timestamp 1669998789
<< deepnwell >>
rect -120 -120 570 590
<< nwell >>
rect 0 0 180 450
<< nsubdiff >>
rect 37 380 143 410
rect 37 60 50 380
rect 130 60 143 380
rect 37 30 143 60
<< nsubdiffcont >>
rect 50 60 130 380
<< metal1 >>
rect 50 380 130 410
rect 50 30 130 60
<< end >>
