magic
tech gf180mcuC
magscale 1 10
timestamp 1669518838
<< metal1 >>
rect 18610 16606 18622 16658
rect 18674 16655 18686 16658
rect 19170 16655 19182 16658
rect 18674 16609 19182 16655
rect 18674 16606 18686 16609
rect 19170 16606 19182 16609
rect 19234 16606 19246 16658
rect 20178 16606 20190 16658
rect 20242 16655 20254 16658
rect 21410 16655 21422 16658
rect 20242 16609 21422 16655
rect 20242 16606 20254 16609
rect 21410 16606 21422 16609
rect 21474 16606 21486 16658
rect 29586 16606 29598 16658
rect 29650 16655 29662 16658
rect 31378 16655 31390 16658
rect 29650 16609 31390 16655
rect 29650 16606 29662 16609
rect 31378 16606 31390 16609
rect 31442 16606 31454 16658
rect 35858 16606 35870 16658
rect 35922 16655 35934 16658
rect 36418 16655 36430 16658
rect 35922 16609 36430 16655
rect 35922 16606 35934 16609
rect 36418 16606 36430 16609
rect 36482 16606 36494 16658
rect 37426 16606 37438 16658
rect 37490 16655 37502 16658
rect 37986 16655 37998 16658
rect 37490 16609 37998 16655
rect 37490 16606 37502 16609
rect 37986 16606 37998 16609
rect 38050 16606 38062 16658
rect 44146 16606 44158 16658
rect 44210 16655 44222 16658
rect 44930 16655 44942 16658
rect 44210 16609 44942 16655
rect 44210 16606 44222 16609
rect 44930 16606 44942 16609
rect 44994 16606 45006 16658
rect 1344 16490 178640 16524
rect 1344 16438 23376 16490
rect 23428 16438 23480 16490
rect 23532 16438 23584 16490
rect 23636 16438 67700 16490
rect 67752 16438 67804 16490
rect 67856 16438 67908 16490
rect 67960 16438 112024 16490
rect 112076 16438 112128 16490
rect 112180 16438 112232 16490
rect 112284 16438 156348 16490
rect 156400 16438 156452 16490
rect 156504 16438 156556 16490
rect 156608 16438 178640 16490
rect 1344 16404 178640 16438
rect 5854 16210 5906 16222
rect 15262 16210 15314 16222
rect 12562 16158 12574 16210
rect 12626 16158 12638 16210
rect 5854 16146 5906 16158
rect 15262 16146 15314 16158
rect 20190 16210 20242 16222
rect 20190 16146 20242 16158
rect 24670 16210 24722 16222
rect 38782 16210 38834 16222
rect 36306 16158 36318 16210
rect 36370 16158 36382 16210
rect 24670 16146 24722 16158
rect 38782 16146 38834 16158
rect 44158 16210 44210 16222
rect 44158 16146 44210 16158
rect 48190 16210 48242 16222
rect 49858 16158 49870 16210
rect 49922 16158 49934 16210
rect 51986 16158 51998 16210
rect 52050 16158 52062 16210
rect 61618 16158 61630 16210
rect 61682 16158 61694 16210
rect 63746 16158 63758 16210
rect 63810 16158 63822 16210
rect 94882 16158 94894 16210
rect 94946 16158 94958 16210
rect 48190 16146 48242 16158
rect 1822 16098 1874 16110
rect 1822 16034 1874 16046
rect 6302 16098 6354 16110
rect 15710 16098 15762 16110
rect 9762 16046 9774 16098
rect 9826 16046 9838 16098
rect 6302 16034 6354 16046
rect 15710 16034 15762 16046
rect 17502 16098 17554 16110
rect 17502 16034 17554 16046
rect 18622 16098 18674 16110
rect 18622 16034 18674 16046
rect 21422 16098 21474 16110
rect 21422 16034 21474 16046
rect 25342 16098 25394 16110
rect 25342 16034 25394 16046
rect 29150 16098 29202 16110
rect 31390 16098 31442 16110
rect 39230 16098 39282 16110
rect 30594 16046 30606 16098
rect 30658 16046 30670 16098
rect 33506 16046 33518 16098
rect 33570 16046 33582 16098
rect 29150 16034 29202 16046
rect 31390 16034 31442 16046
rect 39230 16034 39282 16046
rect 44942 16098 44994 16110
rect 49186 16046 49198 16098
rect 49250 16046 49262 16098
rect 52770 16046 52782 16098
rect 52834 16046 52846 16098
rect 54226 16046 54238 16098
rect 54290 16046 54302 16098
rect 60834 16046 60846 16098
rect 60898 16046 60910 16098
rect 91970 16046 91982 16098
rect 92034 16046 92046 16098
rect 44942 16034 44994 16046
rect 3166 15986 3218 15998
rect 3166 15922 3218 15934
rect 4734 15986 4786 15998
rect 4734 15922 4786 15934
rect 6638 15986 6690 15998
rect 6638 15922 6690 15934
rect 7870 15986 7922 15998
rect 7870 15922 7922 15934
rect 8878 15986 8930 15998
rect 14142 15986 14194 15998
rect 10434 15934 10446 15986
rect 10498 15934 10510 15986
rect 8878 15922 8930 15934
rect 14142 15922 14194 15934
rect 16718 15986 16770 15998
rect 16718 15922 16770 15934
rect 19182 15986 19234 15998
rect 19182 15922 19234 15934
rect 22318 15986 22370 15998
rect 22318 15922 22370 15934
rect 23550 15986 23602 15998
rect 23550 15922 23602 15934
rect 25678 15986 25730 15998
rect 25678 15922 25730 15934
rect 26686 15986 26738 15998
rect 26686 15922 26738 15934
rect 28254 15986 28306 15998
rect 28254 15922 28306 15934
rect 30046 15986 30098 15998
rect 30046 15922 30098 15934
rect 31726 15986 31778 15998
rect 31726 15922 31778 15934
rect 32398 15986 32450 15998
rect 37102 15986 37154 15998
rect 34178 15934 34190 15986
rect 34242 15934 34254 15986
rect 32398 15922 32450 15934
rect 37102 15922 37154 15934
rect 37438 15986 37490 15998
rect 37438 15922 37490 15934
rect 37998 15986 38050 15998
rect 37998 15922 38050 15934
rect 41022 15986 41074 15998
rect 41022 15922 41074 15934
rect 42366 15986 42418 15998
rect 42366 15922 42418 15934
rect 45838 15986 45890 15998
rect 45838 15922 45890 15934
rect 47070 15986 47122 15998
rect 47070 15922 47122 15934
rect 53566 15986 53618 15998
rect 53566 15922 53618 15934
rect 54910 15986 54962 15998
rect 54910 15922 54962 15934
rect 56702 15986 56754 15998
rect 56702 15922 56754 15934
rect 59614 15986 59666 15998
rect 59614 15922 59666 15934
rect 65886 15986 65938 15998
rect 65886 15922 65938 15934
rect 66558 15986 66610 15998
rect 66558 15922 66610 15934
rect 69022 15986 69074 15998
rect 69022 15922 69074 15934
rect 70590 15986 70642 15998
rect 70590 15922 70642 15934
rect 73054 15986 73106 15998
rect 73054 15922 73106 15934
rect 75294 15986 75346 15998
rect 75294 15922 75346 15934
rect 78430 15986 78482 15998
rect 78430 15922 78482 15934
rect 80222 15986 80274 15998
rect 80222 15922 80274 15934
rect 83134 15986 83186 15998
rect 83134 15922 83186 15934
rect 84702 15986 84754 15998
rect 84702 15922 84754 15934
rect 88062 15986 88114 15998
rect 88062 15922 88114 15934
rect 89294 15986 89346 15998
rect 97246 15986 97298 15998
rect 92754 15934 92766 15986
rect 92818 15934 92830 15986
rect 89294 15922 89346 15934
rect 97246 15922 97298 15934
rect 98814 15986 98866 15998
rect 98814 15922 98866 15934
rect 101950 15986 102002 15998
rect 101950 15922 102002 15934
rect 103742 15986 103794 15998
rect 103742 15922 103794 15934
rect 106654 15986 106706 15998
rect 106654 15922 106706 15934
rect 108222 15986 108274 15998
rect 108222 15922 108274 15934
rect 111582 15986 111634 15998
rect 111582 15922 111634 15934
rect 112926 15986 112978 15998
rect 112926 15922 112978 15934
rect 116062 15986 116114 15998
rect 116062 15922 116114 15934
rect 117630 15986 117682 15998
rect 117630 15922 117682 15934
rect 120766 15986 120818 15998
rect 120766 15922 120818 15934
rect 122334 15986 122386 15998
rect 122334 15922 122386 15934
rect 125470 15986 125522 15998
rect 125470 15922 125522 15934
rect 127262 15986 127314 15998
rect 127262 15922 127314 15934
rect 130174 15986 130226 15998
rect 130174 15922 130226 15934
rect 131742 15986 131794 15998
rect 131742 15922 131794 15934
rect 135102 15986 135154 15998
rect 135102 15922 135154 15934
rect 136446 15986 136498 15998
rect 136446 15922 136498 15934
rect 139582 15986 139634 15998
rect 139582 15922 139634 15934
rect 141150 15986 141202 15998
rect 141150 15922 141202 15934
rect 144286 15986 144338 15998
rect 144286 15922 144338 15934
rect 145854 15986 145906 15998
rect 145854 15922 145906 15934
rect 148990 15986 149042 15998
rect 148990 15922 149042 15934
rect 150782 15986 150834 15998
rect 150782 15922 150834 15934
rect 153694 15986 153746 15998
rect 153694 15922 153746 15934
rect 155262 15986 155314 15998
rect 155262 15922 155314 15934
rect 158622 15986 158674 15998
rect 158622 15922 158674 15934
rect 159966 15986 160018 15998
rect 159966 15922 160018 15934
rect 163102 15986 163154 15998
rect 163102 15922 163154 15934
rect 164670 15986 164722 15998
rect 164670 15922 164722 15934
rect 167806 15986 167858 15998
rect 167806 15922 167858 15934
rect 169374 15986 169426 15998
rect 169374 15922 169426 15934
rect 172510 15986 172562 15998
rect 172510 15922 172562 15934
rect 174302 15986 174354 15998
rect 174302 15922 174354 15934
rect 177214 15986 177266 15998
rect 177214 15922 177266 15934
rect 2158 15874 2210 15886
rect 2158 15810 2210 15822
rect 13470 15874 13522 15886
rect 13470 15810 13522 15822
rect 16046 15874 16098 15886
rect 16046 15810 16098 15822
rect 18062 15874 18114 15886
rect 18062 15810 18114 15822
rect 19742 15874 19794 15886
rect 19742 15810 19794 15822
rect 20750 15874 20802 15886
rect 20750 15810 20802 15822
rect 21758 15874 21810 15886
rect 21758 15810 21810 15822
rect 27694 15874 27746 15886
rect 27694 15810 27746 15822
rect 39566 15874 39618 15886
rect 64654 15874 64706 15886
rect 45266 15822 45278 15874
rect 45330 15822 45342 15874
rect 39566 15810 39618 15822
rect 64654 15810 64706 15822
rect 73726 15874 73778 15886
rect 73726 15810 73778 15822
rect 74398 15874 74450 15886
rect 74398 15810 74450 15822
rect 90078 15874 90130 15886
rect 90078 15810 90130 15822
rect 90638 15874 90690 15886
rect 90638 15810 90690 15822
rect 91198 15874 91250 15886
rect 91198 15810 91250 15822
rect 1344 15706 178800 15740
rect 1344 15654 45538 15706
rect 45590 15654 45642 15706
rect 45694 15654 45746 15706
rect 45798 15654 89862 15706
rect 89914 15654 89966 15706
rect 90018 15654 90070 15706
rect 90122 15654 134186 15706
rect 134238 15654 134290 15706
rect 134342 15654 134394 15706
rect 134446 15654 178510 15706
rect 178562 15654 178614 15706
rect 178666 15654 178718 15706
rect 178770 15654 178800 15706
rect 1344 15620 178800 15654
rect 1822 15538 1874 15550
rect 1822 15474 1874 15486
rect 14702 15538 14754 15550
rect 14702 15474 14754 15486
rect 16046 15538 16098 15550
rect 16046 15474 16098 15486
rect 16718 15538 16770 15550
rect 16718 15474 16770 15486
rect 26238 15538 26290 15550
rect 26238 15474 26290 15486
rect 32398 15538 32450 15550
rect 32398 15474 32450 15486
rect 36430 15538 36482 15550
rect 36430 15474 36482 15486
rect 37102 15538 37154 15550
rect 37102 15474 37154 15486
rect 37438 15538 37490 15550
rect 37438 15474 37490 15486
rect 48526 15538 48578 15550
rect 48526 15474 48578 15486
rect 50206 15538 50258 15550
rect 50206 15474 50258 15486
rect 51326 15538 51378 15550
rect 51326 15474 51378 15486
rect 60062 15538 60114 15550
rect 60062 15474 60114 15486
rect 60622 15538 60674 15550
rect 60622 15474 60674 15486
rect 61182 15538 61234 15550
rect 61182 15474 61234 15486
rect 76526 15538 76578 15550
rect 76526 15474 76578 15486
rect 76974 15538 77026 15550
rect 76974 15474 77026 15486
rect 91758 15538 91810 15550
rect 91758 15474 91810 15486
rect 92542 15538 92594 15550
rect 92542 15474 92594 15486
rect 94110 15538 94162 15550
rect 94110 15474 94162 15486
rect 178110 15538 178162 15550
rect 178110 15474 178162 15486
rect 10782 15426 10834 15438
rect 16606 15426 16658 15438
rect 12114 15374 12126 15426
rect 12178 15374 12190 15426
rect 10782 15362 10834 15374
rect 16606 15362 16658 15374
rect 20302 15426 20354 15438
rect 20302 15362 20354 15374
rect 20862 15426 20914 15438
rect 35086 15426 35138 15438
rect 22082 15374 22094 15426
rect 22146 15374 22158 15426
rect 22978 15374 22990 15426
rect 23042 15374 23054 15426
rect 27570 15374 27582 15426
rect 27634 15374 27646 15426
rect 20862 15362 20914 15374
rect 35086 15362 35138 15374
rect 54014 15426 54066 15438
rect 54014 15362 54066 15374
rect 63758 15426 63810 15438
rect 63758 15362 63810 15374
rect 65438 15426 65490 15438
rect 79650 15374 79662 15426
rect 79714 15374 79726 15426
rect 65438 15362 65490 15374
rect 19406 15314 19458 15326
rect 33742 15314 33794 15326
rect 10546 15262 10558 15314
rect 10610 15262 10622 15314
rect 11442 15262 11454 15314
rect 11506 15262 11518 15314
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 26898 15262 26910 15314
rect 26962 15262 26974 15314
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 31714 15262 31726 15314
rect 31778 15262 31790 15314
rect 19406 15250 19458 15262
rect 33742 15250 33794 15262
rect 34190 15314 34242 15326
rect 53566 15314 53618 15326
rect 64654 15314 64706 15326
rect 35858 15262 35870 15314
rect 35922 15262 35934 15314
rect 51986 15262 51998 15314
rect 52050 15262 52062 15314
rect 63186 15262 63198 15314
rect 63250 15262 63262 15314
rect 73602 15262 73614 15314
rect 73666 15262 73678 15314
rect 74834 15262 74846 15314
rect 74898 15262 74910 15314
rect 80434 15262 80446 15314
rect 80498 15262 80510 15314
rect 89506 15262 89518 15314
rect 89570 15262 89582 15314
rect 90738 15262 90750 15314
rect 90802 15262 90814 15314
rect 34190 15250 34242 15262
rect 53566 15250 53618 15262
rect 64654 15250 64706 15262
rect 18510 15202 18562 15214
rect 14242 15150 14254 15202
rect 14306 15150 14318 15202
rect 18510 15138 18562 15150
rect 19742 15202 19794 15214
rect 21758 15202 21810 15214
rect 21186 15150 21198 15202
rect 21250 15150 21262 15202
rect 19742 15138 19794 15150
rect 21758 15138 21810 15150
rect 22654 15202 22706 15214
rect 22654 15138 22706 15150
rect 23550 15202 23602 15214
rect 31054 15202 31106 15214
rect 29698 15150 29710 15202
rect 29762 15150 29774 15202
rect 23550 15138 23602 15150
rect 31054 15138 31106 15150
rect 52670 15202 52722 15214
rect 52670 15138 52722 15150
rect 74174 15202 74226 15214
rect 90078 15202 90130 15214
rect 77522 15150 77534 15202
rect 77586 15150 77598 15202
rect 74174 15138 74226 15150
rect 90078 15138 90130 15150
rect 1344 14922 178640 14956
rect 1344 14870 23376 14922
rect 23428 14870 23480 14922
rect 23532 14870 23584 14922
rect 23636 14870 67700 14922
rect 67752 14870 67804 14922
rect 67856 14870 67908 14922
rect 67960 14870 112024 14922
rect 112076 14870 112128 14922
rect 112180 14870 112232 14922
rect 112284 14870 156348 14922
rect 156400 14870 156452 14922
rect 156504 14870 156556 14922
rect 156608 14870 178640 14922
rect 1344 14836 178640 14870
rect 11006 14642 11058 14654
rect 11006 14578 11058 14590
rect 19518 14642 19570 14654
rect 19518 14578 19570 14590
rect 20526 14642 20578 14654
rect 30046 14642 30098 14654
rect 23426 14590 23438 14642
rect 23490 14590 23502 14642
rect 20526 14578 20578 14590
rect 30046 14578 30098 14590
rect 30382 14642 30434 14654
rect 30382 14578 30434 14590
rect 31166 14642 31218 14654
rect 31166 14578 31218 14590
rect 33182 14642 33234 14654
rect 33182 14578 33234 14590
rect 33742 14642 33794 14654
rect 33742 14578 33794 14590
rect 35086 14642 35138 14654
rect 35086 14578 35138 14590
rect 88958 14642 89010 14654
rect 88958 14578 89010 14590
rect 16830 14530 16882 14542
rect 18958 14530 19010 14542
rect 15362 14478 15374 14530
rect 15426 14478 15438 14530
rect 17490 14478 17502 14530
rect 17554 14478 17566 14530
rect 16830 14466 16882 14478
rect 18958 14466 19010 14478
rect 34190 14530 34242 14542
rect 89854 14530 89906 14542
rect 35858 14478 35870 14530
rect 35922 14478 35934 14530
rect 63186 14478 63198 14530
rect 63250 14478 63262 14530
rect 64530 14478 64542 14530
rect 64594 14478 64606 14530
rect 72706 14478 72718 14530
rect 72770 14478 72782 14530
rect 73938 14478 73950 14530
rect 74002 14478 74014 14530
rect 88386 14478 88398 14530
rect 88450 14478 88462 14530
rect 34190 14466 34242 14478
rect 89854 14466 89906 14478
rect 12574 14418 12626 14430
rect 12574 14354 12626 14366
rect 15934 14418 15986 14430
rect 15934 14354 15986 14366
rect 18062 14418 18114 14430
rect 23214 14418 23266 14430
rect 20850 14366 20862 14418
rect 20914 14366 20926 14418
rect 18062 14354 18114 14366
rect 23214 14354 23266 14366
rect 53678 14418 53730 14430
rect 53678 14354 53730 14366
rect 63758 14418 63810 14430
rect 63758 14354 63810 14366
rect 73278 14418 73330 14430
rect 73278 14354 73330 14366
rect 19966 14306 20018 14318
rect 19966 14242 20018 14254
rect 21870 14306 21922 14318
rect 21870 14242 21922 14254
rect 22654 14306 22706 14318
rect 22654 14242 22706 14254
rect 23998 14306 24050 14318
rect 23998 14242 24050 14254
rect 1344 14138 178800 14172
rect 1344 14086 45538 14138
rect 45590 14086 45642 14138
rect 45694 14086 45746 14138
rect 45798 14086 89862 14138
rect 89914 14086 89966 14138
rect 90018 14086 90070 14138
rect 90122 14086 134186 14138
rect 134238 14086 134290 14138
rect 134342 14086 134394 14138
rect 134446 14086 178510 14138
rect 178562 14086 178614 14138
rect 178666 14086 178718 14138
rect 178770 14086 178800 14138
rect 1344 14052 178800 14086
rect 16606 13970 16658 13982
rect 16606 13906 16658 13918
rect 16942 13970 16994 13982
rect 16942 13906 16994 13918
rect 21298 13806 21310 13858
rect 21362 13806 21374 13858
rect 61630 13746 61682 13758
rect 19282 13694 19294 13746
rect 19346 13694 19358 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 61630 13682 61682 13694
rect 17726 13634 17778 13646
rect 17726 13570 17778 13582
rect 18174 13634 18226 13646
rect 18174 13570 18226 13582
rect 18622 13634 18674 13646
rect 20078 13634 20130 13646
rect 20974 13634 21026 13646
rect 24894 13634 24946 13646
rect 19506 13582 19518 13634
rect 19570 13582 19582 13634
rect 20402 13582 20414 13634
rect 20466 13582 20478 13634
rect 23762 13582 23774 13634
rect 23826 13582 23838 13634
rect 18622 13570 18674 13582
rect 20078 13570 20130 13582
rect 20974 13570 21026 13582
rect 24894 13570 24946 13582
rect 61742 13522 61794 13534
rect 61742 13458 61794 13470
rect 1344 13354 178640 13388
rect 1344 13302 23376 13354
rect 23428 13302 23480 13354
rect 23532 13302 23584 13354
rect 23636 13302 67700 13354
rect 67752 13302 67804 13354
rect 67856 13302 67908 13354
rect 67960 13302 112024 13354
rect 112076 13302 112128 13354
rect 112180 13302 112232 13354
rect 112284 13302 156348 13354
rect 156400 13302 156452 13354
rect 156504 13302 156556 13354
rect 156608 13302 178640 13354
rect 1344 13268 178640 13302
rect 26350 13186 26402 13198
rect 26350 13122 26402 13134
rect 63198 13186 63250 13198
rect 63198 13122 63250 13134
rect 18734 13074 18786 13086
rect 19630 13074 19682 13086
rect 24782 13074 24834 13086
rect 25566 13074 25618 13086
rect 18946 13022 18958 13074
rect 19010 13022 19022 13074
rect 19842 13022 19854 13074
rect 19906 13022 19918 13074
rect 20850 13022 20862 13074
rect 20914 13022 20926 13074
rect 22754 13022 22766 13074
rect 22818 13022 22830 13074
rect 24994 13022 25006 13074
rect 25058 13022 25070 13074
rect 18734 13010 18786 13022
rect 19630 13010 19682 13022
rect 24782 13010 24834 13022
rect 25566 13010 25618 13022
rect 16370 12910 16382 12962
rect 16434 12910 16446 12962
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 17166 12850 17218 12862
rect 17166 12786 17218 12798
rect 20526 12850 20578 12862
rect 20526 12786 20578 12798
rect 26462 12850 26514 12862
rect 26462 12786 26514 12798
rect 40238 12850 40290 12862
rect 40238 12786 40290 12798
rect 40798 12850 40850 12862
rect 40798 12786 40850 12798
rect 63086 12850 63138 12862
rect 63086 12786 63138 12798
rect 40910 12738 40962 12750
rect 40910 12674 40962 12686
rect 61742 12738 61794 12750
rect 61742 12674 61794 12686
rect 62414 12738 62466 12750
rect 62414 12674 62466 12686
rect 1344 12570 178800 12604
rect 1344 12518 45538 12570
rect 45590 12518 45642 12570
rect 45694 12518 45746 12570
rect 45798 12518 89862 12570
rect 89914 12518 89966 12570
rect 90018 12518 90070 12570
rect 90122 12518 134186 12570
rect 134238 12518 134290 12570
rect 134342 12518 134394 12570
rect 134446 12518 178510 12570
rect 178562 12518 178614 12570
rect 178666 12518 178718 12570
rect 178770 12518 178800 12570
rect 1344 12484 178800 12518
rect 17726 12402 17778 12414
rect 17726 12338 17778 12350
rect 19294 12402 19346 12414
rect 19294 12338 19346 12350
rect 20974 12402 21026 12414
rect 20974 12338 21026 12350
rect 23662 12402 23714 12414
rect 23662 12338 23714 12350
rect 24558 12402 24610 12414
rect 27134 12402 27186 12414
rect 26226 12350 26238 12402
rect 26290 12350 26302 12402
rect 26786 12350 26798 12402
rect 26850 12350 26862 12402
rect 24558 12338 24610 12350
rect 27134 12338 27186 12350
rect 39230 12402 39282 12414
rect 39230 12338 39282 12350
rect 60958 12402 61010 12414
rect 60958 12338 61010 12350
rect 62302 12402 62354 12414
rect 62302 12338 62354 12350
rect 19406 12290 19458 12302
rect 16930 12238 16942 12290
rect 16994 12238 17006 12290
rect 18498 12238 18510 12290
rect 18562 12238 18574 12290
rect 19406 12226 19458 12238
rect 19966 12290 20018 12302
rect 22654 12290 22706 12302
rect 25678 12290 25730 12302
rect 20290 12238 20302 12290
rect 20354 12238 20366 12290
rect 22978 12238 22990 12290
rect 23042 12238 23054 12290
rect 19966 12226 20018 12238
rect 22654 12226 22706 12238
rect 25678 12226 25730 12238
rect 27694 12290 27746 12302
rect 27694 12226 27746 12238
rect 39342 12290 39394 12302
rect 39342 12226 39394 12238
rect 39902 12290 39954 12302
rect 39902 12226 39954 12238
rect 40574 12290 40626 12302
rect 40574 12226 40626 12238
rect 41582 12290 41634 12302
rect 41582 12226 41634 12238
rect 60286 12290 60338 12302
rect 60286 12226 60338 12238
rect 61518 12290 61570 12302
rect 61518 12226 61570 12238
rect 63198 12290 63250 12302
rect 63198 12226 63250 12238
rect 63870 12290 63922 12302
rect 63870 12226 63922 12238
rect 16158 12178 16210 12190
rect 16158 12114 16210 12126
rect 16606 12178 16658 12190
rect 16606 12114 16658 12126
rect 18174 12178 18226 12190
rect 22082 12126 22094 12178
rect 22146 12126 22158 12178
rect 23650 12126 23662 12178
rect 23714 12126 23726 12178
rect 18174 12114 18226 12126
rect 20862 12066 20914 12078
rect 20862 12002 20914 12014
rect 21758 12066 21810 12078
rect 21758 12002 21810 12014
rect 24446 12066 24498 12078
rect 24446 12002 24498 12014
rect 25902 11954 25954 11966
rect 25902 11890 25954 11902
rect 60174 11954 60226 11966
rect 60174 11890 60226 11902
rect 1344 11786 178640 11820
rect 1344 11734 23376 11786
rect 23428 11734 23480 11786
rect 23532 11734 23584 11786
rect 23636 11734 67700 11786
rect 67752 11734 67804 11786
rect 67856 11734 67908 11786
rect 67960 11734 112024 11786
rect 112076 11734 112128 11786
rect 112180 11734 112232 11786
rect 112284 11734 156348 11786
rect 156400 11734 156452 11786
rect 156504 11734 156556 11786
rect 156608 11734 178640 11786
rect 1344 11700 178640 11734
rect 25790 11618 25842 11630
rect 25790 11554 25842 11566
rect 26462 11618 26514 11630
rect 26462 11554 26514 11566
rect 39342 11618 39394 11630
rect 39342 11554 39394 11566
rect 40014 11618 40066 11630
rect 40014 11554 40066 11566
rect 42142 11618 42194 11630
rect 42142 11554 42194 11566
rect 51774 11618 51826 11630
rect 51774 11554 51826 11566
rect 60510 11618 60562 11630
rect 60510 11554 60562 11566
rect 61406 11618 61458 11630
rect 61406 11554 61458 11566
rect 62974 11618 63026 11630
rect 62974 11554 63026 11566
rect 63646 11618 63698 11630
rect 63646 11554 63698 11566
rect 17278 11506 17330 11518
rect 17278 11442 17330 11454
rect 17838 11506 17890 11518
rect 18734 11506 18786 11518
rect 19630 11506 19682 11518
rect 52446 11506 52498 11518
rect 18162 11454 18174 11506
rect 18226 11454 18238 11506
rect 18946 11454 18958 11506
rect 19010 11454 19022 11506
rect 19842 11454 19854 11506
rect 19906 11454 19918 11506
rect 22082 11454 22094 11506
rect 22146 11454 22158 11506
rect 22978 11454 22990 11506
rect 23042 11454 23054 11506
rect 23874 11454 23886 11506
rect 23938 11454 23950 11506
rect 17838 11442 17890 11454
rect 18734 11442 18786 11454
rect 19630 11442 19682 11454
rect 52446 11442 52498 11454
rect 53454 11506 53506 11518
rect 53454 11442 53506 11454
rect 26574 11394 26626 11406
rect 25890 11342 25902 11394
rect 25954 11342 25966 11394
rect 26574 11330 26626 11342
rect 40126 11394 40178 11406
rect 40126 11330 40178 11342
rect 51886 11394 51938 11406
rect 51886 11330 51938 11342
rect 60622 11394 60674 11406
rect 60622 11330 60674 11342
rect 61518 11394 61570 11406
rect 61518 11330 61570 11342
rect 63086 11394 63138 11406
rect 63086 11330 63138 11342
rect 63758 11394 63810 11406
rect 63758 11330 63810 11342
rect 20526 11282 20578 11294
rect 20526 11218 20578 11230
rect 21758 11282 21810 11294
rect 21758 11218 21810 11230
rect 22654 11282 22706 11294
rect 22654 11218 22706 11230
rect 23550 11282 23602 11294
rect 23550 11218 23602 11230
rect 39454 11282 39506 11294
rect 39454 11218 39506 11230
rect 40686 11282 40738 11294
rect 40686 11218 40738 11230
rect 41470 11282 41522 11294
rect 41470 11218 41522 11230
rect 42030 11282 42082 11294
rect 42030 11218 42082 11230
rect 20638 11170 20690 11182
rect 20638 11106 20690 11118
rect 24334 11170 24386 11182
rect 24334 11106 24386 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 42702 11170 42754 11182
rect 42702 11106 42754 11118
rect 62078 11170 62130 11182
rect 62078 11106 62130 11118
rect 1344 11002 178800 11036
rect 1344 10950 45538 11002
rect 45590 10950 45642 11002
rect 45694 10950 45746 11002
rect 45798 10950 89862 11002
rect 89914 10950 89966 11002
rect 90018 10950 90070 11002
rect 90122 10950 134186 11002
rect 134238 10950 134290 11002
rect 134342 10950 134394 11002
rect 134446 10950 178510 11002
rect 178562 10950 178614 11002
rect 178666 10950 178718 11002
rect 178770 10950 178800 11002
rect 1344 10916 178800 10950
rect 18062 10834 18114 10846
rect 18062 10770 18114 10782
rect 18510 10834 18562 10846
rect 18510 10770 18562 10782
rect 19182 10834 19234 10846
rect 19182 10770 19234 10782
rect 20974 10834 21026 10846
rect 20974 10770 21026 10782
rect 39790 10834 39842 10846
rect 39790 10770 39842 10782
rect 40462 10834 40514 10846
rect 40462 10770 40514 10782
rect 52334 10834 52386 10846
rect 52334 10770 52386 10782
rect 61854 10834 61906 10846
rect 61854 10770 61906 10782
rect 20302 10722 20354 10734
rect 39902 10722 39954 10734
rect 19954 10670 19966 10722
rect 20018 10670 20030 10722
rect 22082 10670 22094 10722
rect 22146 10670 22158 10722
rect 22978 10670 22990 10722
rect 23042 10670 23054 10722
rect 20302 10658 20354 10670
rect 39902 10658 39954 10670
rect 40574 10722 40626 10734
rect 40574 10658 40626 10670
rect 41582 10722 41634 10734
rect 41582 10658 41634 10670
rect 52446 10722 52498 10734
rect 52446 10658 52498 10670
rect 61966 10722 62018 10734
rect 61966 10658 62018 10670
rect 22654 10610 22706 10622
rect 21858 10558 21870 10610
rect 21922 10558 21934 10610
rect 22654 10546 22706 10558
rect 23438 10610 23490 10622
rect 23438 10546 23490 10558
rect 24110 10610 24162 10622
rect 24110 10546 24162 10558
rect 24558 10610 24610 10622
rect 24558 10546 24610 10558
rect 19070 10498 19122 10510
rect 19070 10434 19122 10446
rect 20862 10498 20914 10510
rect 20862 10434 20914 10446
rect 1344 10218 178640 10252
rect 1344 10166 23376 10218
rect 23428 10166 23480 10218
rect 23532 10166 23584 10218
rect 23636 10166 67700 10218
rect 67752 10166 67804 10218
rect 67856 10166 67908 10218
rect 67960 10166 112024 10218
rect 112076 10166 112128 10218
rect 112180 10166 112232 10218
rect 112284 10166 156348 10218
rect 156400 10166 156452 10218
rect 156504 10166 156556 10218
rect 156608 10166 178640 10218
rect 1344 10132 178640 10166
rect 40462 10050 40514 10062
rect 40462 9986 40514 9998
rect 19070 9938 19122 9950
rect 19070 9874 19122 9886
rect 19518 9938 19570 9950
rect 19518 9874 19570 9886
rect 19966 9938 20018 9950
rect 23326 9938 23378 9950
rect 20850 9886 20862 9938
rect 20914 9886 20926 9938
rect 19966 9874 20018 9886
rect 23326 9874 23378 9886
rect 23774 9938 23826 9950
rect 23774 9874 23826 9886
rect 20526 9826 20578 9838
rect 20526 9762 20578 9774
rect 40574 9826 40626 9838
rect 40574 9762 40626 9774
rect 21646 9714 21698 9726
rect 21646 9650 21698 9662
rect 22542 9714 22594 9726
rect 22542 9650 22594 9662
rect 21758 9602 21810 9614
rect 21758 9538 21810 9550
rect 22654 9602 22706 9614
rect 22654 9538 22706 9550
rect 24222 9602 24274 9614
rect 24222 9538 24274 9550
rect 1344 9434 178800 9468
rect 1344 9382 45538 9434
rect 45590 9382 45642 9434
rect 45694 9382 45746 9434
rect 45798 9382 89862 9434
rect 89914 9382 89966 9434
rect 90018 9382 90070 9434
rect 90122 9382 134186 9434
rect 134238 9382 134290 9434
rect 134342 9382 134394 9434
rect 134446 9382 178510 9434
rect 178562 9382 178614 9434
rect 178666 9382 178718 9434
rect 178770 9382 178800 9434
rect 1344 9348 178800 9382
rect 20414 9266 20466 9278
rect 20414 9202 20466 9214
rect 22766 9266 22818 9278
rect 22766 9202 22818 9214
rect 93886 9266 93938 9278
rect 93886 9202 93938 9214
rect 94446 9266 94498 9278
rect 94446 9202 94498 9214
rect 21310 9154 21362 9166
rect 22206 9154 22258 9166
rect 20962 9102 20974 9154
rect 21026 9102 21038 9154
rect 21858 9102 21870 9154
rect 21922 9102 21934 9154
rect 21310 9090 21362 9102
rect 22206 9090 22258 9102
rect 23102 9154 23154 9166
rect 94770 9102 94782 9154
rect 94834 9102 94846 9154
rect 95890 9102 95902 9154
rect 95954 9102 95966 9154
rect 23102 9090 23154 9102
rect 95566 9042 95618 9054
rect 95566 8978 95618 8990
rect 1344 8650 178640 8684
rect 1344 8598 23376 8650
rect 23428 8598 23480 8650
rect 23532 8598 23584 8650
rect 23636 8598 67700 8650
rect 67752 8598 67804 8650
rect 67856 8598 67908 8650
rect 67960 8598 112024 8650
rect 112076 8598 112128 8650
rect 112180 8598 112232 8650
rect 112284 8598 156348 8650
rect 156400 8598 156452 8650
rect 156504 8598 156556 8650
rect 156608 8598 178640 8650
rect 1344 8564 178640 8598
rect 22542 8370 22594 8382
rect 22542 8306 22594 8318
rect 95342 8370 95394 8382
rect 95342 8306 95394 8318
rect 21646 8034 21698 8046
rect 21646 7970 21698 7982
rect 22094 8034 22146 8046
rect 22094 7970 22146 7982
rect 1344 7866 178800 7900
rect 1344 7814 45538 7866
rect 45590 7814 45642 7866
rect 45694 7814 45746 7866
rect 45798 7814 89862 7866
rect 89914 7814 89966 7866
rect 90018 7814 90070 7866
rect 90122 7814 134186 7866
rect 134238 7814 134290 7866
rect 134342 7814 134394 7866
rect 134446 7814 178510 7866
rect 178562 7814 178614 7866
rect 178666 7814 178718 7866
rect 178770 7814 178800 7866
rect 1344 7780 178800 7814
rect 1344 7082 178640 7116
rect 1344 7030 23376 7082
rect 23428 7030 23480 7082
rect 23532 7030 23584 7082
rect 23636 7030 67700 7082
rect 67752 7030 67804 7082
rect 67856 7030 67908 7082
rect 67960 7030 112024 7082
rect 112076 7030 112128 7082
rect 112180 7030 112232 7082
rect 112284 7030 156348 7082
rect 156400 7030 156452 7082
rect 156504 7030 156556 7082
rect 156608 7030 178640 7082
rect 1344 6996 178640 7030
rect 1344 6298 178800 6332
rect 1344 6246 45538 6298
rect 45590 6246 45642 6298
rect 45694 6246 45746 6298
rect 45798 6246 89862 6298
rect 89914 6246 89966 6298
rect 90018 6246 90070 6298
rect 90122 6246 134186 6298
rect 134238 6246 134290 6298
rect 134342 6246 134394 6298
rect 134446 6246 178510 6298
rect 178562 6246 178614 6298
rect 178666 6246 178718 6298
rect 178770 6246 178800 6298
rect 1344 6212 178800 6246
rect 1344 5514 178640 5548
rect 1344 5462 23376 5514
rect 23428 5462 23480 5514
rect 23532 5462 23584 5514
rect 23636 5462 67700 5514
rect 67752 5462 67804 5514
rect 67856 5462 67908 5514
rect 67960 5462 112024 5514
rect 112076 5462 112128 5514
rect 112180 5462 112232 5514
rect 112284 5462 156348 5514
rect 156400 5462 156452 5514
rect 156504 5462 156556 5514
rect 156608 5462 178640 5514
rect 1344 5428 178640 5462
rect 1344 4730 178800 4764
rect 1344 4678 45538 4730
rect 45590 4678 45642 4730
rect 45694 4678 45746 4730
rect 45798 4678 89862 4730
rect 89914 4678 89966 4730
rect 90018 4678 90070 4730
rect 90122 4678 134186 4730
rect 134238 4678 134290 4730
rect 134342 4678 134394 4730
rect 134446 4678 178510 4730
rect 178562 4678 178614 4730
rect 178666 4678 178718 4730
rect 178770 4678 178800 4730
rect 1344 4644 178800 4678
rect 1344 3946 178640 3980
rect 1344 3894 23376 3946
rect 23428 3894 23480 3946
rect 23532 3894 23584 3946
rect 23636 3894 67700 3946
rect 67752 3894 67804 3946
rect 67856 3894 67908 3946
rect 67960 3894 112024 3946
rect 112076 3894 112128 3946
rect 112180 3894 112232 3946
rect 112284 3894 156348 3946
rect 156400 3894 156452 3946
rect 156504 3894 156556 3946
rect 156608 3894 178640 3946
rect 1344 3860 178640 3894
rect 7310 3330 7362 3342
rect 7310 3266 7362 3278
rect 10670 3330 10722 3342
rect 10670 3266 10722 3278
rect 13582 3330 13634 3342
rect 13582 3266 13634 3278
rect 15150 3330 15202 3342
rect 15150 3266 15202 3278
rect 17502 3330 17554 3342
rect 17502 3266 17554 3278
rect 19630 3330 19682 3342
rect 19630 3266 19682 3278
rect 21422 3330 21474 3342
rect 21422 3266 21474 3278
rect 22990 3330 23042 3342
rect 22990 3266 23042 3278
rect 25342 3330 25394 3342
rect 25342 3266 25394 3278
rect 26350 3330 26402 3342
rect 26350 3266 26402 3278
rect 28030 3330 28082 3342
rect 28030 3266 28082 3278
rect 29710 3330 29762 3342
rect 29710 3266 29762 3278
rect 31390 3330 31442 3342
rect 31390 3266 31442 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 34750 3330 34802 3342
rect 34750 3266 34802 3278
rect 37102 3330 37154 3342
rect 37102 3266 37154 3278
rect 38110 3330 38162 3342
rect 38110 3266 38162 3278
rect 39790 3330 39842 3342
rect 39790 3266 39842 3278
rect 41470 3330 41522 3342
rect 41470 3266 41522 3278
rect 43150 3330 43202 3342
rect 43150 3266 43202 3278
rect 44942 3330 44994 3342
rect 44942 3266 44994 3278
rect 46510 3330 46562 3342
rect 46510 3266 46562 3278
rect 48862 3330 48914 3342
rect 48862 3266 48914 3278
rect 49870 3330 49922 3342
rect 49870 3266 49922 3278
rect 51550 3330 51602 3342
rect 51550 3266 51602 3278
rect 53230 3330 53282 3342
rect 53230 3266 53282 3278
rect 54910 3330 54962 3342
rect 54910 3266 54962 3278
rect 56702 3330 56754 3342
rect 56702 3266 56754 3278
rect 58270 3330 58322 3342
rect 58270 3266 58322 3278
rect 60622 3330 60674 3342
rect 60622 3266 60674 3278
rect 61630 3330 61682 3342
rect 61630 3266 61682 3278
rect 63310 3330 63362 3342
rect 63310 3266 63362 3278
rect 64990 3330 65042 3342
rect 64990 3266 65042 3278
rect 66110 3330 66162 3342
rect 66110 3266 66162 3278
rect 68462 3330 68514 3342
rect 68462 3266 68514 3278
rect 69470 3330 69522 3342
rect 69470 3266 69522 3278
rect 71150 3330 71202 3342
rect 71150 3266 71202 3278
rect 72830 3330 72882 3342
rect 72830 3266 72882 3278
rect 74510 3330 74562 3342
rect 74510 3266 74562 3278
rect 76302 3330 76354 3342
rect 76302 3266 76354 3278
rect 77870 3330 77922 3342
rect 77870 3266 77922 3278
rect 80222 3330 80274 3342
rect 80222 3266 80274 3278
rect 81230 3330 81282 3342
rect 81230 3266 81282 3278
rect 82910 3330 82962 3342
rect 82910 3266 82962 3278
rect 84590 3330 84642 3342
rect 84590 3266 84642 3278
rect 86270 3330 86322 3342
rect 86270 3266 86322 3278
rect 88062 3330 88114 3342
rect 88062 3266 88114 3278
rect 89630 3330 89682 3342
rect 89630 3266 89682 3278
rect 91982 3330 92034 3342
rect 91982 3266 92034 3278
rect 92990 3330 93042 3342
rect 92990 3266 93042 3278
rect 94670 3330 94722 3342
rect 94670 3266 94722 3278
rect 96350 3330 96402 3342
rect 96350 3266 96402 3278
rect 98030 3330 98082 3342
rect 98030 3266 98082 3278
rect 99822 3330 99874 3342
rect 99822 3266 99874 3278
rect 101390 3330 101442 3342
rect 101390 3266 101442 3278
rect 103742 3330 103794 3342
rect 103742 3266 103794 3278
rect 104750 3330 104802 3342
rect 104750 3266 104802 3278
rect 106430 3330 106482 3342
rect 106430 3266 106482 3278
rect 108110 3330 108162 3342
rect 108110 3266 108162 3278
rect 109790 3330 109842 3342
rect 109790 3266 109842 3278
rect 111582 3330 111634 3342
rect 111582 3266 111634 3278
rect 113150 3330 113202 3342
rect 113150 3266 113202 3278
rect 115502 3330 115554 3342
rect 115502 3266 115554 3278
rect 116510 3330 116562 3342
rect 116510 3266 116562 3278
rect 118190 3330 118242 3342
rect 118190 3266 118242 3278
rect 123342 3330 123394 3342
rect 123342 3266 123394 3278
rect 124910 3330 124962 3342
rect 124910 3266 124962 3278
rect 127262 3330 127314 3342
rect 127262 3266 127314 3278
rect 128270 3330 128322 3342
rect 128270 3266 128322 3278
rect 129950 3330 130002 3342
rect 129950 3266 130002 3278
rect 131630 3330 131682 3342
rect 131630 3266 131682 3278
rect 133310 3330 133362 3342
rect 133310 3266 133362 3278
rect 135102 3330 135154 3342
rect 135102 3266 135154 3278
rect 136670 3330 136722 3342
rect 136670 3266 136722 3278
rect 139022 3330 139074 3342
rect 139022 3266 139074 3278
rect 140030 3330 140082 3342
rect 140030 3266 140082 3278
rect 141710 3330 141762 3342
rect 141710 3266 141762 3278
rect 143390 3330 143442 3342
rect 143390 3266 143442 3278
rect 145070 3330 145122 3342
rect 145070 3266 145122 3278
rect 146862 3330 146914 3342
rect 146862 3266 146914 3278
rect 148430 3330 148482 3342
rect 148430 3266 148482 3278
rect 150782 3330 150834 3342
rect 150782 3266 150834 3278
rect 151790 3330 151842 3342
rect 151790 3266 151842 3278
rect 153470 3330 153522 3342
rect 153470 3266 153522 3278
rect 155150 3330 155202 3342
rect 155150 3266 155202 3278
rect 156830 3330 156882 3342
rect 156830 3266 156882 3278
rect 158622 3330 158674 3342
rect 158622 3266 158674 3278
rect 160190 3330 160242 3342
rect 160190 3266 160242 3278
rect 162542 3330 162594 3342
rect 162542 3266 162594 3278
rect 163550 3330 163602 3342
rect 163550 3266 163602 3278
rect 165230 3330 165282 3342
rect 165230 3266 165282 3278
rect 166910 3330 166962 3342
rect 166910 3266 166962 3278
rect 168590 3330 168642 3342
rect 168590 3266 168642 3278
rect 170382 3330 170434 3342
rect 170382 3266 170434 3278
rect 171950 3330 172002 3342
rect 171950 3266 172002 3278
rect 173070 3330 173122 3342
rect 173070 3266 173122 3278
rect 174302 3330 174354 3342
rect 174302 3266 174354 3278
rect 174974 3330 175026 3342
rect 174974 3266 175026 3278
rect 1344 3162 178800 3196
rect 1344 3110 45538 3162
rect 45590 3110 45642 3162
rect 45694 3110 45746 3162
rect 45798 3110 89862 3162
rect 89914 3110 89966 3162
rect 90018 3110 90070 3162
rect 90122 3110 134186 3162
rect 134238 3110 134290 3162
rect 134342 3110 134394 3162
rect 134446 3110 178510 3162
rect 178562 3110 178614 3162
rect 178666 3110 178718 3162
rect 178770 3110 178800 3162
rect 1344 3076 178800 3110
rect 67554 1710 67566 1762
rect 67618 1759 67630 1762
rect 68450 1759 68462 1762
rect 67618 1713 68462 1759
rect 67618 1710 67630 1713
rect 68450 1710 68462 1713
rect 68514 1710 68526 1762
rect 79314 1710 79326 1762
rect 79378 1759 79390 1762
rect 80210 1759 80222 1762
rect 79378 1713 80222 1759
rect 79378 1710 79390 1713
rect 80210 1710 80222 1713
rect 80274 1710 80286 1762
rect 91074 1710 91086 1762
rect 91138 1759 91150 1762
rect 91970 1759 91982 1762
rect 91138 1713 91982 1759
rect 91138 1710 91150 1713
rect 91970 1710 91982 1713
rect 92034 1710 92046 1762
rect 102834 1710 102846 1762
rect 102898 1759 102910 1762
rect 103730 1759 103742 1762
rect 102898 1713 103742 1759
rect 102898 1710 102910 1713
rect 103730 1710 103742 1713
rect 103794 1710 103806 1762
rect 114594 1710 114606 1762
rect 114658 1759 114670 1762
rect 115490 1759 115502 1762
rect 114658 1713 115502 1759
rect 114658 1710 114670 1713
rect 115490 1710 115502 1713
rect 115554 1710 115566 1762
rect 126354 1710 126366 1762
rect 126418 1759 126430 1762
rect 127250 1759 127262 1762
rect 126418 1713 127262 1759
rect 126418 1710 126430 1713
rect 127250 1710 127262 1713
rect 127314 1710 127326 1762
rect 138114 1710 138126 1762
rect 138178 1759 138190 1762
rect 139010 1759 139022 1762
rect 138178 1713 139022 1759
rect 138178 1710 138190 1713
rect 139010 1710 139022 1713
rect 139074 1710 139086 1762
rect 149874 1710 149886 1762
rect 149938 1759 149950 1762
rect 150770 1759 150782 1762
rect 149938 1713 150782 1759
rect 149938 1710 149950 1713
rect 150770 1710 150782 1713
rect 150834 1710 150846 1762
rect 161634 1710 161646 1762
rect 161698 1759 161710 1762
rect 162530 1759 162542 1762
rect 161698 1713 162542 1759
rect 161698 1710 161710 1713
rect 162530 1710 162542 1713
rect 162594 1710 162606 1762
rect 173394 1710 173406 1762
rect 173458 1759 173470 1762
rect 174290 1759 174302 1762
rect 173458 1713 174302 1759
rect 173458 1710 173470 1713
rect 174290 1710 174302 1713
rect 174354 1710 174366 1762
<< via1 >>
rect 18622 16606 18674 16658
rect 19182 16606 19234 16658
rect 20190 16606 20242 16658
rect 21422 16606 21474 16658
rect 29598 16606 29650 16658
rect 31390 16606 31442 16658
rect 35870 16606 35922 16658
rect 36430 16606 36482 16658
rect 37438 16606 37490 16658
rect 37998 16606 38050 16658
rect 44158 16606 44210 16658
rect 44942 16606 44994 16658
rect 23376 16438 23428 16490
rect 23480 16438 23532 16490
rect 23584 16438 23636 16490
rect 67700 16438 67752 16490
rect 67804 16438 67856 16490
rect 67908 16438 67960 16490
rect 112024 16438 112076 16490
rect 112128 16438 112180 16490
rect 112232 16438 112284 16490
rect 156348 16438 156400 16490
rect 156452 16438 156504 16490
rect 156556 16438 156608 16490
rect 5854 16158 5906 16210
rect 12574 16158 12626 16210
rect 15262 16158 15314 16210
rect 20190 16158 20242 16210
rect 24670 16158 24722 16210
rect 36318 16158 36370 16210
rect 38782 16158 38834 16210
rect 44158 16158 44210 16210
rect 48190 16158 48242 16210
rect 49870 16158 49922 16210
rect 51998 16158 52050 16210
rect 61630 16158 61682 16210
rect 63758 16158 63810 16210
rect 94894 16158 94946 16210
rect 1822 16046 1874 16098
rect 6302 16046 6354 16098
rect 9774 16046 9826 16098
rect 15710 16046 15762 16098
rect 17502 16046 17554 16098
rect 18622 16046 18674 16098
rect 21422 16046 21474 16098
rect 25342 16046 25394 16098
rect 29150 16046 29202 16098
rect 30606 16046 30658 16098
rect 31390 16046 31442 16098
rect 33518 16046 33570 16098
rect 39230 16046 39282 16098
rect 44942 16046 44994 16098
rect 49198 16046 49250 16098
rect 52782 16046 52834 16098
rect 54238 16046 54290 16098
rect 60846 16046 60898 16098
rect 91982 16046 92034 16098
rect 3166 15934 3218 15986
rect 4734 15934 4786 15986
rect 6638 15934 6690 15986
rect 7870 15934 7922 15986
rect 8878 15934 8930 15986
rect 10446 15934 10498 15986
rect 14142 15934 14194 15986
rect 16718 15934 16770 15986
rect 19182 15934 19234 15986
rect 22318 15934 22370 15986
rect 23550 15934 23602 15986
rect 25678 15934 25730 15986
rect 26686 15934 26738 15986
rect 28254 15934 28306 15986
rect 30046 15934 30098 15986
rect 31726 15934 31778 15986
rect 32398 15934 32450 15986
rect 34190 15934 34242 15986
rect 37102 15934 37154 15986
rect 37438 15934 37490 15986
rect 37998 15934 38050 15986
rect 41022 15934 41074 15986
rect 42366 15934 42418 15986
rect 45838 15934 45890 15986
rect 47070 15934 47122 15986
rect 53566 15934 53618 15986
rect 54910 15934 54962 15986
rect 56702 15934 56754 15986
rect 59614 15934 59666 15986
rect 65886 15934 65938 15986
rect 66558 15934 66610 15986
rect 69022 15934 69074 15986
rect 70590 15934 70642 15986
rect 73054 15934 73106 15986
rect 75294 15934 75346 15986
rect 78430 15934 78482 15986
rect 80222 15934 80274 15986
rect 83134 15934 83186 15986
rect 84702 15934 84754 15986
rect 88062 15934 88114 15986
rect 89294 15934 89346 15986
rect 92766 15934 92818 15986
rect 97246 15934 97298 15986
rect 98814 15934 98866 15986
rect 101950 15934 102002 15986
rect 103742 15934 103794 15986
rect 106654 15934 106706 15986
rect 108222 15934 108274 15986
rect 111582 15934 111634 15986
rect 112926 15934 112978 15986
rect 116062 15934 116114 15986
rect 117630 15934 117682 15986
rect 120766 15934 120818 15986
rect 122334 15934 122386 15986
rect 125470 15934 125522 15986
rect 127262 15934 127314 15986
rect 130174 15934 130226 15986
rect 131742 15934 131794 15986
rect 135102 15934 135154 15986
rect 136446 15934 136498 15986
rect 139582 15934 139634 15986
rect 141150 15934 141202 15986
rect 144286 15934 144338 15986
rect 145854 15934 145906 15986
rect 148990 15934 149042 15986
rect 150782 15934 150834 15986
rect 153694 15934 153746 15986
rect 155262 15934 155314 15986
rect 158622 15934 158674 15986
rect 159966 15934 160018 15986
rect 163102 15934 163154 15986
rect 164670 15934 164722 15986
rect 167806 15934 167858 15986
rect 169374 15934 169426 15986
rect 172510 15934 172562 15986
rect 174302 15934 174354 15986
rect 177214 15934 177266 15986
rect 2158 15822 2210 15874
rect 13470 15822 13522 15874
rect 16046 15822 16098 15874
rect 18062 15822 18114 15874
rect 19742 15822 19794 15874
rect 20750 15822 20802 15874
rect 21758 15822 21810 15874
rect 27694 15822 27746 15874
rect 39566 15822 39618 15874
rect 45278 15822 45330 15874
rect 64654 15822 64706 15874
rect 73726 15822 73778 15874
rect 74398 15822 74450 15874
rect 90078 15822 90130 15874
rect 90638 15822 90690 15874
rect 91198 15822 91250 15874
rect 45538 15654 45590 15706
rect 45642 15654 45694 15706
rect 45746 15654 45798 15706
rect 89862 15654 89914 15706
rect 89966 15654 90018 15706
rect 90070 15654 90122 15706
rect 134186 15654 134238 15706
rect 134290 15654 134342 15706
rect 134394 15654 134446 15706
rect 178510 15654 178562 15706
rect 178614 15654 178666 15706
rect 178718 15654 178770 15706
rect 1822 15486 1874 15538
rect 14702 15486 14754 15538
rect 16046 15486 16098 15538
rect 16718 15486 16770 15538
rect 26238 15486 26290 15538
rect 32398 15486 32450 15538
rect 36430 15486 36482 15538
rect 37102 15486 37154 15538
rect 37438 15486 37490 15538
rect 48526 15486 48578 15538
rect 50206 15486 50258 15538
rect 51326 15486 51378 15538
rect 60062 15486 60114 15538
rect 60622 15486 60674 15538
rect 61182 15486 61234 15538
rect 76526 15486 76578 15538
rect 76974 15486 77026 15538
rect 91758 15486 91810 15538
rect 92542 15486 92594 15538
rect 94110 15486 94162 15538
rect 178110 15486 178162 15538
rect 10782 15374 10834 15426
rect 12126 15374 12178 15426
rect 16606 15374 16658 15426
rect 20302 15374 20354 15426
rect 20862 15374 20914 15426
rect 22094 15374 22146 15426
rect 22990 15374 23042 15426
rect 27582 15374 27634 15426
rect 35086 15374 35138 15426
rect 54014 15374 54066 15426
rect 63758 15374 63810 15426
rect 65438 15374 65490 15426
rect 79662 15374 79714 15426
rect 10558 15262 10610 15314
rect 11454 15262 11506 15314
rect 17726 15262 17778 15314
rect 19406 15262 19458 15314
rect 26910 15262 26962 15314
rect 30494 15262 30546 15314
rect 31726 15262 31778 15314
rect 33742 15262 33794 15314
rect 34190 15262 34242 15314
rect 35870 15262 35922 15314
rect 51998 15262 52050 15314
rect 53566 15262 53618 15314
rect 63198 15262 63250 15314
rect 64654 15262 64706 15314
rect 73614 15262 73666 15314
rect 74846 15262 74898 15314
rect 80446 15262 80498 15314
rect 89518 15262 89570 15314
rect 90750 15262 90802 15314
rect 14254 15150 14306 15202
rect 18510 15150 18562 15202
rect 19742 15150 19794 15202
rect 21198 15150 21250 15202
rect 21758 15150 21810 15202
rect 22654 15150 22706 15202
rect 23550 15150 23602 15202
rect 29710 15150 29762 15202
rect 31054 15150 31106 15202
rect 52670 15150 52722 15202
rect 74174 15150 74226 15202
rect 77534 15150 77586 15202
rect 90078 15150 90130 15202
rect 23376 14870 23428 14922
rect 23480 14870 23532 14922
rect 23584 14870 23636 14922
rect 67700 14870 67752 14922
rect 67804 14870 67856 14922
rect 67908 14870 67960 14922
rect 112024 14870 112076 14922
rect 112128 14870 112180 14922
rect 112232 14870 112284 14922
rect 156348 14870 156400 14922
rect 156452 14870 156504 14922
rect 156556 14870 156608 14922
rect 11006 14590 11058 14642
rect 19518 14590 19570 14642
rect 20526 14590 20578 14642
rect 23438 14590 23490 14642
rect 30046 14590 30098 14642
rect 30382 14590 30434 14642
rect 31166 14590 31218 14642
rect 33182 14590 33234 14642
rect 33742 14590 33794 14642
rect 35086 14590 35138 14642
rect 88958 14590 89010 14642
rect 15374 14478 15426 14530
rect 16830 14478 16882 14530
rect 17502 14478 17554 14530
rect 18958 14478 19010 14530
rect 34190 14478 34242 14530
rect 35870 14478 35922 14530
rect 63198 14478 63250 14530
rect 64542 14478 64594 14530
rect 72718 14478 72770 14530
rect 73950 14478 74002 14530
rect 88398 14478 88450 14530
rect 89854 14478 89906 14530
rect 12574 14366 12626 14418
rect 15934 14366 15986 14418
rect 18062 14366 18114 14418
rect 20862 14366 20914 14418
rect 23214 14366 23266 14418
rect 53678 14366 53730 14418
rect 63758 14366 63810 14418
rect 73278 14366 73330 14418
rect 19966 14254 20018 14306
rect 21870 14254 21922 14306
rect 22654 14254 22706 14306
rect 23998 14254 24050 14306
rect 45538 14086 45590 14138
rect 45642 14086 45694 14138
rect 45746 14086 45798 14138
rect 89862 14086 89914 14138
rect 89966 14086 90018 14138
rect 90070 14086 90122 14138
rect 134186 14086 134238 14138
rect 134290 14086 134342 14138
rect 134394 14086 134446 14138
rect 178510 14086 178562 14138
rect 178614 14086 178666 14138
rect 178718 14086 178770 14138
rect 16606 13918 16658 13970
rect 16942 13918 16994 13970
rect 21310 13806 21362 13858
rect 19294 13694 19346 13746
rect 21870 13694 21922 13746
rect 61630 13694 61682 13746
rect 17726 13582 17778 13634
rect 18174 13582 18226 13634
rect 18622 13582 18674 13634
rect 19518 13582 19570 13634
rect 20078 13582 20130 13634
rect 20414 13582 20466 13634
rect 20974 13582 21026 13634
rect 23774 13582 23826 13634
rect 24894 13582 24946 13634
rect 61742 13470 61794 13522
rect 23376 13302 23428 13354
rect 23480 13302 23532 13354
rect 23584 13302 23636 13354
rect 67700 13302 67752 13354
rect 67804 13302 67856 13354
rect 67908 13302 67960 13354
rect 112024 13302 112076 13354
rect 112128 13302 112180 13354
rect 112232 13302 112284 13354
rect 156348 13302 156400 13354
rect 156452 13302 156504 13354
rect 156556 13302 156608 13354
rect 26350 13134 26402 13186
rect 63198 13134 63250 13186
rect 18734 13022 18786 13074
rect 18958 13022 19010 13074
rect 19630 13022 19682 13074
rect 19854 13022 19906 13074
rect 20862 13022 20914 13074
rect 22766 13022 22818 13074
rect 24782 13022 24834 13074
rect 25006 13022 25058 13074
rect 25566 13022 25618 13074
rect 16382 12910 16434 12962
rect 17838 12910 17890 12962
rect 21870 12910 21922 12962
rect 17166 12798 17218 12850
rect 20526 12798 20578 12850
rect 26462 12798 26514 12850
rect 40238 12798 40290 12850
rect 40798 12798 40850 12850
rect 63086 12798 63138 12850
rect 40910 12686 40962 12738
rect 61742 12686 61794 12738
rect 62414 12686 62466 12738
rect 45538 12518 45590 12570
rect 45642 12518 45694 12570
rect 45746 12518 45798 12570
rect 89862 12518 89914 12570
rect 89966 12518 90018 12570
rect 90070 12518 90122 12570
rect 134186 12518 134238 12570
rect 134290 12518 134342 12570
rect 134394 12518 134446 12570
rect 178510 12518 178562 12570
rect 178614 12518 178666 12570
rect 178718 12518 178770 12570
rect 17726 12350 17778 12402
rect 19294 12350 19346 12402
rect 20974 12350 21026 12402
rect 23662 12350 23714 12402
rect 24558 12350 24610 12402
rect 26238 12350 26290 12402
rect 26798 12350 26850 12402
rect 27134 12350 27186 12402
rect 39230 12350 39282 12402
rect 60958 12350 61010 12402
rect 62302 12350 62354 12402
rect 16942 12238 16994 12290
rect 18510 12238 18562 12290
rect 19406 12238 19458 12290
rect 19966 12238 20018 12290
rect 20302 12238 20354 12290
rect 22654 12238 22706 12290
rect 22990 12238 23042 12290
rect 25678 12238 25730 12290
rect 27694 12238 27746 12290
rect 39342 12238 39394 12290
rect 39902 12238 39954 12290
rect 40574 12238 40626 12290
rect 41582 12238 41634 12290
rect 60286 12238 60338 12290
rect 61518 12238 61570 12290
rect 63198 12238 63250 12290
rect 63870 12238 63922 12290
rect 16158 12126 16210 12178
rect 16606 12126 16658 12178
rect 18174 12126 18226 12178
rect 22094 12126 22146 12178
rect 23662 12126 23714 12178
rect 20862 12014 20914 12066
rect 21758 12014 21810 12066
rect 24446 12014 24498 12066
rect 25902 11902 25954 11954
rect 60174 11902 60226 11954
rect 23376 11734 23428 11786
rect 23480 11734 23532 11786
rect 23584 11734 23636 11786
rect 67700 11734 67752 11786
rect 67804 11734 67856 11786
rect 67908 11734 67960 11786
rect 112024 11734 112076 11786
rect 112128 11734 112180 11786
rect 112232 11734 112284 11786
rect 156348 11734 156400 11786
rect 156452 11734 156504 11786
rect 156556 11734 156608 11786
rect 25790 11566 25842 11618
rect 26462 11566 26514 11618
rect 39342 11566 39394 11618
rect 40014 11566 40066 11618
rect 42142 11566 42194 11618
rect 51774 11566 51826 11618
rect 60510 11566 60562 11618
rect 61406 11566 61458 11618
rect 62974 11566 63026 11618
rect 63646 11566 63698 11618
rect 17278 11454 17330 11506
rect 17838 11454 17890 11506
rect 18174 11454 18226 11506
rect 18734 11454 18786 11506
rect 18958 11454 19010 11506
rect 19630 11454 19682 11506
rect 19854 11454 19906 11506
rect 22094 11454 22146 11506
rect 22990 11454 23042 11506
rect 23886 11454 23938 11506
rect 52446 11454 52498 11506
rect 53454 11454 53506 11506
rect 25902 11342 25954 11394
rect 26574 11342 26626 11394
rect 40126 11342 40178 11394
rect 51886 11342 51938 11394
rect 60622 11342 60674 11394
rect 61518 11342 61570 11394
rect 63086 11342 63138 11394
rect 63758 11342 63810 11394
rect 20526 11230 20578 11282
rect 21758 11230 21810 11282
rect 22654 11230 22706 11282
rect 23550 11230 23602 11282
rect 39454 11230 39506 11282
rect 40686 11230 40738 11282
rect 41470 11230 41522 11282
rect 42030 11230 42082 11282
rect 20638 11118 20690 11170
rect 24334 11118 24386 11170
rect 24782 11118 24834 11170
rect 42702 11118 42754 11170
rect 62078 11118 62130 11170
rect 45538 10950 45590 11002
rect 45642 10950 45694 11002
rect 45746 10950 45798 11002
rect 89862 10950 89914 11002
rect 89966 10950 90018 11002
rect 90070 10950 90122 11002
rect 134186 10950 134238 11002
rect 134290 10950 134342 11002
rect 134394 10950 134446 11002
rect 178510 10950 178562 11002
rect 178614 10950 178666 11002
rect 178718 10950 178770 11002
rect 18062 10782 18114 10834
rect 18510 10782 18562 10834
rect 19182 10782 19234 10834
rect 20974 10782 21026 10834
rect 39790 10782 39842 10834
rect 40462 10782 40514 10834
rect 52334 10782 52386 10834
rect 61854 10782 61906 10834
rect 19966 10670 20018 10722
rect 20302 10670 20354 10722
rect 22094 10670 22146 10722
rect 22990 10670 23042 10722
rect 39902 10670 39954 10722
rect 40574 10670 40626 10722
rect 41582 10670 41634 10722
rect 52446 10670 52498 10722
rect 61966 10670 62018 10722
rect 21870 10558 21922 10610
rect 22654 10558 22706 10610
rect 23438 10558 23490 10610
rect 24110 10558 24162 10610
rect 24558 10558 24610 10610
rect 19070 10446 19122 10498
rect 20862 10446 20914 10498
rect 23376 10166 23428 10218
rect 23480 10166 23532 10218
rect 23584 10166 23636 10218
rect 67700 10166 67752 10218
rect 67804 10166 67856 10218
rect 67908 10166 67960 10218
rect 112024 10166 112076 10218
rect 112128 10166 112180 10218
rect 112232 10166 112284 10218
rect 156348 10166 156400 10218
rect 156452 10166 156504 10218
rect 156556 10166 156608 10218
rect 40462 9998 40514 10050
rect 19070 9886 19122 9938
rect 19518 9886 19570 9938
rect 19966 9886 20018 9938
rect 20862 9886 20914 9938
rect 23326 9886 23378 9938
rect 23774 9886 23826 9938
rect 20526 9774 20578 9826
rect 40574 9774 40626 9826
rect 21646 9662 21698 9714
rect 22542 9662 22594 9714
rect 21758 9550 21810 9602
rect 22654 9550 22706 9602
rect 24222 9550 24274 9602
rect 45538 9382 45590 9434
rect 45642 9382 45694 9434
rect 45746 9382 45798 9434
rect 89862 9382 89914 9434
rect 89966 9382 90018 9434
rect 90070 9382 90122 9434
rect 134186 9382 134238 9434
rect 134290 9382 134342 9434
rect 134394 9382 134446 9434
rect 178510 9382 178562 9434
rect 178614 9382 178666 9434
rect 178718 9382 178770 9434
rect 20414 9214 20466 9266
rect 22766 9214 22818 9266
rect 93886 9214 93938 9266
rect 94446 9214 94498 9266
rect 20974 9102 21026 9154
rect 21310 9102 21362 9154
rect 21870 9102 21922 9154
rect 22206 9102 22258 9154
rect 23102 9102 23154 9154
rect 94782 9102 94834 9154
rect 95902 9102 95954 9154
rect 95566 8990 95618 9042
rect 23376 8598 23428 8650
rect 23480 8598 23532 8650
rect 23584 8598 23636 8650
rect 67700 8598 67752 8650
rect 67804 8598 67856 8650
rect 67908 8598 67960 8650
rect 112024 8598 112076 8650
rect 112128 8598 112180 8650
rect 112232 8598 112284 8650
rect 156348 8598 156400 8650
rect 156452 8598 156504 8650
rect 156556 8598 156608 8650
rect 22542 8318 22594 8370
rect 95342 8318 95394 8370
rect 21646 7982 21698 8034
rect 22094 7982 22146 8034
rect 45538 7814 45590 7866
rect 45642 7814 45694 7866
rect 45746 7814 45798 7866
rect 89862 7814 89914 7866
rect 89966 7814 90018 7866
rect 90070 7814 90122 7866
rect 134186 7814 134238 7866
rect 134290 7814 134342 7866
rect 134394 7814 134446 7866
rect 178510 7814 178562 7866
rect 178614 7814 178666 7866
rect 178718 7814 178770 7866
rect 23376 7030 23428 7082
rect 23480 7030 23532 7082
rect 23584 7030 23636 7082
rect 67700 7030 67752 7082
rect 67804 7030 67856 7082
rect 67908 7030 67960 7082
rect 112024 7030 112076 7082
rect 112128 7030 112180 7082
rect 112232 7030 112284 7082
rect 156348 7030 156400 7082
rect 156452 7030 156504 7082
rect 156556 7030 156608 7082
rect 45538 6246 45590 6298
rect 45642 6246 45694 6298
rect 45746 6246 45798 6298
rect 89862 6246 89914 6298
rect 89966 6246 90018 6298
rect 90070 6246 90122 6298
rect 134186 6246 134238 6298
rect 134290 6246 134342 6298
rect 134394 6246 134446 6298
rect 178510 6246 178562 6298
rect 178614 6246 178666 6298
rect 178718 6246 178770 6298
rect 23376 5462 23428 5514
rect 23480 5462 23532 5514
rect 23584 5462 23636 5514
rect 67700 5462 67752 5514
rect 67804 5462 67856 5514
rect 67908 5462 67960 5514
rect 112024 5462 112076 5514
rect 112128 5462 112180 5514
rect 112232 5462 112284 5514
rect 156348 5462 156400 5514
rect 156452 5462 156504 5514
rect 156556 5462 156608 5514
rect 45538 4678 45590 4730
rect 45642 4678 45694 4730
rect 45746 4678 45798 4730
rect 89862 4678 89914 4730
rect 89966 4678 90018 4730
rect 90070 4678 90122 4730
rect 134186 4678 134238 4730
rect 134290 4678 134342 4730
rect 134394 4678 134446 4730
rect 178510 4678 178562 4730
rect 178614 4678 178666 4730
rect 178718 4678 178770 4730
rect 23376 3894 23428 3946
rect 23480 3894 23532 3946
rect 23584 3894 23636 3946
rect 67700 3894 67752 3946
rect 67804 3894 67856 3946
rect 67908 3894 67960 3946
rect 112024 3894 112076 3946
rect 112128 3894 112180 3946
rect 112232 3894 112284 3946
rect 156348 3894 156400 3946
rect 156452 3894 156504 3946
rect 156556 3894 156608 3946
rect 7310 3278 7362 3330
rect 10670 3278 10722 3330
rect 13582 3278 13634 3330
rect 15150 3278 15202 3330
rect 17502 3278 17554 3330
rect 19630 3278 19682 3330
rect 21422 3278 21474 3330
rect 22990 3278 23042 3330
rect 25342 3278 25394 3330
rect 26350 3278 26402 3330
rect 28030 3278 28082 3330
rect 29710 3278 29762 3330
rect 31390 3278 31442 3330
rect 33182 3278 33234 3330
rect 34750 3278 34802 3330
rect 37102 3278 37154 3330
rect 38110 3278 38162 3330
rect 39790 3278 39842 3330
rect 41470 3278 41522 3330
rect 43150 3278 43202 3330
rect 44942 3278 44994 3330
rect 46510 3278 46562 3330
rect 48862 3278 48914 3330
rect 49870 3278 49922 3330
rect 51550 3278 51602 3330
rect 53230 3278 53282 3330
rect 54910 3278 54962 3330
rect 56702 3278 56754 3330
rect 58270 3278 58322 3330
rect 60622 3278 60674 3330
rect 61630 3278 61682 3330
rect 63310 3278 63362 3330
rect 64990 3278 65042 3330
rect 66110 3278 66162 3330
rect 68462 3278 68514 3330
rect 69470 3278 69522 3330
rect 71150 3278 71202 3330
rect 72830 3278 72882 3330
rect 74510 3278 74562 3330
rect 76302 3278 76354 3330
rect 77870 3278 77922 3330
rect 80222 3278 80274 3330
rect 81230 3278 81282 3330
rect 82910 3278 82962 3330
rect 84590 3278 84642 3330
rect 86270 3278 86322 3330
rect 88062 3278 88114 3330
rect 89630 3278 89682 3330
rect 91982 3278 92034 3330
rect 92990 3278 93042 3330
rect 94670 3278 94722 3330
rect 96350 3278 96402 3330
rect 98030 3278 98082 3330
rect 99822 3278 99874 3330
rect 101390 3278 101442 3330
rect 103742 3278 103794 3330
rect 104750 3278 104802 3330
rect 106430 3278 106482 3330
rect 108110 3278 108162 3330
rect 109790 3278 109842 3330
rect 111582 3278 111634 3330
rect 113150 3278 113202 3330
rect 115502 3278 115554 3330
rect 116510 3278 116562 3330
rect 118190 3278 118242 3330
rect 123342 3278 123394 3330
rect 124910 3278 124962 3330
rect 127262 3278 127314 3330
rect 128270 3278 128322 3330
rect 129950 3278 130002 3330
rect 131630 3278 131682 3330
rect 133310 3278 133362 3330
rect 135102 3278 135154 3330
rect 136670 3278 136722 3330
rect 139022 3278 139074 3330
rect 140030 3278 140082 3330
rect 141710 3278 141762 3330
rect 143390 3278 143442 3330
rect 145070 3278 145122 3330
rect 146862 3278 146914 3330
rect 148430 3278 148482 3330
rect 150782 3278 150834 3330
rect 151790 3278 151842 3330
rect 153470 3278 153522 3330
rect 155150 3278 155202 3330
rect 156830 3278 156882 3330
rect 158622 3278 158674 3330
rect 160190 3278 160242 3330
rect 162542 3278 162594 3330
rect 163550 3278 163602 3330
rect 165230 3278 165282 3330
rect 166910 3278 166962 3330
rect 168590 3278 168642 3330
rect 170382 3278 170434 3330
rect 171950 3278 172002 3330
rect 173070 3278 173122 3330
rect 174302 3278 174354 3330
rect 174974 3278 175026 3330
rect 45538 3110 45590 3162
rect 45642 3110 45694 3162
rect 45746 3110 45798 3162
rect 89862 3110 89914 3162
rect 89966 3110 90018 3162
rect 90070 3110 90122 3162
rect 134186 3110 134238 3162
rect 134290 3110 134342 3162
rect 134394 3110 134446 3162
rect 178510 3110 178562 3162
rect 178614 3110 178666 3162
rect 178718 3110 178770 3162
rect 67566 1710 67618 1762
rect 68462 1710 68514 1762
rect 79326 1710 79378 1762
rect 80222 1710 80274 1762
rect 91086 1710 91138 1762
rect 91982 1710 92034 1762
rect 102846 1710 102898 1762
rect 103742 1710 103794 1762
rect 114606 1710 114658 1762
rect 115502 1710 115554 1762
rect 126366 1710 126418 1762
rect 127262 1710 127314 1762
rect 138126 1710 138178 1762
rect 139022 1710 139074 1762
rect 149886 1710 149938 1762
rect 150782 1710 150834 1762
rect 161646 1710 161698 1762
rect 162542 1710 162594 1762
rect 173406 1710 173458 1762
rect 174302 1710 174354 1762
<< metal2 >>
rect 1344 19200 1456 20000
rect 2912 19200 3024 20000
rect 4480 19200 4592 20000
rect 6048 19200 6160 20000
rect 7616 19200 7728 20000
rect 9184 19200 9296 20000
rect 10752 19200 10864 20000
rect 12320 19200 12432 20000
rect 13888 19200 14000 20000
rect 15456 19200 15568 20000
rect 17024 19200 17136 20000
rect 18592 19200 18704 20000
rect 20160 19200 20272 20000
rect 21728 19200 21840 20000
rect 23296 19200 23408 20000
rect 24864 19200 24976 20000
rect 26432 19200 26544 20000
rect 28000 19200 28112 20000
rect 29568 19200 29680 20000
rect 31136 19200 31248 20000
rect 32704 19200 32816 20000
rect 34272 19200 34384 20000
rect 35840 19200 35952 20000
rect 37408 19200 37520 20000
rect 38976 19200 39088 20000
rect 40544 19200 40656 20000
rect 42112 19200 42224 20000
rect 43680 19200 43792 20000
rect 45248 19200 45360 20000
rect 46816 19200 46928 20000
rect 48384 19200 48496 20000
rect 49952 19200 50064 20000
rect 51520 19200 51632 20000
rect 53088 19200 53200 20000
rect 54656 19200 54768 20000
rect 56224 19200 56336 20000
rect 57792 19200 57904 20000
rect 59360 19200 59472 20000
rect 60928 19200 61040 20000
rect 62496 19200 62608 20000
rect 64064 19200 64176 20000
rect 65632 19200 65744 20000
rect 67200 19200 67312 20000
rect 68768 19200 68880 20000
rect 70336 19200 70448 20000
rect 71904 19200 72016 20000
rect 73472 19200 73584 20000
rect 75040 19200 75152 20000
rect 76608 19200 76720 20000
rect 78176 19200 78288 20000
rect 79744 19200 79856 20000
rect 81312 19200 81424 20000
rect 82880 19200 82992 20000
rect 84448 19200 84560 20000
rect 86016 19200 86128 20000
rect 87584 19200 87696 20000
rect 89152 19200 89264 20000
rect 90720 19200 90832 20000
rect 92288 19200 92400 20000
rect 93856 19200 93968 20000
rect 95424 19200 95536 20000
rect 96992 19200 97104 20000
rect 98560 19200 98672 20000
rect 100128 19200 100240 20000
rect 101696 19200 101808 20000
rect 103264 19200 103376 20000
rect 104832 19200 104944 20000
rect 106400 19200 106512 20000
rect 107968 19200 108080 20000
rect 109536 19200 109648 20000
rect 111104 19200 111216 20000
rect 112672 19200 112784 20000
rect 114240 19200 114352 20000
rect 115808 19200 115920 20000
rect 117376 19200 117488 20000
rect 118944 19200 119056 20000
rect 120512 19200 120624 20000
rect 122080 19200 122192 20000
rect 123648 19200 123760 20000
rect 125216 19200 125328 20000
rect 126784 19200 126896 20000
rect 128352 19200 128464 20000
rect 129920 19200 130032 20000
rect 131488 19200 131600 20000
rect 133056 19200 133168 20000
rect 134624 19200 134736 20000
rect 136192 19200 136304 20000
rect 137760 19200 137872 20000
rect 139328 19200 139440 20000
rect 140896 19200 141008 20000
rect 142464 19200 142576 20000
rect 144032 19200 144144 20000
rect 145600 19200 145712 20000
rect 147168 19200 147280 20000
rect 148736 19200 148848 20000
rect 150304 19200 150416 20000
rect 151872 19200 151984 20000
rect 153440 19200 153552 20000
rect 155008 19200 155120 20000
rect 156576 19200 156688 20000
rect 158144 19200 158256 20000
rect 159712 19200 159824 20000
rect 161280 19200 161392 20000
rect 162848 19200 162960 20000
rect 164416 19200 164528 20000
rect 165984 19200 166096 20000
rect 167552 19200 167664 20000
rect 169120 19200 169232 20000
rect 170688 19200 170800 20000
rect 172256 19200 172368 20000
rect 173824 19200 173936 20000
rect 175392 19200 175504 20000
rect 176960 19200 177072 20000
rect 178528 19200 178640 20000
rect 1372 16548 1428 19200
rect 1372 16492 1876 16548
rect 1820 16098 1876 16492
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1820 15538 1876 16046
rect 2940 15988 2996 19200
rect 3164 15988 3220 15998
rect 2940 15986 3220 15988
rect 2940 15934 3166 15986
rect 3218 15934 3220 15986
rect 2940 15932 3220 15934
rect 4508 15988 4564 19200
rect 5852 16212 5908 16222
rect 6076 16212 6132 19200
rect 5852 16210 6356 16212
rect 5852 16158 5854 16210
rect 5906 16158 6356 16210
rect 5852 16156 6356 16158
rect 5852 16146 5908 16156
rect 6300 16098 6356 16156
rect 6300 16046 6302 16098
rect 6354 16046 6356 16098
rect 6300 16034 6356 16046
rect 4732 15988 4788 15998
rect 4508 15986 4788 15988
rect 4508 15934 4734 15986
rect 4786 15934 4788 15986
rect 4508 15932 4788 15934
rect 3164 15922 3220 15932
rect 4732 15922 4788 15932
rect 6636 15988 6692 15998
rect 7644 15988 7700 19200
rect 7868 15988 7924 15998
rect 7644 15986 7924 15988
rect 7644 15934 7870 15986
rect 7922 15934 7924 15986
rect 7644 15932 7924 15934
rect 6636 15894 6692 15932
rect 7868 15922 7924 15932
rect 8876 15988 8932 15998
rect 9212 15988 9268 19200
rect 10780 16324 10836 19200
rect 10556 16268 10836 16324
rect 8876 15986 9268 15988
rect 8876 15934 8878 15986
rect 8930 15934 9268 15986
rect 8876 15932 9268 15934
rect 9772 16098 9828 16110
rect 9772 16046 9774 16098
rect 9826 16046 9828 16098
rect 8876 15922 8932 15932
rect 2156 15876 2212 15886
rect 2156 15782 2212 15820
rect 9772 15652 9828 16046
rect 10444 15988 10500 15998
rect 10444 15894 10500 15932
rect 9772 15586 9828 15596
rect 1820 15486 1822 15538
rect 1874 15486 1876 15538
rect 1820 15474 1876 15486
rect 10556 15316 10612 16268
rect 11452 15652 11508 15662
rect 10780 15428 10836 15438
rect 10780 15334 10836 15372
rect 10556 15314 10724 15316
rect 10556 15262 10558 15314
rect 10610 15262 10724 15314
rect 10556 15260 10724 15262
rect 10556 15250 10612 15260
rect 10668 14756 10724 15260
rect 11452 15314 11508 15596
rect 12124 15428 12180 15438
rect 12124 15334 12180 15372
rect 11452 15262 11454 15314
rect 11506 15262 11508 15314
rect 11452 15250 11508 15262
rect 10668 14700 11060 14756
rect 11004 14642 11060 14700
rect 11004 14590 11006 14642
rect 11058 14590 11060 14642
rect 11004 14578 11060 14590
rect 12348 14420 12404 19200
rect 12572 16212 12628 16222
rect 12572 16118 12628 16156
rect 13916 15988 13972 19200
rect 15260 16212 15316 16222
rect 15484 16212 15540 19200
rect 17052 16660 17108 19200
rect 16716 16604 17108 16660
rect 18620 16658 18676 19200
rect 18620 16606 18622 16658
rect 18674 16606 18676 16658
rect 15260 16210 15764 16212
rect 15260 16158 15262 16210
rect 15314 16158 15764 16210
rect 15260 16156 15764 16158
rect 15260 16146 15316 16156
rect 15708 16098 15764 16156
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 16034 15764 16046
rect 14140 15988 14196 15998
rect 13916 15986 14196 15988
rect 13916 15934 14142 15986
rect 14194 15934 14196 15986
rect 13916 15932 14196 15934
rect 14140 15922 14196 15932
rect 16716 15986 16772 16604
rect 18620 16594 18676 16606
rect 19180 16658 19236 16670
rect 19180 16606 19182 16658
rect 19234 16606 19236 16658
rect 17724 16212 17780 16222
rect 16716 15934 16718 15986
rect 16770 15934 16772 15986
rect 16716 15922 16772 15934
rect 16828 16100 16884 16110
rect 13468 15874 13524 15886
rect 13468 15822 13470 15874
rect 13522 15822 13524 15874
rect 13468 15652 13524 15822
rect 15932 15876 15988 15886
rect 13468 15586 13524 15596
rect 14700 15652 14756 15662
rect 14700 15538 14756 15596
rect 14700 15486 14702 15538
rect 14754 15486 14756 15538
rect 14700 15474 14756 15486
rect 15932 15540 15988 15820
rect 16044 15874 16100 15886
rect 16044 15822 16046 15874
rect 16098 15822 16100 15874
rect 16044 15764 16100 15822
rect 16044 15698 16100 15708
rect 16044 15540 16100 15550
rect 15932 15538 16100 15540
rect 15932 15486 16046 15538
rect 16098 15486 16100 15538
rect 15932 15484 16100 15486
rect 16044 15428 16100 15484
rect 16716 15540 16772 15550
rect 16716 15446 16772 15484
rect 16044 15362 16100 15372
rect 16604 15428 16660 15438
rect 16604 15334 16660 15372
rect 14252 15204 14308 15214
rect 14252 15110 14308 15148
rect 15372 15204 15428 15214
rect 15372 14530 15428 15148
rect 15372 14478 15374 14530
rect 15426 14478 15428 14530
rect 12572 14420 12628 14430
rect 12348 14418 12628 14420
rect 12348 14366 12574 14418
rect 12626 14366 12628 14418
rect 12348 14364 12628 14366
rect 12572 14354 12628 14364
rect 15372 12964 15428 14478
rect 16828 14530 16884 16044
rect 17500 16100 17556 16110
rect 17500 16006 17556 16044
rect 17724 15314 17780 16156
rect 18620 16100 18676 16110
rect 18620 16006 18676 16044
rect 19180 15986 19236 16606
rect 20188 16658 20244 19200
rect 20188 16606 20190 16658
rect 20242 16606 20244 16658
rect 20188 16210 20244 16606
rect 20188 16158 20190 16210
rect 20242 16158 20244 16210
rect 20188 16146 20244 16158
rect 21420 16658 21476 16670
rect 21420 16606 21422 16658
rect 21474 16606 21476 16658
rect 19180 15934 19182 15986
rect 19234 15934 19236 15986
rect 19180 15922 19236 15934
rect 19404 16100 19460 16110
rect 18060 15874 18116 15886
rect 18060 15822 18062 15874
rect 18114 15822 18116 15874
rect 18060 15540 18116 15822
rect 18060 15474 18116 15484
rect 19404 15876 19460 16044
rect 21420 16098 21476 16606
rect 21420 16046 21422 16098
rect 21474 16046 21476 16098
rect 21420 16034 21476 16046
rect 21756 16100 21812 19200
rect 23324 17444 23380 19200
rect 23212 17388 23380 17444
rect 21756 16034 21812 16044
rect 22316 16100 22372 16110
rect 22316 15986 22372 16044
rect 22316 15934 22318 15986
rect 22370 15934 22372 15986
rect 22316 15922 22372 15934
rect 23212 15988 23268 17388
rect 23374 16492 23638 16502
rect 23430 16436 23478 16492
rect 23534 16436 23582 16492
rect 23374 16426 23638 16436
rect 24668 16212 24724 16222
rect 24892 16212 24948 19200
rect 25676 16212 25732 16222
rect 24668 16210 25396 16212
rect 24668 16158 24670 16210
rect 24722 16158 25396 16210
rect 24668 16156 25396 16158
rect 24668 16146 24724 16156
rect 25340 16098 25396 16156
rect 25340 16046 25342 16098
rect 25394 16046 25396 16098
rect 25340 16034 25396 16046
rect 23548 15988 23604 15998
rect 23212 15986 23604 15988
rect 23212 15934 23550 15986
rect 23602 15934 23604 15986
rect 23212 15932 23604 15934
rect 23548 15922 23604 15932
rect 25676 15986 25732 16156
rect 25676 15934 25678 15986
rect 25730 15934 25732 15986
rect 25676 15922 25732 15934
rect 26460 15988 26516 19200
rect 27692 16100 27748 16110
rect 26684 15988 26740 15998
rect 26460 15986 26740 15988
rect 26460 15934 26686 15986
rect 26738 15934 26740 15986
rect 26460 15932 26740 15934
rect 26684 15922 26740 15932
rect 19740 15876 19796 15886
rect 19404 15874 19796 15876
rect 19404 15822 19742 15874
rect 19794 15822 19796 15874
rect 19404 15820 19796 15822
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 16828 14478 16830 14530
rect 16882 14478 16884 14530
rect 15932 14420 15988 14430
rect 15932 14326 15988 14364
rect 16604 13972 16660 13982
rect 16828 13972 16884 14478
rect 17500 14532 17556 14542
rect 17724 14532 17780 15262
rect 19404 15314 19460 15820
rect 19740 15810 19796 15820
rect 20748 15874 20804 15886
rect 21756 15876 21812 15886
rect 20748 15822 20750 15874
rect 20802 15822 20804 15874
rect 20300 15428 20356 15438
rect 20748 15428 20804 15822
rect 21644 15874 21812 15876
rect 21644 15822 21758 15874
rect 21810 15822 21812 15874
rect 21644 15820 21812 15822
rect 20860 15428 20916 15438
rect 20300 15426 20916 15428
rect 20300 15374 20302 15426
rect 20354 15374 20862 15426
rect 20914 15374 20916 15426
rect 20300 15372 20916 15374
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 18508 15204 18564 15214
rect 18508 15110 18564 15148
rect 19404 14644 19460 15262
rect 19740 15316 19796 15326
rect 19740 15202 19796 15260
rect 20300 15316 20356 15372
rect 20300 15250 20356 15260
rect 19740 15150 19742 15202
rect 19794 15150 19796 15202
rect 19516 14644 19572 14654
rect 17500 14530 17780 14532
rect 17500 14478 17502 14530
rect 17554 14478 17780 14530
rect 17500 14476 17780 14478
rect 18956 14642 19572 14644
rect 18956 14590 19518 14642
rect 19570 14590 19572 14642
rect 18956 14588 19572 14590
rect 18956 14530 19012 14588
rect 18956 14478 18958 14530
rect 19010 14478 19012 14530
rect 17500 14466 17556 14476
rect 18956 14466 19012 14478
rect 18060 14420 18116 14430
rect 16940 13972 16996 13982
rect 16604 13970 16996 13972
rect 16604 13918 16606 13970
rect 16658 13918 16942 13970
rect 16994 13918 16996 13970
rect 16604 13916 16996 13918
rect 16604 13906 16660 13916
rect 16940 13524 16996 13916
rect 18060 13860 18116 14364
rect 19516 14308 19572 14588
rect 19516 14242 19572 14252
rect 18060 13794 18116 13804
rect 18956 13860 19012 13870
rect 16940 13458 16996 13468
rect 17724 13636 17780 13646
rect 18172 13636 18228 13646
rect 18620 13636 18676 13646
rect 17724 13634 18676 13636
rect 17724 13582 17726 13634
rect 17778 13582 18174 13634
rect 18226 13582 18622 13634
rect 18674 13582 18676 13634
rect 17724 13580 18676 13582
rect 16380 12964 16436 12974
rect 15372 12962 16436 12964
rect 15372 12910 16382 12962
rect 16434 12910 16436 12962
rect 15372 12908 16436 12910
rect 16380 12898 16436 12908
rect 17164 12850 17220 12862
rect 17164 12798 17166 12850
rect 17218 12798 17220 12850
rect 16940 12292 16996 12302
rect 16940 12198 16996 12236
rect 17164 12292 17220 12798
rect 17724 12402 17780 13580
rect 18172 13570 18228 13580
rect 17836 13412 17892 13422
rect 17836 12962 17892 13356
rect 18620 13076 18676 13580
rect 18956 13188 19012 13804
rect 19292 13748 19348 13758
rect 19292 13654 19348 13692
rect 19740 13748 19796 15150
rect 20524 14642 20580 15372
rect 20860 15362 20916 15372
rect 20524 14590 20526 14642
rect 20578 14590 20580 14642
rect 20524 14578 20580 14590
rect 21196 15204 21252 15214
rect 20860 14420 20916 14430
rect 21196 14420 21252 15148
rect 20860 14418 21252 14420
rect 20860 14366 20862 14418
rect 20914 14366 21252 14418
rect 20860 14364 21252 14366
rect 20860 14354 20916 14364
rect 19740 13682 19796 13692
rect 19964 14306 20020 14318
rect 19964 14254 19966 14306
rect 20018 14254 20020 14306
rect 19516 13636 19572 13646
rect 19516 13542 19572 13580
rect 19964 13636 20020 14254
rect 20300 13748 20356 13758
rect 20076 13636 20132 13646
rect 19964 13634 20132 13636
rect 19964 13582 20078 13634
rect 20130 13582 20132 13634
rect 19964 13580 20132 13582
rect 18732 13076 18788 13086
rect 18620 13020 18732 13076
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 18732 12944 18788 13020
rect 18956 13074 19012 13132
rect 18956 13022 18958 13074
rect 19010 13022 19012 13074
rect 18956 13010 19012 13022
rect 19292 13524 19348 13534
rect 17836 12898 17892 12910
rect 17724 12350 17726 12402
rect 17778 12350 17780 12402
rect 17724 12338 17780 12350
rect 19292 12402 19348 13468
rect 19292 12350 19294 12402
rect 19346 12350 19348 12402
rect 18508 12292 18564 12302
rect 17164 12226 17220 12236
rect 18284 12236 18508 12292
rect 16156 12180 16212 12190
rect 16604 12180 16660 12190
rect 16156 12178 16604 12180
rect 16156 12126 16158 12178
rect 16210 12126 16604 12178
rect 16156 12124 16604 12126
rect 16156 12114 16212 12124
rect 16604 12048 16660 12124
rect 17276 12180 17332 12190
rect 17276 11508 17332 12124
rect 18172 12180 18228 12190
rect 18172 12086 18228 12124
rect 17276 11376 17332 11452
rect 17836 11508 17892 11518
rect 17836 11414 17892 11452
rect 18060 11508 18116 11518
rect 18060 10834 18116 11452
rect 18172 11508 18228 11518
rect 18284 11508 18340 12236
rect 18508 12198 18564 12236
rect 18956 12292 19012 12302
rect 18172 11506 18340 11508
rect 18172 11454 18174 11506
rect 18226 11454 18340 11506
rect 18172 11452 18340 11454
rect 18508 11508 18564 11518
rect 18172 11442 18228 11452
rect 18060 10782 18062 10834
rect 18114 10782 18116 10834
rect 18060 10770 18116 10782
rect 18508 10834 18564 11452
rect 18732 11508 18788 11518
rect 18732 11414 18788 11452
rect 18956 11508 19012 12236
rect 19292 12292 19348 12350
rect 19292 12226 19348 12236
rect 19404 13412 19460 13422
rect 19404 12290 19460 13356
rect 19852 13188 19908 13198
rect 19628 13076 19684 13086
rect 19628 12982 19684 13020
rect 19852 13074 19908 13132
rect 19852 13022 19854 13074
rect 19906 13022 19908 13074
rect 19852 12740 19908 13022
rect 19852 12674 19908 12684
rect 19964 13076 20020 13580
rect 20076 13570 20132 13580
rect 19964 12852 20020 13020
rect 20188 12852 20244 12862
rect 19964 12796 20188 12852
rect 19404 12238 19406 12290
rect 19458 12238 19460 12290
rect 19404 12226 19460 12238
rect 19852 12292 19908 12302
rect 19628 11508 19684 11518
rect 18956 11506 19236 11508
rect 18956 11454 18958 11506
rect 19010 11454 19236 11506
rect 18956 11452 19236 11454
rect 18956 11442 19012 11452
rect 18508 10782 18510 10834
rect 18562 10782 18564 10834
rect 18508 10770 18564 10782
rect 19180 10834 19236 11452
rect 19628 11414 19684 11452
rect 19852 11506 19908 12236
rect 19964 12290 20020 12796
rect 20188 12786 20244 12796
rect 20300 12516 20356 13692
rect 20412 13636 20468 13646
rect 20412 13634 20580 13636
rect 20412 13582 20414 13634
rect 20466 13582 20580 13634
rect 20412 13580 20580 13582
rect 20412 13570 20468 13580
rect 19964 12238 19966 12290
rect 20018 12238 20020 12290
rect 19964 12226 20020 12238
rect 20188 12460 20356 12516
rect 20412 13412 20468 13422
rect 19852 11454 19854 11506
rect 19906 11454 19908 11506
rect 19180 10782 19182 10834
rect 19234 10782 19236 10834
rect 19180 10770 19236 10782
rect 19852 11172 19908 11454
rect 19852 10724 19908 11116
rect 20188 11284 20244 12460
rect 20300 12292 20356 12302
rect 20300 12198 20356 12236
rect 20412 11284 20468 13356
rect 20524 13076 20580 13580
rect 20972 13634 21028 13646
rect 20972 13582 20974 13634
rect 21026 13582 21028 13634
rect 20972 13524 21028 13582
rect 20972 13458 21028 13468
rect 21196 13636 21252 14364
rect 21196 13188 21252 13580
rect 21196 13122 21252 13132
rect 21308 14644 21364 14654
rect 21308 13858 21364 14588
rect 21644 14532 21700 15820
rect 21756 15810 21812 15820
rect 27692 15874 27748 16044
rect 28028 15988 28084 19200
rect 29596 16658 29652 19200
rect 29596 16606 29598 16658
rect 29650 16606 29652 16658
rect 29596 16594 29652 16606
rect 29148 16100 29204 16110
rect 29148 16006 29204 16044
rect 30380 16100 30436 16110
rect 28252 15988 28308 15998
rect 28028 15986 28308 15988
rect 28028 15934 28254 15986
rect 28306 15934 28308 15986
rect 28028 15932 28308 15934
rect 28252 15922 28308 15932
rect 30044 15988 30100 15998
rect 30044 15986 30212 15988
rect 30044 15934 30046 15986
rect 30098 15934 30212 15986
rect 30044 15932 30212 15934
rect 30044 15922 30100 15932
rect 27692 15822 27694 15874
rect 27746 15822 27748 15874
rect 26236 15764 26292 15774
rect 26236 15538 26292 15708
rect 27580 15764 27636 15774
rect 26236 15486 26238 15538
rect 26290 15486 26292 15538
rect 26236 15474 26292 15486
rect 26908 15652 26964 15662
rect 22092 15428 22148 15438
rect 22092 15334 22148 15372
rect 22988 15428 23044 15438
rect 21644 14466 21700 14476
rect 21756 15202 21812 15214
rect 21756 15150 21758 15202
rect 21810 15150 21812 15202
rect 21756 14420 21812 15150
rect 21756 14354 21812 14364
rect 22652 15202 22708 15214
rect 22652 15150 22654 15202
rect 22706 15150 22708 15202
rect 21868 14308 21924 14318
rect 21868 14214 21924 14252
rect 22652 14306 22708 15150
rect 22652 14254 22654 14306
rect 22706 14254 22708 14306
rect 21308 13806 21310 13858
rect 21362 13806 21364 13858
rect 20860 13076 20916 13114
rect 21308 13076 21364 13806
rect 20580 13020 20692 13076
rect 20524 13010 20580 13020
rect 20524 12852 20580 12862
rect 20524 12758 20580 12796
rect 20636 12740 20692 13020
rect 20916 13020 21028 13076
rect 20860 13010 20916 13020
rect 20636 12674 20692 12684
rect 20860 12852 20916 12862
rect 20860 12068 20916 12796
rect 20972 12402 21028 13020
rect 21308 13010 21364 13020
rect 21868 13746 21924 13758
rect 21868 13694 21870 13746
rect 21922 13694 21924 13746
rect 21868 13412 21924 13694
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12292 21028 12350
rect 20972 12226 21028 12236
rect 21868 12962 21924 13356
rect 21868 12910 21870 12962
rect 21922 12910 21924 12962
rect 21868 12292 21924 12910
rect 21868 12226 21924 12236
rect 22652 12292 22708 14254
rect 22988 14644 23044 15372
rect 26908 15314 26964 15596
rect 27580 15426 27636 15708
rect 27580 15374 27582 15426
rect 27634 15374 27636 15426
rect 27580 15362 27636 15374
rect 26908 15262 26910 15314
rect 26962 15262 26964 15314
rect 26908 15250 26964 15262
rect 23548 15202 23604 15214
rect 23548 15150 23550 15202
rect 23602 15150 23604 15202
rect 23548 15092 23604 15150
rect 27692 15204 27748 15822
rect 30044 15652 30100 15662
rect 27692 15138 27748 15148
rect 29708 15204 29764 15214
rect 29708 15110 29764 15148
rect 22764 13748 22820 13758
rect 22764 13074 22820 13692
rect 22764 13022 22766 13074
rect 22818 13022 22820 13074
rect 22764 13010 22820 13022
rect 22988 13076 23044 14588
rect 23212 15036 23604 15092
rect 25564 15092 25620 15102
rect 23212 14420 23268 15036
rect 23374 14924 23638 14934
rect 23430 14868 23478 14924
rect 23534 14868 23582 14924
rect 23374 14858 23638 14868
rect 23436 14644 23492 14654
rect 23436 14550 23492 14588
rect 23212 14326 23268 14364
rect 23996 14420 24052 14430
rect 23996 14306 24052 14364
rect 23996 14254 23998 14306
rect 24050 14254 24052 14306
rect 23772 13634 23828 13646
rect 23772 13582 23774 13634
rect 23826 13582 23828 13634
rect 23772 13524 23828 13582
rect 23374 13356 23638 13366
rect 23430 13300 23478 13356
rect 23534 13300 23582 13356
rect 23374 13290 23638 13300
rect 22652 12198 22708 12236
rect 22988 12290 23044 13020
rect 23660 13076 23716 13086
rect 23660 12402 23716 13020
rect 23660 12350 23662 12402
rect 23714 12350 23716 12402
rect 23660 12338 23716 12350
rect 22988 12238 22990 12290
rect 23042 12238 23044 12290
rect 22092 12180 22148 12190
rect 20860 11974 20916 12012
rect 21756 12068 21812 12078
rect 20524 11284 20580 11294
rect 20412 11282 20580 11284
rect 20412 11230 20526 11282
rect 20578 11230 20580 11282
rect 20412 11228 20580 11230
rect 19964 10724 20020 10734
rect 19852 10722 20020 10724
rect 19852 10670 19966 10722
rect 20018 10670 20020 10722
rect 19852 10668 20020 10670
rect 19964 10658 20020 10668
rect 19068 10498 19124 10510
rect 19068 10446 19070 10498
rect 19122 10446 19124 10498
rect 19068 9940 19124 10446
rect 20188 10500 20244 11228
rect 20300 10724 20356 10734
rect 20524 10724 20580 11228
rect 21756 11282 21812 12012
rect 21756 11230 21758 11282
rect 21810 11230 21812 11282
rect 20636 11172 20692 11182
rect 20636 11078 20692 11116
rect 20972 11172 21028 11182
rect 20300 10722 20580 10724
rect 20300 10670 20302 10722
rect 20354 10670 20580 10722
rect 20300 10668 20580 10670
rect 20972 10834 21028 11116
rect 20972 10782 20974 10834
rect 21026 10782 21028 10834
rect 20300 10658 20356 10668
rect 19516 9940 19572 9950
rect 19068 9938 19572 9940
rect 19068 9886 19070 9938
rect 19122 9886 19518 9938
rect 19570 9886 19572 9938
rect 19068 9884 19572 9886
rect 19068 9874 19124 9884
rect 19516 9828 19572 9884
rect 19964 9940 20020 9950
rect 19964 9846 20020 9884
rect 19516 9762 19572 9772
rect 20188 9828 20244 10444
rect 20860 10500 20916 10510
rect 20860 10406 20916 10444
rect 20860 9940 20916 9950
rect 20972 9940 21028 10782
rect 21756 10612 21812 11230
rect 22092 11506 22148 12124
rect 22092 11454 22094 11506
rect 22146 11454 22148 11506
rect 22092 10722 22148 11454
rect 22988 11506 23044 12238
rect 23660 12180 23716 12190
rect 23772 12180 23828 13468
rect 23996 13524 24052 14254
rect 25564 14308 25620 15036
rect 30044 14642 30100 15596
rect 30156 15428 30212 15932
rect 30156 15362 30212 15372
rect 30044 14590 30046 14642
rect 30098 14590 30100 14642
rect 30044 14578 30100 14590
rect 30380 15316 30436 16044
rect 30604 16098 30660 16110
rect 30604 16046 30606 16098
rect 30658 16046 30660 16098
rect 30380 14642 30436 15260
rect 30492 15316 30548 15326
rect 30604 15316 30660 16046
rect 31164 15540 31220 19200
rect 31388 16658 31444 16670
rect 31388 16606 31390 16658
rect 31442 16606 31444 16658
rect 31388 16100 31444 16606
rect 31164 15474 31220 15484
rect 31276 16098 31444 16100
rect 31276 16046 31390 16098
rect 31442 16046 31444 16098
rect 31276 16044 31444 16046
rect 30492 15314 30660 15316
rect 30492 15262 30494 15314
rect 30546 15262 30660 15314
rect 30492 15260 30660 15262
rect 30492 15204 30548 15260
rect 30492 15138 30548 15148
rect 31052 15204 31108 15214
rect 30380 14590 30382 14642
rect 30434 14590 30436 14642
rect 30380 14578 30436 14590
rect 24892 13636 24948 13646
rect 23996 13458 24052 13468
rect 24780 13634 24948 13636
rect 24780 13582 24894 13634
rect 24946 13582 24948 13634
rect 24780 13580 24948 13582
rect 24780 13524 24836 13580
rect 24892 13570 24948 13580
rect 24556 13188 24612 13198
rect 24556 12402 24612 13132
rect 24780 13074 24836 13468
rect 24780 13022 24782 13074
rect 24834 13022 24836 13074
rect 24780 13010 24836 13022
rect 25004 13076 25060 13086
rect 24556 12350 24558 12402
rect 24610 12350 24612 12402
rect 24556 12338 24612 12350
rect 23660 12178 23828 12180
rect 23660 12126 23662 12178
rect 23714 12126 23828 12178
rect 23660 12124 23828 12126
rect 23660 12114 23716 12124
rect 23374 11788 23638 11798
rect 23430 11732 23478 11788
rect 23534 11732 23582 11788
rect 23374 11722 23638 11732
rect 23772 11620 23828 12124
rect 24444 12066 24500 12078
rect 24444 12014 24446 12066
rect 24498 12014 24500 12066
rect 22988 11454 22990 11506
rect 23042 11454 23044 11506
rect 22092 10670 22094 10722
rect 22146 10670 22148 10722
rect 22092 10658 22148 10670
rect 22652 11282 22708 11294
rect 22652 11230 22654 11282
rect 22706 11230 22708 11282
rect 21868 10612 21924 10622
rect 21756 10556 21868 10612
rect 20860 9938 21028 9940
rect 20860 9886 20862 9938
rect 20914 9886 21028 9938
rect 20860 9884 21028 9886
rect 20860 9874 20916 9884
rect 20188 9762 20244 9772
rect 20524 9828 20580 9838
rect 20412 9268 20468 9278
rect 20524 9268 20580 9772
rect 20412 9266 20580 9268
rect 20412 9214 20414 9266
rect 20466 9214 20580 9266
rect 20412 9212 20580 9214
rect 20412 9202 20468 9212
rect 20524 9156 20580 9212
rect 20524 9090 20580 9100
rect 20972 9604 21028 9884
rect 21868 9940 21924 10556
rect 22652 10612 22708 11230
rect 22988 10722 23044 11454
rect 23548 11564 23828 11620
rect 23884 11620 23940 11630
rect 23548 11284 23604 11564
rect 23884 11506 23940 11564
rect 23884 11454 23886 11506
rect 23938 11454 23940 11506
rect 23884 11442 23940 11454
rect 22988 10670 22990 10722
rect 23042 10670 23044 10722
rect 22988 10658 23044 10670
rect 23436 11282 23604 11284
rect 23436 11230 23550 11282
rect 23602 11230 23604 11282
rect 23436 11228 23604 11230
rect 22652 10518 22708 10556
rect 23436 10612 23492 11228
rect 23548 11218 23604 11228
rect 24332 11172 24388 11182
rect 23436 10518 23492 10556
rect 24108 11170 24388 11172
rect 24108 11118 24334 11170
rect 24386 11118 24388 11170
rect 24108 11116 24388 11118
rect 24108 10612 24164 11116
rect 24332 11106 24388 11116
rect 24444 11172 24500 12014
rect 25004 11620 25060 13020
rect 25564 13074 25620 14252
rect 26348 13188 26404 13198
rect 26348 13094 26404 13132
rect 31052 13188 31108 15148
rect 31164 14644 31220 14654
rect 31276 14644 31332 16044
rect 31388 16034 31444 16044
rect 31724 16436 31780 16446
rect 31724 15986 31780 16380
rect 31724 15934 31726 15986
rect 31778 15934 31780 15986
rect 31724 15922 31780 15934
rect 32396 15988 32452 15998
rect 32732 15988 32788 19200
rect 32396 15986 32788 15988
rect 32396 15934 32398 15986
rect 32450 15934 32788 15986
rect 32396 15932 32788 15934
rect 33516 16098 33572 16110
rect 33516 16046 33518 16098
rect 33570 16046 33572 16098
rect 32396 15922 32452 15932
rect 33516 15876 33572 16046
rect 34188 15988 34244 15998
rect 33516 15810 33572 15820
rect 34076 15986 34244 15988
rect 34076 15934 34190 15986
rect 34242 15934 34244 15986
rect 34076 15932 34244 15934
rect 32396 15540 32452 15550
rect 32396 15446 32452 15484
rect 31724 15316 31780 15326
rect 31724 15222 31780 15260
rect 33740 15316 33796 15326
rect 31164 14642 31332 14644
rect 31164 14590 31166 14642
rect 31218 14590 31332 14642
rect 31164 14588 31332 14590
rect 33180 14644 33236 14654
rect 31164 14578 31220 14588
rect 33180 14550 33236 14588
rect 33740 14642 33796 15260
rect 33740 14590 33742 14642
rect 33794 14590 33796 14642
rect 33740 14578 33796 14590
rect 34076 14644 34132 15932
rect 34188 15922 34244 15932
rect 34076 14578 34132 14588
rect 34188 15316 34244 15326
rect 34188 14530 34244 15260
rect 34300 15092 34356 19200
rect 35868 16658 35924 19200
rect 35868 16606 35870 16658
rect 35922 16606 35924 16658
rect 35868 16594 35924 16606
rect 36428 16658 36484 16670
rect 36428 16606 36430 16658
rect 36482 16606 36484 16658
rect 36316 16210 36372 16222
rect 36316 16158 36318 16210
rect 36370 16158 36372 16210
rect 35084 15428 35140 15438
rect 35084 15334 35140 15372
rect 35868 15316 35924 15326
rect 36316 15316 36372 16158
rect 36428 15538 36484 16606
rect 37436 16658 37492 19200
rect 37436 16606 37438 16658
rect 37490 16606 37492 16658
rect 37436 16594 37492 16606
rect 37996 16658 38052 16670
rect 37996 16606 37998 16658
rect 38050 16606 38052 16658
rect 36428 15486 36430 15538
rect 36482 15486 36484 15538
rect 36428 15474 36484 15486
rect 37100 15986 37156 15998
rect 37100 15934 37102 15986
rect 37154 15934 37156 15986
rect 37100 15538 37156 15934
rect 37436 15988 37492 15998
rect 37436 15894 37492 15932
rect 37996 15986 38052 16606
rect 38780 16212 38836 16222
rect 39004 16212 39060 19200
rect 40572 17668 40628 19200
rect 40572 17612 41076 17668
rect 38780 16210 39284 16212
rect 38780 16158 38782 16210
rect 38834 16158 39284 16210
rect 38780 16156 39284 16158
rect 38780 16146 38836 16156
rect 39228 16098 39284 16156
rect 39228 16046 39230 16098
rect 39282 16046 39284 16098
rect 39228 16034 39284 16046
rect 37996 15934 37998 15986
rect 38050 15934 38052 15986
rect 37996 15922 38052 15934
rect 41020 15986 41076 17612
rect 41020 15934 41022 15986
rect 41074 15934 41076 15986
rect 41020 15922 41076 15934
rect 42140 15988 42196 19200
rect 43708 17108 43764 19200
rect 43708 17052 44212 17108
rect 44156 16658 44212 17052
rect 44156 16606 44158 16658
rect 44210 16606 44212 16658
rect 44156 16210 44212 16606
rect 44156 16158 44158 16210
rect 44210 16158 44212 16210
rect 44156 16146 44212 16158
rect 44940 16658 44996 16670
rect 44940 16606 44942 16658
rect 44994 16606 44996 16658
rect 44940 16098 44996 16606
rect 44940 16046 44942 16098
rect 44994 16046 44996 16098
rect 44940 16034 44996 16046
rect 45276 16100 45332 19200
rect 45276 16034 45332 16044
rect 45836 16100 45892 16110
rect 42364 15988 42420 15998
rect 42140 15986 42420 15988
rect 42140 15934 42366 15986
rect 42418 15934 42420 15986
rect 42140 15932 42420 15934
rect 42364 15922 42420 15932
rect 45836 15986 45892 16044
rect 45836 15934 45838 15986
rect 45890 15934 45892 15986
rect 45836 15922 45892 15934
rect 46844 15988 46900 19200
rect 48188 16212 48244 16222
rect 48188 16118 48244 16156
rect 49868 16212 49924 16222
rect 49868 16118 49924 16156
rect 48524 16100 48580 16110
rect 47068 15988 47124 15998
rect 46844 15986 47124 15988
rect 46844 15934 47070 15986
rect 47122 15934 47124 15986
rect 46844 15932 47124 15934
rect 47068 15922 47124 15932
rect 39564 15874 39620 15886
rect 39564 15822 39566 15874
rect 39618 15822 39620 15874
rect 37100 15486 37102 15538
rect 37154 15486 37156 15538
rect 35868 15314 36372 15316
rect 35868 15262 35870 15314
rect 35922 15262 36372 15314
rect 35868 15260 36372 15262
rect 34300 15026 34356 15036
rect 35084 15204 35140 15214
rect 34188 14478 34190 14530
rect 34242 14478 34244 14530
rect 35084 14644 35140 15148
rect 35084 14512 35140 14588
rect 35868 14530 35924 15260
rect 37100 15092 37156 15486
rect 37436 15764 37492 15774
rect 37436 15538 37492 15708
rect 37436 15486 37438 15538
rect 37490 15486 37492 15538
rect 37436 15474 37492 15486
rect 39564 15540 39620 15822
rect 45276 15876 45332 15886
rect 45276 15782 45332 15820
rect 48524 15876 48580 16044
rect 49196 16100 49252 16110
rect 49196 16006 49252 16044
rect 45536 15708 45800 15718
rect 45592 15652 45640 15708
rect 45696 15652 45744 15708
rect 45536 15642 45800 15652
rect 39564 15474 39620 15484
rect 48524 15538 48580 15820
rect 48524 15486 48526 15538
rect 48578 15486 48580 15538
rect 48524 15474 48580 15486
rect 49980 15540 50036 19200
rect 50204 15540 50260 15550
rect 49980 15538 50260 15540
rect 49980 15486 50206 15538
rect 50258 15486 50260 15538
rect 49980 15484 50260 15486
rect 50204 15474 50260 15484
rect 51324 15540 51380 15550
rect 51548 15540 51604 19200
rect 51324 15538 51604 15540
rect 51324 15486 51326 15538
rect 51378 15486 51604 15538
rect 51324 15484 51604 15486
rect 51996 16210 52052 16222
rect 51996 16158 51998 16210
rect 52050 16158 52052 16210
rect 51996 16100 52052 16158
rect 51324 15474 51380 15484
rect 51996 15314 52052 16044
rect 52780 16100 52836 16110
rect 54236 16100 54292 16110
rect 52780 16006 52836 16044
rect 54124 16098 54292 16100
rect 54124 16046 54238 16098
rect 54290 16046 54292 16098
rect 54124 16044 54292 16046
rect 53564 15988 53620 15998
rect 53452 15986 53620 15988
rect 53452 15934 53566 15986
rect 53618 15934 53620 15986
rect 53452 15932 53620 15934
rect 52668 15652 52724 15662
rect 51996 15262 51998 15314
rect 52050 15262 52052 15314
rect 51996 15250 52052 15262
rect 52108 15428 52164 15438
rect 37100 15026 37156 15036
rect 34188 14466 34244 14478
rect 35868 14478 35870 14530
rect 35922 14478 35924 14530
rect 35868 14466 35924 14478
rect 39228 14644 39284 14654
rect 31052 13122 31108 13132
rect 25564 13022 25566 13074
rect 25618 13022 25620 13074
rect 25564 12292 25620 13022
rect 26460 12852 26516 12862
rect 26460 12850 26852 12852
rect 26460 12798 26462 12850
rect 26514 12798 26852 12850
rect 26460 12796 26852 12798
rect 26460 12786 26516 12796
rect 26236 12404 26292 12414
rect 26236 12310 26292 12348
rect 25676 12292 25732 12302
rect 25564 12290 25732 12292
rect 25564 12238 25678 12290
rect 25730 12238 25732 12290
rect 25564 12236 25732 12238
rect 25676 12226 25732 12236
rect 25900 11954 25956 11966
rect 25900 11902 25902 11954
rect 25954 11902 25956 11954
rect 25004 11554 25060 11564
rect 25788 11620 25844 11630
rect 25900 11620 25956 11902
rect 25788 11618 25956 11620
rect 25788 11566 25790 11618
rect 25842 11566 25956 11618
rect 25788 11564 25956 11566
rect 26460 11620 26516 11630
rect 25788 11554 25844 11564
rect 26460 11526 26516 11564
rect 25900 11396 25956 11406
rect 25900 11302 25956 11340
rect 26572 11394 26628 12796
rect 26796 12402 26852 12796
rect 26796 12350 26798 12402
rect 26850 12350 26852 12402
rect 26796 12338 26852 12350
rect 27132 12404 27188 12414
rect 27132 12310 27188 12348
rect 39228 12402 39284 14588
rect 45536 14140 45800 14150
rect 45592 14084 45640 14140
rect 45696 14084 45744 14140
rect 45536 14074 45800 14084
rect 40236 12852 40292 12862
rect 40236 12758 40292 12796
rect 40796 12852 40852 12862
rect 40796 12758 40852 12796
rect 39228 12350 39230 12402
rect 39282 12350 39284 12402
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 26572 11330 26628 11342
rect 27692 12290 27748 12302
rect 27692 12238 27694 12290
rect 27746 12238 27748 12290
rect 27692 11396 27748 12238
rect 39228 11620 39284 12350
rect 40908 12738 40964 12750
rect 40908 12686 40910 12738
rect 40962 12686 40964 12738
rect 39340 12292 39396 12302
rect 39900 12292 39956 12302
rect 39340 12290 39956 12292
rect 39340 12238 39342 12290
rect 39394 12238 39902 12290
rect 39954 12238 39956 12290
rect 39340 12236 39956 12238
rect 39340 12226 39396 12236
rect 39900 12226 39956 12236
rect 40124 12292 40180 12302
rect 39340 11620 39396 11630
rect 39228 11564 39340 11620
rect 39340 11488 39396 11564
rect 39788 11620 39844 11630
rect 27692 11330 27748 11340
rect 39452 11284 39508 11294
rect 39452 11190 39508 11228
rect 24780 11172 24836 11182
rect 24444 11170 24836 11172
rect 24444 11118 24782 11170
rect 24834 11118 24836 11170
rect 24444 11116 24836 11118
rect 24108 10518 24164 10556
rect 23374 10220 23638 10230
rect 23430 10164 23478 10220
rect 23534 10164 23582 10220
rect 23374 10154 23638 10164
rect 21868 9874 21924 9884
rect 22764 9940 22820 9950
rect 20972 9154 21028 9548
rect 21644 9714 21700 9726
rect 21644 9662 21646 9714
rect 21698 9662 21700 9714
rect 20972 9102 20974 9154
rect 21026 9102 21028 9154
rect 20972 9090 21028 9102
rect 21308 9156 21364 9166
rect 21308 9062 21364 9100
rect 21644 9156 21700 9662
rect 22540 9714 22596 9726
rect 22540 9662 22542 9714
rect 22594 9662 22596 9714
rect 21756 9604 21812 9614
rect 21756 9156 21812 9548
rect 21868 9156 21924 9166
rect 21756 9154 21924 9156
rect 21756 9102 21870 9154
rect 21922 9102 21924 9154
rect 21756 9100 21924 9102
rect 21644 9090 21700 9100
rect 21868 9090 21924 9100
rect 22204 9156 22260 9166
rect 22204 8428 22260 9100
rect 22092 8372 22260 8428
rect 22540 9156 22596 9662
rect 22652 9604 22708 9614
rect 22652 9510 22708 9548
rect 22764 9266 22820 9884
rect 23324 9940 23380 9950
rect 23324 9846 23380 9884
rect 23772 9940 23828 9950
rect 23772 9846 23828 9884
rect 22764 9214 22766 9266
rect 22818 9214 22820 9266
rect 22764 9202 22820 9214
rect 24220 9604 24276 9614
rect 24444 9604 24500 11116
rect 24780 11106 24836 11116
rect 39788 10836 39844 11564
rect 40012 11620 40068 11630
rect 40012 11526 40068 11564
rect 40124 11394 40180 12236
rect 40124 11342 40126 11394
rect 40178 11342 40180 11394
rect 40124 11330 40180 11342
rect 40572 12290 40628 12302
rect 40572 12238 40574 12290
rect 40626 12238 40628 12290
rect 39788 10704 39844 10780
rect 40460 10836 40516 10846
rect 39900 10724 39956 10734
rect 39900 10630 39956 10668
rect 24556 10612 24612 10622
rect 24556 10518 24612 10556
rect 40460 10050 40516 10780
rect 40572 10722 40628 12238
rect 40908 11620 40964 12686
rect 45536 12572 45800 12582
rect 45592 12516 45640 12572
rect 45696 12516 45744 12572
rect 45536 12506 45800 12516
rect 41580 12292 41636 12302
rect 41580 12198 41636 12236
rect 52108 11732 52164 15372
rect 40908 11554 40964 11564
rect 42140 11620 42196 11630
rect 42140 11526 42196 11564
rect 51772 11620 51828 11630
rect 52108 11620 52164 11676
rect 51772 11618 52164 11620
rect 51772 11566 51774 11618
rect 51826 11566 52164 11618
rect 51772 11564 52164 11566
rect 52668 15202 52724 15596
rect 53452 15428 53508 15932
rect 53564 15922 53620 15932
rect 53452 15362 53508 15372
rect 54012 15426 54068 15438
rect 54012 15374 54014 15426
rect 54066 15374 54068 15426
rect 53564 15316 53620 15326
rect 54012 15316 54068 15374
rect 53564 15314 54068 15316
rect 53564 15262 53566 15314
rect 53618 15262 54068 15314
rect 53564 15260 54068 15262
rect 53564 15250 53620 15260
rect 54124 15204 54180 16044
rect 54236 16034 54292 16044
rect 54684 15988 54740 19200
rect 56252 17668 56308 19200
rect 56252 17612 56756 17668
rect 54908 15988 54964 15998
rect 54684 15986 54964 15988
rect 54684 15934 54910 15986
rect 54962 15934 54964 15986
rect 54684 15932 54964 15934
rect 54908 15922 54964 15932
rect 56700 15986 56756 17612
rect 56700 15934 56702 15986
rect 56754 15934 56756 15986
rect 56700 15922 56756 15934
rect 59388 15988 59444 19200
rect 60620 16436 60676 16446
rect 60060 16212 60116 16222
rect 59612 15988 59668 15998
rect 59388 15986 59668 15988
rect 59388 15934 59614 15986
rect 59666 15934 59668 15986
rect 59388 15932 59668 15934
rect 59612 15922 59668 15932
rect 60060 15538 60116 16156
rect 60060 15486 60062 15538
rect 60114 15486 60116 15538
rect 60060 15474 60116 15486
rect 60620 15538 60676 16380
rect 60844 16212 60900 16222
rect 60844 16098 60900 16156
rect 60844 16046 60846 16098
rect 60898 16046 60900 16098
rect 60844 16034 60900 16046
rect 60620 15486 60622 15538
rect 60674 15486 60676 15538
rect 60620 15474 60676 15486
rect 60956 15540 61012 19200
rect 61628 16436 61684 16446
rect 61628 16210 61684 16380
rect 63756 16212 63812 16222
rect 61628 16158 61630 16210
rect 61682 16158 61684 16210
rect 61628 16146 61684 16158
rect 63196 16210 63812 16212
rect 63196 16158 63758 16210
rect 63810 16158 63812 16210
rect 63196 16156 63812 16158
rect 61180 15540 61236 15550
rect 60956 15538 61236 15540
rect 60956 15486 61182 15538
rect 61234 15486 61236 15538
rect 60956 15484 61236 15486
rect 61180 15474 61236 15484
rect 52668 15150 52670 15202
rect 52722 15150 52724 15202
rect 51772 11554 51828 11564
rect 52444 11506 52500 11518
rect 52444 11454 52446 11506
rect 52498 11454 52500 11506
rect 51884 11396 51940 11406
rect 51884 11302 51940 11340
rect 40684 11284 40740 11294
rect 40684 11190 40740 11228
rect 41468 11284 41524 11294
rect 41468 11190 41524 11228
rect 42028 11284 42084 11294
rect 42028 11190 42084 11228
rect 52332 11284 52388 11294
rect 42700 11170 42756 11182
rect 42700 11118 42702 11170
rect 42754 11118 42756 11170
rect 40572 10670 40574 10722
rect 40626 10670 40628 10722
rect 40572 10658 40628 10670
rect 41580 10724 41636 10734
rect 41580 10630 41636 10668
rect 40460 9998 40462 10050
rect 40514 9998 40516 10050
rect 40460 9986 40516 9998
rect 40572 10388 40628 10398
rect 40572 9826 40628 10332
rect 42700 10388 42756 11118
rect 45536 11004 45800 11014
rect 45592 10948 45640 11004
rect 45696 10948 45744 11004
rect 45536 10938 45800 10948
rect 52332 10834 52388 11228
rect 52332 10782 52334 10834
rect 52386 10782 52388 10834
rect 52332 10770 52388 10782
rect 52444 10722 52500 11454
rect 52668 11284 52724 15150
rect 53676 15148 54180 15204
rect 63196 15314 63252 16156
rect 63756 16146 63812 16156
rect 64092 16100 64148 19200
rect 64092 16034 64148 16044
rect 65660 15988 65716 19200
rect 68796 16660 68852 19200
rect 68796 16604 69076 16660
rect 67698 16492 67962 16502
rect 67754 16436 67802 16492
rect 67858 16436 67906 16492
rect 67698 16426 67962 16436
rect 66556 16100 66612 16110
rect 65884 15988 65940 15998
rect 65660 15986 65940 15988
rect 65660 15934 65886 15986
rect 65938 15934 65940 15986
rect 65660 15932 65940 15934
rect 65884 15922 65940 15932
rect 66556 15986 66612 16044
rect 66556 15934 66558 15986
rect 66610 15934 66612 15986
rect 66556 15922 66612 15934
rect 69020 15986 69076 16604
rect 69020 15934 69022 15986
rect 69074 15934 69076 15986
rect 69020 15922 69076 15934
rect 70364 15988 70420 19200
rect 73500 17668 73556 19200
rect 73052 17612 73556 17668
rect 70588 15988 70644 15998
rect 70364 15986 70644 15988
rect 70364 15934 70590 15986
rect 70642 15934 70644 15986
rect 70364 15932 70644 15934
rect 70588 15922 70644 15932
rect 73052 15986 73108 17612
rect 73052 15934 73054 15986
rect 73106 15934 73108 15986
rect 73052 15922 73108 15934
rect 75068 15988 75124 19200
rect 76524 16212 76580 16222
rect 75292 15988 75348 15998
rect 75068 15986 75348 15988
rect 75068 15934 75294 15986
rect 75346 15934 75348 15986
rect 75068 15932 75348 15934
rect 75292 15922 75348 15932
rect 64652 15876 64708 15886
rect 64540 15874 64708 15876
rect 64540 15822 64654 15874
rect 64706 15822 64708 15874
rect 64540 15820 64708 15822
rect 63196 15262 63198 15314
rect 63250 15262 63252 15314
rect 53676 14418 53732 15148
rect 63196 14530 63252 15262
rect 63756 15652 63812 15662
rect 63756 15426 63812 15596
rect 63756 15374 63758 15426
rect 63810 15374 63812 15426
rect 63756 15204 63812 15374
rect 63756 15138 63812 15148
rect 63196 14478 63198 14530
rect 63250 14478 63252 14530
rect 63196 14466 63252 14478
rect 64540 14530 64596 15820
rect 64652 15810 64708 15820
rect 73724 15876 73780 15886
rect 73724 15874 74004 15876
rect 73724 15822 73726 15874
rect 73778 15822 74004 15874
rect 73724 15820 74004 15822
rect 73724 15810 73780 15820
rect 65436 15426 65492 15438
rect 65436 15374 65438 15426
rect 65490 15374 65492 15426
rect 64652 15316 64708 15326
rect 65436 15316 65492 15374
rect 64652 15314 65492 15316
rect 64652 15262 64654 15314
rect 64706 15262 65492 15314
rect 64652 15260 65492 15262
rect 72716 15316 72772 15326
rect 64652 15250 64708 15260
rect 67698 14924 67962 14934
rect 67754 14868 67802 14924
rect 67858 14868 67906 14924
rect 67698 14858 67962 14868
rect 64540 14478 64542 14530
rect 64594 14478 64596 14530
rect 64540 14466 64596 14478
rect 72716 14530 72772 15260
rect 73612 15316 73668 15326
rect 73612 15222 73668 15260
rect 72716 14478 72718 14530
rect 72770 14478 72772 14530
rect 72716 14466 72772 14478
rect 73948 14530 74004 15820
rect 74396 15874 74452 15886
rect 74396 15822 74398 15874
rect 74450 15822 74452 15874
rect 74396 15316 74452 15822
rect 76524 15538 76580 16156
rect 76524 15486 76526 15538
rect 76578 15486 76580 15538
rect 74844 15316 74900 15326
rect 74396 15314 74900 15316
rect 74396 15262 74846 15314
rect 74898 15262 74900 15314
rect 74396 15260 74900 15262
rect 74844 15250 74900 15260
rect 74172 15204 74228 15214
rect 74172 14644 74228 15148
rect 76524 15204 76580 15486
rect 76972 15988 77028 15998
rect 78204 15988 78260 19200
rect 79772 17668 79828 19200
rect 79772 17612 80276 17668
rect 78428 15988 78484 15998
rect 78204 15986 78484 15988
rect 78204 15934 78430 15986
rect 78482 15934 78484 15986
rect 78204 15932 78484 15934
rect 76972 15538 77028 15932
rect 78428 15922 78484 15932
rect 80220 15986 80276 17612
rect 80220 15934 80222 15986
rect 80274 15934 80276 15986
rect 80220 15922 80276 15934
rect 82908 15988 82964 19200
rect 83132 15988 83188 15998
rect 82908 15986 83188 15988
rect 82908 15934 83134 15986
rect 83186 15934 83188 15986
rect 82908 15932 83188 15934
rect 84476 15988 84532 19200
rect 87612 17668 87668 19200
rect 87612 17612 88116 17668
rect 84700 15988 84756 15998
rect 84476 15986 84756 15988
rect 84476 15934 84702 15986
rect 84754 15934 84756 15986
rect 84476 15932 84756 15934
rect 83132 15922 83188 15932
rect 84700 15922 84756 15932
rect 88060 15986 88116 17612
rect 88060 15934 88062 15986
rect 88114 15934 88116 15986
rect 88060 15922 88116 15934
rect 89180 15988 89236 19200
rect 92316 16660 92372 19200
rect 92316 16604 92596 16660
rect 91196 16100 91252 16110
rect 89292 15988 89348 15998
rect 89180 15986 89348 15988
rect 89180 15934 89294 15986
rect 89346 15934 89348 15986
rect 89180 15932 89348 15934
rect 89292 15922 89348 15932
rect 90076 15876 90132 15914
rect 90076 15810 90132 15820
rect 90636 15874 90692 15886
rect 90636 15822 90638 15874
rect 90690 15822 90692 15874
rect 89860 15708 90124 15718
rect 89916 15652 89964 15708
rect 90020 15652 90068 15708
rect 89860 15642 90124 15652
rect 76972 15486 76974 15538
rect 77026 15486 77028 15538
rect 76972 15428 77028 15486
rect 76972 15362 77028 15372
rect 79660 15428 79716 15438
rect 79660 15334 79716 15372
rect 76524 15138 76580 15148
rect 77532 15316 77588 15326
rect 77532 15202 77588 15260
rect 77532 15150 77534 15202
rect 77586 15150 77588 15202
rect 77532 15138 77588 15150
rect 80444 15314 80500 15326
rect 80444 15262 80446 15314
rect 80498 15262 80500 15314
rect 80444 15204 80500 15262
rect 80444 15138 80500 15148
rect 89516 15316 89572 15326
rect 74172 14578 74228 14588
rect 88956 14644 89012 14654
rect 88956 14550 89012 14588
rect 73948 14478 73950 14530
rect 74002 14478 74004 14530
rect 73948 14466 74004 14478
rect 88396 14532 88452 14542
rect 88396 14438 88452 14476
rect 89516 14532 89572 15260
rect 90076 15204 90132 15214
rect 89516 14466 89572 14476
rect 89740 15202 90132 15204
rect 89740 15150 90078 15202
rect 90130 15150 90132 15202
rect 89740 15148 90132 15150
rect 53676 14366 53678 14418
rect 53730 14366 53732 14418
rect 53676 14354 53732 14366
rect 63308 14420 63364 14430
rect 61628 13748 61684 13758
rect 60956 13746 61684 13748
rect 60956 13694 61630 13746
rect 61682 13694 61684 13746
rect 60956 13692 61684 13694
rect 60620 12740 60676 12750
rect 60284 12292 60340 12302
rect 60284 12198 60340 12236
rect 60172 11954 60228 11966
rect 60172 11902 60174 11954
rect 60226 11902 60228 11954
rect 60172 11620 60228 11902
rect 60172 11554 60228 11564
rect 60508 11620 60564 11630
rect 60508 11526 60564 11564
rect 53452 11506 53508 11518
rect 53452 11454 53454 11506
rect 53506 11454 53508 11506
rect 53452 11396 53508 11454
rect 53452 11330 53508 11340
rect 60620 11394 60676 12684
rect 60956 12402 61012 13692
rect 61628 13682 61684 13692
rect 61740 13524 61796 13534
rect 61740 13430 61796 13468
rect 63308 13524 63364 14364
rect 63756 14420 63812 14430
rect 63756 14326 63812 14364
rect 73276 14420 73332 14430
rect 73276 14326 73332 14364
rect 89740 14420 89796 15148
rect 90076 15138 90132 15148
rect 89852 14532 89908 14542
rect 90636 14532 90692 15822
rect 90748 15876 90804 15886
rect 90748 15314 90804 15820
rect 90748 15262 90750 15314
rect 90802 15262 90804 15314
rect 90748 15250 90804 15262
rect 91196 15874 91252 16044
rect 91980 16100 92036 16110
rect 91980 16006 92036 16044
rect 91196 15822 91198 15874
rect 91250 15822 91252 15874
rect 91196 15204 91252 15822
rect 91756 15988 91812 15998
rect 91756 15540 91812 15932
rect 91756 15408 91812 15484
rect 92540 15538 92596 16604
rect 92764 15988 92820 15998
rect 92764 15894 92820 15932
rect 92540 15486 92542 15538
rect 92594 15486 92596 15538
rect 92540 15474 92596 15486
rect 93884 15540 93940 19200
rect 94892 16210 94948 16222
rect 94892 16158 94894 16210
rect 94946 16158 94948 16210
rect 94108 15540 94164 15550
rect 93884 15538 94164 15540
rect 93884 15486 94110 15538
rect 94162 15486 94164 15538
rect 93884 15484 94164 15486
rect 94108 15474 94164 15484
rect 94892 15316 94948 16158
rect 97020 15988 97076 19200
rect 97244 15988 97300 15998
rect 97020 15986 97300 15988
rect 97020 15934 97246 15986
rect 97298 15934 97300 15986
rect 97020 15932 97300 15934
rect 98588 15988 98644 19200
rect 98812 15988 98868 15998
rect 98588 15986 98868 15988
rect 98588 15934 98814 15986
rect 98866 15934 98868 15986
rect 98588 15932 98868 15934
rect 101724 15988 101780 19200
rect 103292 17668 103348 19200
rect 103292 17612 103796 17668
rect 101948 15988 102004 15998
rect 101724 15986 102004 15988
rect 101724 15934 101950 15986
rect 102002 15934 102004 15986
rect 101724 15932 102004 15934
rect 97244 15922 97300 15932
rect 98812 15922 98868 15932
rect 101948 15922 102004 15932
rect 103740 15986 103796 17612
rect 103740 15934 103742 15986
rect 103794 15934 103796 15986
rect 103740 15922 103796 15934
rect 106428 15988 106484 19200
rect 106652 15988 106708 15998
rect 106428 15986 106708 15988
rect 106428 15934 106654 15986
rect 106706 15934 106708 15986
rect 106428 15932 106708 15934
rect 107996 15988 108052 19200
rect 111132 17668 111188 19200
rect 111132 17612 111636 17668
rect 108220 15988 108276 15998
rect 107996 15986 108276 15988
rect 107996 15934 108222 15986
rect 108274 15934 108276 15986
rect 107996 15932 108276 15934
rect 106652 15922 106708 15932
rect 108220 15922 108276 15932
rect 111580 15986 111636 17612
rect 112022 16492 112286 16502
rect 112078 16436 112126 16492
rect 112182 16436 112230 16492
rect 112022 16426 112286 16436
rect 111580 15934 111582 15986
rect 111634 15934 111636 15986
rect 111580 15922 111636 15934
rect 112700 15988 112756 19200
rect 115836 16660 115892 19200
rect 115836 16604 116116 16660
rect 112924 15988 112980 15998
rect 112700 15986 112980 15988
rect 112700 15934 112926 15986
rect 112978 15934 112980 15986
rect 112700 15932 112980 15934
rect 112924 15922 112980 15932
rect 116060 15986 116116 16604
rect 116060 15934 116062 15986
rect 116114 15934 116116 15986
rect 116060 15922 116116 15934
rect 117404 15988 117460 19200
rect 117628 15988 117684 15998
rect 117404 15986 117684 15988
rect 117404 15934 117630 15986
rect 117682 15934 117684 15986
rect 117404 15932 117684 15934
rect 120540 15988 120596 19200
rect 120764 15988 120820 15998
rect 120540 15986 120820 15988
rect 120540 15934 120766 15986
rect 120818 15934 120820 15986
rect 120540 15932 120820 15934
rect 122108 15988 122164 19200
rect 122332 15988 122388 15998
rect 122108 15986 122388 15988
rect 122108 15934 122334 15986
rect 122386 15934 122388 15986
rect 122108 15932 122388 15934
rect 125244 15988 125300 19200
rect 126812 17668 126868 19200
rect 126812 17612 127316 17668
rect 125468 15988 125524 15998
rect 125244 15986 125524 15988
rect 125244 15934 125470 15986
rect 125522 15934 125524 15986
rect 125244 15932 125524 15934
rect 117628 15922 117684 15932
rect 120764 15922 120820 15932
rect 122332 15922 122388 15932
rect 125468 15922 125524 15932
rect 127260 15986 127316 17612
rect 127260 15934 127262 15986
rect 127314 15934 127316 15986
rect 127260 15922 127316 15934
rect 129948 15988 130004 19200
rect 130172 15988 130228 15998
rect 129948 15986 130228 15988
rect 129948 15934 130174 15986
rect 130226 15934 130228 15986
rect 129948 15932 130228 15934
rect 131516 15988 131572 19200
rect 134652 17668 134708 19200
rect 134652 17612 135156 17668
rect 131740 15988 131796 15998
rect 131516 15986 131796 15988
rect 131516 15934 131742 15986
rect 131794 15934 131796 15986
rect 131516 15932 131796 15934
rect 130172 15922 130228 15932
rect 131740 15922 131796 15932
rect 135100 15986 135156 17612
rect 135100 15934 135102 15986
rect 135154 15934 135156 15986
rect 135100 15922 135156 15934
rect 136220 15988 136276 19200
rect 139356 16660 139412 19200
rect 139356 16604 139636 16660
rect 136444 15988 136500 15998
rect 136220 15986 136500 15988
rect 136220 15934 136446 15986
rect 136498 15934 136500 15986
rect 136220 15932 136500 15934
rect 136444 15922 136500 15932
rect 139580 15986 139636 16604
rect 139580 15934 139582 15986
rect 139634 15934 139636 15986
rect 139580 15922 139636 15934
rect 140924 15988 140980 19200
rect 141148 15988 141204 15998
rect 140924 15986 141204 15988
rect 140924 15934 141150 15986
rect 141202 15934 141204 15986
rect 140924 15932 141204 15934
rect 144060 15988 144116 19200
rect 144284 15988 144340 15998
rect 144060 15986 144340 15988
rect 144060 15934 144286 15986
rect 144338 15934 144340 15986
rect 144060 15932 144340 15934
rect 145628 15988 145684 19200
rect 145852 15988 145908 15998
rect 145628 15986 145908 15988
rect 145628 15934 145854 15986
rect 145906 15934 145908 15986
rect 145628 15932 145908 15934
rect 148764 15988 148820 19200
rect 150332 17668 150388 19200
rect 150332 17612 150836 17668
rect 148988 15988 149044 15998
rect 148764 15986 149044 15988
rect 148764 15934 148990 15986
rect 149042 15934 149044 15986
rect 148764 15932 149044 15934
rect 141148 15922 141204 15932
rect 144284 15922 144340 15932
rect 145852 15922 145908 15932
rect 148988 15922 149044 15932
rect 150780 15986 150836 17612
rect 150780 15934 150782 15986
rect 150834 15934 150836 15986
rect 150780 15922 150836 15934
rect 153468 15988 153524 19200
rect 153692 15988 153748 15998
rect 153468 15986 153748 15988
rect 153468 15934 153694 15986
rect 153746 15934 153748 15986
rect 153468 15932 153748 15934
rect 155036 15988 155092 19200
rect 158172 17668 158228 19200
rect 158172 17612 158676 17668
rect 156346 16492 156610 16502
rect 156402 16436 156450 16492
rect 156506 16436 156554 16492
rect 156346 16426 156610 16436
rect 155260 15988 155316 15998
rect 155036 15986 155316 15988
rect 155036 15934 155262 15986
rect 155314 15934 155316 15986
rect 155036 15932 155316 15934
rect 153692 15922 153748 15932
rect 155260 15922 155316 15932
rect 158620 15986 158676 17612
rect 158620 15934 158622 15986
rect 158674 15934 158676 15986
rect 158620 15922 158676 15934
rect 159740 15988 159796 19200
rect 162876 16660 162932 19200
rect 162876 16604 163156 16660
rect 159964 15988 160020 15998
rect 159740 15986 160020 15988
rect 159740 15934 159966 15986
rect 160018 15934 160020 15986
rect 159740 15932 160020 15934
rect 159964 15922 160020 15932
rect 163100 15986 163156 16604
rect 163100 15934 163102 15986
rect 163154 15934 163156 15986
rect 163100 15922 163156 15934
rect 164444 15988 164500 19200
rect 164668 15988 164724 15998
rect 164444 15986 164724 15988
rect 164444 15934 164670 15986
rect 164722 15934 164724 15986
rect 164444 15932 164724 15934
rect 167580 15988 167636 19200
rect 167804 15988 167860 15998
rect 167580 15986 167860 15988
rect 167580 15934 167806 15986
rect 167858 15934 167860 15986
rect 167580 15932 167860 15934
rect 169148 15988 169204 19200
rect 169372 15988 169428 15998
rect 169148 15986 169428 15988
rect 169148 15934 169374 15986
rect 169426 15934 169428 15986
rect 169148 15932 169428 15934
rect 172284 15988 172340 19200
rect 173852 17668 173908 19200
rect 173852 17612 174356 17668
rect 172508 15988 172564 15998
rect 172284 15986 172564 15988
rect 172284 15934 172510 15986
rect 172562 15934 172564 15986
rect 172284 15932 172564 15934
rect 164668 15922 164724 15932
rect 167804 15922 167860 15932
rect 169372 15922 169428 15932
rect 172508 15922 172564 15932
rect 174300 15986 174356 17612
rect 174300 15934 174302 15986
rect 174354 15934 174356 15986
rect 174300 15922 174356 15934
rect 176988 15988 177044 19200
rect 178556 17444 178612 19200
rect 178108 17388 178612 17444
rect 177212 15988 177268 15998
rect 176988 15986 177268 15988
rect 176988 15934 177214 15986
rect 177266 15934 177268 15986
rect 176988 15932 177268 15934
rect 177212 15922 177268 15932
rect 134184 15708 134448 15718
rect 134240 15652 134288 15708
rect 134344 15652 134392 15708
rect 134184 15642 134448 15652
rect 178108 15538 178164 17388
rect 178508 15708 178772 15718
rect 178564 15652 178612 15708
rect 178668 15652 178716 15708
rect 178508 15642 178772 15652
rect 178108 15486 178110 15538
rect 178162 15486 178164 15538
rect 178108 15474 178164 15486
rect 94892 15250 94948 15260
rect 91196 15138 91252 15148
rect 112022 14924 112286 14934
rect 112078 14868 112126 14924
rect 112182 14868 112230 14924
rect 112022 14858 112286 14868
rect 156346 14924 156610 14934
rect 156402 14868 156450 14924
rect 156506 14868 156554 14924
rect 156346 14858 156610 14868
rect 89852 14530 90692 14532
rect 89852 14478 89854 14530
rect 89906 14478 90692 14530
rect 89852 14476 90692 14478
rect 93884 14644 93940 14654
rect 89852 14466 89908 14476
rect 63196 13188 63252 13198
rect 63308 13188 63364 13468
rect 67698 13356 67962 13366
rect 67754 13300 67802 13356
rect 67858 13300 67906 13356
rect 67698 13290 67962 13300
rect 63196 13186 63364 13188
rect 63196 13134 63198 13186
rect 63250 13134 63364 13186
rect 63196 13132 63364 13134
rect 63084 12852 63140 12862
rect 62524 12850 63140 12852
rect 62524 12798 63086 12850
rect 63138 12798 63140 12850
rect 62524 12796 63140 12798
rect 60956 12350 60958 12402
rect 61010 12350 61012 12402
rect 60956 12338 61012 12350
rect 61740 12738 61796 12750
rect 61740 12686 61742 12738
rect 61794 12686 61796 12738
rect 61516 12290 61572 12302
rect 61516 12238 61518 12290
rect 61570 12238 61572 12290
rect 61404 11620 61460 11630
rect 61404 11526 61460 11564
rect 60620 11342 60622 11394
rect 60674 11342 60676 11394
rect 60620 11330 60676 11342
rect 61516 11394 61572 12238
rect 61740 12292 61796 12686
rect 62412 12740 62468 12750
rect 62412 12646 62468 12684
rect 62300 12404 62356 12414
rect 62524 12404 62580 12796
rect 63084 12786 63140 12796
rect 63196 12516 63252 13132
rect 62300 12402 62580 12404
rect 62300 12350 62302 12402
rect 62354 12350 62580 12402
rect 62300 12348 62580 12350
rect 62972 12460 63252 12516
rect 62300 12338 62356 12348
rect 61740 12226 61796 12236
rect 61516 11342 61518 11394
rect 61570 11342 61572 11394
rect 61516 11330 61572 11342
rect 61852 11620 61908 11630
rect 52668 11218 52724 11228
rect 61852 10834 61908 11564
rect 62972 11620 63028 12460
rect 62972 11488 63028 11564
rect 63196 12290 63252 12302
rect 63868 12292 63924 12302
rect 63196 12238 63198 12290
rect 63250 12238 63252 12290
rect 63084 11396 63140 11406
rect 63196 11396 63252 12238
rect 63756 12290 63924 12292
rect 63756 12238 63870 12290
rect 63922 12238 63924 12290
rect 63756 12236 63924 12238
rect 63644 11620 63700 11630
rect 63644 11526 63700 11564
rect 63084 11394 63252 11396
rect 63084 11342 63086 11394
rect 63138 11342 63252 11394
rect 63084 11340 63252 11342
rect 63756 11394 63812 12236
rect 63868 12226 63924 12236
rect 67698 11788 67962 11798
rect 67754 11732 67802 11788
rect 67858 11732 67906 11788
rect 67698 11722 67962 11732
rect 63756 11342 63758 11394
rect 63810 11342 63812 11394
rect 63084 11330 63140 11340
rect 63756 11330 63812 11342
rect 61852 10782 61854 10834
rect 61906 10782 61908 10834
rect 61852 10770 61908 10782
rect 62076 11170 62132 11182
rect 62076 11118 62078 11170
rect 62130 11118 62132 11170
rect 52444 10670 52446 10722
rect 52498 10670 52500 10722
rect 52444 10658 52500 10670
rect 61964 10724 62020 10734
rect 62076 10724 62132 11118
rect 61964 10722 62132 10724
rect 61964 10670 61966 10722
rect 62018 10670 62132 10722
rect 61964 10668 62132 10670
rect 61964 10658 62020 10668
rect 42700 10322 42756 10332
rect 67698 10220 67962 10230
rect 67754 10164 67802 10220
rect 67858 10164 67906 10220
rect 67698 10154 67962 10164
rect 40572 9774 40574 9826
rect 40626 9774 40628 9826
rect 40572 9762 40628 9774
rect 24220 9602 24500 9604
rect 24220 9550 24222 9602
rect 24274 9550 24500 9602
rect 24220 9548 24500 9550
rect 21644 8036 21700 8046
rect 22092 8036 22148 8372
rect 22540 8370 22596 9100
rect 23100 9156 23156 9166
rect 23100 9062 23156 9100
rect 24220 9156 24276 9548
rect 45536 9436 45800 9446
rect 45592 9380 45640 9436
rect 45696 9380 45744 9436
rect 45536 9370 45800 9380
rect 24220 9090 24276 9100
rect 89740 9044 89796 14364
rect 89860 14140 90124 14150
rect 89916 14084 89964 14140
rect 90020 14084 90068 14140
rect 89860 14074 90124 14084
rect 89860 12572 90124 12582
rect 89916 12516 89964 12572
rect 90020 12516 90068 12572
rect 89860 12506 90124 12516
rect 89860 11004 90124 11014
rect 89916 10948 89964 11004
rect 90020 10948 90068 11004
rect 89860 10938 90124 10948
rect 89860 9436 90124 9446
rect 89916 9380 89964 9436
rect 90020 9380 90068 9436
rect 89860 9370 90124 9380
rect 93884 9268 93940 14588
rect 134184 14140 134448 14150
rect 134240 14084 134288 14140
rect 134344 14084 134392 14140
rect 134184 14074 134448 14084
rect 178508 14140 178772 14150
rect 178564 14084 178612 14140
rect 178668 14084 178716 14140
rect 178508 14074 178772 14084
rect 112022 13356 112286 13366
rect 112078 13300 112126 13356
rect 112182 13300 112230 13356
rect 112022 13290 112286 13300
rect 156346 13356 156610 13366
rect 156402 13300 156450 13356
rect 156506 13300 156554 13356
rect 156346 13290 156610 13300
rect 134184 12572 134448 12582
rect 134240 12516 134288 12572
rect 134344 12516 134392 12572
rect 134184 12506 134448 12516
rect 178508 12572 178772 12582
rect 178564 12516 178612 12572
rect 178668 12516 178716 12572
rect 178508 12506 178772 12516
rect 112022 11788 112286 11798
rect 112078 11732 112126 11788
rect 112182 11732 112230 11788
rect 112022 11722 112286 11732
rect 156346 11788 156610 11798
rect 156402 11732 156450 11788
rect 156506 11732 156554 11788
rect 156346 11722 156610 11732
rect 134184 11004 134448 11014
rect 134240 10948 134288 11004
rect 134344 10948 134392 11004
rect 134184 10938 134448 10948
rect 178508 11004 178772 11014
rect 178564 10948 178612 11004
rect 178668 10948 178716 11004
rect 178508 10938 178772 10948
rect 112022 10220 112286 10230
rect 112078 10164 112126 10220
rect 112182 10164 112230 10220
rect 112022 10154 112286 10164
rect 156346 10220 156610 10230
rect 156402 10164 156450 10220
rect 156506 10164 156554 10220
rect 156346 10154 156610 10164
rect 134184 9436 134448 9446
rect 134240 9380 134288 9436
rect 134344 9380 134392 9436
rect 134184 9370 134448 9380
rect 178508 9436 178772 9446
rect 178564 9380 178612 9436
rect 178668 9380 178716 9436
rect 178508 9370 178772 9380
rect 93884 9136 93940 9212
rect 94444 9268 94500 9278
rect 94444 9174 94500 9212
rect 94780 9154 94836 9166
rect 89740 8978 89796 8988
rect 94780 9102 94782 9154
rect 94834 9102 94836 9154
rect 23374 8652 23638 8662
rect 23430 8596 23478 8652
rect 23534 8596 23582 8652
rect 23374 8586 23638 8596
rect 67698 8652 67962 8662
rect 67754 8596 67802 8652
rect 67858 8596 67906 8652
rect 67698 8586 67962 8596
rect 22540 8318 22542 8370
rect 22594 8318 22596 8370
rect 22540 8306 22596 8318
rect 21644 8034 22148 8036
rect 21644 7982 21646 8034
rect 21698 7982 22094 8034
rect 22146 7982 22148 8034
rect 21644 7980 22148 7982
rect 21644 7970 21700 7980
rect 22092 7970 22148 7980
rect 45536 7868 45800 7878
rect 45592 7812 45640 7868
rect 45696 7812 45744 7868
rect 45536 7802 45800 7812
rect 89860 7868 90124 7878
rect 89916 7812 89964 7868
rect 90020 7812 90068 7868
rect 89860 7802 90124 7812
rect 23374 7084 23638 7094
rect 23430 7028 23478 7084
rect 23534 7028 23582 7084
rect 23374 7018 23638 7028
rect 67698 7084 67962 7094
rect 67754 7028 67802 7084
rect 67858 7028 67906 7084
rect 67698 7018 67962 7028
rect 45536 6300 45800 6310
rect 45592 6244 45640 6300
rect 45696 6244 45744 6300
rect 45536 6234 45800 6244
rect 89860 6300 90124 6310
rect 89916 6244 89964 6300
rect 90020 6244 90068 6300
rect 89860 6234 90124 6244
rect 23374 5516 23638 5526
rect 23430 5460 23478 5516
rect 23534 5460 23582 5516
rect 23374 5450 23638 5460
rect 67698 5516 67962 5526
rect 67754 5460 67802 5516
rect 67858 5460 67906 5516
rect 67698 5450 67962 5460
rect 45536 4732 45800 4742
rect 45592 4676 45640 4732
rect 45696 4676 45744 4732
rect 45536 4666 45800 4676
rect 89860 4732 90124 4742
rect 89916 4676 89964 4732
rect 90020 4676 90068 4732
rect 89860 4666 90124 4676
rect 94780 4340 94836 9102
rect 95900 9154 95956 9166
rect 95900 9102 95902 9154
rect 95954 9102 95956 9154
rect 95340 9044 95396 9054
rect 95340 8370 95396 8988
rect 95564 9044 95620 9054
rect 95564 8950 95620 8988
rect 95340 8318 95342 8370
rect 95394 8318 95396 8370
rect 95340 8306 95396 8318
rect 94780 4274 94836 4284
rect 95900 4228 95956 9102
rect 112022 8652 112286 8662
rect 112078 8596 112126 8652
rect 112182 8596 112230 8652
rect 112022 8586 112286 8596
rect 156346 8652 156610 8662
rect 156402 8596 156450 8652
rect 156506 8596 156554 8652
rect 156346 8586 156610 8596
rect 134184 7868 134448 7878
rect 134240 7812 134288 7868
rect 134344 7812 134392 7868
rect 134184 7802 134448 7812
rect 178508 7868 178772 7878
rect 178564 7812 178612 7868
rect 178668 7812 178716 7868
rect 178508 7802 178772 7812
rect 112022 7084 112286 7094
rect 112078 7028 112126 7084
rect 112182 7028 112230 7084
rect 112022 7018 112286 7028
rect 156346 7084 156610 7094
rect 156402 7028 156450 7084
rect 156506 7028 156554 7084
rect 156346 7018 156610 7028
rect 134184 6300 134448 6310
rect 134240 6244 134288 6300
rect 134344 6244 134392 6300
rect 134184 6234 134448 6244
rect 178508 6300 178772 6310
rect 178564 6244 178612 6300
rect 178668 6244 178716 6300
rect 178508 6234 178772 6244
rect 112022 5516 112286 5526
rect 112078 5460 112126 5516
rect 112182 5460 112230 5516
rect 112022 5450 112286 5460
rect 156346 5516 156610 5526
rect 156402 5460 156450 5516
rect 156506 5460 156554 5516
rect 156346 5450 156610 5460
rect 134184 4732 134448 4742
rect 134240 4676 134288 4732
rect 134344 4676 134392 4732
rect 134184 4666 134448 4676
rect 178508 4732 178772 4742
rect 178564 4676 178612 4732
rect 178668 4676 178716 4732
rect 178508 4666 178772 4676
rect 95900 4162 95956 4172
rect 119644 4340 119700 4350
rect 23374 3948 23638 3958
rect 23430 3892 23478 3948
rect 23534 3892 23582 3948
rect 23374 3882 23638 3892
rect 67698 3948 67962 3958
rect 67754 3892 67802 3948
rect 67858 3892 67906 3948
rect 67698 3882 67962 3892
rect 112022 3948 112286 3958
rect 112078 3892 112126 3948
rect 112182 3892 112230 3948
rect 112022 3882 112286 3892
rect 7308 3332 7364 3342
rect 10668 3332 10724 3342
rect 7084 3330 7364 3332
rect 7084 3278 7310 3330
rect 7362 3278 7364 3330
rect 7084 3276 7364 3278
rect 7084 800 7140 3276
rect 7308 3266 7364 3276
rect 10444 3330 10724 3332
rect 10444 3278 10670 3330
rect 10722 3278 10724 3330
rect 10444 3276 10724 3278
rect 10444 800 10500 3276
rect 10668 3266 10724 3276
rect 12684 3332 12740 3342
rect 12684 800 12740 3276
rect 13580 3332 13636 3342
rect 15148 3332 15204 3342
rect 17500 3332 17556 3342
rect 19628 3332 19684 3342
rect 21420 3332 21476 3342
rect 22988 3332 23044 3342
rect 13580 3238 13636 3276
rect 14924 3330 15204 3332
rect 14924 3278 15150 3330
rect 15202 3278 15204 3330
rect 14924 3276 15204 3278
rect 14924 800 14980 3276
rect 15148 3266 15204 3276
rect 17164 3330 17556 3332
rect 17164 3278 17502 3330
rect 17554 3278 17556 3330
rect 17164 3276 17556 3278
rect 17164 800 17220 3276
rect 17500 3266 17556 3276
rect 19404 3330 19684 3332
rect 19404 3278 19630 3330
rect 19682 3278 19684 3330
rect 19404 3276 19684 3278
rect 19404 800 19460 3276
rect 19628 3266 19684 3276
rect 21084 3330 21476 3332
rect 21084 3278 21422 3330
rect 21474 3278 21476 3330
rect 21084 3276 21476 3278
rect 21084 800 21140 3276
rect 21420 3266 21476 3276
rect 22764 3330 23044 3332
rect 22764 3278 22990 3330
rect 23042 3278 23044 3330
rect 22764 3276 23044 3278
rect 22764 800 22820 3276
rect 22988 3266 23044 3276
rect 24444 3332 24500 3342
rect 24444 800 24500 3276
rect 25340 3332 25396 3342
rect 26348 3332 26404 3342
rect 28028 3332 28084 3342
rect 29708 3332 29764 3342
rect 31388 3332 31444 3342
rect 33180 3332 33236 3342
rect 34748 3332 34804 3342
rect 25340 3238 25396 3276
rect 26124 3330 26404 3332
rect 26124 3278 26350 3330
rect 26402 3278 26404 3330
rect 26124 3276 26404 3278
rect 26124 800 26180 3276
rect 26348 3266 26404 3276
rect 27804 3330 28084 3332
rect 27804 3278 28030 3330
rect 28082 3278 28084 3330
rect 27804 3276 28084 3278
rect 27804 800 27860 3276
rect 28028 3266 28084 3276
rect 29484 3330 29764 3332
rect 29484 3278 29710 3330
rect 29762 3278 29764 3330
rect 29484 3276 29764 3278
rect 29484 800 29540 3276
rect 29708 3266 29764 3276
rect 31164 3330 31444 3332
rect 31164 3278 31390 3330
rect 31442 3278 31444 3330
rect 31164 3276 31444 3278
rect 31164 800 31220 3276
rect 31388 3266 31444 3276
rect 32844 3330 33236 3332
rect 32844 3278 33182 3330
rect 33234 3278 33236 3330
rect 32844 3276 33236 3278
rect 32844 800 32900 3276
rect 33180 3266 33236 3276
rect 34524 3330 34804 3332
rect 34524 3278 34750 3330
rect 34802 3278 34804 3330
rect 34524 3276 34804 3278
rect 34524 800 34580 3276
rect 34748 3266 34804 3276
rect 36204 3332 36260 3342
rect 36204 800 36260 3276
rect 37100 3332 37156 3342
rect 38108 3332 38164 3342
rect 39788 3332 39844 3342
rect 41468 3332 41524 3342
rect 43148 3332 43204 3342
rect 44940 3332 44996 3342
rect 46508 3332 46564 3342
rect 37100 3238 37156 3276
rect 37884 3330 38164 3332
rect 37884 3278 38110 3330
rect 38162 3278 38164 3330
rect 37884 3276 38164 3278
rect 37884 800 37940 3276
rect 38108 3266 38164 3276
rect 39564 3330 39844 3332
rect 39564 3278 39790 3330
rect 39842 3278 39844 3330
rect 39564 3276 39844 3278
rect 39564 800 39620 3276
rect 39788 3266 39844 3276
rect 41244 3330 41524 3332
rect 41244 3278 41470 3330
rect 41522 3278 41524 3330
rect 41244 3276 41524 3278
rect 41244 800 41300 3276
rect 41468 3266 41524 3276
rect 42924 3330 43204 3332
rect 42924 3278 43150 3330
rect 43202 3278 43204 3330
rect 42924 3276 43204 3278
rect 42924 800 42980 3276
rect 43148 3266 43204 3276
rect 44604 3330 44996 3332
rect 44604 3278 44942 3330
rect 44994 3278 44996 3330
rect 44604 3276 44996 3278
rect 44604 800 44660 3276
rect 44940 3266 44996 3276
rect 46284 3330 46564 3332
rect 46284 3278 46510 3330
rect 46562 3278 46564 3330
rect 46284 3276 46564 3278
rect 45536 3164 45800 3174
rect 45592 3108 45640 3164
rect 45696 3108 45744 3164
rect 45536 3098 45800 3108
rect 46284 800 46340 3276
rect 46508 3266 46564 3276
rect 47964 3332 48020 3342
rect 47964 800 48020 3276
rect 48860 3332 48916 3342
rect 49868 3332 49924 3342
rect 51548 3332 51604 3342
rect 53228 3332 53284 3342
rect 54908 3332 54964 3342
rect 56700 3332 56756 3342
rect 58268 3332 58324 3342
rect 48860 3238 48916 3276
rect 49644 3330 49924 3332
rect 49644 3278 49870 3330
rect 49922 3278 49924 3330
rect 49644 3276 49924 3278
rect 49644 800 49700 3276
rect 49868 3266 49924 3276
rect 51324 3330 51604 3332
rect 51324 3278 51550 3330
rect 51602 3278 51604 3330
rect 51324 3276 51604 3278
rect 51324 800 51380 3276
rect 51548 3266 51604 3276
rect 53004 3330 53284 3332
rect 53004 3278 53230 3330
rect 53282 3278 53284 3330
rect 53004 3276 53284 3278
rect 53004 800 53060 3276
rect 53228 3266 53284 3276
rect 54684 3330 54964 3332
rect 54684 3278 54910 3330
rect 54962 3278 54964 3330
rect 54684 3276 54964 3278
rect 54684 800 54740 3276
rect 54908 3266 54964 3276
rect 56364 3330 56756 3332
rect 56364 3278 56702 3330
rect 56754 3278 56756 3330
rect 56364 3276 56756 3278
rect 56364 800 56420 3276
rect 56700 3266 56756 3276
rect 58044 3330 58324 3332
rect 58044 3278 58270 3330
rect 58322 3278 58324 3330
rect 58044 3276 58324 3278
rect 58044 800 58100 3276
rect 58268 3266 58324 3276
rect 59724 3332 59780 3342
rect 59724 800 59780 3276
rect 60620 3332 60676 3342
rect 61628 3332 61684 3342
rect 63308 3332 63364 3342
rect 64988 3332 65044 3342
rect 66108 3332 66164 3342
rect 60620 3238 60676 3276
rect 61404 3330 61684 3332
rect 61404 3278 61630 3330
rect 61682 3278 61684 3330
rect 61404 3276 61684 3278
rect 61404 800 61460 3276
rect 61628 3266 61684 3276
rect 63084 3330 63364 3332
rect 63084 3278 63310 3330
rect 63362 3278 63364 3330
rect 63084 3276 63364 3278
rect 63084 800 63140 3276
rect 63308 3266 63364 3276
rect 64764 3330 65044 3332
rect 64764 3278 64990 3330
rect 65042 3278 65044 3330
rect 64764 3276 65044 3278
rect 64764 800 64820 3276
rect 64988 3266 65044 3276
rect 65884 3330 66164 3332
rect 65884 3278 66110 3330
rect 66162 3278 66164 3330
rect 65884 3276 66164 3278
rect 65884 800 65940 3276
rect 66108 3266 66164 3276
rect 68460 3330 68516 3342
rect 69468 3332 69524 3342
rect 71148 3332 71204 3342
rect 72828 3332 72884 3342
rect 74508 3332 74564 3342
rect 76300 3332 76356 3342
rect 77868 3332 77924 3342
rect 68460 3278 68462 3330
rect 68514 3278 68516 3330
rect 67564 1762 67620 1774
rect 67564 1710 67566 1762
rect 67618 1710 67620 1762
rect 67564 800 67620 1710
rect 68460 1762 68516 3278
rect 68460 1710 68462 1762
rect 68514 1710 68516 1762
rect 68460 1698 68516 1710
rect 69244 3330 69524 3332
rect 69244 3278 69470 3330
rect 69522 3278 69524 3330
rect 69244 3276 69524 3278
rect 69244 800 69300 3276
rect 69468 3266 69524 3276
rect 70924 3330 71204 3332
rect 70924 3278 71150 3330
rect 71202 3278 71204 3330
rect 70924 3276 71204 3278
rect 70924 800 70980 3276
rect 71148 3266 71204 3276
rect 72604 3330 72884 3332
rect 72604 3278 72830 3330
rect 72882 3278 72884 3330
rect 72604 3276 72884 3278
rect 72604 800 72660 3276
rect 72828 3266 72884 3276
rect 74284 3330 74564 3332
rect 74284 3278 74510 3330
rect 74562 3278 74564 3330
rect 74284 3276 74564 3278
rect 74284 800 74340 3276
rect 74508 3266 74564 3276
rect 75964 3330 76356 3332
rect 75964 3278 76302 3330
rect 76354 3278 76356 3330
rect 75964 3276 76356 3278
rect 75964 800 76020 3276
rect 76300 3266 76356 3276
rect 77644 3330 77924 3332
rect 77644 3278 77870 3330
rect 77922 3278 77924 3330
rect 77644 3276 77924 3278
rect 77644 800 77700 3276
rect 77868 3266 77924 3276
rect 80220 3330 80276 3342
rect 81228 3332 81284 3342
rect 82908 3332 82964 3342
rect 84588 3332 84644 3342
rect 86268 3332 86324 3342
rect 88060 3332 88116 3342
rect 89628 3332 89684 3342
rect 80220 3278 80222 3330
rect 80274 3278 80276 3330
rect 79324 1762 79380 1774
rect 79324 1710 79326 1762
rect 79378 1710 79380 1762
rect 79324 800 79380 1710
rect 80220 1762 80276 3278
rect 80220 1710 80222 1762
rect 80274 1710 80276 1762
rect 80220 1698 80276 1710
rect 81004 3330 81284 3332
rect 81004 3278 81230 3330
rect 81282 3278 81284 3330
rect 81004 3276 81284 3278
rect 81004 800 81060 3276
rect 81228 3266 81284 3276
rect 82684 3330 82964 3332
rect 82684 3278 82910 3330
rect 82962 3278 82964 3330
rect 82684 3276 82964 3278
rect 82684 800 82740 3276
rect 82908 3266 82964 3276
rect 84364 3330 84644 3332
rect 84364 3278 84590 3330
rect 84642 3278 84644 3330
rect 84364 3276 84644 3278
rect 84364 800 84420 3276
rect 84588 3266 84644 3276
rect 86044 3330 86324 3332
rect 86044 3278 86270 3330
rect 86322 3278 86324 3330
rect 86044 3276 86324 3278
rect 86044 800 86100 3276
rect 86268 3266 86324 3276
rect 87724 3330 88116 3332
rect 87724 3278 88062 3330
rect 88114 3278 88116 3330
rect 87724 3276 88116 3278
rect 87724 800 87780 3276
rect 88060 3266 88116 3276
rect 89404 3330 89684 3332
rect 89404 3278 89630 3330
rect 89682 3278 89684 3330
rect 89404 3276 89684 3278
rect 89404 800 89460 3276
rect 89628 3266 89684 3276
rect 91980 3330 92036 3342
rect 92988 3332 93044 3342
rect 94668 3332 94724 3342
rect 96348 3332 96404 3342
rect 98028 3332 98084 3342
rect 99820 3332 99876 3342
rect 101388 3332 101444 3342
rect 91980 3278 91982 3330
rect 92034 3278 92036 3330
rect 89860 3164 90124 3174
rect 89916 3108 89964 3164
rect 90020 3108 90068 3164
rect 89860 3098 90124 3108
rect 91084 1762 91140 1774
rect 91084 1710 91086 1762
rect 91138 1710 91140 1762
rect 91084 800 91140 1710
rect 91980 1762 92036 3278
rect 91980 1710 91982 1762
rect 92034 1710 92036 1762
rect 91980 1698 92036 1710
rect 92764 3330 93044 3332
rect 92764 3278 92990 3330
rect 93042 3278 93044 3330
rect 92764 3276 93044 3278
rect 92764 800 92820 3276
rect 92988 3266 93044 3276
rect 94444 3330 94724 3332
rect 94444 3278 94670 3330
rect 94722 3278 94724 3330
rect 94444 3276 94724 3278
rect 94444 800 94500 3276
rect 94668 3266 94724 3276
rect 96124 3330 96404 3332
rect 96124 3278 96350 3330
rect 96402 3278 96404 3330
rect 96124 3276 96404 3278
rect 96124 800 96180 3276
rect 96348 3266 96404 3276
rect 97804 3330 98084 3332
rect 97804 3278 98030 3330
rect 98082 3278 98084 3330
rect 97804 3276 98084 3278
rect 97804 800 97860 3276
rect 98028 3266 98084 3276
rect 99484 3330 99876 3332
rect 99484 3278 99822 3330
rect 99874 3278 99876 3330
rect 99484 3276 99876 3278
rect 99484 800 99540 3276
rect 99820 3266 99876 3276
rect 101164 3330 101444 3332
rect 101164 3278 101390 3330
rect 101442 3278 101444 3330
rect 101164 3276 101444 3278
rect 101164 800 101220 3276
rect 101388 3266 101444 3276
rect 103740 3330 103796 3342
rect 104748 3332 104804 3342
rect 106428 3332 106484 3342
rect 108108 3332 108164 3342
rect 109788 3332 109844 3342
rect 111580 3332 111636 3342
rect 113148 3332 113204 3342
rect 103740 3278 103742 3330
rect 103794 3278 103796 3330
rect 102844 1762 102900 1774
rect 102844 1710 102846 1762
rect 102898 1710 102900 1762
rect 102844 800 102900 1710
rect 103740 1762 103796 3278
rect 103740 1710 103742 1762
rect 103794 1710 103796 1762
rect 103740 1698 103796 1710
rect 104524 3330 104804 3332
rect 104524 3278 104750 3330
rect 104802 3278 104804 3330
rect 104524 3276 104804 3278
rect 104524 800 104580 3276
rect 104748 3266 104804 3276
rect 106204 3330 106484 3332
rect 106204 3278 106430 3330
rect 106482 3278 106484 3330
rect 106204 3276 106484 3278
rect 106204 800 106260 3276
rect 106428 3266 106484 3276
rect 107884 3330 108164 3332
rect 107884 3278 108110 3330
rect 108162 3278 108164 3330
rect 107884 3276 108164 3278
rect 107884 800 107940 3276
rect 108108 3266 108164 3276
rect 109564 3330 109844 3332
rect 109564 3278 109790 3330
rect 109842 3278 109844 3330
rect 109564 3276 109844 3278
rect 109564 800 109620 3276
rect 109788 3266 109844 3276
rect 111244 3330 111636 3332
rect 111244 3278 111582 3330
rect 111634 3278 111636 3330
rect 111244 3276 111636 3278
rect 111244 800 111300 3276
rect 111580 3266 111636 3276
rect 112924 3330 113204 3332
rect 112924 3278 113150 3330
rect 113202 3278 113204 3330
rect 112924 3276 113204 3278
rect 112924 800 112980 3276
rect 113148 3266 113204 3276
rect 115500 3330 115556 3342
rect 116508 3332 116564 3342
rect 118188 3332 118244 3342
rect 115500 3278 115502 3330
rect 115554 3278 115556 3330
rect 114604 1762 114660 1774
rect 114604 1710 114606 1762
rect 114658 1710 114660 1762
rect 114604 800 114660 1710
rect 115500 1762 115556 3278
rect 115500 1710 115502 1762
rect 115554 1710 115556 1762
rect 115500 1698 115556 1710
rect 116284 3330 116564 3332
rect 116284 3278 116510 3330
rect 116562 3278 116564 3330
rect 116284 3276 116564 3278
rect 116284 800 116340 3276
rect 116508 3266 116564 3276
rect 117964 3330 118244 3332
rect 117964 3278 118190 3330
rect 118242 3278 118244 3330
rect 117964 3276 118244 3278
rect 117964 800 118020 3276
rect 118188 3266 118244 3276
rect 119644 800 119700 4284
rect 121324 4228 121380 4238
rect 121324 800 121380 4172
rect 156346 3948 156610 3958
rect 156402 3892 156450 3948
rect 156506 3892 156554 3948
rect 156346 3882 156610 3892
rect 123340 3332 123396 3342
rect 124908 3332 124964 3342
rect 123004 3330 123396 3332
rect 123004 3278 123342 3330
rect 123394 3278 123396 3330
rect 123004 3276 123396 3278
rect 123004 800 123060 3276
rect 123340 3266 123396 3276
rect 124684 3330 124964 3332
rect 124684 3278 124910 3330
rect 124962 3278 124964 3330
rect 124684 3276 124964 3278
rect 124684 800 124740 3276
rect 124908 3266 124964 3276
rect 127260 3330 127316 3342
rect 128268 3332 128324 3342
rect 129948 3332 130004 3342
rect 131628 3332 131684 3342
rect 133308 3332 133364 3342
rect 135100 3332 135156 3342
rect 136668 3332 136724 3342
rect 127260 3278 127262 3330
rect 127314 3278 127316 3330
rect 126364 1762 126420 1774
rect 126364 1710 126366 1762
rect 126418 1710 126420 1762
rect 126364 800 126420 1710
rect 127260 1762 127316 3278
rect 127260 1710 127262 1762
rect 127314 1710 127316 1762
rect 127260 1698 127316 1710
rect 128044 3330 128324 3332
rect 128044 3278 128270 3330
rect 128322 3278 128324 3330
rect 128044 3276 128324 3278
rect 128044 800 128100 3276
rect 128268 3266 128324 3276
rect 129724 3330 130004 3332
rect 129724 3278 129950 3330
rect 130002 3278 130004 3330
rect 129724 3276 130004 3278
rect 129724 800 129780 3276
rect 129948 3266 130004 3276
rect 131404 3330 131684 3332
rect 131404 3278 131630 3330
rect 131682 3278 131684 3330
rect 131404 3276 131684 3278
rect 131404 800 131460 3276
rect 131628 3266 131684 3276
rect 133084 3330 133364 3332
rect 133084 3278 133310 3330
rect 133362 3278 133364 3330
rect 133084 3276 133364 3278
rect 133084 800 133140 3276
rect 133308 3266 133364 3276
rect 134764 3330 135156 3332
rect 134764 3278 135102 3330
rect 135154 3278 135156 3330
rect 134764 3276 135156 3278
rect 134184 3164 134448 3174
rect 134240 3108 134288 3164
rect 134344 3108 134392 3164
rect 134184 3098 134448 3108
rect 134764 800 134820 3276
rect 135100 3266 135156 3276
rect 136444 3330 136724 3332
rect 136444 3278 136670 3330
rect 136722 3278 136724 3330
rect 136444 3276 136724 3278
rect 136444 800 136500 3276
rect 136668 3266 136724 3276
rect 139020 3330 139076 3342
rect 140028 3332 140084 3342
rect 141708 3332 141764 3342
rect 143388 3332 143444 3342
rect 145068 3332 145124 3342
rect 146860 3332 146916 3342
rect 148428 3332 148484 3342
rect 139020 3278 139022 3330
rect 139074 3278 139076 3330
rect 138124 1762 138180 1774
rect 138124 1710 138126 1762
rect 138178 1710 138180 1762
rect 138124 800 138180 1710
rect 139020 1762 139076 3278
rect 139020 1710 139022 1762
rect 139074 1710 139076 1762
rect 139020 1698 139076 1710
rect 139804 3330 140084 3332
rect 139804 3278 140030 3330
rect 140082 3278 140084 3330
rect 139804 3276 140084 3278
rect 139804 800 139860 3276
rect 140028 3266 140084 3276
rect 141484 3330 141764 3332
rect 141484 3278 141710 3330
rect 141762 3278 141764 3330
rect 141484 3276 141764 3278
rect 141484 800 141540 3276
rect 141708 3266 141764 3276
rect 143164 3330 143444 3332
rect 143164 3278 143390 3330
rect 143442 3278 143444 3330
rect 143164 3276 143444 3278
rect 143164 800 143220 3276
rect 143388 3266 143444 3276
rect 144844 3330 145124 3332
rect 144844 3278 145070 3330
rect 145122 3278 145124 3330
rect 144844 3276 145124 3278
rect 144844 800 144900 3276
rect 145068 3266 145124 3276
rect 146524 3330 146916 3332
rect 146524 3278 146862 3330
rect 146914 3278 146916 3330
rect 146524 3276 146916 3278
rect 146524 800 146580 3276
rect 146860 3266 146916 3276
rect 148204 3330 148484 3332
rect 148204 3278 148430 3330
rect 148482 3278 148484 3330
rect 148204 3276 148484 3278
rect 148204 800 148260 3276
rect 148428 3266 148484 3276
rect 150780 3330 150836 3342
rect 151788 3332 151844 3342
rect 153468 3332 153524 3342
rect 155148 3332 155204 3342
rect 156828 3332 156884 3342
rect 158620 3332 158676 3342
rect 160188 3332 160244 3342
rect 150780 3278 150782 3330
rect 150834 3278 150836 3330
rect 149884 1762 149940 1774
rect 149884 1710 149886 1762
rect 149938 1710 149940 1762
rect 149884 800 149940 1710
rect 150780 1762 150836 3278
rect 150780 1710 150782 1762
rect 150834 1710 150836 1762
rect 150780 1698 150836 1710
rect 151564 3330 151844 3332
rect 151564 3278 151790 3330
rect 151842 3278 151844 3330
rect 151564 3276 151844 3278
rect 151564 800 151620 3276
rect 151788 3266 151844 3276
rect 153244 3330 153524 3332
rect 153244 3278 153470 3330
rect 153522 3278 153524 3330
rect 153244 3276 153524 3278
rect 153244 800 153300 3276
rect 153468 3266 153524 3276
rect 154924 3330 155204 3332
rect 154924 3278 155150 3330
rect 155202 3278 155204 3330
rect 154924 3276 155204 3278
rect 154924 800 154980 3276
rect 155148 3266 155204 3276
rect 156604 3330 156884 3332
rect 156604 3278 156830 3330
rect 156882 3278 156884 3330
rect 156604 3276 156884 3278
rect 156604 800 156660 3276
rect 156828 3266 156884 3276
rect 158284 3330 158676 3332
rect 158284 3278 158622 3330
rect 158674 3278 158676 3330
rect 158284 3276 158676 3278
rect 158284 800 158340 3276
rect 158620 3266 158676 3276
rect 159964 3330 160244 3332
rect 159964 3278 160190 3330
rect 160242 3278 160244 3330
rect 159964 3276 160244 3278
rect 159964 800 160020 3276
rect 160188 3266 160244 3276
rect 162540 3330 162596 3342
rect 163548 3332 163604 3342
rect 165228 3332 165284 3342
rect 166908 3332 166964 3342
rect 168588 3332 168644 3342
rect 170380 3332 170436 3342
rect 171948 3332 172004 3342
rect 173068 3332 173124 3342
rect 162540 3278 162542 3330
rect 162594 3278 162596 3330
rect 161644 1762 161700 1774
rect 161644 1710 161646 1762
rect 161698 1710 161700 1762
rect 161644 800 161700 1710
rect 162540 1762 162596 3278
rect 162540 1710 162542 1762
rect 162594 1710 162596 1762
rect 162540 1698 162596 1710
rect 163324 3330 163604 3332
rect 163324 3278 163550 3330
rect 163602 3278 163604 3330
rect 163324 3276 163604 3278
rect 163324 800 163380 3276
rect 163548 3266 163604 3276
rect 165004 3330 165284 3332
rect 165004 3278 165230 3330
rect 165282 3278 165284 3330
rect 165004 3276 165284 3278
rect 165004 800 165060 3276
rect 165228 3266 165284 3276
rect 166684 3330 166964 3332
rect 166684 3278 166910 3330
rect 166962 3278 166964 3330
rect 166684 3276 166964 3278
rect 166684 800 166740 3276
rect 166908 3266 166964 3276
rect 168364 3330 168644 3332
rect 168364 3278 168590 3330
rect 168642 3278 168644 3330
rect 168364 3276 168644 3278
rect 168364 800 168420 3276
rect 168588 3266 168644 3276
rect 170044 3330 170436 3332
rect 170044 3278 170382 3330
rect 170434 3278 170436 3330
rect 170044 3276 170436 3278
rect 170044 800 170100 3276
rect 170380 3266 170436 3276
rect 171724 3330 172004 3332
rect 171724 3278 171950 3330
rect 172002 3278 172004 3330
rect 171724 3276 172004 3278
rect 171724 800 171780 3276
rect 171948 3266 172004 3276
rect 172844 3330 173124 3332
rect 172844 3278 173070 3330
rect 173122 3278 173124 3330
rect 172844 3276 173124 3278
rect 172844 800 172900 3276
rect 173068 3266 173124 3276
rect 173964 3332 174020 3342
rect 173404 1762 173460 1774
rect 173404 1710 173406 1762
rect 173458 1710 173460 1762
rect 173404 800 173460 1710
rect 173964 800 174020 3276
rect 174300 3330 174356 3342
rect 174300 3278 174302 3330
rect 174354 3278 174356 3330
rect 174300 1762 174356 3278
rect 174972 3332 175028 3342
rect 174972 3238 175028 3276
rect 178508 3164 178772 3174
rect 178564 3108 178612 3164
rect 178668 3108 178716 3164
rect 178508 3098 178772 3108
rect 174300 1710 174302 1762
rect 174354 1710 174356 1762
rect 174300 1698 174356 1710
rect 5936 0 6048 800
rect 6496 0 6608 800
rect 7056 0 7168 800
rect 7616 0 7728 800
rect 8176 0 8288 800
rect 8736 0 8848 800
rect 9296 0 9408 800
rect 9856 0 9968 800
rect 10416 0 10528 800
rect 10976 0 11088 800
rect 11536 0 11648 800
rect 12096 0 12208 800
rect 12656 0 12768 800
rect 13216 0 13328 800
rect 13776 0 13888 800
rect 14336 0 14448 800
rect 14896 0 15008 800
rect 15456 0 15568 800
rect 16016 0 16128 800
rect 16576 0 16688 800
rect 17136 0 17248 800
rect 17696 0 17808 800
rect 18256 0 18368 800
rect 18816 0 18928 800
rect 19376 0 19488 800
rect 19936 0 20048 800
rect 20496 0 20608 800
rect 21056 0 21168 800
rect 21616 0 21728 800
rect 22176 0 22288 800
rect 22736 0 22848 800
rect 23296 0 23408 800
rect 23856 0 23968 800
rect 24416 0 24528 800
rect 24976 0 25088 800
rect 25536 0 25648 800
rect 26096 0 26208 800
rect 26656 0 26768 800
rect 27216 0 27328 800
rect 27776 0 27888 800
rect 28336 0 28448 800
rect 28896 0 29008 800
rect 29456 0 29568 800
rect 30016 0 30128 800
rect 30576 0 30688 800
rect 31136 0 31248 800
rect 31696 0 31808 800
rect 32256 0 32368 800
rect 32816 0 32928 800
rect 33376 0 33488 800
rect 33936 0 34048 800
rect 34496 0 34608 800
rect 35056 0 35168 800
rect 35616 0 35728 800
rect 36176 0 36288 800
rect 36736 0 36848 800
rect 37296 0 37408 800
rect 37856 0 37968 800
rect 38416 0 38528 800
rect 38976 0 39088 800
rect 39536 0 39648 800
rect 40096 0 40208 800
rect 40656 0 40768 800
rect 41216 0 41328 800
rect 41776 0 41888 800
rect 42336 0 42448 800
rect 42896 0 43008 800
rect 43456 0 43568 800
rect 44016 0 44128 800
rect 44576 0 44688 800
rect 45136 0 45248 800
rect 45696 0 45808 800
rect 46256 0 46368 800
rect 46816 0 46928 800
rect 47376 0 47488 800
rect 47936 0 48048 800
rect 48496 0 48608 800
rect 49056 0 49168 800
rect 49616 0 49728 800
rect 50176 0 50288 800
rect 50736 0 50848 800
rect 51296 0 51408 800
rect 51856 0 51968 800
rect 52416 0 52528 800
rect 52976 0 53088 800
rect 53536 0 53648 800
rect 54096 0 54208 800
rect 54656 0 54768 800
rect 55216 0 55328 800
rect 55776 0 55888 800
rect 56336 0 56448 800
rect 56896 0 57008 800
rect 57456 0 57568 800
rect 58016 0 58128 800
rect 58576 0 58688 800
rect 59136 0 59248 800
rect 59696 0 59808 800
rect 60256 0 60368 800
rect 60816 0 60928 800
rect 61376 0 61488 800
rect 61936 0 62048 800
rect 62496 0 62608 800
rect 63056 0 63168 800
rect 63616 0 63728 800
rect 64176 0 64288 800
rect 64736 0 64848 800
rect 65296 0 65408 800
rect 65856 0 65968 800
rect 66416 0 66528 800
rect 66976 0 67088 800
rect 67536 0 67648 800
rect 68096 0 68208 800
rect 68656 0 68768 800
rect 69216 0 69328 800
rect 69776 0 69888 800
rect 70336 0 70448 800
rect 70896 0 71008 800
rect 71456 0 71568 800
rect 72016 0 72128 800
rect 72576 0 72688 800
rect 73136 0 73248 800
rect 73696 0 73808 800
rect 74256 0 74368 800
rect 74816 0 74928 800
rect 75376 0 75488 800
rect 75936 0 76048 800
rect 76496 0 76608 800
rect 77056 0 77168 800
rect 77616 0 77728 800
rect 78176 0 78288 800
rect 78736 0 78848 800
rect 79296 0 79408 800
rect 79856 0 79968 800
rect 80416 0 80528 800
rect 80976 0 81088 800
rect 81536 0 81648 800
rect 82096 0 82208 800
rect 82656 0 82768 800
rect 83216 0 83328 800
rect 83776 0 83888 800
rect 84336 0 84448 800
rect 84896 0 85008 800
rect 85456 0 85568 800
rect 86016 0 86128 800
rect 86576 0 86688 800
rect 87136 0 87248 800
rect 87696 0 87808 800
rect 88256 0 88368 800
rect 88816 0 88928 800
rect 89376 0 89488 800
rect 89936 0 90048 800
rect 90496 0 90608 800
rect 91056 0 91168 800
rect 91616 0 91728 800
rect 92176 0 92288 800
rect 92736 0 92848 800
rect 93296 0 93408 800
rect 93856 0 93968 800
rect 94416 0 94528 800
rect 94976 0 95088 800
rect 95536 0 95648 800
rect 96096 0 96208 800
rect 96656 0 96768 800
rect 97216 0 97328 800
rect 97776 0 97888 800
rect 98336 0 98448 800
rect 98896 0 99008 800
rect 99456 0 99568 800
rect 100016 0 100128 800
rect 100576 0 100688 800
rect 101136 0 101248 800
rect 101696 0 101808 800
rect 102256 0 102368 800
rect 102816 0 102928 800
rect 103376 0 103488 800
rect 103936 0 104048 800
rect 104496 0 104608 800
rect 105056 0 105168 800
rect 105616 0 105728 800
rect 106176 0 106288 800
rect 106736 0 106848 800
rect 107296 0 107408 800
rect 107856 0 107968 800
rect 108416 0 108528 800
rect 108976 0 109088 800
rect 109536 0 109648 800
rect 110096 0 110208 800
rect 110656 0 110768 800
rect 111216 0 111328 800
rect 111776 0 111888 800
rect 112336 0 112448 800
rect 112896 0 113008 800
rect 113456 0 113568 800
rect 114016 0 114128 800
rect 114576 0 114688 800
rect 115136 0 115248 800
rect 115696 0 115808 800
rect 116256 0 116368 800
rect 116816 0 116928 800
rect 117376 0 117488 800
rect 117936 0 118048 800
rect 118496 0 118608 800
rect 119056 0 119168 800
rect 119616 0 119728 800
rect 120176 0 120288 800
rect 120736 0 120848 800
rect 121296 0 121408 800
rect 121856 0 121968 800
rect 122416 0 122528 800
rect 122976 0 123088 800
rect 123536 0 123648 800
rect 124096 0 124208 800
rect 124656 0 124768 800
rect 125216 0 125328 800
rect 125776 0 125888 800
rect 126336 0 126448 800
rect 126896 0 127008 800
rect 127456 0 127568 800
rect 128016 0 128128 800
rect 128576 0 128688 800
rect 129136 0 129248 800
rect 129696 0 129808 800
rect 130256 0 130368 800
rect 130816 0 130928 800
rect 131376 0 131488 800
rect 131936 0 132048 800
rect 132496 0 132608 800
rect 133056 0 133168 800
rect 133616 0 133728 800
rect 134176 0 134288 800
rect 134736 0 134848 800
rect 135296 0 135408 800
rect 135856 0 135968 800
rect 136416 0 136528 800
rect 136976 0 137088 800
rect 137536 0 137648 800
rect 138096 0 138208 800
rect 138656 0 138768 800
rect 139216 0 139328 800
rect 139776 0 139888 800
rect 140336 0 140448 800
rect 140896 0 141008 800
rect 141456 0 141568 800
rect 142016 0 142128 800
rect 142576 0 142688 800
rect 143136 0 143248 800
rect 143696 0 143808 800
rect 144256 0 144368 800
rect 144816 0 144928 800
rect 145376 0 145488 800
rect 145936 0 146048 800
rect 146496 0 146608 800
rect 147056 0 147168 800
rect 147616 0 147728 800
rect 148176 0 148288 800
rect 148736 0 148848 800
rect 149296 0 149408 800
rect 149856 0 149968 800
rect 150416 0 150528 800
rect 150976 0 151088 800
rect 151536 0 151648 800
rect 152096 0 152208 800
rect 152656 0 152768 800
rect 153216 0 153328 800
rect 153776 0 153888 800
rect 154336 0 154448 800
rect 154896 0 155008 800
rect 155456 0 155568 800
rect 156016 0 156128 800
rect 156576 0 156688 800
rect 157136 0 157248 800
rect 157696 0 157808 800
rect 158256 0 158368 800
rect 158816 0 158928 800
rect 159376 0 159488 800
rect 159936 0 160048 800
rect 160496 0 160608 800
rect 161056 0 161168 800
rect 161616 0 161728 800
rect 162176 0 162288 800
rect 162736 0 162848 800
rect 163296 0 163408 800
rect 163856 0 163968 800
rect 164416 0 164528 800
rect 164976 0 165088 800
rect 165536 0 165648 800
rect 166096 0 166208 800
rect 166656 0 166768 800
rect 167216 0 167328 800
rect 167776 0 167888 800
rect 168336 0 168448 800
rect 168896 0 169008 800
rect 169456 0 169568 800
rect 170016 0 170128 800
rect 170576 0 170688 800
rect 171136 0 171248 800
rect 171696 0 171808 800
rect 172256 0 172368 800
rect 172816 0 172928 800
rect 173376 0 173488 800
rect 173936 0 174048 800
<< via2 >>
rect 6636 15986 6692 15988
rect 6636 15934 6638 15986
rect 6638 15934 6690 15986
rect 6690 15934 6692 15986
rect 6636 15932 6692 15934
rect 2156 15874 2212 15876
rect 2156 15822 2158 15874
rect 2158 15822 2210 15874
rect 2210 15822 2212 15874
rect 2156 15820 2212 15822
rect 10444 15986 10500 15988
rect 10444 15934 10446 15986
rect 10446 15934 10498 15986
rect 10498 15934 10500 15986
rect 10444 15932 10500 15934
rect 9772 15596 9828 15652
rect 11452 15596 11508 15652
rect 10780 15426 10836 15428
rect 10780 15374 10782 15426
rect 10782 15374 10834 15426
rect 10834 15374 10836 15426
rect 10780 15372 10836 15374
rect 12124 15426 12180 15428
rect 12124 15374 12126 15426
rect 12126 15374 12178 15426
rect 12178 15374 12180 15426
rect 12124 15372 12180 15374
rect 12572 16210 12628 16212
rect 12572 16158 12574 16210
rect 12574 16158 12626 16210
rect 12626 16158 12628 16210
rect 12572 16156 12628 16158
rect 17724 16156 17780 16212
rect 16828 16044 16884 16100
rect 15932 15820 15988 15876
rect 13468 15596 13524 15652
rect 14700 15596 14756 15652
rect 16044 15708 16100 15764
rect 16716 15538 16772 15540
rect 16716 15486 16718 15538
rect 16718 15486 16770 15538
rect 16770 15486 16772 15538
rect 16716 15484 16772 15486
rect 16044 15372 16100 15428
rect 16604 15426 16660 15428
rect 16604 15374 16606 15426
rect 16606 15374 16658 15426
rect 16658 15374 16660 15426
rect 16604 15372 16660 15374
rect 14252 15202 14308 15204
rect 14252 15150 14254 15202
rect 14254 15150 14306 15202
rect 14306 15150 14308 15202
rect 14252 15148 14308 15150
rect 15372 15148 15428 15204
rect 17500 16098 17556 16100
rect 17500 16046 17502 16098
rect 17502 16046 17554 16098
rect 17554 16046 17556 16098
rect 17500 16044 17556 16046
rect 18620 16098 18676 16100
rect 18620 16046 18622 16098
rect 18622 16046 18674 16098
rect 18674 16046 18676 16098
rect 18620 16044 18676 16046
rect 19404 16044 19460 16100
rect 18060 15484 18116 15540
rect 21756 16044 21812 16100
rect 22316 16044 22372 16100
rect 23374 16490 23430 16492
rect 23374 16438 23376 16490
rect 23376 16438 23428 16490
rect 23428 16438 23430 16490
rect 23374 16436 23430 16438
rect 23478 16490 23534 16492
rect 23478 16438 23480 16490
rect 23480 16438 23532 16490
rect 23532 16438 23534 16490
rect 23478 16436 23534 16438
rect 23582 16490 23638 16492
rect 23582 16438 23584 16490
rect 23584 16438 23636 16490
rect 23636 16438 23638 16490
rect 23582 16436 23638 16438
rect 25676 16156 25732 16212
rect 27692 16044 27748 16100
rect 15932 14418 15988 14420
rect 15932 14366 15934 14418
rect 15934 14366 15986 14418
rect 15986 14366 15988 14418
rect 15932 14364 15988 14366
rect 18508 15202 18564 15204
rect 18508 15150 18510 15202
rect 18510 15150 18562 15202
rect 18562 15150 18564 15202
rect 18508 15148 18564 15150
rect 19740 15260 19796 15316
rect 20300 15260 20356 15316
rect 18060 14418 18116 14420
rect 18060 14366 18062 14418
rect 18062 14366 18114 14418
rect 18114 14366 18116 14418
rect 18060 14364 18116 14366
rect 19516 14252 19572 14308
rect 18060 13804 18116 13860
rect 18956 13804 19012 13860
rect 16940 13468 16996 13524
rect 16940 12290 16996 12292
rect 16940 12238 16942 12290
rect 16942 12238 16994 12290
rect 16994 12238 16996 12290
rect 16940 12236 16996 12238
rect 17836 13356 17892 13412
rect 19292 13746 19348 13748
rect 19292 13694 19294 13746
rect 19294 13694 19346 13746
rect 19346 13694 19348 13746
rect 19292 13692 19348 13694
rect 21196 15202 21252 15204
rect 21196 15150 21198 15202
rect 21198 15150 21250 15202
rect 21250 15150 21252 15202
rect 21196 15148 21252 15150
rect 19740 13692 19796 13748
rect 19516 13634 19572 13636
rect 19516 13582 19518 13634
rect 19518 13582 19570 13634
rect 19570 13582 19572 13634
rect 19516 13580 19572 13582
rect 20300 13692 20356 13748
rect 18956 13132 19012 13188
rect 18732 13074 18788 13076
rect 18732 13022 18734 13074
rect 18734 13022 18786 13074
rect 18786 13022 18788 13074
rect 18732 13020 18788 13022
rect 19292 13468 19348 13524
rect 17164 12236 17220 12292
rect 18508 12290 18564 12292
rect 18508 12238 18510 12290
rect 18510 12238 18562 12290
rect 18562 12238 18564 12290
rect 18508 12236 18564 12238
rect 16604 12178 16660 12180
rect 16604 12126 16606 12178
rect 16606 12126 16658 12178
rect 16658 12126 16660 12178
rect 16604 12124 16660 12126
rect 17276 12124 17332 12180
rect 18172 12178 18228 12180
rect 18172 12126 18174 12178
rect 18174 12126 18226 12178
rect 18226 12126 18228 12178
rect 18172 12124 18228 12126
rect 17276 11506 17332 11508
rect 17276 11454 17278 11506
rect 17278 11454 17330 11506
rect 17330 11454 17332 11506
rect 17276 11452 17332 11454
rect 17836 11506 17892 11508
rect 17836 11454 17838 11506
rect 17838 11454 17890 11506
rect 17890 11454 17892 11506
rect 17836 11452 17892 11454
rect 18060 11452 18116 11508
rect 18956 12236 19012 12292
rect 18508 11452 18564 11508
rect 18732 11506 18788 11508
rect 18732 11454 18734 11506
rect 18734 11454 18786 11506
rect 18786 11454 18788 11506
rect 18732 11452 18788 11454
rect 19292 12236 19348 12292
rect 19404 13356 19460 13412
rect 19852 13132 19908 13188
rect 19628 13074 19684 13076
rect 19628 13022 19630 13074
rect 19630 13022 19682 13074
rect 19682 13022 19684 13074
rect 19628 13020 19684 13022
rect 19852 12684 19908 12740
rect 19964 13020 20020 13076
rect 20188 12796 20244 12852
rect 19852 12236 19908 12292
rect 19628 11506 19684 11508
rect 19628 11454 19630 11506
rect 19630 11454 19682 11506
rect 19682 11454 19684 11506
rect 19628 11452 19684 11454
rect 20412 13356 20468 13412
rect 19852 11116 19908 11172
rect 20300 12290 20356 12292
rect 20300 12238 20302 12290
rect 20302 12238 20354 12290
rect 20354 12238 20356 12290
rect 20300 12236 20356 12238
rect 20188 11228 20244 11284
rect 20972 13468 21028 13524
rect 21196 13580 21252 13636
rect 21196 13132 21252 13188
rect 21308 14588 21364 14644
rect 29148 16098 29204 16100
rect 29148 16046 29150 16098
rect 29150 16046 29202 16098
rect 29202 16046 29204 16098
rect 29148 16044 29204 16046
rect 30380 16044 30436 16100
rect 26236 15708 26292 15764
rect 27580 15708 27636 15764
rect 26908 15596 26964 15652
rect 22092 15426 22148 15428
rect 22092 15374 22094 15426
rect 22094 15374 22146 15426
rect 22146 15374 22148 15426
rect 22092 15372 22148 15374
rect 22988 15426 23044 15428
rect 22988 15374 22990 15426
rect 22990 15374 23042 15426
rect 23042 15374 23044 15426
rect 22988 15372 23044 15374
rect 21644 14476 21700 14532
rect 21756 14364 21812 14420
rect 21868 14306 21924 14308
rect 21868 14254 21870 14306
rect 21870 14254 21922 14306
rect 21922 14254 21924 14306
rect 21868 14252 21924 14254
rect 20524 13020 20580 13076
rect 20524 12850 20580 12852
rect 20524 12798 20526 12850
rect 20526 12798 20578 12850
rect 20578 12798 20580 12850
rect 20524 12796 20580 12798
rect 20860 13074 20916 13076
rect 20860 13022 20862 13074
rect 20862 13022 20914 13074
rect 20914 13022 20916 13074
rect 20860 13020 20916 13022
rect 20636 12684 20692 12740
rect 20860 12796 20916 12852
rect 21308 13020 21364 13076
rect 21868 13356 21924 13412
rect 20972 12236 21028 12292
rect 21868 12236 21924 12292
rect 30044 15596 30100 15652
rect 27692 15148 27748 15204
rect 29708 15202 29764 15204
rect 29708 15150 29710 15202
rect 29710 15150 29762 15202
rect 29762 15150 29764 15202
rect 29708 15148 29764 15150
rect 22988 14588 23044 14644
rect 22764 13692 22820 13748
rect 25564 15036 25620 15092
rect 23374 14922 23430 14924
rect 23374 14870 23376 14922
rect 23376 14870 23428 14922
rect 23428 14870 23430 14922
rect 23374 14868 23430 14870
rect 23478 14922 23534 14924
rect 23478 14870 23480 14922
rect 23480 14870 23532 14922
rect 23532 14870 23534 14922
rect 23478 14868 23534 14870
rect 23582 14922 23638 14924
rect 23582 14870 23584 14922
rect 23584 14870 23636 14922
rect 23636 14870 23638 14922
rect 23582 14868 23638 14870
rect 23436 14642 23492 14644
rect 23436 14590 23438 14642
rect 23438 14590 23490 14642
rect 23490 14590 23492 14642
rect 23436 14588 23492 14590
rect 23212 14418 23268 14420
rect 23212 14366 23214 14418
rect 23214 14366 23266 14418
rect 23266 14366 23268 14418
rect 23212 14364 23268 14366
rect 23996 14364 24052 14420
rect 23772 13468 23828 13524
rect 23374 13354 23430 13356
rect 23374 13302 23376 13354
rect 23376 13302 23428 13354
rect 23428 13302 23430 13354
rect 23374 13300 23430 13302
rect 23478 13354 23534 13356
rect 23478 13302 23480 13354
rect 23480 13302 23532 13354
rect 23532 13302 23534 13354
rect 23478 13300 23534 13302
rect 23582 13354 23638 13356
rect 23582 13302 23584 13354
rect 23584 13302 23636 13354
rect 23636 13302 23638 13354
rect 23582 13300 23638 13302
rect 22988 13020 23044 13076
rect 22652 12290 22708 12292
rect 22652 12238 22654 12290
rect 22654 12238 22706 12290
rect 22706 12238 22708 12290
rect 22652 12236 22708 12238
rect 23660 13020 23716 13076
rect 22092 12178 22148 12180
rect 22092 12126 22094 12178
rect 22094 12126 22146 12178
rect 22146 12126 22148 12178
rect 22092 12124 22148 12126
rect 20860 12066 20916 12068
rect 20860 12014 20862 12066
rect 20862 12014 20914 12066
rect 20914 12014 20916 12066
rect 20860 12012 20916 12014
rect 21756 12066 21812 12068
rect 21756 12014 21758 12066
rect 21758 12014 21810 12066
rect 21810 12014 21812 12066
rect 21756 12012 21812 12014
rect 20636 11170 20692 11172
rect 20636 11118 20638 11170
rect 20638 11118 20690 11170
rect 20690 11118 20692 11170
rect 20636 11116 20692 11118
rect 20972 11116 21028 11172
rect 20188 10444 20244 10500
rect 19964 9938 20020 9940
rect 19964 9886 19966 9938
rect 19966 9886 20018 9938
rect 20018 9886 20020 9938
rect 19964 9884 20020 9886
rect 19516 9772 19572 9828
rect 20860 10498 20916 10500
rect 20860 10446 20862 10498
rect 20862 10446 20914 10498
rect 20914 10446 20916 10498
rect 20860 10444 20916 10446
rect 30156 15372 30212 15428
rect 30380 15260 30436 15316
rect 31164 15484 31220 15540
rect 30492 15148 30548 15204
rect 31052 15202 31108 15204
rect 31052 15150 31054 15202
rect 31054 15150 31106 15202
rect 31106 15150 31108 15202
rect 31052 15148 31108 15150
rect 25564 14252 25620 14308
rect 23996 13468 24052 13524
rect 24780 13468 24836 13524
rect 24556 13132 24612 13188
rect 25004 13074 25060 13076
rect 25004 13022 25006 13074
rect 25006 13022 25058 13074
rect 25058 13022 25060 13074
rect 25004 13020 25060 13022
rect 23374 11786 23430 11788
rect 23374 11734 23376 11786
rect 23376 11734 23428 11786
rect 23428 11734 23430 11786
rect 23374 11732 23430 11734
rect 23478 11786 23534 11788
rect 23478 11734 23480 11786
rect 23480 11734 23532 11786
rect 23532 11734 23534 11786
rect 23478 11732 23534 11734
rect 23582 11786 23638 11788
rect 23582 11734 23584 11786
rect 23584 11734 23636 11786
rect 23636 11734 23638 11786
rect 23582 11732 23638 11734
rect 21868 10610 21924 10612
rect 21868 10558 21870 10610
rect 21870 10558 21922 10610
rect 21922 10558 21924 10610
rect 21868 10556 21924 10558
rect 20188 9772 20244 9828
rect 20524 9826 20580 9828
rect 20524 9774 20526 9826
rect 20526 9774 20578 9826
rect 20578 9774 20580 9826
rect 20524 9772 20580 9774
rect 20524 9100 20580 9156
rect 23884 11564 23940 11620
rect 22652 10610 22708 10612
rect 22652 10558 22654 10610
rect 22654 10558 22706 10610
rect 22706 10558 22708 10610
rect 22652 10556 22708 10558
rect 23436 10610 23492 10612
rect 23436 10558 23438 10610
rect 23438 10558 23490 10610
rect 23490 10558 23492 10610
rect 23436 10556 23492 10558
rect 26348 13186 26404 13188
rect 26348 13134 26350 13186
rect 26350 13134 26402 13186
rect 26402 13134 26404 13186
rect 26348 13132 26404 13134
rect 31724 16380 31780 16436
rect 33516 15820 33572 15876
rect 32396 15538 32452 15540
rect 32396 15486 32398 15538
rect 32398 15486 32450 15538
rect 32450 15486 32452 15538
rect 32396 15484 32452 15486
rect 31724 15314 31780 15316
rect 31724 15262 31726 15314
rect 31726 15262 31778 15314
rect 31778 15262 31780 15314
rect 31724 15260 31780 15262
rect 33740 15314 33796 15316
rect 33740 15262 33742 15314
rect 33742 15262 33794 15314
rect 33794 15262 33796 15314
rect 33740 15260 33796 15262
rect 33180 14642 33236 14644
rect 33180 14590 33182 14642
rect 33182 14590 33234 14642
rect 33234 14590 33236 14642
rect 33180 14588 33236 14590
rect 34076 14588 34132 14644
rect 34188 15314 34244 15316
rect 34188 15262 34190 15314
rect 34190 15262 34242 15314
rect 34242 15262 34244 15314
rect 34188 15260 34244 15262
rect 35084 15426 35140 15428
rect 35084 15374 35086 15426
rect 35086 15374 35138 15426
rect 35138 15374 35140 15426
rect 35084 15372 35140 15374
rect 37436 15986 37492 15988
rect 37436 15934 37438 15986
rect 37438 15934 37490 15986
rect 37490 15934 37492 15986
rect 37436 15932 37492 15934
rect 45276 16044 45332 16100
rect 45836 16044 45892 16100
rect 48188 16210 48244 16212
rect 48188 16158 48190 16210
rect 48190 16158 48242 16210
rect 48242 16158 48244 16210
rect 48188 16156 48244 16158
rect 49868 16210 49924 16212
rect 49868 16158 49870 16210
rect 49870 16158 49922 16210
rect 49922 16158 49924 16210
rect 49868 16156 49924 16158
rect 48524 16044 48580 16100
rect 34300 15036 34356 15092
rect 35084 15148 35140 15204
rect 35084 14642 35140 14644
rect 35084 14590 35086 14642
rect 35086 14590 35138 14642
rect 35138 14590 35140 14642
rect 35084 14588 35140 14590
rect 37436 15708 37492 15764
rect 45276 15874 45332 15876
rect 45276 15822 45278 15874
rect 45278 15822 45330 15874
rect 45330 15822 45332 15874
rect 45276 15820 45332 15822
rect 49196 16098 49252 16100
rect 49196 16046 49198 16098
rect 49198 16046 49250 16098
rect 49250 16046 49252 16098
rect 49196 16044 49252 16046
rect 48524 15820 48580 15876
rect 45536 15706 45592 15708
rect 45536 15654 45538 15706
rect 45538 15654 45590 15706
rect 45590 15654 45592 15706
rect 45536 15652 45592 15654
rect 45640 15706 45696 15708
rect 45640 15654 45642 15706
rect 45642 15654 45694 15706
rect 45694 15654 45696 15706
rect 45640 15652 45696 15654
rect 45744 15706 45800 15708
rect 45744 15654 45746 15706
rect 45746 15654 45798 15706
rect 45798 15654 45800 15706
rect 45744 15652 45800 15654
rect 39564 15484 39620 15540
rect 51996 16044 52052 16100
rect 52780 16098 52836 16100
rect 52780 16046 52782 16098
rect 52782 16046 52834 16098
rect 52834 16046 52836 16098
rect 52780 16044 52836 16046
rect 52668 15596 52724 15652
rect 52108 15372 52164 15428
rect 37100 15036 37156 15092
rect 39228 14588 39284 14644
rect 31052 13132 31108 13188
rect 26236 12402 26292 12404
rect 26236 12350 26238 12402
rect 26238 12350 26290 12402
rect 26290 12350 26292 12402
rect 26236 12348 26292 12350
rect 25004 11564 25060 11620
rect 26460 11618 26516 11620
rect 26460 11566 26462 11618
rect 26462 11566 26514 11618
rect 26514 11566 26516 11618
rect 26460 11564 26516 11566
rect 25900 11394 25956 11396
rect 25900 11342 25902 11394
rect 25902 11342 25954 11394
rect 25954 11342 25956 11394
rect 25900 11340 25956 11342
rect 27132 12402 27188 12404
rect 27132 12350 27134 12402
rect 27134 12350 27186 12402
rect 27186 12350 27188 12402
rect 27132 12348 27188 12350
rect 45536 14138 45592 14140
rect 45536 14086 45538 14138
rect 45538 14086 45590 14138
rect 45590 14086 45592 14138
rect 45536 14084 45592 14086
rect 45640 14138 45696 14140
rect 45640 14086 45642 14138
rect 45642 14086 45694 14138
rect 45694 14086 45696 14138
rect 45640 14084 45696 14086
rect 45744 14138 45800 14140
rect 45744 14086 45746 14138
rect 45746 14086 45798 14138
rect 45798 14086 45800 14138
rect 45744 14084 45800 14086
rect 40236 12850 40292 12852
rect 40236 12798 40238 12850
rect 40238 12798 40290 12850
rect 40290 12798 40292 12850
rect 40236 12796 40292 12798
rect 40796 12850 40852 12852
rect 40796 12798 40798 12850
rect 40798 12798 40850 12850
rect 40850 12798 40852 12850
rect 40796 12796 40852 12798
rect 40124 12236 40180 12292
rect 39340 11618 39396 11620
rect 39340 11566 39342 11618
rect 39342 11566 39394 11618
rect 39394 11566 39396 11618
rect 39340 11564 39396 11566
rect 39788 11564 39844 11620
rect 27692 11340 27748 11396
rect 39452 11282 39508 11284
rect 39452 11230 39454 11282
rect 39454 11230 39506 11282
rect 39506 11230 39508 11282
rect 39452 11228 39508 11230
rect 24108 10610 24164 10612
rect 24108 10558 24110 10610
rect 24110 10558 24162 10610
rect 24162 10558 24164 10610
rect 24108 10556 24164 10558
rect 23374 10218 23430 10220
rect 23374 10166 23376 10218
rect 23376 10166 23428 10218
rect 23428 10166 23430 10218
rect 23374 10164 23430 10166
rect 23478 10218 23534 10220
rect 23478 10166 23480 10218
rect 23480 10166 23532 10218
rect 23532 10166 23534 10218
rect 23478 10164 23534 10166
rect 23582 10218 23638 10220
rect 23582 10166 23584 10218
rect 23584 10166 23636 10218
rect 23636 10166 23638 10218
rect 23582 10164 23638 10166
rect 21868 9884 21924 9940
rect 22764 9884 22820 9940
rect 20972 9548 21028 9604
rect 21308 9154 21364 9156
rect 21308 9102 21310 9154
rect 21310 9102 21362 9154
rect 21362 9102 21364 9154
rect 21308 9100 21364 9102
rect 21644 9100 21700 9156
rect 21756 9602 21812 9604
rect 21756 9550 21758 9602
rect 21758 9550 21810 9602
rect 21810 9550 21812 9602
rect 21756 9548 21812 9550
rect 22204 9154 22260 9156
rect 22204 9102 22206 9154
rect 22206 9102 22258 9154
rect 22258 9102 22260 9154
rect 22204 9100 22260 9102
rect 22652 9602 22708 9604
rect 22652 9550 22654 9602
rect 22654 9550 22706 9602
rect 22706 9550 22708 9602
rect 22652 9548 22708 9550
rect 23324 9938 23380 9940
rect 23324 9886 23326 9938
rect 23326 9886 23378 9938
rect 23378 9886 23380 9938
rect 23324 9884 23380 9886
rect 23772 9938 23828 9940
rect 23772 9886 23774 9938
rect 23774 9886 23826 9938
rect 23826 9886 23828 9938
rect 23772 9884 23828 9886
rect 40012 11618 40068 11620
rect 40012 11566 40014 11618
rect 40014 11566 40066 11618
rect 40066 11566 40068 11618
rect 40012 11564 40068 11566
rect 39788 10834 39844 10836
rect 39788 10782 39790 10834
rect 39790 10782 39842 10834
rect 39842 10782 39844 10834
rect 39788 10780 39844 10782
rect 40460 10834 40516 10836
rect 40460 10782 40462 10834
rect 40462 10782 40514 10834
rect 40514 10782 40516 10834
rect 40460 10780 40516 10782
rect 39900 10722 39956 10724
rect 39900 10670 39902 10722
rect 39902 10670 39954 10722
rect 39954 10670 39956 10722
rect 39900 10668 39956 10670
rect 24556 10610 24612 10612
rect 24556 10558 24558 10610
rect 24558 10558 24610 10610
rect 24610 10558 24612 10610
rect 24556 10556 24612 10558
rect 45536 12570 45592 12572
rect 45536 12518 45538 12570
rect 45538 12518 45590 12570
rect 45590 12518 45592 12570
rect 45536 12516 45592 12518
rect 45640 12570 45696 12572
rect 45640 12518 45642 12570
rect 45642 12518 45694 12570
rect 45694 12518 45696 12570
rect 45640 12516 45696 12518
rect 45744 12570 45800 12572
rect 45744 12518 45746 12570
rect 45746 12518 45798 12570
rect 45798 12518 45800 12570
rect 45744 12516 45800 12518
rect 41580 12290 41636 12292
rect 41580 12238 41582 12290
rect 41582 12238 41634 12290
rect 41634 12238 41636 12290
rect 41580 12236 41636 12238
rect 52108 11676 52164 11732
rect 40908 11564 40964 11620
rect 42140 11618 42196 11620
rect 42140 11566 42142 11618
rect 42142 11566 42194 11618
rect 42194 11566 42196 11618
rect 42140 11564 42196 11566
rect 53452 15372 53508 15428
rect 60620 16380 60676 16436
rect 60060 16156 60116 16212
rect 60844 16156 60900 16212
rect 61628 16380 61684 16436
rect 51884 11394 51940 11396
rect 51884 11342 51886 11394
rect 51886 11342 51938 11394
rect 51938 11342 51940 11394
rect 51884 11340 51940 11342
rect 40684 11282 40740 11284
rect 40684 11230 40686 11282
rect 40686 11230 40738 11282
rect 40738 11230 40740 11282
rect 40684 11228 40740 11230
rect 41468 11282 41524 11284
rect 41468 11230 41470 11282
rect 41470 11230 41522 11282
rect 41522 11230 41524 11282
rect 41468 11228 41524 11230
rect 42028 11282 42084 11284
rect 42028 11230 42030 11282
rect 42030 11230 42082 11282
rect 42082 11230 42084 11282
rect 42028 11228 42084 11230
rect 52332 11228 52388 11284
rect 41580 10722 41636 10724
rect 41580 10670 41582 10722
rect 41582 10670 41634 10722
rect 41634 10670 41636 10722
rect 41580 10668 41636 10670
rect 40572 10332 40628 10388
rect 45536 11002 45592 11004
rect 45536 10950 45538 11002
rect 45538 10950 45590 11002
rect 45590 10950 45592 11002
rect 45536 10948 45592 10950
rect 45640 11002 45696 11004
rect 45640 10950 45642 11002
rect 45642 10950 45694 11002
rect 45694 10950 45696 11002
rect 45640 10948 45696 10950
rect 45744 11002 45800 11004
rect 45744 10950 45746 11002
rect 45746 10950 45798 11002
rect 45798 10950 45800 11002
rect 45744 10948 45800 10950
rect 64092 16044 64148 16100
rect 67698 16490 67754 16492
rect 67698 16438 67700 16490
rect 67700 16438 67752 16490
rect 67752 16438 67754 16490
rect 67698 16436 67754 16438
rect 67802 16490 67858 16492
rect 67802 16438 67804 16490
rect 67804 16438 67856 16490
rect 67856 16438 67858 16490
rect 67802 16436 67858 16438
rect 67906 16490 67962 16492
rect 67906 16438 67908 16490
rect 67908 16438 67960 16490
rect 67960 16438 67962 16490
rect 67906 16436 67962 16438
rect 66556 16044 66612 16100
rect 76524 16156 76580 16212
rect 63756 15596 63812 15652
rect 63756 15148 63812 15204
rect 72716 15260 72772 15316
rect 67698 14922 67754 14924
rect 67698 14870 67700 14922
rect 67700 14870 67752 14922
rect 67752 14870 67754 14922
rect 67698 14868 67754 14870
rect 67802 14922 67858 14924
rect 67802 14870 67804 14922
rect 67804 14870 67856 14922
rect 67856 14870 67858 14922
rect 67802 14868 67858 14870
rect 67906 14922 67962 14924
rect 67906 14870 67908 14922
rect 67908 14870 67960 14922
rect 67960 14870 67962 14922
rect 67906 14868 67962 14870
rect 73612 15314 73668 15316
rect 73612 15262 73614 15314
rect 73614 15262 73666 15314
rect 73666 15262 73668 15314
rect 73612 15260 73668 15262
rect 74172 15202 74228 15204
rect 74172 15150 74174 15202
rect 74174 15150 74226 15202
rect 74226 15150 74228 15202
rect 74172 15148 74228 15150
rect 76972 15932 77028 15988
rect 91196 16044 91252 16100
rect 90076 15874 90132 15876
rect 90076 15822 90078 15874
rect 90078 15822 90130 15874
rect 90130 15822 90132 15874
rect 90076 15820 90132 15822
rect 89860 15706 89916 15708
rect 89860 15654 89862 15706
rect 89862 15654 89914 15706
rect 89914 15654 89916 15706
rect 89860 15652 89916 15654
rect 89964 15706 90020 15708
rect 89964 15654 89966 15706
rect 89966 15654 90018 15706
rect 90018 15654 90020 15706
rect 89964 15652 90020 15654
rect 90068 15706 90124 15708
rect 90068 15654 90070 15706
rect 90070 15654 90122 15706
rect 90122 15654 90124 15706
rect 90068 15652 90124 15654
rect 76972 15372 77028 15428
rect 79660 15426 79716 15428
rect 79660 15374 79662 15426
rect 79662 15374 79714 15426
rect 79714 15374 79716 15426
rect 79660 15372 79716 15374
rect 76524 15148 76580 15204
rect 77532 15260 77588 15316
rect 80444 15148 80500 15204
rect 89516 15314 89572 15316
rect 89516 15262 89518 15314
rect 89518 15262 89570 15314
rect 89570 15262 89572 15314
rect 89516 15260 89572 15262
rect 74172 14588 74228 14644
rect 88956 14642 89012 14644
rect 88956 14590 88958 14642
rect 88958 14590 89010 14642
rect 89010 14590 89012 14642
rect 88956 14588 89012 14590
rect 88396 14530 88452 14532
rect 88396 14478 88398 14530
rect 88398 14478 88450 14530
rect 88450 14478 88452 14530
rect 88396 14476 88452 14478
rect 89516 14476 89572 14532
rect 63308 14364 63364 14420
rect 60620 12684 60676 12740
rect 60284 12290 60340 12292
rect 60284 12238 60286 12290
rect 60286 12238 60338 12290
rect 60338 12238 60340 12290
rect 60284 12236 60340 12238
rect 60172 11564 60228 11620
rect 60508 11618 60564 11620
rect 60508 11566 60510 11618
rect 60510 11566 60562 11618
rect 60562 11566 60564 11618
rect 60508 11564 60564 11566
rect 53452 11340 53508 11396
rect 61740 13522 61796 13524
rect 61740 13470 61742 13522
rect 61742 13470 61794 13522
rect 61794 13470 61796 13522
rect 61740 13468 61796 13470
rect 63756 14418 63812 14420
rect 63756 14366 63758 14418
rect 63758 14366 63810 14418
rect 63810 14366 63812 14418
rect 63756 14364 63812 14366
rect 73276 14418 73332 14420
rect 73276 14366 73278 14418
rect 73278 14366 73330 14418
rect 73330 14366 73332 14418
rect 73276 14364 73332 14366
rect 90748 15820 90804 15876
rect 91980 16098 92036 16100
rect 91980 16046 91982 16098
rect 91982 16046 92034 16098
rect 92034 16046 92036 16098
rect 91980 16044 92036 16046
rect 91756 15932 91812 15988
rect 91756 15538 91812 15540
rect 91756 15486 91758 15538
rect 91758 15486 91810 15538
rect 91810 15486 91812 15538
rect 91756 15484 91812 15486
rect 92764 15986 92820 15988
rect 92764 15934 92766 15986
rect 92766 15934 92818 15986
rect 92818 15934 92820 15986
rect 92764 15932 92820 15934
rect 112022 16490 112078 16492
rect 112022 16438 112024 16490
rect 112024 16438 112076 16490
rect 112076 16438 112078 16490
rect 112022 16436 112078 16438
rect 112126 16490 112182 16492
rect 112126 16438 112128 16490
rect 112128 16438 112180 16490
rect 112180 16438 112182 16490
rect 112126 16436 112182 16438
rect 112230 16490 112286 16492
rect 112230 16438 112232 16490
rect 112232 16438 112284 16490
rect 112284 16438 112286 16490
rect 112230 16436 112286 16438
rect 156346 16490 156402 16492
rect 156346 16438 156348 16490
rect 156348 16438 156400 16490
rect 156400 16438 156402 16490
rect 156346 16436 156402 16438
rect 156450 16490 156506 16492
rect 156450 16438 156452 16490
rect 156452 16438 156504 16490
rect 156504 16438 156506 16490
rect 156450 16436 156506 16438
rect 156554 16490 156610 16492
rect 156554 16438 156556 16490
rect 156556 16438 156608 16490
rect 156608 16438 156610 16490
rect 156554 16436 156610 16438
rect 134184 15706 134240 15708
rect 134184 15654 134186 15706
rect 134186 15654 134238 15706
rect 134238 15654 134240 15706
rect 134184 15652 134240 15654
rect 134288 15706 134344 15708
rect 134288 15654 134290 15706
rect 134290 15654 134342 15706
rect 134342 15654 134344 15706
rect 134288 15652 134344 15654
rect 134392 15706 134448 15708
rect 134392 15654 134394 15706
rect 134394 15654 134446 15706
rect 134446 15654 134448 15706
rect 134392 15652 134448 15654
rect 178508 15706 178564 15708
rect 178508 15654 178510 15706
rect 178510 15654 178562 15706
rect 178562 15654 178564 15706
rect 178508 15652 178564 15654
rect 178612 15706 178668 15708
rect 178612 15654 178614 15706
rect 178614 15654 178666 15706
rect 178666 15654 178668 15706
rect 178612 15652 178668 15654
rect 178716 15706 178772 15708
rect 178716 15654 178718 15706
rect 178718 15654 178770 15706
rect 178770 15654 178772 15706
rect 178716 15652 178772 15654
rect 94892 15260 94948 15316
rect 91196 15148 91252 15204
rect 112022 14922 112078 14924
rect 112022 14870 112024 14922
rect 112024 14870 112076 14922
rect 112076 14870 112078 14922
rect 112022 14868 112078 14870
rect 112126 14922 112182 14924
rect 112126 14870 112128 14922
rect 112128 14870 112180 14922
rect 112180 14870 112182 14922
rect 112126 14868 112182 14870
rect 112230 14922 112286 14924
rect 112230 14870 112232 14922
rect 112232 14870 112284 14922
rect 112284 14870 112286 14922
rect 112230 14868 112286 14870
rect 156346 14922 156402 14924
rect 156346 14870 156348 14922
rect 156348 14870 156400 14922
rect 156400 14870 156402 14922
rect 156346 14868 156402 14870
rect 156450 14922 156506 14924
rect 156450 14870 156452 14922
rect 156452 14870 156504 14922
rect 156504 14870 156506 14922
rect 156450 14868 156506 14870
rect 156554 14922 156610 14924
rect 156554 14870 156556 14922
rect 156556 14870 156608 14922
rect 156608 14870 156610 14922
rect 156554 14868 156610 14870
rect 93884 14588 93940 14644
rect 89740 14364 89796 14420
rect 63308 13468 63364 13524
rect 67698 13354 67754 13356
rect 67698 13302 67700 13354
rect 67700 13302 67752 13354
rect 67752 13302 67754 13354
rect 67698 13300 67754 13302
rect 67802 13354 67858 13356
rect 67802 13302 67804 13354
rect 67804 13302 67856 13354
rect 67856 13302 67858 13354
rect 67802 13300 67858 13302
rect 67906 13354 67962 13356
rect 67906 13302 67908 13354
rect 67908 13302 67960 13354
rect 67960 13302 67962 13354
rect 67906 13300 67962 13302
rect 61404 11618 61460 11620
rect 61404 11566 61406 11618
rect 61406 11566 61458 11618
rect 61458 11566 61460 11618
rect 61404 11564 61460 11566
rect 62412 12738 62468 12740
rect 62412 12686 62414 12738
rect 62414 12686 62466 12738
rect 62466 12686 62468 12738
rect 62412 12684 62468 12686
rect 61740 12236 61796 12292
rect 61852 11564 61908 11620
rect 52668 11228 52724 11284
rect 62972 11618 63028 11620
rect 62972 11566 62974 11618
rect 62974 11566 63026 11618
rect 63026 11566 63028 11618
rect 62972 11564 63028 11566
rect 63644 11618 63700 11620
rect 63644 11566 63646 11618
rect 63646 11566 63698 11618
rect 63698 11566 63700 11618
rect 63644 11564 63700 11566
rect 67698 11786 67754 11788
rect 67698 11734 67700 11786
rect 67700 11734 67752 11786
rect 67752 11734 67754 11786
rect 67698 11732 67754 11734
rect 67802 11786 67858 11788
rect 67802 11734 67804 11786
rect 67804 11734 67856 11786
rect 67856 11734 67858 11786
rect 67802 11732 67858 11734
rect 67906 11786 67962 11788
rect 67906 11734 67908 11786
rect 67908 11734 67960 11786
rect 67960 11734 67962 11786
rect 67906 11732 67962 11734
rect 42700 10332 42756 10388
rect 67698 10218 67754 10220
rect 67698 10166 67700 10218
rect 67700 10166 67752 10218
rect 67752 10166 67754 10218
rect 67698 10164 67754 10166
rect 67802 10218 67858 10220
rect 67802 10166 67804 10218
rect 67804 10166 67856 10218
rect 67856 10166 67858 10218
rect 67802 10164 67858 10166
rect 67906 10218 67962 10220
rect 67906 10166 67908 10218
rect 67908 10166 67960 10218
rect 67960 10166 67962 10218
rect 67906 10164 67962 10166
rect 22540 9100 22596 9156
rect 23100 9154 23156 9156
rect 23100 9102 23102 9154
rect 23102 9102 23154 9154
rect 23154 9102 23156 9154
rect 23100 9100 23156 9102
rect 45536 9434 45592 9436
rect 45536 9382 45538 9434
rect 45538 9382 45590 9434
rect 45590 9382 45592 9434
rect 45536 9380 45592 9382
rect 45640 9434 45696 9436
rect 45640 9382 45642 9434
rect 45642 9382 45694 9434
rect 45694 9382 45696 9434
rect 45640 9380 45696 9382
rect 45744 9434 45800 9436
rect 45744 9382 45746 9434
rect 45746 9382 45798 9434
rect 45798 9382 45800 9434
rect 45744 9380 45800 9382
rect 24220 9100 24276 9156
rect 89860 14138 89916 14140
rect 89860 14086 89862 14138
rect 89862 14086 89914 14138
rect 89914 14086 89916 14138
rect 89860 14084 89916 14086
rect 89964 14138 90020 14140
rect 89964 14086 89966 14138
rect 89966 14086 90018 14138
rect 90018 14086 90020 14138
rect 89964 14084 90020 14086
rect 90068 14138 90124 14140
rect 90068 14086 90070 14138
rect 90070 14086 90122 14138
rect 90122 14086 90124 14138
rect 90068 14084 90124 14086
rect 89860 12570 89916 12572
rect 89860 12518 89862 12570
rect 89862 12518 89914 12570
rect 89914 12518 89916 12570
rect 89860 12516 89916 12518
rect 89964 12570 90020 12572
rect 89964 12518 89966 12570
rect 89966 12518 90018 12570
rect 90018 12518 90020 12570
rect 89964 12516 90020 12518
rect 90068 12570 90124 12572
rect 90068 12518 90070 12570
rect 90070 12518 90122 12570
rect 90122 12518 90124 12570
rect 90068 12516 90124 12518
rect 89860 11002 89916 11004
rect 89860 10950 89862 11002
rect 89862 10950 89914 11002
rect 89914 10950 89916 11002
rect 89860 10948 89916 10950
rect 89964 11002 90020 11004
rect 89964 10950 89966 11002
rect 89966 10950 90018 11002
rect 90018 10950 90020 11002
rect 89964 10948 90020 10950
rect 90068 11002 90124 11004
rect 90068 10950 90070 11002
rect 90070 10950 90122 11002
rect 90122 10950 90124 11002
rect 90068 10948 90124 10950
rect 89860 9434 89916 9436
rect 89860 9382 89862 9434
rect 89862 9382 89914 9434
rect 89914 9382 89916 9434
rect 89860 9380 89916 9382
rect 89964 9434 90020 9436
rect 89964 9382 89966 9434
rect 89966 9382 90018 9434
rect 90018 9382 90020 9434
rect 89964 9380 90020 9382
rect 90068 9434 90124 9436
rect 90068 9382 90070 9434
rect 90070 9382 90122 9434
rect 90122 9382 90124 9434
rect 90068 9380 90124 9382
rect 134184 14138 134240 14140
rect 134184 14086 134186 14138
rect 134186 14086 134238 14138
rect 134238 14086 134240 14138
rect 134184 14084 134240 14086
rect 134288 14138 134344 14140
rect 134288 14086 134290 14138
rect 134290 14086 134342 14138
rect 134342 14086 134344 14138
rect 134288 14084 134344 14086
rect 134392 14138 134448 14140
rect 134392 14086 134394 14138
rect 134394 14086 134446 14138
rect 134446 14086 134448 14138
rect 134392 14084 134448 14086
rect 178508 14138 178564 14140
rect 178508 14086 178510 14138
rect 178510 14086 178562 14138
rect 178562 14086 178564 14138
rect 178508 14084 178564 14086
rect 178612 14138 178668 14140
rect 178612 14086 178614 14138
rect 178614 14086 178666 14138
rect 178666 14086 178668 14138
rect 178612 14084 178668 14086
rect 178716 14138 178772 14140
rect 178716 14086 178718 14138
rect 178718 14086 178770 14138
rect 178770 14086 178772 14138
rect 178716 14084 178772 14086
rect 112022 13354 112078 13356
rect 112022 13302 112024 13354
rect 112024 13302 112076 13354
rect 112076 13302 112078 13354
rect 112022 13300 112078 13302
rect 112126 13354 112182 13356
rect 112126 13302 112128 13354
rect 112128 13302 112180 13354
rect 112180 13302 112182 13354
rect 112126 13300 112182 13302
rect 112230 13354 112286 13356
rect 112230 13302 112232 13354
rect 112232 13302 112284 13354
rect 112284 13302 112286 13354
rect 112230 13300 112286 13302
rect 156346 13354 156402 13356
rect 156346 13302 156348 13354
rect 156348 13302 156400 13354
rect 156400 13302 156402 13354
rect 156346 13300 156402 13302
rect 156450 13354 156506 13356
rect 156450 13302 156452 13354
rect 156452 13302 156504 13354
rect 156504 13302 156506 13354
rect 156450 13300 156506 13302
rect 156554 13354 156610 13356
rect 156554 13302 156556 13354
rect 156556 13302 156608 13354
rect 156608 13302 156610 13354
rect 156554 13300 156610 13302
rect 134184 12570 134240 12572
rect 134184 12518 134186 12570
rect 134186 12518 134238 12570
rect 134238 12518 134240 12570
rect 134184 12516 134240 12518
rect 134288 12570 134344 12572
rect 134288 12518 134290 12570
rect 134290 12518 134342 12570
rect 134342 12518 134344 12570
rect 134288 12516 134344 12518
rect 134392 12570 134448 12572
rect 134392 12518 134394 12570
rect 134394 12518 134446 12570
rect 134446 12518 134448 12570
rect 134392 12516 134448 12518
rect 178508 12570 178564 12572
rect 178508 12518 178510 12570
rect 178510 12518 178562 12570
rect 178562 12518 178564 12570
rect 178508 12516 178564 12518
rect 178612 12570 178668 12572
rect 178612 12518 178614 12570
rect 178614 12518 178666 12570
rect 178666 12518 178668 12570
rect 178612 12516 178668 12518
rect 178716 12570 178772 12572
rect 178716 12518 178718 12570
rect 178718 12518 178770 12570
rect 178770 12518 178772 12570
rect 178716 12516 178772 12518
rect 112022 11786 112078 11788
rect 112022 11734 112024 11786
rect 112024 11734 112076 11786
rect 112076 11734 112078 11786
rect 112022 11732 112078 11734
rect 112126 11786 112182 11788
rect 112126 11734 112128 11786
rect 112128 11734 112180 11786
rect 112180 11734 112182 11786
rect 112126 11732 112182 11734
rect 112230 11786 112286 11788
rect 112230 11734 112232 11786
rect 112232 11734 112284 11786
rect 112284 11734 112286 11786
rect 112230 11732 112286 11734
rect 156346 11786 156402 11788
rect 156346 11734 156348 11786
rect 156348 11734 156400 11786
rect 156400 11734 156402 11786
rect 156346 11732 156402 11734
rect 156450 11786 156506 11788
rect 156450 11734 156452 11786
rect 156452 11734 156504 11786
rect 156504 11734 156506 11786
rect 156450 11732 156506 11734
rect 156554 11786 156610 11788
rect 156554 11734 156556 11786
rect 156556 11734 156608 11786
rect 156608 11734 156610 11786
rect 156554 11732 156610 11734
rect 134184 11002 134240 11004
rect 134184 10950 134186 11002
rect 134186 10950 134238 11002
rect 134238 10950 134240 11002
rect 134184 10948 134240 10950
rect 134288 11002 134344 11004
rect 134288 10950 134290 11002
rect 134290 10950 134342 11002
rect 134342 10950 134344 11002
rect 134288 10948 134344 10950
rect 134392 11002 134448 11004
rect 134392 10950 134394 11002
rect 134394 10950 134446 11002
rect 134446 10950 134448 11002
rect 134392 10948 134448 10950
rect 178508 11002 178564 11004
rect 178508 10950 178510 11002
rect 178510 10950 178562 11002
rect 178562 10950 178564 11002
rect 178508 10948 178564 10950
rect 178612 11002 178668 11004
rect 178612 10950 178614 11002
rect 178614 10950 178666 11002
rect 178666 10950 178668 11002
rect 178612 10948 178668 10950
rect 178716 11002 178772 11004
rect 178716 10950 178718 11002
rect 178718 10950 178770 11002
rect 178770 10950 178772 11002
rect 178716 10948 178772 10950
rect 112022 10218 112078 10220
rect 112022 10166 112024 10218
rect 112024 10166 112076 10218
rect 112076 10166 112078 10218
rect 112022 10164 112078 10166
rect 112126 10218 112182 10220
rect 112126 10166 112128 10218
rect 112128 10166 112180 10218
rect 112180 10166 112182 10218
rect 112126 10164 112182 10166
rect 112230 10218 112286 10220
rect 112230 10166 112232 10218
rect 112232 10166 112284 10218
rect 112284 10166 112286 10218
rect 112230 10164 112286 10166
rect 156346 10218 156402 10220
rect 156346 10166 156348 10218
rect 156348 10166 156400 10218
rect 156400 10166 156402 10218
rect 156346 10164 156402 10166
rect 156450 10218 156506 10220
rect 156450 10166 156452 10218
rect 156452 10166 156504 10218
rect 156504 10166 156506 10218
rect 156450 10164 156506 10166
rect 156554 10218 156610 10220
rect 156554 10166 156556 10218
rect 156556 10166 156608 10218
rect 156608 10166 156610 10218
rect 156554 10164 156610 10166
rect 134184 9434 134240 9436
rect 134184 9382 134186 9434
rect 134186 9382 134238 9434
rect 134238 9382 134240 9434
rect 134184 9380 134240 9382
rect 134288 9434 134344 9436
rect 134288 9382 134290 9434
rect 134290 9382 134342 9434
rect 134342 9382 134344 9434
rect 134288 9380 134344 9382
rect 134392 9434 134448 9436
rect 134392 9382 134394 9434
rect 134394 9382 134446 9434
rect 134446 9382 134448 9434
rect 134392 9380 134448 9382
rect 178508 9434 178564 9436
rect 178508 9382 178510 9434
rect 178510 9382 178562 9434
rect 178562 9382 178564 9434
rect 178508 9380 178564 9382
rect 178612 9434 178668 9436
rect 178612 9382 178614 9434
rect 178614 9382 178666 9434
rect 178666 9382 178668 9434
rect 178612 9380 178668 9382
rect 178716 9434 178772 9436
rect 178716 9382 178718 9434
rect 178718 9382 178770 9434
rect 178770 9382 178772 9434
rect 178716 9380 178772 9382
rect 93884 9266 93940 9268
rect 93884 9214 93886 9266
rect 93886 9214 93938 9266
rect 93938 9214 93940 9266
rect 93884 9212 93940 9214
rect 94444 9266 94500 9268
rect 94444 9214 94446 9266
rect 94446 9214 94498 9266
rect 94498 9214 94500 9266
rect 94444 9212 94500 9214
rect 89740 8988 89796 9044
rect 23374 8650 23430 8652
rect 23374 8598 23376 8650
rect 23376 8598 23428 8650
rect 23428 8598 23430 8650
rect 23374 8596 23430 8598
rect 23478 8650 23534 8652
rect 23478 8598 23480 8650
rect 23480 8598 23532 8650
rect 23532 8598 23534 8650
rect 23478 8596 23534 8598
rect 23582 8650 23638 8652
rect 23582 8598 23584 8650
rect 23584 8598 23636 8650
rect 23636 8598 23638 8650
rect 23582 8596 23638 8598
rect 67698 8650 67754 8652
rect 67698 8598 67700 8650
rect 67700 8598 67752 8650
rect 67752 8598 67754 8650
rect 67698 8596 67754 8598
rect 67802 8650 67858 8652
rect 67802 8598 67804 8650
rect 67804 8598 67856 8650
rect 67856 8598 67858 8650
rect 67802 8596 67858 8598
rect 67906 8650 67962 8652
rect 67906 8598 67908 8650
rect 67908 8598 67960 8650
rect 67960 8598 67962 8650
rect 67906 8596 67962 8598
rect 45536 7866 45592 7868
rect 45536 7814 45538 7866
rect 45538 7814 45590 7866
rect 45590 7814 45592 7866
rect 45536 7812 45592 7814
rect 45640 7866 45696 7868
rect 45640 7814 45642 7866
rect 45642 7814 45694 7866
rect 45694 7814 45696 7866
rect 45640 7812 45696 7814
rect 45744 7866 45800 7868
rect 45744 7814 45746 7866
rect 45746 7814 45798 7866
rect 45798 7814 45800 7866
rect 45744 7812 45800 7814
rect 89860 7866 89916 7868
rect 89860 7814 89862 7866
rect 89862 7814 89914 7866
rect 89914 7814 89916 7866
rect 89860 7812 89916 7814
rect 89964 7866 90020 7868
rect 89964 7814 89966 7866
rect 89966 7814 90018 7866
rect 90018 7814 90020 7866
rect 89964 7812 90020 7814
rect 90068 7866 90124 7868
rect 90068 7814 90070 7866
rect 90070 7814 90122 7866
rect 90122 7814 90124 7866
rect 90068 7812 90124 7814
rect 23374 7082 23430 7084
rect 23374 7030 23376 7082
rect 23376 7030 23428 7082
rect 23428 7030 23430 7082
rect 23374 7028 23430 7030
rect 23478 7082 23534 7084
rect 23478 7030 23480 7082
rect 23480 7030 23532 7082
rect 23532 7030 23534 7082
rect 23478 7028 23534 7030
rect 23582 7082 23638 7084
rect 23582 7030 23584 7082
rect 23584 7030 23636 7082
rect 23636 7030 23638 7082
rect 23582 7028 23638 7030
rect 67698 7082 67754 7084
rect 67698 7030 67700 7082
rect 67700 7030 67752 7082
rect 67752 7030 67754 7082
rect 67698 7028 67754 7030
rect 67802 7082 67858 7084
rect 67802 7030 67804 7082
rect 67804 7030 67856 7082
rect 67856 7030 67858 7082
rect 67802 7028 67858 7030
rect 67906 7082 67962 7084
rect 67906 7030 67908 7082
rect 67908 7030 67960 7082
rect 67960 7030 67962 7082
rect 67906 7028 67962 7030
rect 45536 6298 45592 6300
rect 45536 6246 45538 6298
rect 45538 6246 45590 6298
rect 45590 6246 45592 6298
rect 45536 6244 45592 6246
rect 45640 6298 45696 6300
rect 45640 6246 45642 6298
rect 45642 6246 45694 6298
rect 45694 6246 45696 6298
rect 45640 6244 45696 6246
rect 45744 6298 45800 6300
rect 45744 6246 45746 6298
rect 45746 6246 45798 6298
rect 45798 6246 45800 6298
rect 45744 6244 45800 6246
rect 89860 6298 89916 6300
rect 89860 6246 89862 6298
rect 89862 6246 89914 6298
rect 89914 6246 89916 6298
rect 89860 6244 89916 6246
rect 89964 6298 90020 6300
rect 89964 6246 89966 6298
rect 89966 6246 90018 6298
rect 90018 6246 90020 6298
rect 89964 6244 90020 6246
rect 90068 6298 90124 6300
rect 90068 6246 90070 6298
rect 90070 6246 90122 6298
rect 90122 6246 90124 6298
rect 90068 6244 90124 6246
rect 23374 5514 23430 5516
rect 23374 5462 23376 5514
rect 23376 5462 23428 5514
rect 23428 5462 23430 5514
rect 23374 5460 23430 5462
rect 23478 5514 23534 5516
rect 23478 5462 23480 5514
rect 23480 5462 23532 5514
rect 23532 5462 23534 5514
rect 23478 5460 23534 5462
rect 23582 5514 23638 5516
rect 23582 5462 23584 5514
rect 23584 5462 23636 5514
rect 23636 5462 23638 5514
rect 23582 5460 23638 5462
rect 67698 5514 67754 5516
rect 67698 5462 67700 5514
rect 67700 5462 67752 5514
rect 67752 5462 67754 5514
rect 67698 5460 67754 5462
rect 67802 5514 67858 5516
rect 67802 5462 67804 5514
rect 67804 5462 67856 5514
rect 67856 5462 67858 5514
rect 67802 5460 67858 5462
rect 67906 5514 67962 5516
rect 67906 5462 67908 5514
rect 67908 5462 67960 5514
rect 67960 5462 67962 5514
rect 67906 5460 67962 5462
rect 45536 4730 45592 4732
rect 45536 4678 45538 4730
rect 45538 4678 45590 4730
rect 45590 4678 45592 4730
rect 45536 4676 45592 4678
rect 45640 4730 45696 4732
rect 45640 4678 45642 4730
rect 45642 4678 45694 4730
rect 45694 4678 45696 4730
rect 45640 4676 45696 4678
rect 45744 4730 45800 4732
rect 45744 4678 45746 4730
rect 45746 4678 45798 4730
rect 45798 4678 45800 4730
rect 45744 4676 45800 4678
rect 89860 4730 89916 4732
rect 89860 4678 89862 4730
rect 89862 4678 89914 4730
rect 89914 4678 89916 4730
rect 89860 4676 89916 4678
rect 89964 4730 90020 4732
rect 89964 4678 89966 4730
rect 89966 4678 90018 4730
rect 90018 4678 90020 4730
rect 89964 4676 90020 4678
rect 90068 4730 90124 4732
rect 90068 4678 90070 4730
rect 90070 4678 90122 4730
rect 90122 4678 90124 4730
rect 90068 4676 90124 4678
rect 95340 8988 95396 9044
rect 95564 9042 95620 9044
rect 95564 8990 95566 9042
rect 95566 8990 95618 9042
rect 95618 8990 95620 9042
rect 95564 8988 95620 8990
rect 94780 4284 94836 4340
rect 112022 8650 112078 8652
rect 112022 8598 112024 8650
rect 112024 8598 112076 8650
rect 112076 8598 112078 8650
rect 112022 8596 112078 8598
rect 112126 8650 112182 8652
rect 112126 8598 112128 8650
rect 112128 8598 112180 8650
rect 112180 8598 112182 8650
rect 112126 8596 112182 8598
rect 112230 8650 112286 8652
rect 112230 8598 112232 8650
rect 112232 8598 112284 8650
rect 112284 8598 112286 8650
rect 112230 8596 112286 8598
rect 156346 8650 156402 8652
rect 156346 8598 156348 8650
rect 156348 8598 156400 8650
rect 156400 8598 156402 8650
rect 156346 8596 156402 8598
rect 156450 8650 156506 8652
rect 156450 8598 156452 8650
rect 156452 8598 156504 8650
rect 156504 8598 156506 8650
rect 156450 8596 156506 8598
rect 156554 8650 156610 8652
rect 156554 8598 156556 8650
rect 156556 8598 156608 8650
rect 156608 8598 156610 8650
rect 156554 8596 156610 8598
rect 134184 7866 134240 7868
rect 134184 7814 134186 7866
rect 134186 7814 134238 7866
rect 134238 7814 134240 7866
rect 134184 7812 134240 7814
rect 134288 7866 134344 7868
rect 134288 7814 134290 7866
rect 134290 7814 134342 7866
rect 134342 7814 134344 7866
rect 134288 7812 134344 7814
rect 134392 7866 134448 7868
rect 134392 7814 134394 7866
rect 134394 7814 134446 7866
rect 134446 7814 134448 7866
rect 134392 7812 134448 7814
rect 178508 7866 178564 7868
rect 178508 7814 178510 7866
rect 178510 7814 178562 7866
rect 178562 7814 178564 7866
rect 178508 7812 178564 7814
rect 178612 7866 178668 7868
rect 178612 7814 178614 7866
rect 178614 7814 178666 7866
rect 178666 7814 178668 7866
rect 178612 7812 178668 7814
rect 178716 7866 178772 7868
rect 178716 7814 178718 7866
rect 178718 7814 178770 7866
rect 178770 7814 178772 7866
rect 178716 7812 178772 7814
rect 112022 7082 112078 7084
rect 112022 7030 112024 7082
rect 112024 7030 112076 7082
rect 112076 7030 112078 7082
rect 112022 7028 112078 7030
rect 112126 7082 112182 7084
rect 112126 7030 112128 7082
rect 112128 7030 112180 7082
rect 112180 7030 112182 7082
rect 112126 7028 112182 7030
rect 112230 7082 112286 7084
rect 112230 7030 112232 7082
rect 112232 7030 112284 7082
rect 112284 7030 112286 7082
rect 112230 7028 112286 7030
rect 156346 7082 156402 7084
rect 156346 7030 156348 7082
rect 156348 7030 156400 7082
rect 156400 7030 156402 7082
rect 156346 7028 156402 7030
rect 156450 7082 156506 7084
rect 156450 7030 156452 7082
rect 156452 7030 156504 7082
rect 156504 7030 156506 7082
rect 156450 7028 156506 7030
rect 156554 7082 156610 7084
rect 156554 7030 156556 7082
rect 156556 7030 156608 7082
rect 156608 7030 156610 7082
rect 156554 7028 156610 7030
rect 134184 6298 134240 6300
rect 134184 6246 134186 6298
rect 134186 6246 134238 6298
rect 134238 6246 134240 6298
rect 134184 6244 134240 6246
rect 134288 6298 134344 6300
rect 134288 6246 134290 6298
rect 134290 6246 134342 6298
rect 134342 6246 134344 6298
rect 134288 6244 134344 6246
rect 134392 6298 134448 6300
rect 134392 6246 134394 6298
rect 134394 6246 134446 6298
rect 134446 6246 134448 6298
rect 134392 6244 134448 6246
rect 178508 6298 178564 6300
rect 178508 6246 178510 6298
rect 178510 6246 178562 6298
rect 178562 6246 178564 6298
rect 178508 6244 178564 6246
rect 178612 6298 178668 6300
rect 178612 6246 178614 6298
rect 178614 6246 178666 6298
rect 178666 6246 178668 6298
rect 178612 6244 178668 6246
rect 178716 6298 178772 6300
rect 178716 6246 178718 6298
rect 178718 6246 178770 6298
rect 178770 6246 178772 6298
rect 178716 6244 178772 6246
rect 112022 5514 112078 5516
rect 112022 5462 112024 5514
rect 112024 5462 112076 5514
rect 112076 5462 112078 5514
rect 112022 5460 112078 5462
rect 112126 5514 112182 5516
rect 112126 5462 112128 5514
rect 112128 5462 112180 5514
rect 112180 5462 112182 5514
rect 112126 5460 112182 5462
rect 112230 5514 112286 5516
rect 112230 5462 112232 5514
rect 112232 5462 112284 5514
rect 112284 5462 112286 5514
rect 112230 5460 112286 5462
rect 156346 5514 156402 5516
rect 156346 5462 156348 5514
rect 156348 5462 156400 5514
rect 156400 5462 156402 5514
rect 156346 5460 156402 5462
rect 156450 5514 156506 5516
rect 156450 5462 156452 5514
rect 156452 5462 156504 5514
rect 156504 5462 156506 5514
rect 156450 5460 156506 5462
rect 156554 5514 156610 5516
rect 156554 5462 156556 5514
rect 156556 5462 156608 5514
rect 156608 5462 156610 5514
rect 156554 5460 156610 5462
rect 134184 4730 134240 4732
rect 134184 4678 134186 4730
rect 134186 4678 134238 4730
rect 134238 4678 134240 4730
rect 134184 4676 134240 4678
rect 134288 4730 134344 4732
rect 134288 4678 134290 4730
rect 134290 4678 134342 4730
rect 134342 4678 134344 4730
rect 134288 4676 134344 4678
rect 134392 4730 134448 4732
rect 134392 4678 134394 4730
rect 134394 4678 134446 4730
rect 134446 4678 134448 4730
rect 134392 4676 134448 4678
rect 178508 4730 178564 4732
rect 178508 4678 178510 4730
rect 178510 4678 178562 4730
rect 178562 4678 178564 4730
rect 178508 4676 178564 4678
rect 178612 4730 178668 4732
rect 178612 4678 178614 4730
rect 178614 4678 178666 4730
rect 178666 4678 178668 4730
rect 178612 4676 178668 4678
rect 178716 4730 178772 4732
rect 178716 4678 178718 4730
rect 178718 4678 178770 4730
rect 178770 4678 178772 4730
rect 178716 4676 178772 4678
rect 95900 4172 95956 4228
rect 119644 4284 119700 4340
rect 23374 3946 23430 3948
rect 23374 3894 23376 3946
rect 23376 3894 23428 3946
rect 23428 3894 23430 3946
rect 23374 3892 23430 3894
rect 23478 3946 23534 3948
rect 23478 3894 23480 3946
rect 23480 3894 23532 3946
rect 23532 3894 23534 3946
rect 23478 3892 23534 3894
rect 23582 3946 23638 3948
rect 23582 3894 23584 3946
rect 23584 3894 23636 3946
rect 23636 3894 23638 3946
rect 23582 3892 23638 3894
rect 67698 3946 67754 3948
rect 67698 3894 67700 3946
rect 67700 3894 67752 3946
rect 67752 3894 67754 3946
rect 67698 3892 67754 3894
rect 67802 3946 67858 3948
rect 67802 3894 67804 3946
rect 67804 3894 67856 3946
rect 67856 3894 67858 3946
rect 67802 3892 67858 3894
rect 67906 3946 67962 3948
rect 67906 3894 67908 3946
rect 67908 3894 67960 3946
rect 67960 3894 67962 3946
rect 67906 3892 67962 3894
rect 112022 3946 112078 3948
rect 112022 3894 112024 3946
rect 112024 3894 112076 3946
rect 112076 3894 112078 3946
rect 112022 3892 112078 3894
rect 112126 3946 112182 3948
rect 112126 3894 112128 3946
rect 112128 3894 112180 3946
rect 112180 3894 112182 3946
rect 112126 3892 112182 3894
rect 112230 3946 112286 3948
rect 112230 3894 112232 3946
rect 112232 3894 112284 3946
rect 112284 3894 112286 3946
rect 112230 3892 112286 3894
rect 12684 3276 12740 3332
rect 13580 3330 13636 3332
rect 13580 3278 13582 3330
rect 13582 3278 13634 3330
rect 13634 3278 13636 3330
rect 13580 3276 13636 3278
rect 24444 3276 24500 3332
rect 25340 3330 25396 3332
rect 25340 3278 25342 3330
rect 25342 3278 25394 3330
rect 25394 3278 25396 3330
rect 25340 3276 25396 3278
rect 36204 3276 36260 3332
rect 37100 3330 37156 3332
rect 37100 3278 37102 3330
rect 37102 3278 37154 3330
rect 37154 3278 37156 3330
rect 37100 3276 37156 3278
rect 45536 3162 45592 3164
rect 45536 3110 45538 3162
rect 45538 3110 45590 3162
rect 45590 3110 45592 3162
rect 45536 3108 45592 3110
rect 45640 3162 45696 3164
rect 45640 3110 45642 3162
rect 45642 3110 45694 3162
rect 45694 3110 45696 3162
rect 45640 3108 45696 3110
rect 45744 3162 45800 3164
rect 45744 3110 45746 3162
rect 45746 3110 45798 3162
rect 45798 3110 45800 3162
rect 45744 3108 45800 3110
rect 47964 3276 48020 3332
rect 48860 3330 48916 3332
rect 48860 3278 48862 3330
rect 48862 3278 48914 3330
rect 48914 3278 48916 3330
rect 48860 3276 48916 3278
rect 59724 3276 59780 3332
rect 60620 3330 60676 3332
rect 60620 3278 60622 3330
rect 60622 3278 60674 3330
rect 60674 3278 60676 3330
rect 60620 3276 60676 3278
rect 89860 3162 89916 3164
rect 89860 3110 89862 3162
rect 89862 3110 89914 3162
rect 89914 3110 89916 3162
rect 89860 3108 89916 3110
rect 89964 3162 90020 3164
rect 89964 3110 89966 3162
rect 89966 3110 90018 3162
rect 90018 3110 90020 3162
rect 89964 3108 90020 3110
rect 90068 3162 90124 3164
rect 90068 3110 90070 3162
rect 90070 3110 90122 3162
rect 90122 3110 90124 3162
rect 90068 3108 90124 3110
rect 121324 4172 121380 4228
rect 156346 3946 156402 3948
rect 156346 3894 156348 3946
rect 156348 3894 156400 3946
rect 156400 3894 156402 3946
rect 156346 3892 156402 3894
rect 156450 3946 156506 3948
rect 156450 3894 156452 3946
rect 156452 3894 156504 3946
rect 156504 3894 156506 3946
rect 156450 3892 156506 3894
rect 156554 3946 156610 3948
rect 156554 3894 156556 3946
rect 156556 3894 156608 3946
rect 156608 3894 156610 3946
rect 156554 3892 156610 3894
rect 134184 3162 134240 3164
rect 134184 3110 134186 3162
rect 134186 3110 134238 3162
rect 134238 3110 134240 3162
rect 134184 3108 134240 3110
rect 134288 3162 134344 3164
rect 134288 3110 134290 3162
rect 134290 3110 134342 3162
rect 134342 3110 134344 3162
rect 134288 3108 134344 3110
rect 134392 3162 134448 3164
rect 134392 3110 134394 3162
rect 134394 3110 134446 3162
rect 134446 3110 134448 3162
rect 134392 3108 134448 3110
rect 173964 3276 174020 3332
rect 174972 3330 175028 3332
rect 174972 3278 174974 3330
rect 174974 3278 175026 3330
rect 175026 3278 175028 3330
rect 174972 3276 175028 3278
rect 178508 3162 178564 3164
rect 178508 3110 178510 3162
rect 178510 3110 178562 3162
rect 178562 3110 178564 3162
rect 178508 3108 178564 3110
rect 178612 3162 178668 3164
rect 178612 3110 178614 3162
rect 178614 3110 178666 3162
rect 178666 3110 178668 3162
rect 178612 3108 178668 3110
rect 178716 3162 178772 3164
rect 178716 3110 178718 3162
rect 178718 3110 178770 3162
rect 178770 3110 178772 3162
rect 178716 3108 178772 3110
<< metal3 >>
rect 23364 16436 23374 16492
rect 23430 16436 23478 16492
rect 23534 16436 23582 16492
rect 23638 16436 23648 16492
rect 67688 16436 67698 16492
rect 67754 16436 67802 16492
rect 67858 16436 67906 16492
rect 67962 16436 67972 16492
rect 112012 16436 112022 16492
rect 112078 16436 112126 16492
rect 112182 16436 112230 16492
rect 112286 16436 112296 16492
rect 156336 16436 156346 16492
rect 156402 16436 156450 16492
rect 156506 16436 156554 16492
rect 156610 16436 156620 16492
rect 31714 16380 31724 16436
rect 31780 16380 60620 16436
rect 60676 16380 61628 16436
rect 61684 16380 61694 16436
rect 12562 16156 12572 16212
rect 12628 16156 17724 16212
rect 17780 16156 17790 16212
rect 25666 16156 25676 16212
rect 25732 16156 48188 16212
rect 48244 16156 49868 16212
rect 49924 16156 49934 16212
rect 50092 16156 60060 16212
rect 60116 16156 60844 16212
rect 60900 16156 76524 16212
rect 76580 16156 76590 16212
rect 50092 16100 50148 16156
rect 16818 16044 16828 16100
rect 16884 16044 17500 16100
rect 17556 16044 18620 16100
rect 18676 16044 19404 16100
rect 19460 16044 19470 16100
rect 21746 16044 21756 16100
rect 21812 16044 22316 16100
rect 22372 16044 22382 16100
rect 27682 16044 27692 16100
rect 27748 16044 29148 16100
rect 29204 16044 30380 16100
rect 30436 16044 30446 16100
rect 45266 16044 45276 16100
rect 45332 16044 45836 16100
rect 45892 16044 45902 16100
rect 48514 16044 48524 16100
rect 48580 16044 49196 16100
rect 49252 16044 50148 16100
rect 51986 16044 51996 16100
rect 52052 16044 52780 16100
rect 52836 16044 52846 16100
rect 64082 16044 64092 16100
rect 64148 16044 66556 16100
rect 66612 16044 66622 16100
rect 91186 16044 91196 16100
rect 91252 16044 91980 16100
rect 92036 16044 92046 16100
rect 6626 15932 6636 15988
rect 6692 15932 10444 15988
rect 10500 15932 10510 15988
rect 37426 15932 37436 15988
rect 37492 15932 76972 15988
rect 77028 15932 77038 15988
rect 91746 15932 91756 15988
rect 91812 15932 92764 15988
rect 92820 15932 92830 15988
rect 2146 15820 2156 15876
rect 2212 15820 15932 15876
rect 15988 15820 15998 15876
rect 31892 15820 33516 15876
rect 33572 15820 45276 15876
rect 45332 15820 48524 15876
rect 48580 15820 48590 15876
rect 90066 15820 90076 15876
rect 90132 15820 90748 15876
rect 90804 15820 90814 15876
rect 16034 15708 16044 15764
rect 16100 15708 26236 15764
rect 26292 15708 27580 15764
rect 27636 15708 27646 15764
rect 31892 15652 31948 15820
rect 37436 15764 37492 15820
rect 37426 15708 37436 15764
rect 37492 15708 37502 15764
rect 45526 15652 45536 15708
rect 45592 15652 45640 15708
rect 45696 15652 45744 15708
rect 45800 15652 45810 15708
rect 89850 15652 89860 15708
rect 89916 15652 89964 15708
rect 90020 15652 90068 15708
rect 90124 15652 90134 15708
rect 134174 15652 134184 15708
rect 134240 15652 134288 15708
rect 134344 15652 134392 15708
rect 134448 15652 134458 15708
rect 178498 15652 178508 15708
rect 178564 15652 178612 15708
rect 178668 15652 178716 15708
rect 178772 15652 178782 15708
rect 9762 15596 9772 15652
rect 9828 15596 11452 15652
rect 11508 15596 13468 15652
rect 13524 15596 14700 15652
rect 14756 15596 26908 15652
rect 26964 15596 30044 15652
rect 30100 15596 31948 15652
rect 52658 15596 52668 15652
rect 52724 15596 63756 15652
rect 63812 15596 63822 15652
rect 16706 15484 16716 15540
rect 16772 15484 18060 15540
rect 18116 15484 18126 15540
rect 31154 15484 31164 15540
rect 31220 15484 32396 15540
rect 32452 15484 32462 15540
rect 39554 15484 39564 15540
rect 39620 15484 91756 15540
rect 91812 15484 91822 15540
rect 10770 15372 10780 15428
rect 10836 15372 12124 15428
rect 12180 15372 12190 15428
rect 16034 15372 16044 15428
rect 16100 15372 16604 15428
rect 16660 15372 16670 15428
rect 22082 15372 22092 15428
rect 22148 15372 22988 15428
rect 23044 15372 30156 15428
rect 30212 15372 35084 15428
rect 35140 15372 52108 15428
rect 52164 15372 53452 15428
rect 53508 15372 53518 15428
rect 76962 15372 76972 15428
rect 77028 15372 79660 15428
rect 79716 15372 79726 15428
rect 19730 15260 19740 15316
rect 19796 15260 20300 15316
rect 20356 15260 20366 15316
rect 30370 15260 30380 15316
rect 30436 15260 31724 15316
rect 31780 15260 33740 15316
rect 33796 15260 34188 15316
rect 34244 15260 34254 15316
rect 72706 15260 72716 15316
rect 72772 15260 73612 15316
rect 73668 15260 77532 15316
rect 77588 15260 77598 15316
rect 89506 15260 89516 15316
rect 89572 15260 94892 15316
rect 94948 15260 94958 15316
rect 14242 15148 14252 15204
rect 14308 15148 15372 15204
rect 15428 15148 15438 15204
rect 18498 15148 18508 15204
rect 18564 15148 21196 15204
rect 21252 15148 21262 15204
rect 26796 15148 27692 15204
rect 27748 15148 27758 15204
rect 29698 15148 29708 15204
rect 29764 15148 30492 15204
rect 30548 15148 30558 15204
rect 31042 15148 31052 15204
rect 31108 15148 35084 15204
rect 35140 15148 35150 15204
rect 63746 15148 63756 15204
rect 63812 15148 74172 15204
rect 74228 15148 74238 15204
rect 76514 15148 76524 15204
rect 76580 15148 80444 15204
rect 80500 15148 91196 15204
rect 91252 15148 91262 15204
rect 26796 15092 26852 15148
rect 25554 15036 25564 15092
rect 25620 15036 26852 15092
rect 34290 15036 34300 15092
rect 34356 15036 37100 15092
rect 37156 15036 37166 15092
rect 23364 14868 23374 14924
rect 23430 14868 23478 14924
rect 23534 14868 23582 14924
rect 23638 14868 23648 14924
rect 67688 14868 67698 14924
rect 67754 14868 67802 14924
rect 67858 14868 67906 14924
rect 67962 14868 67972 14924
rect 112012 14868 112022 14924
rect 112078 14868 112126 14924
rect 112182 14868 112230 14924
rect 112286 14868 112296 14924
rect 156336 14868 156346 14924
rect 156402 14868 156450 14924
rect 156506 14868 156554 14924
rect 156610 14868 156620 14924
rect 21298 14588 21308 14644
rect 21364 14588 22988 14644
rect 23044 14588 23436 14644
rect 23492 14588 23502 14644
rect 31892 14588 33180 14644
rect 33236 14588 34076 14644
rect 34132 14588 34142 14644
rect 35074 14588 35084 14644
rect 35140 14588 39228 14644
rect 39284 14588 39294 14644
rect 74162 14588 74172 14644
rect 74228 14588 88956 14644
rect 89012 14588 93884 14644
rect 93940 14588 93950 14644
rect 31892 14532 31948 14588
rect 21634 14476 21644 14532
rect 21700 14476 31948 14532
rect 88386 14476 88396 14532
rect 88452 14476 89516 14532
rect 89572 14476 89582 14532
rect 15922 14364 15932 14420
rect 15988 14364 18060 14420
rect 18116 14364 18126 14420
rect 21746 14364 21756 14420
rect 21812 14364 23212 14420
rect 23268 14364 23996 14420
rect 24052 14364 24062 14420
rect 63298 14364 63308 14420
rect 63364 14364 63756 14420
rect 63812 14364 73276 14420
rect 73332 14364 89740 14420
rect 89796 14364 89806 14420
rect 19506 14252 19516 14308
rect 19572 14252 21868 14308
rect 21924 14252 25564 14308
rect 25620 14252 25630 14308
rect 45526 14084 45536 14140
rect 45592 14084 45640 14140
rect 45696 14084 45744 14140
rect 45800 14084 45810 14140
rect 89850 14084 89860 14140
rect 89916 14084 89964 14140
rect 90020 14084 90068 14140
rect 90124 14084 90134 14140
rect 134174 14084 134184 14140
rect 134240 14084 134288 14140
rect 134344 14084 134392 14140
rect 134448 14084 134458 14140
rect 178498 14084 178508 14140
rect 178564 14084 178612 14140
rect 178668 14084 178716 14140
rect 178772 14084 178782 14140
rect 18050 13804 18060 13860
rect 18116 13804 18956 13860
rect 19012 13804 19022 13860
rect 19282 13692 19292 13748
rect 19348 13692 19740 13748
rect 19796 13692 20300 13748
rect 20356 13692 22764 13748
rect 22820 13692 22830 13748
rect 19292 13580 19516 13636
rect 19572 13580 21196 13636
rect 21252 13580 21262 13636
rect 19292 13524 19348 13580
rect 16930 13468 16940 13524
rect 16996 13468 17892 13524
rect 19282 13468 19292 13524
rect 19348 13468 19358 13524
rect 20962 13468 20972 13524
rect 21028 13468 21038 13524
rect 23762 13468 23772 13524
rect 23828 13468 23996 13524
rect 24052 13468 24780 13524
rect 24836 13468 24846 13524
rect 61730 13468 61740 13524
rect 61796 13468 63308 13524
rect 63364 13468 63374 13524
rect 17836 13412 17892 13468
rect 20972 13412 21028 13468
rect 17826 13356 17836 13412
rect 17892 13356 17902 13412
rect 19394 13356 19404 13412
rect 19460 13356 20412 13412
rect 20468 13356 21868 13412
rect 21924 13356 21934 13412
rect 23364 13300 23374 13356
rect 23430 13300 23478 13356
rect 23534 13300 23582 13356
rect 23638 13300 23648 13356
rect 67688 13300 67698 13356
rect 67754 13300 67802 13356
rect 67858 13300 67906 13356
rect 67962 13300 67972 13356
rect 112012 13300 112022 13356
rect 112078 13300 112126 13356
rect 112182 13300 112230 13356
rect 112286 13300 112296 13356
rect 156336 13300 156346 13356
rect 156402 13300 156450 13356
rect 156506 13300 156554 13356
rect 156610 13300 156620 13356
rect 18946 13132 18956 13188
rect 19012 13132 19852 13188
rect 19908 13132 19918 13188
rect 21186 13132 21196 13188
rect 21252 13132 24556 13188
rect 24612 13132 26348 13188
rect 26404 13132 31052 13188
rect 31108 13132 31118 13188
rect 18722 13020 18732 13076
rect 18788 13020 19628 13076
rect 19684 13020 19964 13076
rect 20020 13020 20030 13076
rect 20514 13020 20524 13076
rect 20580 13020 20860 13076
rect 20916 13020 21308 13076
rect 21364 13020 21374 13076
rect 22978 13020 22988 13076
rect 23044 13020 23660 13076
rect 23716 13020 25004 13076
rect 25060 13020 25070 13076
rect 20178 12796 20188 12852
rect 20244 12796 20524 12852
rect 20580 12796 20860 12852
rect 20916 12796 20926 12852
rect 40226 12796 40236 12852
rect 40292 12796 40796 12852
rect 40852 12796 40862 12852
rect 19842 12684 19852 12740
rect 19908 12684 20636 12740
rect 20692 12684 20702 12740
rect 60610 12684 60620 12740
rect 60676 12684 62412 12740
rect 62468 12684 62478 12740
rect 45526 12516 45536 12572
rect 45592 12516 45640 12572
rect 45696 12516 45744 12572
rect 45800 12516 45810 12572
rect 89850 12516 89860 12572
rect 89916 12516 89964 12572
rect 90020 12516 90068 12572
rect 90124 12516 90134 12572
rect 134174 12516 134184 12572
rect 134240 12516 134288 12572
rect 134344 12516 134392 12572
rect 134448 12516 134458 12572
rect 178498 12516 178508 12572
rect 178564 12516 178612 12572
rect 178668 12516 178716 12572
rect 178772 12516 178782 12572
rect 26226 12348 26236 12404
rect 26292 12348 27132 12404
rect 27188 12348 27198 12404
rect 16930 12236 16940 12292
rect 16996 12236 17164 12292
rect 17220 12236 18508 12292
rect 18564 12236 18956 12292
rect 19012 12236 19292 12292
rect 19348 12236 19852 12292
rect 19908 12236 19918 12292
rect 20290 12236 20300 12292
rect 20356 12236 20972 12292
rect 21028 12236 21038 12292
rect 21858 12236 21868 12292
rect 21924 12236 22652 12292
rect 22708 12236 22718 12292
rect 40114 12236 40124 12292
rect 40180 12236 41580 12292
rect 41636 12236 41646 12292
rect 60274 12236 60284 12292
rect 60340 12236 61740 12292
rect 61796 12236 61806 12292
rect 20972 12180 21028 12236
rect 16594 12124 16604 12180
rect 16660 12124 17276 12180
rect 17332 12124 18172 12180
rect 18228 12124 18238 12180
rect 20972 12124 22092 12180
rect 22148 12124 22158 12180
rect 20850 12012 20860 12068
rect 20916 12012 21756 12068
rect 21812 12012 21822 12068
rect 23364 11732 23374 11788
rect 23430 11732 23478 11788
rect 23534 11732 23582 11788
rect 23638 11732 23648 11788
rect 67688 11732 67698 11788
rect 67754 11732 67802 11788
rect 67858 11732 67906 11788
rect 67962 11732 67972 11788
rect 112012 11732 112022 11788
rect 112078 11732 112126 11788
rect 112182 11732 112230 11788
rect 112286 11732 112296 11788
rect 156336 11732 156346 11788
rect 156402 11732 156450 11788
rect 156506 11732 156554 11788
rect 156610 11732 156620 11788
rect 52098 11676 52108 11732
rect 52164 11676 60228 11732
rect 60172 11620 60228 11676
rect 23874 11564 23884 11620
rect 23940 11564 25004 11620
rect 25060 11564 26460 11620
rect 26516 11564 26526 11620
rect 39330 11564 39340 11620
rect 39396 11564 39788 11620
rect 39844 11564 40012 11620
rect 40068 11564 40908 11620
rect 40964 11564 42140 11620
rect 42196 11564 43708 11620
rect 60162 11564 60172 11620
rect 60228 11564 60508 11620
rect 60564 11564 61404 11620
rect 61460 11564 61852 11620
rect 61908 11564 62972 11620
rect 63028 11564 63644 11620
rect 63700 11564 63710 11620
rect 17266 11452 17276 11508
rect 17332 11452 17836 11508
rect 17892 11452 18060 11508
rect 18116 11452 18508 11508
rect 18564 11452 18732 11508
rect 18788 11452 19628 11508
rect 19684 11452 20188 11508
rect 20132 11228 20188 11452
rect 25890 11340 25900 11396
rect 25956 11340 27692 11396
rect 27748 11340 27758 11396
rect 43652 11284 43708 11564
rect 51874 11340 51884 11396
rect 51940 11340 53452 11396
rect 53508 11340 53518 11396
rect 20244 11228 20254 11284
rect 39442 11228 39452 11284
rect 39508 11228 40684 11284
rect 40740 11228 40750 11284
rect 41458 11228 41468 11284
rect 41524 11228 42028 11284
rect 42084 11228 42094 11284
rect 43652 11228 52332 11284
rect 52388 11228 52668 11284
rect 52724 11228 52734 11284
rect 19842 11116 19852 11172
rect 19908 11116 20636 11172
rect 20692 11116 20972 11172
rect 21028 11116 21038 11172
rect 45526 10948 45536 11004
rect 45592 10948 45640 11004
rect 45696 10948 45744 11004
rect 45800 10948 45810 11004
rect 89850 10948 89860 11004
rect 89916 10948 89964 11004
rect 90020 10948 90068 11004
rect 90124 10948 90134 11004
rect 134174 10948 134184 11004
rect 134240 10948 134288 11004
rect 134344 10948 134392 11004
rect 134448 10948 134458 11004
rect 178498 10948 178508 11004
rect 178564 10948 178612 11004
rect 178668 10948 178716 11004
rect 178772 10948 178782 11004
rect 39778 10780 39788 10836
rect 39844 10780 40460 10836
rect 40516 10780 40526 10836
rect 39890 10668 39900 10724
rect 39956 10668 41580 10724
rect 41636 10668 41646 10724
rect 21858 10556 21868 10612
rect 21924 10556 22652 10612
rect 22708 10556 23436 10612
rect 23492 10556 24108 10612
rect 24164 10556 24556 10612
rect 24612 10556 24622 10612
rect 20178 10444 20188 10500
rect 20244 10444 20860 10500
rect 20916 10444 20926 10500
rect 40562 10332 40572 10388
rect 40628 10332 42700 10388
rect 42756 10332 42766 10388
rect 23364 10164 23374 10220
rect 23430 10164 23478 10220
rect 23534 10164 23582 10220
rect 23638 10164 23648 10220
rect 67688 10164 67698 10220
rect 67754 10164 67802 10220
rect 67858 10164 67906 10220
rect 67962 10164 67972 10220
rect 112012 10164 112022 10220
rect 112078 10164 112126 10220
rect 112182 10164 112230 10220
rect 112286 10164 112296 10220
rect 156336 10164 156346 10220
rect 156402 10164 156450 10220
rect 156506 10164 156554 10220
rect 156610 10164 156620 10220
rect 19954 9884 19964 9940
rect 20020 9884 21868 9940
rect 21924 9884 22764 9940
rect 22820 9884 23324 9940
rect 23380 9884 23772 9940
rect 23828 9884 23838 9940
rect 19506 9772 19516 9828
rect 19572 9772 20188 9828
rect 20244 9772 20524 9828
rect 20580 9772 20590 9828
rect 20962 9548 20972 9604
rect 21028 9548 21756 9604
rect 21812 9548 22652 9604
rect 22708 9548 22718 9604
rect 45526 9380 45536 9436
rect 45592 9380 45640 9436
rect 45696 9380 45744 9436
rect 45800 9380 45810 9436
rect 89850 9380 89860 9436
rect 89916 9380 89964 9436
rect 90020 9380 90068 9436
rect 90124 9380 90134 9436
rect 134174 9380 134184 9436
rect 134240 9380 134288 9436
rect 134344 9380 134392 9436
rect 134448 9380 134458 9436
rect 178498 9380 178508 9436
rect 178564 9380 178612 9436
rect 178668 9380 178716 9436
rect 178772 9380 178782 9436
rect 93874 9212 93884 9268
rect 93940 9212 94444 9268
rect 94500 9212 94510 9268
rect 20514 9100 20524 9156
rect 20580 9100 21308 9156
rect 21364 9100 21644 9156
rect 21700 9100 22204 9156
rect 22260 9100 22540 9156
rect 22596 9100 23100 9156
rect 23156 9100 24220 9156
rect 24276 9100 24286 9156
rect 89730 8988 89740 9044
rect 89796 8988 95340 9044
rect 95396 8988 95564 9044
rect 95620 8988 95630 9044
rect 23364 8596 23374 8652
rect 23430 8596 23478 8652
rect 23534 8596 23582 8652
rect 23638 8596 23648 8652
rect 67688 8596 67698 8652
rect 67754 8596 67802 8652
rect 67858 8596 67906 8652
rect 67962 8596 67972 8652
rect 112012 8596 112022 8652
rect 112078 8596 112126 8652
rect 112182 8596 112230 8652
rect 112286 8596 112296 8652
rect 156336 8596 156346 8652
rect 156402 8596 156450 8652
rect 156506 8596 156554 8652
rect 156610 8596 156620 8652
rect 45526 7812 45536 7868
rect 45592 7812 45640 7868
rect 45696 7812 45744 7868
rect 45800 7812 45810 7868
rect 89850 7812 89860 7868
rect 89916 7812 89964 7868
rect 90020 7812 90068 7868
rect 90124 7812 90134 7868
rect 134174 7812 134184 7868
rect 134240 7812 134288 7868
rect 134344 7812 134392 7868
rect 134448 7812 134458 7868
rect 178498 7812 178508 7868
rect 178564 7812 178612 7868
rect 178668 7812 178716 7868
rect 178772 7812 178782 7868
rect 23364 7028 23374 7084
rect 23430 7028 23478 7084
rect 23534 7028 23582 7084
rect 23638 7028 23648 7084
rect 67688 7028 67698 7084
rect 67754 7028 67802 7084
rect 67858 7028 67906 7084
rect 67962 7028 67972 7084
rect 112012 7028 112022 7084
rect 112078 7028 112126 7084
rect 112182 7028 112230 7084
rect 112286 7028 112296 7084
rect 156336 7028 156346 7084
rect 156402 7028 156450 7084
rect 156506 7028 156554 7084
rect 156610 7028 156620 7084
rect 45526 6244 45536 6300
rect 45592 6244 45640 6300
rect 45696 6244 45744 6300
rect 45800 6244 45810 6300
rect 89850 6244 89860 6300
rect 89916 6244 89964 6300
rect 90020 6244 90068 6300
rect 90124 6244 90134 6300
rect 134174 6244 134184 6300
rect 134240 6244 134288 6300
rect 134344 6244 134392 6300
rect 134448 6244 134458 6300
rect 178498 6244 178508 6300
rect 178564 6244 178612 6300
rect 178668 6244 178716 6300
rect 178772 6244 178782 6300
rect 23364 5460 23374 5516
rect 23430 5460 23478 5516
rect 23534 5460 23582 5516
rect 23638 5460 23648 5516
rect 67688 5460 67698 5516
rect 67754 5460 67802 5516
rect 67858 5460 67906 5516
rect 67962 5460 67972 5516
rect 112012 5460 112022 5516
rect 112078 5460 112126 5516
rect 112182 5460 112230 5516
rect 112286 5460 112296 5516
rect 156336 5460 156346 5516
rect 156402 5460 156450 5516
rect 156506 5460 156554 5516
rect 156610 5460 156620 5516
rect 45526 4676 45536 4732
rect 45592 4676 45640 4732
rect 45696 4676 45744 4732
rect 45800 4676 45810 4732
rect 89850 4676 89860 4732
rect 89916 4676 89964 4732
rect 90020 4676 90068 4732
rect 90124 4676 90134 4732
rect 134174 4676 134184 4732
rect 134240 4676 134288 4732
rect 134344 4676 134392 4732
rect 134448 4676 134458 4732
rect 178498 4676 178508 4732
rect 178564 4676 178612 4732
rect 178668 4676 178716 4732
rect 178772 4676 178782 4732
rect 94770 4284 94780 4340
rect 94836 4284 119644 4340
rect 119700 4284 119710 4340
rect 95890 4172 95900 4228
rect 95956 4172 121324 4228
rect 121380 4172 121390 4228
rect 23364 3892 23374 3948
rect 23430 3892 23478 3948
rect 23534 3892 23582 3948
rect 23638 3892 23648 3948
rect 67688 3892 67698 3948
rect 67754 3892 67802 3948
rect 67858 3892 67906 3948
rect 67962 3892 67972 3948
rect 112012 3892 112022 3948
rect 112078 3892 112126 3948
rect 112182 3892 112230 3948
rect 112286 3892 112296 3948
rect 156336 3892 156346 3948
rect 156402 3892 156450 3948
rect 156506 3892 156554 3948
rect 156610 3892 156620 3948
rect 12674 3276 12684 3332
rect 12740 3276 13580 3332
rect 13636 3276 13646 3332
rect 24434 3276 24444 3332
rect 24500 3276 25340 3332
rect 25396 3276 25406 3332
rect 36194 3276 36204 3332
rect 36260 3276 37100 3332
rect 37156 3276 37166 3332
rect 47954 3276 47964 3332
rect 48020 3276 48860 3332
rect 48916 3276 48926 3332
rect 59714 3276 59724 3332
rect 59780 3276 60620 3332
rect 60676 3276 60686 3332
rect 173954 3276 173964 3332
rect 174020 3276 174972 3332
rect 175028 3276 175038 3332
rect 45526 3108 45536 3164
rect 45592 3108 45640 3164
rect 45696 3108 45744 3164
rect 45800 3108 45810 3164
rect 89850 3108 89860 3164
rect 89916 3108 89964 3164
rect 90020 3108 90068 3164
rect 90124 3108 90134 3164
rect 134174 3108 134184 3164
rect 134240 3108 134288 3164
rect 134344 3108 134392 3164
rect 134448 3108 134458 3164
rect 178498 3108 178508 3164
rect 178564 3108 178612 3164
rect 178668 3108 178716 3164
rect 178772 3108 178782 3164
<< via3 >>
rect 23374 16436 23430 16492
rect 23478 16436 23534 16492
rect 23582 16436 23638 16492
rect 67698 16436 67754 16492
rect 67802 16436 67858 16492
rect 67906 16436 67962 16492
rect 112022 16436 112078 16492
rect 112126 16436 112182 16492
rect 112230 16436 112286 16492
rect 156346 16436 156402 16492
rect 156450 16436 156506 16492
rect 156554 16436 156610 16492
rect 45536 15652 45592 15708
rect 45640 15652 45696 15708
rect 45744 15652 45800 15708
rect 89860 15652 89916 15708
rect 89964 15652 90020 15708
rect 90068 15652 90124 15708
rect 134184 15652 134240 15708
rect 134288 15652 134344 15708
rect 134392 15652 134448 15708
rect 178508 15652 178564 15708
rect 178612 15652 178668 15708
rect 178716 15652 178772 15708
rect 23374 14868 23430 14924
rect 23478 14868 23534 14924
rect 23582 14868 23638 14924
rect 67698 14868 67754 14924
rect 67802 14868 67858 14924
rect 67906 14868 67962 14924
rect 112022 14868 112078 14924
rect 112126 14868 112182 14924
rect 112230 14868 112286 14924
rect 156346 14868 156402 14924
rect 156450 14868 156506 14924
rect 156554 14868 156610 14924
rect 45536 14084 45592 14140
rect 45640 14084 45696 14140
rect 45744 14084 45800 14140
rect 89860 14084 89916 14140
rect 89964 14084 90020 14140
rect 90068 14084 90124 14140
rect 134184 14084 134240 14140
rect 134288 14084 134344 14140
rect 134392 14084 134448 14140
rect 178508 14084 178564 14140
rect 178612 14084 178668 14140
rect 178716 14084 178772 14140
rect 23374 13300 23430 13356
rect 23478 13300 23534 13356
rect 23582 13300 23638 13356
rect 67698 13300 67754 13356
rect 67802 13300 67858 13356
rect 67906 13300 67962 13356
rect 112022 13300 112078 13356
rect 112126 13300 112182 13356
rect 112230 13300 112286 13356
rect 156346 13300 156402 13356
rect 156450 13300 156506 13356
rect 156554 13300 156610 13356
rect 45536 12516 45592 12572
rect 45640 12516 45696 12572
rect 45744 12516 45800 12572
rect 89860 12516 89916 12572
rect 89964 12516 90020 12572
rect 90068 12516 90124 12572
rect 134184 12516 134240 12572
rect 134288 12516 134344 12572
rect 134392 12516 134448 12572
rect 178508 12516 178564 12572
rect 178612 12516 178668 12572
rect 178716 12516 178772 12572
rect 23374 11732 23430 11788
rect 23478 11732 23534 11788
rect 23582 11732 23638 11788
rect 67698 11732 67754 11788
rect 67802 11732 67858 11788
rect 67906 11732 67962 11788
rect 112022 11732 112078 11788
rect 112126 11732 112182 11788
rect 112230 11732 112286 11788
rect 156346 11732 156402 11788
rect 156450 11732 156506 11788
rect 156554 11732 156610 11788
rect 45536 10948 45592 11004
rect 45640 10948 45696 11004
rect 45744 10948 45800 11004
rect 89860 10948 89916 11004
rect 89964 10948 90020 11004
rect 90068 10948 90124 11004
rect 134184 10948 134240 11004
rect 134288 10948 134344 11004
rect 134392 10948 134448 11004
rect 178508 10948 178564 11004
rect 178612 10948 178668 11004
rect 178716 10948 178772 11004
rect 23374 10164 23430 10220
rect 23478 10164 23534 10220
rect 23582 10164 23638 10220
rect 67698 10164 67754 10220
rect 67802 10164 67858 10220
rect 67906 10164 67962 10220
rect 112022 10164 112078 10220
rect 112126 10164 112182 10220
rect 112230 10164 112286 10220
rect 156346 10164 156402 10220
rect 156450 10164 156506 10220
rect 156554 10164 156610 10220
rect 45536 9380 45592 9436
rect 45640 9380 45696 9436
rect 45744 9380 45800 9436
rect 89860 9380 89916 9436
rect 89964 9380 90020 9436
rect 90068 9380 90124 9436
rect 134184 9380 134240 9436
rect 134288 9380 134344 9436
rect 134392 9380 134448 9436
rect 178508 9380 178564 9436
rect 178612 9380 178668 9436
rect 178716 9380 178772 9436
rect 23374 8596 23430 8652
rect 23478 8596 23534 8652
rect 23582 8596 23638 8652
rect 67698 8596 67754 8652
rect 67802 8596 67858 8652
rect 67906 8596 67962 8652
rect 112022 8596 112078 8652
rect 112126 8596 112182 8652
rect 112230 8596 112286 8652
rect 156346 8596 156402 8652
rect 156450 8596 156506 8652
rect 156554 8596 156610 8652
rect 45536 7812 45592 7868
rect 45640 7812 45696 7868
rect 45744 7812 45800 7868
rect 89860 7812 89916 7868
rect 89964 7812 90020 7868
rect 90068 7812 90124 7868
rect 134184 7812 134240 7868
rect 134288 7812 134344 7868
rect 134392 7812 134448 7868
rect 178508 7812 178564 7868
rect 178612 7812 178668 7868
rect 178716 7812 178772 7868
rect 23374 7028 23430 7084
rect 23478 7028 23534 7084
rect 23582 7028 23638 7084
rect 67698 7028 67754 7084
rect 67802 7028 67858 7084
rect 67906 7028 67962 7084
rect 112022 7028 112078 7084
rect 112126 7028 112182 7084
rect 112230 7028 112286 7084
rect 156346 7028 156402 7084
rect 156450 7028 156506 7084
rect 156554 7028 156610 7084
rect 45536 6244 45592 6300
rect 45640 6244 45696 6300
rect 45744 6244 45800 6300
rect 89860 6244 89916 6300
rect 89964 6244 90020 6300
rect 90068 6244 90124 6300
rect 134184 6244 134240 6300
rect 134288 6244 134344 6300
rect 134392 6244 134448 6300
rect 178508 6244 178564 6300
rect 178612 6244 178668 6300
rect 178716 6244 178772 6300
rect 23374 5460 23430 5516
rect 23478 5460 23534 5516
rect 23582 5460 23638 5516
rect 67698 5460 67754 5516
rect 67802 5460 67858 5516
rect 67906 5460 67962 5516
rect 112022 5460 112078 5516
rect 112126 5460 112182 5516
rect 112230 5460 112286 5516
rect 156346 5460 156402 5516
rect 156450 5460 156506 5516
rect 156554 5460 156610 5516
rect 45536 4676 45592 4732
rect 45640 4676 45696 4732
rect 45744 4676 45800 4732
rect 89860 4676 89916 4732
rect 89964 4676 90020 4732
rect 90068 4676 90124 4732
rect 134184 4676 134240 4732
rect 134288 4676 134344 4732
rect 134392 4676 134448 4732
rect 178508 4676 178564 4732
rect 178612 4676 178668 4732
rect 178716 4676 178772 4732
rect 23374 3892 23430 3948
rect 23478 3892 23534 3948
rect 23582 3892 23638 3948
rect 67698 3892 67754 3948
rect 67802 3892 67858 3948
rect 67906 3892 67962 3948
rect 112022 3892 112078 3948
rect 112126 3892 112182 3948
rect 112230 3892 112286 3948
rect 156346 3892 156402 3948
rect 156450 3892 156506 3948
rect 156554 3892 156610 3948
rect 45536 3108 45592 3164
rect 45640 3108 45696 3164
rect 45744 3108 45800 3164
rect 89860 3108 89916 3164
rect 89964 3108 90020 3164
rect 90068 3108 90124 3164
rect 134184 3108 134240 3164
rect 134288 3108 134344 3164
rect 134392 3108 134448 3164
rect 178508 3108 178564 3164
rect 178612 3108 178668 3164
rect 178716 3108 178772 3164
<< metal4 >>
rect 23346 16492 23666 16524
rect 23346 16436 23374 16492
rect 23430 16436 23478 16492
rect 23534 16436 23582 16492
rect 23638 16436 23666 16492
rect 23346 14924 23666 16436
rect 23346 14868 23374 14924
rect 23430 14868 23478 14924
rect 23534 14868 23582 14924
rect 23638 14868 23666 14924
rect 23346 13356 23666 14868
rect 23346 13300 23374 13356
rect 23430 13300 23478 13356
rect 23534 13300 23582 13356
rect 23638 13300 23666 13356
rect 23346 11788 23666 13300
rect 23346 11732 23374 11788
rect 23430 11732 23478 11788
rect 23534 11732 23582 11788
rect 23638 11732 23666 11788
rect 23346 10220 23666 11732
rect 23346 10164 23374 10220
rect 23430 10164 23478 10220
rect 23534 10164 23582 10220
rect 23638 10164 23666 10220
rect 23346 8652 23666 10164
rect 23346 8596 23374 8652
rect 23430 8596 23478 8652
rect 23534 8596 23582 8652
rect 23638 8596 23666 8652
rect 23346 7084 23666 8596
rect 23346 7028 23374 7084
rect 23430 7028 23478 7084
rect 23534 7028 23582 7084
rect 23638 7028 23666 7084
rect 23346 5516 23666 7028
rect 23346 5460 23374 5516
rect 23430 5460 23478 5516
rect 23534 5460 23582 5516
rect 23638 5460 23666 5516
rect 23346 3948 23666 5460
rect 23346 3892 23374 3948
rect 23430 3892 23478 3948
rect 23534 3892 23582 3948
rect 23638 3892 23666 3948
rect 23346 3076 23666 3892
rect 45508 15708 45828 16524
rect 45508 15652 45536 15708
rect 45592 15652 45640 15708
rect 45696 15652 45744 15708
rect 45800 15652 45828 15708
rect 45508 14140 45828 15652
rect 45508 14084 45536 14140
rect 45592 14084 45640 14140
rect 45696 14084 45744 14140
rect 45800 14084 45828 14140
rect 45508 12572 45828 14084
rect 45508 12516 45536 12572
rect 45592 12516 45640 12572
rect 45696 12516 45744 12572
rect 45800 12516 45828 12572
rect 45508 11004 45828 12516
rect 45508 10948 45536 11004
rect 45592 10948 45640 11004
rect 45696 10948 45744 11004
rect 45800 10948 45828 11004
rect 45508 9436 45828 10948
rect 45508 9380 45536 9436
rect 45592 9380 45640 9436
rect 45696 9380 45744 9436
rect 45800 9380 45828 9436
rect 45508 7868 45828 9380
rect 45508 7812 45536 7868
rect 45592 7812 45640 7868
rect 45696 7812 45744 7868
rect 45800 7812 45828 7868
rect 45508 6300 45828 7812
rect 45508 6244 45536 6300
rect 45592 6244 45640 6300
rect 45696 6244 45744 6300
rect 45800 6244 45828 6300
rect 45508 4732 45828 6244
rect 45508 4676 45536 4732
rect 45592 4676 45640 4732
rect 45696 4676 45744 4732
rect 45800 4676 45828 4732
rect 45508 3164 45828 4676
rect 45508 3108 45536 3164
rect 45592 3108 45640 3164
rect 45696 3108 45744 3164
rect 45800 3108 45828 3164
rect 45508 3076 45828 3108
rect 67670 16492 67990 16524
rect 67670 16436 67698 16492
rect 67754 16436 67802 16492
rect 67858 16436 67906 16492
rect 67962 16436 67990 16492
rect 67670 14924 67990 16436
rect 67670 14868 67698 14924
rect 67754 14868 67802 14924
rect 67858 14868 67906 14924
rect 67962 14868 67990 14924
rect 67670 13356 67990 14868
rect 67670 13300 67698 13356
rect 67754 13300 67802 13356
rect 67858 13300 67906 13356
rect 67962 13300 67990 13356
rect 67670 11788 67990 13300
rect 67670 11732 67698 11788
rect 67754 11732 67802 11788
rect 67858 11732 67906 11788
rect 67962 11732 67990 11788
rect 67670 10220 67990 11732
rect 67670 10164 67698 10220
rect 67754 10164 67802 10220
rect 67858 10164 67906 10220
rect 67962 10164 67990 10220
rect 67670 8652 67990 10164
rect 67670 8596 67698 8652
rect 67754 8596 67802 8652
rect 67858 8596 67906 8652
rect 67962 8596 67990 8652
rect 67670 7084 67990 8596
rect 67670 7028 67698 7084
rect 67754 7028 67802 7084
rect 67858 7028 67906 7084
rect 67962 7028 67990 7084
rect 67670 5516 67990 7028
rect 67670 5460 67698 5516
rect 67754 5460 67802 5516
rect 67858 5460 67906 5516
rect 67962 5460 67990 5516
rect 67670 3948 67990 5460
rect 67670 3892 67698 3948
rect 67754 3892 67802 3948
rect 67858 3892 67906 3948
rect 67962 3892 67990 3948
rect 67670 3076 67990 3892
rect 89832 15708 90152 16524
rect 89832 15652 89860 15708
rect 89916 15652 89964 15708
rect 90020 15652 90068 15708
rect 90124 15652 90152 15708
rect 89832 14140 90152 15652
rect 89832 14084 89860 14140
rect 89916 14084 89964 14140
rect 90020 14084 90068 14140
rect 90124 14084 90152 14140
rect 89832 12572 90152 14084
rect 89832 12516 89860 12572
rect 89916 12516 89964 12572
rect 90020 12516 90068 12572
rect 90124 12516 90152 12572
rect 89832 11004 90152 12516
rect 89832 10948 89860 11004
rect 89916 10948 89964 11004
rect 90020 10948 90068 11004
rect 90124 10948 90152 11004
rect 89832 9436 90152 10948
rect 89832 9380 89860 9436
rect 89916 9380 89964 9436
rect 90020 9380 90068 9436
rect 90124 9380 90152 9436
rect 89832 7868 90152 9380
rect 89832 7812 89860 7868
rect 89916 7812 89964 7868
rect 90020 7812 90068 7868
rect 90124 7812 90152 7868
rect 89832 6300 90152 7812
rect 89832 6244 89860 6300
rect 89916 6244 89964 6300
rect 90020 6244 90068 6300
rect 90124 6244 90152 6300
rect 89832 4732 90152 6244
rect 89832 4676 89860 4732
rect 89916 4676 89964 4732
rect 90020 4676 90068 4732
rect 90124 4676 90152 4732
rect 89832 3164 90152 4676
rect 89832 3108 89860 3164
rect 89916 3108 89964 3164
rect 90020 3108 90068 3164
rect 90124 3108 90152 3164
rect 89832 3076 90152 3108
rect 111994 16492 112314 16524
rect 111994 16436 112022 16492
rect 112078 16436 112126 16492
rect 112182 16436 112230 16492
rect 112286 16436 112314 16492
rect 111994 14924 112314 16436
rect 111994 14868 112022 14924
rect 112078 14868 112126 14924
rect 112182 14868 112230 14924
rect 112286 14868 112314 14924
rect 111994 13356 112314 14868
rect 111994 13300 112022 13356
rect 112078 13300 112126 13356
rect 112182 13300 112230 13356
rect 112286 13300 112314 13356
rect 111994 11788 112314 13300
rect 111994 11732 112022 11788
rect 112078 11732 112126 11788
rect 112182 11732 112230 11788
rect 112286 11732 112314 11788
rect 111994 10220 112314 11732
rect 111994 10164 112022 10220
rect 112078 10164 112126 10220
rect 112182 10164 112230 10220
rect 112286 10164 112314 10220
rect 111994 8652 112314 10164
rect 111994 8596 112022 8652
rect 112078 8596 112126 8652
rect 112182 8596 112230 8652
rect 112286 8596 112314 8652
rect 111994 7084 112314 8596
rect 111994 7028 112022 7084
rect 112078 7028 112126 7084
rect 112182 7028 112230 7084
rect 112286 7028 112314 7084
rect 111994 5516 112314 7028
rect 111994 5460 112022 5516
rect 112078 5460 112126 5516
rect 112182 5460 112230 5516
rect 112286 5460 112314 5516
rect 111994 3948 112314 5460
rect 111994 3892 112022 3948
rect 112078 3892 112126 3948
rect 112182 3892 112230 3948
rect 112286 3892 112314 3948
rect 111994 3076 112314 3892
rect 134156 15708 134476 16524
rect 134156 15652 134184 15708
rect 134240 15652 134288 15708
rect 134344 15652 134392 15708
rect 134448 15652 134476 15708
rect 134156 14140 134476 15652
rect 134156 14084 134184 14140
rect 134240 14084 134288 14140
rect 134344 14084 134392 14140
rect 134448 14084 134476 14140
rect 134156 12572 134476 14084
rect 134156 12516 134184 12572
rect 134240 12516 134288 12572
rect 134344 12516 134392 12572
rect 134448 12516 134476 12572
rect 134156 11004 134476 12516
rect 134156 10948 134184 11004
rect 134240 10948 134288 11004
rect 134344 10948 134392 11004
rect 134448 10948 134476 11004
rect 134156 9436 134476 10948
rect 134156 9380 134184 9436
rect 134240 9380 134288 9436
rect 134344 9380 134392 9436
rect 134448 9380 134476 9436
rect 134156 7868 134476 9380
rect 134156 7812 134184 7868
rect 134240 7812 134288 7868
rect 134344 7812 134392 7868
rect 134448 7812 134476 7868
rect 134156 6300 134476 7812
rect 134156 6244 134184 6300
rect 134240 6244 134288 6300
rect 134344 6244 134392 6300
rect 134448 6244 134476 6300
rect 134156 4732 134476 6244
rect 134156 4676 134184 4732
rect 134240 4676 134288 4732
rect 134344 4676 134392 4732
rect 134448 4676 134476 4732
rect 134156 3164 134476 4676
rect 134156 3108 134184 3164
rect 134240 3108 134288 3164
rect 134344 3108 134392 3164
rect 134448 3108 134476 3164
rect 134156 3076 134476 3108
rect 156318 16492 156638 16524
rect 156318 16436 156346 16492
rect 156402 16436 156450 16492
rect 156506 16436 156554 16492
rect 156610 16436 156638 16492
rect 156318 14924 156638 16436
rect 156318 14868 156346 14924
rect 156402 14868 156450 14924
rect 156506 14868 156554 14924
rect 156610 14868 156638 14924
rect 156318 13356 156638 14868
rect 156318 13300 156346 13356
rect 156402 13300 156450 13356
rect 156506 13300 156554 13356
rect 156610 13300 156638 13356
rect 156318 11788 156638 13300
rect 156318 11732 156346 11788
rect 156402 11732 156450 11788
rect 156506 11732 156554 11788
rect 156610 11732 156638 11788
rect 156318 10220 156638 11732
rect 156318 10164 156346 10220
rect 156402 10164 156450 10220
rect 156506 10164 156554 10220
rect 156610 10164 156638 10220
rect 156318 8652 156638 10164
rect 156318 8596 156346 8652
rect 156402 8596 156450 8652
rect 156506 8596 156554 8652
rect 156610 8596 156638 8652
rect 156318 7084 156638 8596
rect 156318 7028 156346 7084
rect 156402 7028 156450 7084
rect 156506 7028 156554 7084
rect 156610 7028 156638 7084
rect 156318 5516 156638 7028
rect 156318 5460 156346 5516
rect 156402 5460 156450 5516
rect 156506 5460 156554 5516
rect 156610 5460 156638 5516
rect 156318 3948 156638 5460
rect 156318 3892 156346 3948
rect 156402 3892 156450 3948
rect 156506 3892 156554 3948
rect 156610 3892 156638 3948
rect 156318 3076 156638 3892
rect 178480 15708 178800 16524
rect 178480 15652 178508 15708
rect 178564 15652 178612 15708
rect 178668 15652 178716 15708
rect 178772 15652 178800 15708
rect 178480 14140 178800 15652
rect 178480 14084 178508 14140
rect 178564 14084 178612 14140
rect 178668 14084 178716 14140
rect 178772 14084 178800 14140
rect 178480 12572 178800 14084
rect 178480 12516 178508 12572
rect 178564 12516 178612 12572
rect 178668 12516 178716 12572
rect 178772 12516 178800 12572
rect 178480 11004 178800 12516
rect 178480 10948 178508 11004
rect 178564 10948 178612 11004
rect 178668 10948 178716 11004
rect 178772 10948 178800 11004
rect 178480 9436 178800 10948
rect 178480 9380 178508 9436
rect 178564 9380 178612 9436
rect 178668 9380 178716 9436
rect 178772 9380 178800 9436
rect 178480 7868 178800 9380
rect 178480 7812 178508 7868
rect 178564 7812 178612 7868
rect 178668 7812 178716 7868
rect 178772 7812 178800 7868
rect 178480 6300 178800 7812
rect 178480 6244 178508 6300
rect 178564 6244 178612 6300
rect 178668 6244 178716 6300
rect 178772 6244 178800 6300
rect 178480 4732 178800 6244
rect 178480 4676 178508 4732
rect 178564 4676 178612 4732
rect 178668 4676 178716 4732
rect 178772 4676 178800 4732
rect 178480 3164 178800 4676
rect 178480 3108 178508 3164
rect 178564 3108 178612 3164
rect 178668 3108 178716 3164
rect 178772 3108 178800 3164
rect 178480 3076 178800 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__030__I pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__A1
timestamp 1667941163
transform 1 0 25536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__CLK
timestamp 1667941163
transform 1 0 13440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__CLK
timestamp 1667941163
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__CLK
timestamp 1667941163
transform -1 0 30128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__D
timestamp 1667941163
transform 1 0 26208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__CLK
timestamp 1667941163
transform 1 0 37408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__D
timestamp 1667941163
transform -1 0 33264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__CLK
timestamp 1667941163
transform 1 0 48496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__D
timestamp 1667941163
transform -1 0 48272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__CLK
timestamp 1667941163
transform 1 0 60032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__D
timestamp 1667941163
transform -1 0 60704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__CLK
timestamp 1667941163
transform 1 0 76496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__D
timestamp 1667941163
transform 1 0 76944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__CLK
timestamp 1667941163
transform 1 0 91168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__D
timestamp 1667941163
transform -1 0 91840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__I
timestamp 1667941163
transform 1 0 93856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I
timestamp 1667941163
transform -1 0 95424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout13_I
timestamp 1667941163
transform 1 0 19488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1667941163
transform -1 0 1904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1667941163
transform -1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1667941163
transform 1 0 10976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1667941163
transform -1 0 15344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1667941163
transform 1 0 20160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1667941163
transform -1 0 24752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1667941163
transform -1 0 31248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1667941163
transform -1 0 37184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1667941163
transform -1 0 38864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1667941163
transform 1 0 44128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[0\].pun_I
timestamp 1667941163
transform 1 0 23296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[0\].pup_I
timestamp 1667941163
transform 1 0 23072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[1\].pun_I
timestamp 1667941163
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[1\].pup_I
timestamp 1667941163
transform 1 0 18480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[2\].pun_I
timestamp 1667941163
transform -1 0 17808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[2\].pup_I
timestamp 1667941163
transform 1 0 24192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[3\].pun_I
timestamp 1667941163
transform 1 0 24304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[4\].pun_I
timestamp 1667941163
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[4\].pup_I
timestamp 1667941163
transform -1 0 21728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[5\].pun_I
timestamp 1667941163
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[5\].pup_I
timestamp 1667941163
transform -1 0 22624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[6\].pun_I
timestamp 1667941163
transform 1 0 23744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[6\].pup_I
timestamp 1667941163
transform -1 0 16240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[7\].pup_I
timestamp 1667941163
transform 1 0 24752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[8\].pup_I
timestamp 1667941163
transform 1 0 19488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[10\].pun_I
timestamp 1667941163
transform -1 0 23632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[10\].pup_I
timestamp 1667941163
transform -1 0 20832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[11\].pun_I
timestamp 1667941163
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[12\].pun_I
timestamp 1667941163
transform 1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[12\].pup_I
timestamp 1667941163
transform -1 0 22176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[13\].pun_I
timestamp 1667941163
transform 1 0 23968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[13\].pup_I
timestamp 1667941163
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[14\].pun_I
timestamp 1667941163
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[14\].pup_I
timestamp 1667941163
transform 1 0 20384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[15\].pun_I
timestamp 1667941163
transform 1 0 23408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[15\].pup_I
timestamp 1667941163
transform 1 0 17248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[16\].pun_I
timestamp 1667941163
transform 1 0 24080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[16\].pup_I
timestamp 1667941163
transform 1 0 20272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[17\].pun_I
timestamp 1667941163
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[17\].pup_I
timestamp 1667941163
transform 1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[18\].pun_I
timestamp 1667941163
transform -1 0 22848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[18\].pup_I
timestamp 1667941163
transform 1 0 18032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[0\].ptrimn_I
timestamp 1667941163
transform 1 0 19712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[0\].ptrimp_I
timestamp 1667941163
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[1\].ptrimn_I
timestamp 1667941163
transform -1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[1\].ptrimp_I
timestamp 1667941163
transform 1 0 16912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[2\].ptrimn_I
timestamp 1667941163
transform 1 0 27664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[2\].ptrimp_I
timestamp 1667941163
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ptrimn_I
timestamp 1667941163
transform 1 0 33712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ptrimp_I
timestamp 1667941163
transform 1 0 33712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 6384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 6832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51
timestamp 1667941163
transform 1 0 7056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56
timestamp 1667941163
transform 1 0 7616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64
timestamp 1667941163
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1667941163
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1667941163
transform 1 0 9408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80
timestamp 1667941163
transform 1 0 10304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 10976 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102
timestamp 1667941163
transform 1 0 12768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1667941163
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112
timestamp 1667941163
transform 1 0 13888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120
timestamp 1667941163
transform 1 0 14784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_126
timestamp 1667941163
transform 1 0 15456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134
timestamp 1667941163
transform 1 0 16352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 16800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1667941163
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_147
timestamp 1667941163
transform 1 0 17808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155
timestamp 1667941163
transform 1 0 18704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159
timestamp 1667941163
transform 1 0 19152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_161
timestamp 1667941163
transform 1 0 19376 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_166
timestamp 1667941163
transform 1 0 19936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_182
timestamp 1667941163
transform 1 0 21728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190
timestamp 1667941163
transform 1 0 22624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_196
timestamp 1667941163
transform 1 0 23296 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_204
timestamp 1667941163
transform 1 0 24192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_208
timestamp 1667941163
transform 1 0 24640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1667941163
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_217
timestamp 1667941163
transform 1 0 25648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_221
timestamp 1667941163
transform 1 0 26096 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_226
timestamp 1667941163
transform 1 0 26656 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_234
timestamp 1667941163
transform 1 0 27552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_236
timestamp 1667941163
transform 1 0 27776 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_241
timestamp 1667941163
transform 1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 29008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 29456 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_256
timestamp 1667941163
transform 1 0 30016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_264
timestamp 1667941163
transform 1 0 30912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_266
timestamp 1667941163
transform 1 0 31136 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_271
timestamp 1667941163
transform 1 0 31696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1667941163
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_287
timestamp 1667941163
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_295
timestamp 1667941163
transform 1 0 34384 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_301
timestamp 1667941163
transform 1 0 35056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_309
timestamp 1667941163
transform 1 0 35952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1667941163
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1667941163
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_322
timestamp 1667941163
transform 1 0 37408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_326
timestamp 1667941163
transform 1 0 37856 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_331
timestamp 1667941163
transform 1 0 38416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_339
timestamp 1667941163
transform 1 0 39312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_341
timestamp 1667941163
transform 1 0 39536 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_346
timestamp 1667941163
transform 1 0 40096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1667941163
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_356
timestamp 1667941163
transform 1 0 41216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_361
timestamp 1667941163
transform 1 0 41776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_369
timestamp 1667941163
transform 1 0 42672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_371
timestamp 1667941163
transform 1 0 42896 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_376
timestamp 1667941163
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1667941163
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1667941163
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_392
timestamp 1667941163
transform 1 0 45248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_400
timestamp 1667941163
transform 1 0 46144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_406
timestamp 1667941163
transform 1 0 46816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_414
timestamp 1667941163
transform 1 0 47712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1667941163
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1667941163
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_427
timestamp 1667941163
transform 1 0 49168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_431
timestamp 1667941163
transform 1 0 49616 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_436
timestamp 1667941163
transform 1 0 50176 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_444
timestamp 1667941163
transform 1 0 51072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_446
timestamp 1667941163
transform 1 0 51296 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_451
timestamp 1667941163
transform 1 0 51856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_457
timestamp 1667941163
transform 1 0 52528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_461
timestamp 1667941163
transform 1 0 52976 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_466
timestamp 1667941163
transform 1 0 53536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_474
timestamp 1667941163
transform 1 0 54432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_476
timestamp 1667941163
transform 1 0 54656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_481
timestamp 1667941163
transform 1 0 55216 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1667941163
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1667941163
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_497
timestamp 1667941163
transform 1 0 57008 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_505
timestamp 1667941163
transform 1 0 57904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_511
timestamp 1667941163
transform 1 0 58576 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_519
timestamp 1667941163
transform 1 0 59472 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_523
timestamp 1667941163
transform 1 0 59920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1667941163
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_532
timestamp 1667941163
transform 1 0 60928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_536
timestamp 1667941163
transform 1 0 61376 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_541
timestamp 1667941163
transform 1 0 61936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_549
timestamp 1667941163
transform 1 0 62832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_551
timestamp 1667941163
transform 1 0 63056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_556
timestamp 1667941163
transform 1 0 63616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_562
timestamp 1667941163
transform 1 0 64288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_566
timestamp 1667941163
transform 1 0 64736 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_571
timestamp 1667941163
transform 1 0 65296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_575
timestamp 1667941163
transform 1 0 65744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_581
timestamp 1667941163
transform 1 0 66416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_589
timestamp 1667941163
transform 1 0 67312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_593
timestamp 1667941163
transform 1 0 67760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1667941163
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_602
timestamp 1667941163
transform 1 0 68768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_606
timestamp 1667941163
transform 1 0 69216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_611
timestamp 1667941163
transform 1 0 69776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_619
timestamp 1667941163
transform 1 0 70672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_621
timestamp 1667941163
transform 1 0 70896 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_626
timestamp 1667941163
transform 1 0 71456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_632
timestamp 1667941163
transform 1 0 72128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_636
timestamp 1667941163
transform 1 0 72576 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_641
timestamp 1667941163
transform 1 0 73136 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_649
timestamp 1667941163
transform 1 0 74032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_651
timestamp 1667941163
transform 1 0 74256 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_656
timestamp 1667941163
transform 1 0 74816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1667941163
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1667941163
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_672
timestamp 1667941163
transform 1 0 76608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_680
timestamp 1667941163
transform 1 0 77504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_686
timestamp 1667941163
transform 1 0 78176 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_694
timestamp 1667941163
transform 1 0 79072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_698
timestamp 1667941163
transform 1 0 79520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1667941163
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_707
timestamp 1667941163
transform 1 0 80528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_711
timestamp 1667941163
transform 1 0 80976 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_716
timestamp 1667941163
transform 1 0 81536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_724
timestamp 1667941163
transform 1 0 82432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_726
timestamp 1667941163
transform 1 0 82656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_731
timestamp 1667941163
transform 1 0 83216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_737
timestamp 1667941163
transform 1 0 83888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_741
timestamp 1667941163
transform 1 0 84336 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_746
timestamp 1667941163
transform 1 0 84896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_754
timestamp 1667941163
transform 1 0 85792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_756
timestamp 1667941163
transform 1 0 86016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_761
timestamp 1667941163
transform 1 0 86576 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_769
timestamp 1667941163
transform 1 0 87472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1667941163
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_777
timestamp 1667941163
transform 1 0 88368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_785
timestamp 1667941163
transform 1 0 89264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_791
timestamp 1667941163
transform 1 0 89936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_799
timestamp 1667941163
transform 1 0 90832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_803
timestamp 1667941163
transform 1 0 91280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1667941163
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_812
timestamp 1667941163
transform 1 0 92288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_816
timestamp 1667941163
transform 1 0 92736 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_821
timestamp 1667941163
transform 1 0 93296 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_829
timestamp 1667941163
transform 1 0 94192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_831
timestamp 1667941163
transform 1 0 94416 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_836
timestamp 1667941163
transform 1 0 94976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_842
timestamp 1667941163
transform 1 0 95648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_846
timestamp 1667941163
transform 1 0 96096 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_851
timestamp 1667941163
transform 1 0 96656 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_859
timestamp 1667941163
transform 1 0 97552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_861
timestamp 1667941163
transform 1 0 97776 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_866
timestamp 1667941163
transform 1 0 98336 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1667941163
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1667941163
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_882
timestamp 1667941163
transform 1 0 100128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_890
timestamp 1667941163
transform 1 0 101024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_896
timestamp 1667941163
transform 1 0 101696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_904
timestamp 1667941163
transform 1 0 102592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_908
timestamp 1667941163
transform 1 0 103040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_912
timestamp 1667941163
transform 1 0 103488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_917
timestamp 1667941163
transform 1 0 104048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_921
timestamp 1667941163
transform 1 0 104496 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_926
timestamp 1667941163
transform 1 0 105056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_934
timestamp 1667941163
transform 1 0 105952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_936
timestamp 1667941163
transform 1 0 106176 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_941
timestamp 1667941163
transform 1 0 106736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_947
timestamp 1667941163
transform 1 0 107408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_951
timestamp 1667941163
transform 1 0 107856 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_956
timestamp 1667941163
transform 1 0 108416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_964
timestamp 1667941163
transform 1 0 109312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_966
timestamp 1667941163
transform 1 0 109536 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_971
timestamp 1667941163
transform 1 0 110096 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1667941163
transform 1 0 110992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1667941163
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_987
timestamp 1667941163
transform 1 0 111888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_995
timestamp 1667941163
transform 1 0 112784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1001
timestamp 1667941163
transform 1 0 113456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1009
timestamp 1667941163
transform 1 0 114352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1013
timestamp 1667941163
transform 1 0 114800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1667941163
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1022
timestamp 1667941163
transform 1 0 115808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1026
timestamp 1667941163
transform 1 0 116256 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1031
timestamp 1667941163
transform 1 0 116816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1039
timestamp 1667941163
transform 1 0 117712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1041
timestamp 1667941163
transform 1 0 117936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1046
timestamp 1667941163
transform 1 0 118496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1052
timestamp 1667941163
transform 1 0 119168 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1667941163
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1667941163
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1092
timestamp 1667941163
transform 1 0 123648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1100
timestamp 1667941163
transform 1 0 124544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1106
timestamp 1667941163
transform 1 0 125216 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1114
timestamp 1667941163
transform 1 0 126112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1118
timestamp 1667941163
transform 1 0 126560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1667941163
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1127
timestamp 1667941163
transform 1 0 127568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1131
timestamp 1667941163
transform 1 0 128016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1136
timestamp 1667941163
transform 1 0 128576 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1144
timestamp 1667941163
transform 1 0 129472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1146
timestamp 1667941163
transform 1 0 129696 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1151
timestamp 1667941163
transform 1 0 130256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1157
timestamp 1667941163
transform 1 0 130928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1161
timestamp 1667941163
transform 1 0 131376 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1166
timestamp 1667941163
transform 1 0 131936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1174
timestamp 1667941163
transform 1 0 132832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1176
timestamp 1667941163
transform 1 0 133056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1181
timestamp 1667941163
transform 1 0 133616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1189
timestamp 1667941163
transform 1 0 134512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1192
timestamp 1667941163
transform 1 0 134848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1197
timestamp 1667941163
transform 1 0 135408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1205
timestamp 1667941163
transform 1 0 136304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1211
timestamp 1667941163
transform 1 0 136976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1219
timestamp 1667941163
transform 1 0 137872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1223
timestamp 1667941163
transform 1 0 138320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1667941163
transform 1 0 138768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1232
timestamp 1667941163
transform 1 0 139328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1236
timestamp 1667941163
transform 1 0 139776 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1241
timestamp 1667941163
transform 1 0 140336 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1249
timestamp 1667941163
transform 1 0 141232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1251
timestamp 1667941163
transform 1 0 141456 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1256
timestamp 1667941163
transform 1 0 142016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1262
timestamp 1667941163
transform 1 0 142688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1266
timestamp 1667941163
transform 1 0 143136 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1271
timestamp 1667941163
transform 1 0 143696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1279
timestamp 1667941163
transform 1 0 144592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1281
timestamp 1667941163
transform 1 0 144816 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1286
timestamp 1667941163
transform 1 0 145376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1294
timestamp 1667941163
transform 1 0 146272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1297
timestamp 1667941163
transform 1 0 146608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1302
timestamp 1667941163
transform 1 0 147168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1310
timestamp 1667941163
transform 1 0 148064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1316
timestamp 1667941163
transform 1 0 148736 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1324
timestamp 1667941163
transform 1 0 149632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1328
timestamp 1667941163
transform 1 0 150080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1332
timestamp 1667941163
transform 1 0 150528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1337
timestamp 1667941163
transform 1 0 151088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1341
timestamp 1667941163
transform 1 0 151536 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1346
timestamp 1667941163
transform 1 0 152096 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1354
timestamp 1667941163
transform 1 0 152992 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1356
timestamp 1667941163
transform 1 0 153216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1361
timestamp 1667941163
transform 1 0 153776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1367
timestamp 1667941163
transform 1 0 154448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1371
timestamp 1667941163
transform 1 0 154896 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1376
timestamp 1667941163
transform 1 0 155456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1384
timestamp 1667941163
transform 1 0 156352 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1386
timestamp 1667941163
transform 1 0 156576 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1391
timestamp 1667941163
transform 1 0 157136 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1399
timestamp 1667941163
transform 1 0 158032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1402
timestamp 1667941163
transform 1 0 158368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1407
timestamp 1667941163
transform 1 0 158928 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1415
timestamp 1667941163
transform 1 0 159824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1421
timestamp 1667941163
transform 1 0 160496 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1429
timestamp 1667941163
transform 1 0 161392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1433
timestamp 1667941163
transform 1 0 161840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1437
timestamp 1667941163
transform 1 0 162288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1442
timestamp 1667941163
transform 1 0 162848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1446
timestamp 1667941163
transform 1 0 163296 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1451
timestamp 1667941163
transform 1 0 163856 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1459
timestamp 1667941163
transform 1 0 164752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1461
timestamp 1667941163
transform 1 0 164976 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1466
timestamp 1667941163
transform 1 0 165536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1472
timestamp 1667941163
transform 1 0 166208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1476
timestamp 1667941163
transform 1 0 166656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1481
timestamp 1667941163
transform 1 0 167216 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1489
timestamp 1667941163
transform 1 0 168112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1491
timestamp 1667941163
transform 1 0 168336 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1496
timestamp 1667941163
transform 1 0 168896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1504
timestamp 1667941163
transform 1 0 169792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1507
timestamp 1667941163
transform 1 0 170128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1512
timestamp 1667941163
transform 1 0 170688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1520
timestamp 1667941163
transform 1 0 171584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1526
timestamp 1667941163
transform 1 0 172256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1530
timestamp 1667941163
transform 1 0 172704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1536
timestamp 1667941163
transform 1 0 173376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1542
timestamp 1667941163
transform 1 0 174048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1547
timestamp 1667941163
transform 1 0 174608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1553
timestamp 1667941163
transform 1 0 175280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1569
timestamp 1667941163
transform 1 0 177072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1573
timestamp 1667941163
transform 1 0 177520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1577
timestamp 1667941163
transform 1 0 177968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1667941163
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1667941163
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1667941163
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1667941163
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1667941163
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1667941163
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1667941163
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1667941163
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1667941163
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1667941163
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1667941163
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1667941163
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428
timestamp 1667941163
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1667941163
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1667941163
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_499
timestamp 1667941163
transform 1 0 57232 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_563
timestamp 1667941163
transform 1 0 64400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1667941163
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_570
timestamp 1667941163
transform 1 0 65184 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_634
timestamp 1667941163
transform 1 0 72352 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1667941163
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_641
timestamp 1667941163
transform 1 0 73136 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_705
timestamp 1667941163
transform 1 0 80304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1667941163
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_712
timestamp 1667941163
transform 1 0 81088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_776
timestamp 1667941163
transform 1 0 88256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1667941163
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_783
timestamp 1667941163
transform 1 0 89040 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_847
timestamp 1667941163
transform 1 0 96208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1667941163
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_854
timestamp 1667941163
transform 1 0 96992 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_918
timestamp 1667941163
transform 1 0 104160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_922
timestamp 1667941163
transform 1 0 104608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_925
timestamp 1667941163
transform 1 0 104944 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_989
timestamp 1667941163
transform 1 0 112112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_993
timestamp 1667941163
transform 1 0 112560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_996
timestamp 1667941163
transform 1 0 112896 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1060
timestamp 1667941163
transform 1 0 120064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1064
timestamp 1667941163
transform 1 0 120512 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1067
timestamp 1667941163
transform 1 0 120848 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1131
timestamp 1667941163
transform 1 0 128016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1135
timestamp 1667941163
transform 1 0 128464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1138
timestamp 1667941163
transform 1 0 128800 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1202
timestamp 1667941163
transform 1 0 135968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1667941163
transform 1 0 136416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1209
timestamp 1667941163
transform 1 0 136752 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1273
timestamp 1667941163
transform 1 0 143920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1277
timestamp 1667941163
transform 1 0 144368 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1280
timestamp 1667941163
transform 1 0 144704 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1344
timestamp 1667941163
transform 1 0 151872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1348
timestamp 1667941163
transform 1 0 152320 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1351
timestamp 1667941163
transform 1 0 152656 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1415
timestamp 1667941163
transform 1 0 159824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1419
timestamp 1667941163
transform 1 0 160272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1422
timestamp 1667941163
transform 1 0 160608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1486
timestamp 1667941163
transform 1 0 167776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1490
timestamp 1667941163
transform 1 0 168224 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1493
timestamp 1667941163
transform 1 0 168560 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1557
timestamp 1667941163
transform 1 0 175728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1561
timestamp 1667941163
transform 1 0 176176 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1564
timestamp 1667941163
transform 1 0 176512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1580
timestamp 1667941163
transform 1 0 178304 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1667941163
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1667941163
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1667941163
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1667941163
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1667941163
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1667941163
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1667941163
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1667941163
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1667941163
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1667941163
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1667941163
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1667941163
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1667941163
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1667941163
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1667941163
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1667941163
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1667941163
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_463
timestamp 1667941163
transform 1 0 53200 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1667941163
transform 1 0 60368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1667941163
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_534
timestamp 1667941163
transform 1 0 61152 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_598
timestamp 1667941163
transform 1 0 68320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1667941163
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_605
timestamp 1667941163
transform 1 0 69104 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_669
timestamp 1667941163
transform 1 0 76272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1667941163
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_676
timestamp 1667941163
transform 1 0 77056 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_740
timestamp 1667941163
transform 1 0 84224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1667941163
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_747
timestamp 1667941163
transform 1 0 85008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_811
timestamp 1667941163
transform 1 0 92176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1667941163
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_818
timestamp 1667941163
transform 1 0 92960 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_882
timestamp 1667941163
transform 1 0 100128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_886
timestamp 1667941163
transform 1 0 100576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_889
timestamp 1667941163
transform 1 0 100912 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_953
timestamp 1667941163
transform 1 0 108080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1667941163
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_960
timestamp 1667941163
transform 1 0 108864 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1024
timestamp 1667941163
transform 1 0 116032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1667941163
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1031
timestamp 1667941163
transform 1 0 116816 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1095
timestamp 1667941163
transform 1 0 123984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1099
timestamp 1667941163
transform 1 0 124432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1102
timestamp 1667941163
transform 1 0 124768 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1166
timestamp 1667941163
transform 1 0 131936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1170
timestamp 1667941163
transform 1 0 132384 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1173
timestamp 1667941163
transform 1 0 132720 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1237
timestamp 1667941163
transform 1 0 139888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1241
timestamp 1667941163
transform 1 0 140336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1244
timestamp 1667941163
transform 1 0 140672 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1308
timestamp 1667941163
transform 1 0 147840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1312
timestamp 1667941163
transform 1 0 148288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1315
timestamp 1667941163
transform 1 0 148624 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1379
timestamp 1667941163
transform 1 0 155792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1383
timestamp 1667941163
transform 1 0 156240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1386
timestamp 1667941163
transform 1 0 156576 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1450
timestamp 1667941163
transform 1 0 163744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1454
timestamp 1667941163
transform 1 0 164192 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1457
timestamp 1667941163
transform 1 0 164528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1521
timestamp 1667941163
transform 1 0 171696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1525
timestamp 1667941163
transform 1 0 172144 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_1528
timestamp 1667941163
transform 1 0 172480 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1560
timestamp 1667941163
transform 1 0 176064 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1576
timestamp 1667941163
transform 1 0 177856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1580
timestamp 1667941163
transform 1 0 178304 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1667941163
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1667941163
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1667941163
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1667941163
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1667941163
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1667941163
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1667941163
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1667941163
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1667941163
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1667941163
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1667941163
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1667941163
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1667941163
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1667941163
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1667941163
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1667941163
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1667941163
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1667941163
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1667941163
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1667941163
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1667941163
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1667941163
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_641
timestamp 1667941163
transform 1 0 73136 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_705
timestamp 1667941163
transform 1 0 80304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1667941163
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_712
timestamp 1667941163
transform 1 0 81088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_776
timestamp 1667941163
transform 1 0 88256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1667941163
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_783
timestamp 1667941163
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_847
timestamp 1667941163
transform 1 0 96208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1667941163
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_854
timestamp 1667941163
transform 1 0 96992 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_918
timestamp 1667941163
transform 1 0 104160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1667941163
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_925
timestamp 1667941163
transform 1 0 104944 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_989
timestamp 1667941163
transform 1 0 112112 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1667941163
transform 1 0 112560 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_996
timestamp 1667941163
transform 1 0 112896 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1060
timestamp 1667941163
transform 1 0 120064 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1064
timestamp 1667941163
transform 1 0 120512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1067
timestamp 1667941163
transform 1 0 120848 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1131
timestamp 1667941163
transform 1 0 128016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1135
timestamp 1667941163
transform 1 0 128464 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1138
timestamp 1667941163
transform 1 0 128800 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1202
timestamp 1667941163
transform 1 0 135968 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1206
timestamp 1667941163
transform 1 0 136416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1209
timestamp 1667941163
transform 1 0 136752 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1273
timestamp 1667941163
transform 1 0 143920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1667941163
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1280
timestamp 1667941163
transform 1 0 144704 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1344
timestamp 1667941163
transform 1 0 151872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1348
timestamp 1667941163
transform 1 0 152320 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1351
timestamp 1667941163
transform 1 0 152656 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1415
timestamp 1667941163
transform 1 0 159824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1419
timestamp 1667941163
transform 1 0 160272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1422
timestamp 1667941163
transform 1 0 160608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1486
timestamp 1667941163
transform 1 0 167776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1490
timestamp 1667941163
transform 1 0 168224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1493
timestamp 1667941163
transform 1 0 168560 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1557
timestamp 1667941163
transform 1 0 175728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1561
timestamp 1667941163
transform 1 0 176176 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1564
timestamp 1667941163
transform 1 0 176512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1580
timestamp 1667941163
transform 1 0 178304 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1667941163
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1667941163
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1667941163
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1667941163
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1667941163
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1667941163
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1667941163
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1667941163
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1667941163
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1667941163
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1667941163
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1667941163
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1667941163
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1667941163
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1667941163
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1667941163
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1667941163
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1667941163
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1667941163
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1667941163
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1667941163
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1667941163
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1667941163
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1667941163
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1667941163
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1667941163
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1667941163
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1667941163
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1667941163
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1667941163
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1667941163
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_818
timestamp 1667941163
transform 1 0 92960 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_882
timestamp 1667941163
transform 1 0 100128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1667941163
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_889
timestamp 1667941163
transform 1 0 100912 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_953
timestamp 1667941163
transform 1 0 108080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1667941163
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_960
timestamp 1667941163
transform 1 0 108864 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1024
timestamp 1667941163
transform 1 0 116032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1028
timestamp 1667941163
transform 1 0 116480 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1031
timestamp 1667941163
transform 1 0 116816 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1095
timestamp 1667941163
transform 1 0 123984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1667941163
transform 1 0 124432 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1102
timestamp 1667941163
transform 1 0 124768 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1166
timestamp 1667941163
transform 1 0 131936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1170
timestamp 1667941163
transform 1 0 132384 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1173
timestamp 1667941163
transform 1 0 132720 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1237
timestamp 1667941163
transform 1 0 139888 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1241
timestamp 1667941163
transform 1 0 140336 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1244
timestamp 1667941163
transform 1 0 140672 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1308
timestamp 1667941163
transform 1 0 147840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1312
timestamp 1667941163
transform 1 0 148288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1315
timestamp 1667941163
transform 1 0 148624 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1379
timestamp 1667941163
transform 1 0 155792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1383
timestamp 1667941163
transform 1 0 156240 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1386
timestamp 1667941163
transform 1 0 156576 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1450
timestamp 1667941163
transform 1 0 163744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1454
timestamp 1667941163
transform 1 0 164192 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1457
timestamp 1667941163
transform 1 0 164528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1521
timestamp 1667941163
transform 1 0 171696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1525
timestamp 1667941163
transform 1 0 172144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1528
timestamp 1667941163
transform 1 0 172480 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1560
timestamp 1667941163
transform 1 0 176064 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1576
timestamp 1667941163
transform 1 0 177856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1580
timestamp 1667941163
transform 1 0 178304 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1667941163
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1667941163
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1667941163
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1667941163
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1667941163
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1667941163
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1667941163
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1667941163
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1667941163
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1667941163
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1667941163
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1667941163
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1667941163
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1667941163
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1667941163
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1667941163
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1667941163
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1667941163
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1667941163
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1667941163
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1667941163
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1667941163
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1667941163
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1667941163
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1667941163
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1667941163
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1667941163
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1667941163
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1667941163
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1667941163
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1667941163
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1667941163
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_854
timestamp 1667941163
transform 1 0 96992 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_918
timestamp 1667941163
transform 1 0 104160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_922
timestamp 1667941163
transform 1 0 104608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_925
timestamp 1667941163
transform 1 0 104944 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1667941163
transform 1 0 112112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1667941163
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_996
timestamp 1667941163
transform 1 0 112896 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1060
timestamp 1667941163
transform 1 0 120064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1064
timestamp 1667941163
transform 1 0 120512 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1067
timestamp 1667941163
transform 1 0 120848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1131
timestamp 1667941163
transform 1 0 128016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1667941163
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1138
timestamp 1667941163
transform 1 0 128800 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1202
timestamp 1667941163
transform 1 0 135968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1667941163
transform 1 0 136416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1209
timestamp 1667941163
transform 1 0 136752 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1273
timestamp 1667941163
transform 1 0 143920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1277
timestamp 1667941163
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1280
timestamp 1667941163
transform 1 0 144704 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1344
timestamp 1667941163
transform 1 0 151872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1348
timestamp 1667941163
transform 1 0 152320 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1351
timestamp 1667941163
transform 1 0 152656 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1415
timestamp 1667941163
transform 1 0 159824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1419
timestamp 1667941163
transform 1 0 160272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1422
timestamp 1667941163
transform 1 0 160608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1486
timestamp 1667941163
transform 1 0 167776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1490
timestamp 1667941163
transform 1 0 168224 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1493
timestamp 1667941163
transform 1 0 168560 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1557
timestamp 1667941163
transform 1 0 175728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1561
timestamp 1667941163
transform 1 0 176176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1564
timestamp 1667941163
transform 1 0 176512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1580
timestamp 1667941163
transform 1 0 178304 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1667941163
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1667941163
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1667941163
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1667941163
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1667941163
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_179
timestamp 1667941163
transform 1 0 21392 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_182
timestamp 1667941163
transform 1 0 21728 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_186
timestamp 1667941163
transform 1 0 22176 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_190
timestamp 1667941163
transform 1 0 22624 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_222
timestamp 1667941163
transform 1 0 26208 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_238
timestamp 1667941163
transform 1 0 28000 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_246
timestamp 1667941163
transform 1 0 28896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1667941163
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1667941163
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1667941163
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1667941163
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1667941163
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1667941163
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1667941163
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1667941163
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1667941163
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1667941163
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1667941163
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1667941163
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1667941163
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1667941163
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1667941163
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1667941163
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1667941163
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1667941163
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1667941163
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1667941163
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1667941163
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1667941163
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1667941163
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1667941163
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_818
timestamp 1667941163
transform 1 0 92960 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_834
timestamp 1667941163
transform 1 0 94752 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_840
timestamp 1667941163
transform 1 0 95424 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_872
timestamp 1667941163
transform 1 0 99008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_880
timestamp 1667941163
transform 1 0 99904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_884
timestamp 1667941163
transform 1 0 100352 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1667941163
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1667941163
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1667941163
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1667941163
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1667941163
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1667941163
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1667941163
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1031
timestamp 1667941163
transform 1 0 116816 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1095
timestamp 1667941163
transform 1 0 123984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1099
timestamp 1667941163
transform 1 0 124432 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1102
timestamp 1667941163
transform 1 0 124768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1166
timestamp 1667941163
transform 1 0 131936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1170
timestamp 1667941163
transform 1 0 132384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1173
timestamp 1667941163
transform 1 0 132720 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1237
timestamp 1667941163
transform 1 0 139888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1241
timestamp 1667941163
transform 1 0 140336 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1244
timestamp 1667941163
transform 1 0 140672 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1308
timestamp 1667941163
transform 1 0 147840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1312
timestamp 1667941163
transform 1 0 148288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1315
timestamp 1667941163
transform 1 0 148624 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1379
timestamp 1667941163
transform 1 0 155792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1383
timestamp 1667941163
transform 1 0 156240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1386
timestamp 1667941163
transform 1 0 156576 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1450
timestamp 1667941163
transform 1 0 163744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1454
timestamp 1667941163
transform 1 0 164192 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1457
timestamp 1667941163
transform 1 0 164528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1521
timestamp 1667941163
transform 1 0 171696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1525
timestamp 1667941163
transform 1 0 172144 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1528
timestamp 1667941163
transform 1 0 172480 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1560
timestamp 1667941163
transform 1 0 176064 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1576
timestamp 1667941163
transform 1 0 177856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1580
timestamp 1667941163
transform 1 0 178304 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1667941163
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1667941163
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_144
timestamp 1667941163
transform 1 0 17472 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_160
timestamp 1667941163
transform 1 0 19264 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_168
timestamp 1667941163
transform 1 0 20160 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_172
timestamp 1667941163
transform 1 0 20608 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_180
timestamp 1667941163
transform 1 0 21504 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_188
timestamp 1667941163
transform 1 0 22400 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_192
timestamp 1667941163
transform 1 0 22848 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_196
timestamp 1667941163
transform 1 0 23296 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1667941163
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1667941163
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1667941163
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1667941163
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1667941163
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1667941163
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1667941163
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1667941163
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1667941163
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1667941163
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1667941163
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1667941163
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1667941163
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1667941163
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1667941163
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1667941163
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1667941163
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1667941163
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1667941163
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1667941163
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1667941163
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1667941163
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1667941163
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1667941163
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1667941163
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_783
timestamp 1667941163
transform 1 0 89040 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_815
timestamp 1667941163
transform 1 0 92624 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_823
timestamp 1667941163
transform 1 0 93520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_825
timestamp 1667941163
transform 1 0 93744 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_828
timestamp 1667941163
transform 1 0 94080 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_836
timestamp 1667941163
transform 1 0 94976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_846
timestamp 1667941163
transform 1 0 96096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_850
timestamp 1667941163
transform 1 0 96544 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1667941163
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1667941163
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1667941163
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1667941163
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1667941163
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1667941163
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_996
timestamp 1667941163
transform 1 0 112896 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1060
timestamp 1667941163
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1667941163
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1067
timestamp 1667941163
transform 1 0 120848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1131
timestamp 1667941163
transform 1 0 128016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1135
timestamp 1667941163
transform 1 0 128464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1138
timestamp 1667941163
transform 1 0 128800 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1667941163
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1667941163
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1667941163
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1667941163
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1667941163
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1280
timestamp 1667941163
transform 1 0 144704 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1344
timestamp 1667941163
transform 1 0 151872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1348
timestamp 1667941163
transform 1 0 152320 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1351
timestamp 1667941163
transform 1 0 152656 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1415
timestamp 1667941163
transform 1 0 159824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1419
timestamp 1667941163
transform 1 0 160272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1422
timestamp 1667941163
transform 1 0 160608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1486
timestamp 1667941163
transform 1 0 167776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1490
timestamp 1667941163
transform 1 0 168224 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1493
timestamp 1667941163
transform 1 0 168560 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1557
timestamp 1667941163
transform 1 0 175728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1561
timestamp 1667941163
transform 1 0 176176 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1564
timestamp 1667941163
transform 1 0 176512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1580
timestamp 1667941163
transform 1 0 178304 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1667941163
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1667941163
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1667941163
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_108
timestamp 1667941163
transform 1 0 13440 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_140
timestamp 1667941163
transform 1 0 17024 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_156
timestamp 1667941163
transform 1 0 18816 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_160
timestamp 1667941163
transform 1 0 19264 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_164
timestamp 1667941163
transform 1 0 19712 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_168
timestamp 1667941163
transform 1 0 20160 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_179
timestamp 1667941163
transform 1 0 21392 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_186
timestamp 1667941163
transform 1 0 22176 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 23072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_198
timestamp 1667941163
transform 1 0 23520 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_202
timestamp 1667941163
transform 1 0 23968 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_206
timestamp 1667941163
transform 1 0 24416 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_238
timestamp 1667941163
transform 1 0 28000 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_246
timestamp 1667941163
transform 1 0 28896 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1667941163
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1667941163
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1667941163
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_321
timestamp 1667941163
transform 1 0 37296 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_337
timestamp 1667941163
transform 1 0 39088 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_345
timestamp 1667941163
transform 1 0 39984 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_347
timestamp 1667941163
transform 1 0 40208 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_352
timestamp 1667941163
transform 1 0 40768 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_384
timestamp 1667941163
transform 1 0 44352 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_388
timestamp 1667941163
transform 1 0 44800 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1667941163
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1667941163
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1667941163
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1667941163
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1667941163
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1667941163
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1667941163
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1667941163
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1667941163
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1667941163
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1667941163
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1667941163
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1667941163
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1667941163
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1667941163
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1667941163
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1667941163
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1667941163
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1667941163
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1667941163
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1667941163
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1667941163
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1667941163
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1667941163
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1667941163
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1667941163
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1667941163
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1031
timestamp 1667941163
transform 1 0 116816 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1095
timestamp 1667941163
transform 1 0 123984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1099
timestamp 1667941163
transform 1 0 124432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1102
timestamp 1667941163
transform 1 0 124768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1166
timestamp 1667941163
transform 1 0 131936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1170
timestamp 1667941163
transform 1 0 132384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1667941163
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1667941163
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1667941163
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1244
timestamp 1667941163
transform 1 0 140672 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1308
timestamp 1667941163
transform 1 0 147840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1312
timestamp 1667941163
transform 1 0 148288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1315
timestamp 1667941163
transform 1 0 148624 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1379
timestamp 1667941163
transform 1 0 155792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1383
timestamp 1667941163
transform 1 0 156240 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1386
timestamp 1667941163
transform 1 0 156576 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1450
timestamp 1667941163
transform 1 0 163744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1454
timestamp 1667941163
transform 1 0 164192 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1457
timestamp 1667941163
transform 1 0 164528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1521
timestamp 1667941163
transform 1 0 171696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1525
timestamp 1667941163
transform 1 0 172144 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1528
timestamp 1667941163
transform 1 0 172480 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_1560
timestamp 1667941163
transform 1 0 176064 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1576
timestamp 1667941163
transform 1 0 177856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1580
timestamp 1667941163
transform 1 0 178304 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1667941163
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1667941163
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_144
timestamp 1667941163
transform 1 0 17472 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_148
timestamp 1667941163
transform 1 0 17920 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_151
timestamp 1667941163
transform 1 0 18256 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_155
timestamp 1667941163
transform 1 0 18704 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_163
timestamp 1667941163
transform 1 0 19600 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_171
timestamp 1667941163
transform 1 0 20496 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_179
timestamp 1667941163
transform 1 0 21392 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_187
timestamp 1667941163
transform 1 0 22288 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_195
timestamp 1667941163
transform 1 0 23184 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_199
timestamp 1667941163
transform 1 0 23632 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_205
timestamp 1667941163
transform 1 0 24304 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_209
timestamp 1667941163
transform 1 0 24752 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1667941163
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1667941163
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1667941163
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_286
timestamp 1667941163
transform 1 0 33376 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_318
timestamp 1667941163
transform 1 0 36960 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_334
timestamp 1667941163
transform 1 0 38752 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_346
timestamp 1667941163
transform 1 0 40096 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_352
timestamp 1667941163
transform 1 0 40768 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1667941163
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1667941163
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_362
timestamp 1667941163
transform 1 0 41888 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_428
timestamp 1667941163
transform 1 0 49280 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_444
timestamp 1667941163
transform 1 0 51072 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_452
timestamp 1667941163
transform 1 0 51968 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_458
timestamp 1667941163
transform 1 0 52640 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_490
timestamp 1667941163
transform 1 0 56224 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_494
timestamp 1667941163
transform 1 0 56672 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1667941163
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_499
timestamp 1667941163
transform 1 0 57232 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_531
timestamp 1667941163
transform 1 0 60816 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_543
timestamp 1667941163
transform 1 0 62160 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_559
timestamp 1667941163
transform 1 0 63952 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1667941163
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1667941163
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1667941163
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1667941163
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1667941163
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1667941163
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1667941163
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1667941163
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1667941163
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1667941163
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1667941163
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1667941163
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1667941163
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1667941163
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1667941163
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1667941163
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1667941163
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1667941163
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1667941163
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_996
timestamp 1667941163
transform 1 0 112896 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1667941163
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1667941163
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1667941163
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1667941163
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1667941163
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1667941163
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1667941163
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1667941163
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1667941163
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1667941163
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1667941163
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1280
timestamp 1667941163
transform 1 0 144704 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1344
timestamp 1667941163
transform 1 0 151872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1348
timestamp 1667941163
transform 1 0 152320 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1351
timestamp 1667941163
transform 1 0 152656 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1415
timestamp 1667941163
transform 1 0 159824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1419
timestamp 1667941163
transform 1 0 160272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1422
timestamp 1667941163
transform 1 0 160608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1486
timestamp 1667941163
transform 1 0 167776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1490
timestamp 1667941163
transform 1 0 168224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1493
timestamp 1667941163
transform 1 0 168560 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1557
timestamp 1667941163
transform 1 0 175728 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1561
timestamp 1667941163
transform 1 0 176176 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_1564
timestamp 1667941163
transform 1 0 176512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1580
timestamp 1667941163
transform 1 0 178304 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1667941163
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1667941163
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1667941163
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_108
timestamp 1667941163
transform 1 0 13440 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_140
timestamp 1667941163
transform 1 0 17024 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_144
timestamp 1667941163
transform 1 0 17472 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_152
timestamp 1667941163
transform 1 0 18368 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_160
timestamp 1667941163
transform 1 0 19264 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_168
timestamp 1667941163
transform 1 0 20160 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_179
timestamp 1667941163
transform 1 0 21392 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_187
timestamp 1667941163
transform 1 0 22288 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_195
timestamp 1667941163
transform 1 0 23184 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_203
timestamp 1667941163
transform 1 0 24080 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_207
timestamp 1667941163
transform 1 0 24528 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_211
timestamp 1667941163
transform 1 0 24976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_221
timestamp 1667941163
transform 1 0 26096 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_227
timestamp 1667941163
transform 1 0 26768 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1667941163
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1667941163
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1667941163
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_321
timestamp 1667941163
transform 1 0 37296 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_337
timestamp 1667941163
transform 1 0 39088 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_342
timestamp 1667941163
transform 1 0 39648 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_348
timestamp 1667941163
transform 1 0 40320 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_354
timestamp 1667941163
transform 1 0 40992 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_360
timestamp 1667941163
transform 1 0 41664 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_366
timestamp 1667941163
transform 1 0 42336 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_372
timestamp 1667941163
transform 1 0 43008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_388
timestamp 1667941163
transform 1 0 44800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_392
timestamp 1667941163
transform 1 0 45248 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_424
timestamp 1667941163
transform 1 0 48832 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_440
timestamp 1667941163
transform 1 0 50624 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_448
timestamp 1667941163
transform 1 0 51520 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_453
timestamp 1667941163
transform 1 0 52080 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_459
timestamp 1667941163
transform 1 0 52752 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1667941163
transform 1 0 53200 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_468
timestamp 1667941163
transform 1 0 53760 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_500
timestamp 1667941163
transform 1 0 57344 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_516
timestamp 1667941163
transform 1 0 59136 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_524
timestamp 1667941163
transform 1 0 60032 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_526
timestamp 1667941163
transform 1 0 60256 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1667941163
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_534
timestamp 1667941163
transform 1 0 61152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_539
timestamp 1667941163
transform 1 0 61712 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_545
timestamp 1667941163
transform 1 0 62384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_553
timestamp 1667941163
transform 1 0 63280 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_559
timestamp 1667941163
transform 1 0 63952 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_591
timestamp 1667941163
transform 1 0 67536 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_599
timestamp 1667941163
transform 1 0 68432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1667941163
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1667941163
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1667941163
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1667941163
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1667941163
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1667941163
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1667941163
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1667941163
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1667941163
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1667941163
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_882
timestamp 1667941163
transform 1 0 100128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1667941163
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1667941163
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1667941163
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1667941163
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1667941163
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1667941163
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1667941163
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1667941163
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1667941163
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1667941163
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1667941163
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1667941163
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1667941163
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1667941163
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1667941163
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1667941163
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1244
timestamp 1667941163
transform 1 0 140672 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1308
timestamp 1667941163
transform 1 0 147840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1312
timestamp 1667941163
transform 1 0 148288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1315
timestamp 1667941163
transform 1 0 148624 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1379
timestamp 1667941163
transform 1 0 155792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1383
timestamp 1667941163
transform 1 0 156240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1386
timestamp 1667941163
transform 1 0 156576 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1450
timestamp 1667941163
transform 1 0 163744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1454
timestamp 1667941163
transform 1 0 164192 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1457
timestamp 1667941163
transform 1 0 164528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1521
timestamp 1667941163
transform 1 0 171696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1525
timestamp 1667941163
transform 1 0 172144 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_1528
timestamp 1667941163
transform 1 0 172480 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_1560
timestamp 1667941163
transform 1 0 176064 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1576
timestamp 1667941163
transform 1 0 177856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1580
timestamp 1667941163
transform 1 0 178304 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1667941163
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_73
timestamp 1667941163
transform 1 0 9520 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_105
timestamp 1667941163
transform 1 0 13104 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_121
timestamp 1667941163
transform 1 0 14896 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_129
timestamp 1667941163
transform 1 0 15792 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_133
timestamp 1667941163
transform 1 0 16240 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1667941163
transform 1 0 17472 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_147
timestamp 1667941163
transform 1 0 17808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_155
timestamp 1667941163
transform 1 0 18704 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_163
timestamp 1667941163
transform 1 0 19600 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_171
timestamp 1667941163
transform 1 0 20496 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_179
timestamp 1667941163
transform 1 0 21392 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_187
timestamp 1667941163
transform 1 0 22288 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_195
timestamp 1667941163
transform 1 0 23184 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_203
timestamp 1667941163
transform 1 0 24080 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_211
timestamp 1667941163
transform 1 0 24976 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1667941163
transform 1 0 25424 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_224
timestamp 1667941163
transform 1 0 26432 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_232
timestamp 1667941163
transform 1 0 27328 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_238
timestamp 1667941163
transform 1 0 28000 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_270
timestamp 1667941163
transform 1 0 31584 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_278
timestamp 1667941163
transform 1 0 32480 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1667941163
transform 1 0 32928 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_286
timestamp 1667941163
transform 1 0 33376 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_318
timestamp 1667941163
transform 1 0 36960 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_334
timestamp 1667941163
transform 1 0 38752 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_336
timestamp 1667941163
transform 1 0 38976 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_341
timestamp 1667941163
transform 1 0 39536 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_347
timestamp 1667941163
transform 1 0 40208 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_353
timestamp 1667941163
transform 1 0 40880 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1667941163
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_362
timestamp 1667941163
transform 1 0 41888 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1667941163
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1667941163
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1667941163
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_499
timestamp 1667941163
transform 1 0 57232 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_515
timestamp 1667941163
transform 1 0 59024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_523
timestamp 1667941163
transform 1 0 59920 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_528
timestamp 1667941163
transform 1 0 60480 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_534
timestamp 1667941163
transform 1 0 61152 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_540
timestamp 1667941163
transform 1 0 61824 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_546
timestamp 1667941163
transform 1 0 62496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_550
timestamp 1667941163
transform 1 0 62944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_555
timestamp 1667941163
transform 1 0 63504 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_561
timestamp 1667941163
transform 1 0 64176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_565
timestamp 1667941163
transform 1 0 64624 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1667941163
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1667941163
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1667941163
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1667941163
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1667941163
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1667941163
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1667941163
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1667941163
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1667941163
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1667941163
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1667941163
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1667941163
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1667941163
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_854
timestamp 1667941163
transform 1 0 96992 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_918
timestamp 1667941163
transform 1 0 104160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1667941163
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1667941163
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1667941163
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1667941163
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1667941163
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1667941163
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1667941163
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1667941163
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1667941163
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1667941163
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1667941163
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1667941163
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1667941163
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1667941163
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1273
timestamp 1667941163
transform 1 0 143920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1667941163
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1280
timestamp 1667941163
transform 1 0 144704 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1344
timestamp 1667941163
transform 1 0 151872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1348
timestamp 1667941163
transform 1 0 152320 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1351
timestamp 1667941163
transform 1 0 152656 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1415
timestamp 1667941163
transform 1 0 159824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1419
timestamp 1667941163
transform 1 0 160272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1422
timestamp 1667941163
transform 1 0 160608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1486
timestamp 1667941163
transform 1 0 167776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1490
timestamp 1667941163
transform 1 0 168224 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1493
timestamp 1667941163
transform 1 0 168560 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1557
timestamp 1667941163
transform 1 0 175728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1561
timestamp 1667941163
transform 1 0 176176 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_1564
timestamp 1667941163
transform 1 0 176512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1580
timestamp 1667941163
transform 1 0 178304 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1667941163
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1667941163
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1667941163
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_108
timestamp 1667941163
transform 1 0 13440 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_124
timestamp 1667941163
transform 1 0 15232 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_132
timestamp 1667941163
transform 1 0 16128 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_150
timestamp 1667941163
transform 1 0 18144 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_160
timestamp 1667941163
transform 1 0 19264 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_168
timestamp 1667941163
transform 1 0 20160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1667941163
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_206
timestamp 1667941163
transform 1 0 24416 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_214
timestamp 1667941163
transform 1 0 25312 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_218
timestamp 1667941163
transform 1 0 25760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_226
timestamp 1667941163
transform 1 0 26656 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_242
timestamp 1667941163
transform 1 0 28448 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_246
timestamp 1667941163
transform 1 0 28896 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1667941163
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1667941163
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1667941163
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_321
timestamp 1667941163
transform 1 0 37296 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_337
timestamp 1667941163
transform 1 0 39088 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_349
timestamp 1667941163
transform 1 0 40432 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_355
timestamp 1667941163
transform 1 0 41104 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_387
timestamp 1667941163
transform 1 0 44688 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1667941163
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1667941163
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1667941163
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1667941163
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1667941163
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1667941163
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1667941163
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_534
timestamp 1667941163
transform 1 0 61152 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_542
timestamp 1667941163
transform 1 0 62048 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_548
timestamp 1667941163
transform 1 0 62720 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_554
timestamp 1667941163
transform 1 0 63392 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_586
timestamp 1667941163
transform 1 0 66976 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1667941163
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1667941163
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1667941163
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1667941163
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1667941163
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1667941163
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1667941163
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1667941163
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1667941163
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1667941163
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1667941163
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1667941163
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1667941163
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_889
timestamp 1667941163
transform 1 0 100912 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_953
timestamp 1667941163
transform 1 0 108080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1667941163
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1667941163
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1667941163
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1667941163
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1667941163
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1667941163
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1667941163
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1667941163
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1667941163
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1667941163
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1667941163
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1667941163
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1667941163
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1244
timestamp 1667941163
transform 1 0 140672 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1308
timestamp 1667941163
transform 1 0 147840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1312
timestamp 1667941163
transform 1 0 148288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1315
timestamp 1667941163
transform 1 0 148624 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1379
timestamp 1667941163
transform 1 0 155792 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1383
timestamp 1667941163
transform 1 0 156240 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1386
timestamp 1667941163
transform 1 0 156576 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1450
timestamp 1667941163
transform 1 0 163744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1454
timestamp 1667941163
transform 1 0 164192 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1457
timestamp 1667941163
transform 1 0 164528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1521
timestamp 1667941163
transform 1 0 171696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1525
timestamp 1667941163
transform 1 0 172144 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_1528
timestamp 1667941163
transform 1 0 172480 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_1560
timestamp 1667941163
transform 1 0 176064 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1576
timestamp 1667941163
transform 1 0 177856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1580
timestamp 1667941163
transform 1 0 178304 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1667941163
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_73
timestamp 1667941163
transform 1 0 9520 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_105
timestamp 1667941163
transform 1 0 13104 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_121
timestamp 1667941163
transform 1 0 14896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_129
timestamp 1667941163
transform 1 0 15792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_133
timestamp 1667941163
transform 1 0 16240 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_137
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_144
timestamp 1667941163
transform 1 0 17472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_148
timestamp 1667941163
transform 1 0 17920 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_152
timestamp 1667941163
transform 1 0 18368 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_156
timestamp 1667941163
transform 1 0 18816 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_164
timestamp 1667941163
transform 1 0 19712 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_172
timestamp 1667941163
transform 1 0 20608 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_180
timestamp 1667941163
transform 1 0 21504 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_208
timestamp 1667941163
transform 1 0 24640 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1667941163
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1667941163
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1667941163
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1667941163
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1667941163
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1667941163
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1667941163
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1667941163
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1667941163
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1667941163
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1667941163
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1667941163
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_499
timestamp 1667941163
transform 1 0 57232 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_531
timestamp 1667941163
transform 1 0 60816 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_535
timestamp 1667941163
transform 1 0 61264 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_541
timestamp 1667941163
transform 1 0 61936 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_557
timestamp 1667941163
transform 1 0 63728 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_565
timestamp 1667941163
transform 1 0 64624 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1667941163
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1667941163
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1667941163
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1667941163
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1667941163
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1667941163
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1667941163
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1667941163
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1667941163
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1667941163
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1667941163
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1667941163
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1667941163
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1667941163
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1667941163
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1667941163
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1667941163
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1667941163
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1667941163
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1667941163
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1667941163
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1667941163
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1667941163
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1667941163
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1667941163
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1667941163
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1667941163
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1667941163
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1667941163
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1667941163
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1667941163
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1280
timestamp 1667941163
transform 1 0 144704 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1344
timestamp 1667941163
transform 1 0 151872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1348
timestamp 1667941163
transform 1 0 152320 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1351
timestamp 1667941163
transform 1 0 152656 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1415
timestamp 1667941163
transform 1 0 159824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1419
timestamp 1667941163
transform 1 0 160272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1422
timestamp 1667941163
transform 1 0 160608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1486
timestamp 1667941163
transform 1 0 167776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1490
timestamp 1667941163
transform 1 0 168224 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1493
timestamp 1667941163
transform 1 0 168560 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1557
timestamp 1667941163
transform 1 0 175728 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1561
timestamp 1667941163
transform 1 0 176176 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_1564
timestamp 1667941163
transform 1 0 176512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1580
timestamp 1667941163
transform 1 0 178304 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1667941163
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_37
timestamp 1667941163
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_69
timestamp 1667941163
transform 1 0 9072 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_85
timestamp 1667941163
transform 1 0 10864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_88
timestamp 1667941163
transform 1 0 11200 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_96
timestamp 1667941163
transform 1 0 12096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_98
timestamp 1667941163
transform 1 0 12320 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_103
timestamp 1667941163
transform 1 0 12880 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_108
timestamp 1667941163
transform 1 0 13440 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_116
timestamp 1667941163
transform 1 0 14336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_120
timestamp 1667941163
transform 1 0 14784 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_139
timestamp 1667941163
transform 1 0 16912 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_158
timestamp 1667941163
transform 1 0 19040 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_164
timestamp 1667941163
transform 1 0 19712 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_168
timestamp 1667941163
transform 1 0 20160 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1667941163
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_179
timestamp 1667941163
transform 1 0 21392 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_181
timestamp 1667941163
transform 1 0 21616 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_192
timestamp 1667941163
transform 1 0 22848 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_200
timestamp 1667941163
transform 1 0 23744 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_204
timestamp 1667941163
transform 1 0 24192 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_236
timestamp 1667941163
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_244
timestamp 1667941163
transform 1 0 28672 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_250
timestamp 1667941163
transform 1 0 29344 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_254
timestamp 1667941163
transform 1 0 29792 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_257
timestamp 1667941163
transform 1 0 30128 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_261
timestamp 1667941163
transform 1 0 30576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_267
timestamp 1667941163
transform 1 0 31248 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_285
timestamp 1667941163
transform 1 0 33264 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_291
timestamp 1667941163
transform 1 0 33936 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_310
timestamp 1667941163
transform 1 0 36064 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1667941163
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1667941163
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1667941163
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1667941163
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1667941163
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1667941163
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1667941163
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_463
timestamp 1667941163
transform 1 0 53200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_469
timestamp 1667941163
transform 1 0 53872 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_501
timestamp 1667941163
transform 1 0 57456 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_517
timestamp 1667941163
transform 1 0 59248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_525
timestamp 1667941163
transform 1 0 60144 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_529
timestamp 1667941163
transform 1 0 60592 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1667941163
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_534
timestamp 1667941163
transform 1 0 61152 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_542
timestamp 1667941163
transform 1 0 62048 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_546
timestamp 1667941163
transform 1 0 62496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_548
timestamp 1667941163
transform 1 0 62720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_566
timestamp 1667941163
transform 1 0 64736 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1667941163
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1667941163
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_605
timestamp 1667941163
transform 1 0 69104 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_621
timestamp 1667941163
transform 1 0 70896 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_629
timestamp 1667941163
transform 1 0 71792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_633
timestamp 1667941163
transform 1 0 72240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_651
timestamp 1667941163
transform 1 0 74256 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_667
timestamp 1667941163
transform 1 0 76048 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_671
timestamp 1667941163
transform 1 0 76496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1667941163
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1667941163
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1667941163
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1667941163
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_747
timestamp 1667941163
transform 1 0 85008 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_763
timestamp 1667941163
transform 1 0 86800 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_771
timestamp 1667941163
transform 1 0 87696 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_773
timestamp 1667941163
transform 1 0 87920 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_791
timestamp 1667941163
transform 1 0 89936 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_807
timestamp 1667941163
transform 1 0 91728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1667941163
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1667941163
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1667941163
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1667941163
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1667941163
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1667941163
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1667941163
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1667941163
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1667941163
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1667941163
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1667941163
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1667941163
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1667941163
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1667941163
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1667941163
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1667941163
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1667941163
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1667941163
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1667941163
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1244
timestamp 1667941163
transform 1 0 140672 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1308
timestamp 1667941163
transform 1 0 147840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1312
timestamp 1667941163
transform 1 0 148288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1315
timestamp 1667941163
transform 1 0 148624 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1379
timestamp 1667941163
transform 1 0 155792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1383
timestamp 1667941163
transform 1 0 156240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1386
timestamp 1667941163
transform 1 0 156576 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1450
timestamp 1667941163
transform 1 0 163744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1454
timestamp 1667941163
transform 1 0 164192 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1457
timestamp 1667941163
transform 1 0 164528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1521
timestamp 1667941163
transform 1 0 171696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1525
timestamp 1667941163
transform 1 0 172144 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_1528
timestamp 1667941163
transform 1 0 172480 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_1560
timestamp 1667941163
transform 1 0 176064 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1576
timestamp 1667941163
transform 1 0 177856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1580
timestamp 1667941163
transform 1 0 178304 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1667941163
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_5
timestamp 1667941163
transform 1 0 1904 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_69
timestamp 1667941163
transform 1 0 9072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_73
timestamp 1667941163
transform 1 0 9520 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_77
timestamp 1667941163
transform 1 0 9968 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_79
timestamp 1667941163
transform 1 0 10192 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_86
timestamp 1667941163
transform 1 0 10976 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_117
timestamp 1667941163
transform 1 0 14448 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_121
timestamp 1667941163
transform 1 0 14896 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_129
timestamp 1667941163
transform 1 0 15792 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_133
timestamp 1667941163
transform 1 0 16240 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_139
timestamp 1667941163
transform 1 0 16912 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_144
timestamp 1667941163
transform 1 0 17472 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_162
timestamp 1667941163
transform 1 0 19488 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 19936 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_168
timestamp 1667941163
transform 1 0 20160 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_171
timestamp 1667941163
transform 1 0 20496 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_179
timestamp 1667941163
transform 1 0 21392 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_187
timestamp 1667941163
transform 1 0 22288 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_195
timestamp 1667941163
transform 1 0 23184 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_199
timestamp 1667941163
transform 1 0 23632 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_207
timestamp 1667941163
transform 1 0 24528 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_211
timestamp 1667941163
transform 1 0 24976 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_215
timestamp 1667941163
transform 1 0 25424 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_219
timestamp 1667941163
transform 1 0 25872 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_221
timestamp 1667941163
transform 1 0 26096 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_224
timestamp 1667941163
transform 1 0 26432 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_255
timestamp 1667941163
transform 1 0 29904 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_274
timestamp 1667941163
transform 1 0 32032 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_280
timestamp 1667941163
transform 1 0 32704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_286
timestamp 1667941163
transform 1 0 33376 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_288
timestamp 1667941163
transform 1 0 33600 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_291
timestamp 1667941163
transform 1 0 33936 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_310
timestamp 1667941163
transform 1 0 36064 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_316
timestamp 1667941163
transform 1 0 36736 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_320
timestamp 1667941163
transform 1 0 37184 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_324
timestamp 1667941163
transform 1 0 37632 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_340
timestamp 1667941163
transform 1 0 39424 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_348
timestamp 1667941163
transform 1 0 40320 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_352
timestamp 1667941163
transform 1 0 40768 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1667941163
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1667941163
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_423
timestamp 1667941163
transform 1 0 48720 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1667941163
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_428
timestamp 1667941163
transform 1 0 49280 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_432
timestamp 1667941163
transform 1 0 49728 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_434
timestamp 1667941163
transform 1 0 49952 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_439
timestamp 1667941163
transform 1 0 50512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_443
timestamp 1667941163
transform 1 0 50960 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_448
timestamp 1667941163
transform 1 0 51520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_467
timestamp 1667941163
transform 1 0 53648 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_473
timestamp 1667941163
transform 1 0 54320 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_489
timestamp 1667941163
transform 1 0 56112 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_499
timestamp 1667941163
transform 1 0 57232 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_515
timestamp 1667941163
transform 1 0 59024 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_523
timestamp 1667941163
transform 1 0 59920 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_526
timestamp 1667941163
transform 1 0 60256 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_530
timestamp 1667941163
transform 1 0 60704 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_532
timestamp 1667941163
transform 1 0 60928 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_537
timestamp 1667941163
transform 1 0 61488 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_545
timestamp 1667941163
transform 1 0 62384 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_566
timestamp 1667941163
transform 1 0 64736 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_570
timestamp 1667941163
transform 1 0 65184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_575
timestamp 1667941163
transform 1 0 65744 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_641
timestamp 1667941163
transform 1 0 73136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_659
timestamp 1667941163
transform 1 0 75152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_667
timestamp 1667941163
transform 1 0 76048 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_673
timestamp 1667941163
transform 1 0 76720 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_677
timestamp 1667941163
transform 1 0 77168 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_708
timestamp 1667941163
transform 1 0 80640 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1667941163
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1667941163
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1667941163
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_783
timestamp 1667941163
transform 1 0 89040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_801
timestamp 1667941163
transform 1 0 91056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_805
timestamp 1667941163
transform 1 0 91504 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_808
timestamp 1667941163
transform 1 0 91840 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_812
timestamp 1667941163
transform 1 0 92288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_817
timestamp 1667941163
transform 1 0 92848 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_825
timestamp 1667941163
transform 1 0 93744 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_831
timestamp 1667941163
transform 1 0 94416 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1667941163
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1667941163
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1667941163
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1667941163
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1667941163
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1667941163
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1667941163
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1667941163
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1667941163
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1667941163
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1667941163
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1667941163
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1667941163
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1667941163
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1667941163
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1667941163
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1667941163
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1667941163
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1273
timestamp 1667941163
transform 1 0 143920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1667941163
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1280
timestamp 1667941163
transform 1 0 144704 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1344
timestamp 1667941163
transform 1 0 151872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1348
timestamp 1667941163
transform 1 0 152320 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1351
timestamp 1667941163
transform 1 0 152656 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1415
timestamp 1667941163
transform 1 0 159824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1419
timestamp 1667941163
transform 1 0 160272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1422
timestamp 1667941163
transform 1 0 160608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1486
timestamp 1667941163
transform 1 0 167776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1490
timestamp 1667941163
transform 1 0 168224 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1493
timestamp 1667941163
transform 1 0 168560 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1557
timestamp 1667941163
transform 1 0 175728 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1561
timestamp 1667941163
transform 1 0 176176 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_1564
timestamp 1667941163
transform 1 0 176512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1572
timestamp 1667941163
transform 1 0 177408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1580
timestamp 1667941163
transform 1 0 178304 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1667941163
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_9
timestamp 1667941163
transform 1 0 2352 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_13
timestamp 1667941163
transform 1 0 2800 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_19
timestamp 1667941163
transform 1 0 3472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_27
timestamp 1667941163
transform 1 0 4368 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_33
timestamp 1667941163
transform 1 0 5040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_37
timestamp 1667941163
transform 1 0 5488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_41
timestamp 1667941163
transform 1 0 5936 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_49
timestamp 1667941163
transform 1 0 6832 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_61
timestamp 1667941163
transform 1 0 8176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_69
timestamp 1667941163
transform 1 0 9072 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_72
timestamp 1667941163
transform 1 0 9408 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_102
timestamp 1667941163
transform 1 0 12768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_104
timestamp 1667941163
transform 1 0 12992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_107
timestamp 1667941163
transform 1 0 13328 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_110
timestamp 1667941163
transform 1 0 13664 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_112
timestamp 1667941163
transform 1 0 13888 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_117
timestamp 1667941163
transform 1 0 14448 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_121
timestamp 1667941163
transform 1 0 14896 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_125
timestamp 1667941163
transform 1 0 15344 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_133
timestamp 1667941163
transform 1 0 16240 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 16912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_142
timestamp 1667941163
transform 1 0 17248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_146
timestamp 1667941163
transform 1 0 17696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_156
timestamp 1667941163
transform 1 0 18816 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_162
timestamp 1667941163
transform 1 0 19488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_166
timestamp 1667941163
transform 1 0 19936 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_170
timestamp 1667941163
transform 1 0 20384 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_174
timestamp 1667941163
transform 1 0 20832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_177
timestamp 1667941163
transform 1 0 21168 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_184
timestamp 1667941163
transform 1 0 21952 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_190
timestamp 1667941163
transform 1 0 22624 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 23072 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_196
timestamp 1667941163
transform 1 0 23296 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_201
timestamp 1667941163
transform 1 0 23856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_205
timestamp 1667941163
transform 1 0 24304 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_209
timestamp 1667941163
transform 1 0 24752 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_212
timestamp 1667941163
transform 1 0 25088 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_219
timestamp 1667941163
transform 1 0 25872 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_223
timestamp 1667941163
transform 1 0 26320 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_229
timestamp 1667941163
transform 1 0 26992 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_233
timestamp 1667941163
transform 1 0 27440 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_237
timestamp 1667941163
transform 1 0 27888 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_243
timestamp 1667941163
transform 1 0 28560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1667941163
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_265
timestamp 1667941163
transform 1 0 31024 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_273
timestamp 1667941163
transform 1 0 31920 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_279
timestamp 1667941163
transform 1 0 32592 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_282
timestamp 1667941163
transform 1 0 32928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_284
timestamp 1667941163
transform 1 0 33152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_314
timestamp 1667941163
transform 1 0 36512 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_317
timestamp 1667941163
transform 1 0 36848 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_324
timestamp 1667941163
transform 1 0 37632 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_330
timestamp 1667941163
transform 1 0 38304 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_332
timestamp 1667941163
transform 1 0 38528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_335
timestamp 1667941163
transform 1 0 38864 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_343
timestamp 1667941163
transform 1 0 39760 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_347
timestamp 1667941163
transform 1 0 40208 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_349
timestamp 1667941163
transform 1 0 40432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_352
timestamp 1667941163
transform 1 0 40768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_357
timestamp 1667941163
transform 1 0 41328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_369
timestamp 1667941163
transform 1 0 42672 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_377
timestamp 1667941163
transform 1 0 43568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_381
timestamp 1667941163
transform 1 0 44016 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_384
timestamp 1667941163
transform 1 0 44352 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_387
timestamp 1667941163
transform 1 0 44688 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_394
timestamp 1667941163
transform 1 0 45472 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_400
timestamp 1667941163
transform 1 0 46144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_404
timestamp 1667941163
transform 1 0 46592 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_406
timestamp 1667941163
transform 1 0 46816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_411
timestamp 1667941163
transform 1 0 47376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_415
timestamp 1667941163
transform 1 0 47824 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_419
timestamp 1667941163
transform 1 0 48272 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_422
timestamp 1667941163
transform 1 0 48608 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_424
timestamp 1667941163
transform 1 0 48832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_454
timestamp 1667941163
transform 1 0 52192 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_457
timestamp 1667941163
transform 1 0 52528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_475
timestamp 1667941163
transform 1 0 54544 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_481
timestamp 1667941163
transform 1 0 55216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_489
timestamp 1667941163
transform 1 0 56112 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_492
timestamp 1667941163
transform 1 0 56448 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_497
timestamp 1667941163
transform 1 0 57008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_513
timestamp 1667941163
transform 1 0 58800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_517
timestamp 1667941163
transform 1 0 59248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_523
timestamp 1667941163
transform 1 0 59920 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_527
timestamp 1667941163
transform 1 0 60368 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_529
timestamp 1667941163
transform 1 0 60592 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_559
timestamp 1667941163
transform 1 0 63952 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_562
timestamp 1667941163
transform 1 0 64288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_568
timestamp 1667941163
transform 1 0 64960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_572
timestamp 1667941163
transform 1 0 65408 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_574
timestamp 1667941163
transform 1 0 65632 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_579
timestamp 1667941163
transform 1 0 66192 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_585
timestamp 1667941163
transform 1 0 66864 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_593
timestamp 1667941163
transform 1 0 67760 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_597
timestamp 1667941163
transform 1 0 68208 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_601
timestamp 1667941163
transform 1 0 68656 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_607
timestamp 1667941163
transform 1 0 69328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_615
timestamp 1667941163
transform 1 0 70224 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_621
timestamp 1667941163
transform 1 0 70896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_629
timestamp 1667941163
transform 1 0 71792 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_632
timestamp 1667941163
transform 1 0 72128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_636
timestamp 1667941163
transform 1 0 72576 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_642
timestamp 1667941163
transform 1 0 73248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_648
timestamp 1667941163
transform 1 0 73920 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_654
timestamp 1667941163
transform 1 0 74592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_658
timestamp 1667941163
transform 1 0 75040 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_663
timestamp 1667941163
transform 1 0 75600 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_667
timestamp 1667941163
transform 1 0 76048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_683
timestamp 1667941163
transform 1 0 77840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_691
timestamp 1667941163
transform 1 0 78736 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_699
timestamp 1667941163
transform 1 0 79632 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_702
timestamp 1667941163
transform 1 0 79968 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_707
timestamp 1667941163
transform 1 0 80528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_723
timestamp 1667941163
transform 1 0 82320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_727
timestamp 1667941163
transform 1 0 82768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_733
timestamp 1667941163
transform 1 0 83440 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_737
timestamp 1667941163
transform 1 0 83888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_741
timestamp 1667941163
transform 1 0 84336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_747
timestamp 1667941163
transform 1 0 85008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_763
timestamp 1667941163
transform 1 0 86800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_767
timestamp 1667941163
transform 1 0 87248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_769
timestamp 1667941163
transform 1 0 87472 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_772
timestamp 1667941163
transform 1 0 87808 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_777
timestamp 1667941163
transform 1 0 88368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_781
timestamp 1667941163
transform 1 0 88816 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_783
timestamp 1667941163
transform 1 0 89040 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_788
timestamp 1667941163
transform 1 0 89600 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_794
timestamp 1667941163
transform 1 0 90272 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_800
timestamp 1667941163
transform 1 0 90944 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_804
timestamp 1667941163
transform 1 0 91392 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_807
timestamp 1667941163
transform 1 0 91728 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_837
timestamp 1667941163
transform 1 0 95088 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_839
timestamp 1667941163
transform 1 0 95312 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_842
timestamp 1667941163
transform 1 0 95648 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_850
timestamp 1667941163
transform 1 0 96544 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_854
timestamp 1667941163
transform 1 0 96992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_859
timestamp 1667941163
transform 1 0 97552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_867
timestamp 1667941163
transform 1 0 98448 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_873
timestamp 1667941163
transform 1 0 99120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_877
timestamp 1667941163
transform 1 0 99568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_893
timestamp 1667941163
transform 1 0 101360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_901
timestamp 1667941163
transform 1 0 102256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_909
timestamp 1667941163
transform 1 0 103152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_912
timestamp 1667941163
transform 1 0 103488 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_917
timestamp 1667941163
transform 1 0 104048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_933
timestamp 1667941163
transform 1 0 105840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_937
timestamp 1667941163
transform 1 0 106288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_943
timestamp 1667941163
transform 1 0 106960 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_947
timestamp 1667941163
transform 1 0 107408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_951
timestamp 1667941163
transform 1 0 107856 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_957
timestamp 1667941163
transform 1 0 108528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_973
timestamp 1667941163
transform 1 0 110320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_977
timestamp 1667941163
transform 1 0 110768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_979
timestamp 1667941163
transform 1 0 110992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_982
timestamp 1667941163
transform 1 0 111328 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_987
timestamp 1667941163
transform 1 0 111888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_999
timestamp 1667941163
transform 1 0 113232 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1017
timestamp 1667941163
transform 1 0 115248 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1021
timestamp 1667941163
transform 1 0 115696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1027
timestamp 1667941163
transform 1 0 116368 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1035
timestamp 1667941163
transform 1 0 117264 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1041
timestamp 1667941163
transform 1 0 117936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1049
timestamp 1667941163
transform 1 0 118832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1052
timestamp 1667941163
transform 1 0 119168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1060
timestamp 1667941163
transform 1 0 120064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1064
timestamp 1667941163
transform 1 0 120512 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1069
timestamp 1667941163
transform 1 0 121072 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1077
timestamp 1667941163
transform 1 0 121968 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1083
timestamp 1667941163
transform 1 0 122640 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1087
timestamp 1667941163
transform 1 0 123088 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1103
timestamp 1667941163
transform 1 0 124880 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1111
timestamp 1667941163
transform 1 0 125776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1119
timestamp 1667941163
transform 1 0 126672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1122
timestamp 1667941163
transform 1 0 127008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1127
timestamp 1667941163
transform 1 0 127568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1143
timestamp 1667941163
transform 1 0 129360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1147
timestamp 1667941163
transform 1 0 129808 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1153
timestamp 1667941163
transform 1 0 130480 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1157
timestamp 1667941163
transform 1 0 130928 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1161
timestamp 1667941163
transform 1 0 131376 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1167
timestamp 1667941163
transform 1 0 132048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1183
timestamp 1667941163
transform 1 0 133840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1187
timestamp 1667941163
transform 1 0 134288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1189
timestamp 1667941163
transform 1 0 134512 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1192
timestamp 1667941163
transform 1 0 134848 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1197
timestamp 1667941163
transform 1 0 135408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1209
timestamp 1667941163
transform 1 0 136752 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1227
timestamp 1667941163
transform 1 0 138768 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1231
timestamp 1667941163
transform 1 0 139216 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1237
timestamp 1667941163
transform 1 0 139888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1245
timestamp 1667941163
transform 1 0 140784 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1251
timestamp 1667941163
transform 1 0 141456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1259
timestamp 1667941163
transform 1 0 142352 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1262
timestamp 1667941163
transform 1 0 142688 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1270
timestamp 1667941163
transform 1 0 143584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1274
timestamp 1667941163
transform 1 0 144032 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1279
timestamp 1667941163
transform 1 0 144592 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1287
timestamp 1667941163
transform 1 0 145488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1293
timestamp 1667941163
transform 1 0 146160 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1297
timestamp 1667941163
transform 1 0 146608 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1313
timestamp 1667941163
transform 1 0 148400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1321
timestamp 1667941163
transform 1 0 149296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1329
timestamp 1667941163
transform 1 0 150192 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1332
timestamp 1667941163
transform 1 0 150528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1337
timestamp 1667941163
transform 1 0 151088 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1353
timestamp 1667941163
transform 1 0 152880 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1357
timestamp 1667941163
transform 1 0 153328 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1363
timestamp 1667941163
transform 1 0 154000 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1367
timestamp 1667941163
transform 1 0 154448 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1371
timestamp 1667941163
transform 1 0 154896 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1377
timestamp 1667941163
transform 1 0 155568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1393
timestamp 1667941163
transform 1 0 157360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1397
timestamp 1667941163
transform 1 0 157808 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1399
timestamp 1667941163
transform 1 0 158032 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1402
timestamp 1667941163
transform 1 0 158368 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1407
timestamp 1667941163
transform 1 0 158928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1419
timestamp 1667941163
transform 1 0 160272 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1437
timestamp 1667941163
transform 1 0 162288 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1441
timestamp 1667941163
transform 1 0 162736 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1447
timestamp 1667941163
transform 1 0 163408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1455
timestamp 1667941163
transform 1 0 164304 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1461
timestamp 1667941163
transform 1 0 164976 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1469
timestamp 1667941163
transform 1 0 165872 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1472
timestamp 1667941163
transform 1 0 166208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1480
timestamp 1667941163
transform 1 0 167104 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1484
timestamp 1667941163
transform 1 0 167552 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1489
timestamp 1667941163
transform 1 0 168112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1497
timestamp 1667941163
transform 1 0 169008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1503
timestamp 1667941163
transform 1 0 169680 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1507
timestamp 1667941163
transform 1 0 170128 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1523
timestamp 1667941163
transform 1 0 171920 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1531
timestamp 1667941163
transform 1 0 172816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1539
timestamp 1667941163
transform 1 0 173712 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1542
timestamp 1667941163
transform 1 0 174048 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1547
timestamp 1667941163
transform 1 0 174608 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1563
timestamp 1667941163
transform 1 0 176400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1567
timestamp 1667941163
transform 1 0 176848 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1573
timestamp 1667941163
transform 1 0 177520 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1577
timestamp 1667941163
transform 1 0 177968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 178640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 178640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 178640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 178640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 178640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 178640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 178640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 178640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 178640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 178640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 178640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 178640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 178640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 178640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 178640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 178640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 178640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1667941163
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1667941163
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1667941163
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1667941163
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1667941163
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1667941163
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1667941163
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1667941163
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1667941163
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1667941163
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1667941163
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1667941163
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1667941163
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1667941163
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1667941163
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1667941163
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1667941163
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1667941163
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1667941163
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1667941163
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1667941163
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1667941163
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1667941163
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1667941163
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1667941163
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1667941163
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1667941163
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1667941163
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1667941163
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1667941163
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1667941163
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1667941163
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1667941163
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1667941163
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1667941163
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1667941163
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1667941163
transform 1 0 150304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1667941163
transform 1 0 154224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1667941163
transform 1 0 158144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1667941163
transform 1 0 162064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1667941163
transform 1 0 165984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1667941163
transform 1 0 169904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1667941163
transform 1 0 173824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1667941163
transform 1 0 177744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1667941163
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_81
timestamp 1667941163
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_82
timestamp 1667941163
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_83
timestamp 1667941163
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1667941163
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1667941163
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1667941163
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1667941163
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1667941163
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1667941163
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1667941163
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1667941163
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1667941163
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1667941163
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1667941163
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1667941163
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1667941163
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1667941163
transform 1 0 152432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1667941163
transform 1 0 160384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1667941163
transform 1 0 168336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1667941163
transform 1 0 176288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1667941163
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1667941163
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1667941163
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1667941163
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1667941163
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1667941163
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1667941163
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1667941163
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1667941163
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1667941163
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1667941163
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1667941163
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1667941163
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1667941163
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1667941163
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1667941163
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1667941163
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1667941163
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1667941163
transform 1 0 148400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1667941163
transform 1 0 156352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1667941163
transform 1 0 164304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1667941163
transform 1 0 172256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1667941163
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1667941163
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1667941163
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1667941163
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1667941163
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1667941163
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1667941163
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1667941163
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1667941163
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1667941163
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1667941163
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1667941163
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1667941163
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1667941163
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1667941163
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1667941163
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1667941163
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1667941163
transform 1 0 152432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1667941163
transform 1 0 160384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1667941163
transform 1 0 168336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1667941163
transform 1 0 176288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1667941163
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1667941163
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1667941163
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1667941163
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1667941163
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1667941163
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1667941163
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1667941163
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1667941163
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1667941163
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1667941163
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1667941163
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1667941163
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1667941163
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1667941163
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1667941163
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1667941163
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1667941163
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 148400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 156352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 164304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 172256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 152432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 160384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 168336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 176288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 148400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 156352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 164304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 172256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 152432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 160384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 168336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 176288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 148400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 156352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 164304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 172256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 152432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 160384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 168336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 176288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1667941163
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1667941163
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1667941163
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1667941163
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1667941163
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1667941163
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1667941163
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1667941163
transform 1 0 148400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1667941163
transform 1 0 156352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1667941163
transform 1 0 164304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1667941163
transform 1 0 172256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1667941163
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1667941163
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1667941163
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1667941163
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1667941163
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1667941163
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1667941163
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1667941163
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1667941163
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1667941163
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1667941163
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1667941163
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1667941163
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1667941163
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1667941163
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1667941163
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1667941163
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1667941163
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1667941163
transform 1 0 152432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1667941163
transform 1 0 160384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1667941163
transform 1 0 168336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1667941163
transform 1 0 176288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1667941163
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1667941163
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1667941163
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1667941163
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1667941163
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1667941163
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1667941163
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1667941163
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1667941163
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1667941163
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1667941163
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1667941163
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1667941163
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1667941163
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1667941163
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1667941163
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1667941163
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1667941163
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1667941163
transform 1 0 148400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1667941163
transform 1 0 156352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1667941163
transform 1 0 164304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1667941163
transform 1 0 172256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1667941163
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1667941163
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1667941163
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1667941163
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1667941163
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1667941163
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1667941163
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1667941163
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1667941163
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1667941163
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1667941163
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1667941163
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1667941163
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1667941163
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1667941163
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1667941163
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1667941163
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1667941163
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1667941163
transform 1 0 152432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1667941163
transform 1 0 160384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1667941163
transform 1 0 168336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1667941163
transform 1 0 176288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1667941163
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1667941163
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1667941163
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1667941163
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1667941163
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1667941163
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1667941163
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1667941163
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1667941163
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1667941163
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1667941163
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1667941163
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1667941163
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1667941163
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1667941163
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1667941163
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1667941163
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1667941163
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1667941163
transform 1 0 148400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1667941163
transform 1 0 156352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1667941163
transform 1 0 164304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1667941163
transform 1 0 172256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1667941163
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1667941163
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1667941163
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1667941163
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1667941163
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1667941163
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1667941163
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1667941163
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1667941163
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1667941163
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1667941163
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1667941163
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1667941163
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1667941163
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1667941163
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1667941163
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1667941163
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1667941163
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1667941163
transform 1 0 152432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1667941163
transform 1 0 160384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1667941163
transform 1 0 168336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1667941163
transform 1 0 176288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1667941163
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1667941163
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1667941163
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1667941163
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1667941163
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1667941163
transform 1 0 24864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1667941163
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1667941163
transform 1 0 32704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1667941163
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1667941163
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1667941163
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1667941163
transform 1 0 48384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1667941163
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1667941163
transform 1 0 56224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1667941163
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1667941163
transform 1 0 64064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1667941163
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1667941163
transform 1 0 71904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1667941163
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1667941163
transform 1 0 79744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1667941163
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1667941163
transform 1 0 87584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1667941163
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1667941163
transform 1 0 95424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1667941163
transform 1 0 99344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1667941163
transform 1 0 103264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1667941163
transform 1 0 107184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1667941163
transform 1 0 111104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1667941163
transform 1 0 115024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1667941163
transform 1 0 118944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1667941163
transform 1 0 122864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1667941163
transform 1 0 126784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1667941163
transform 1 0 130704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1667941163
transform 1 0 134624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1667941163
transform 1 0 138544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1667941163
transform 1 0 142464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1667941163
transform 1 0 146384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1667941163
transform 1 0 150304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1667941163
transform 1 0 154224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1667941163
transform 1 0 158144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1667941163
transform 1 0 162064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1667941163
transform 1 0 165984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1667941163
transform 1 0 169904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1667941163
transform 1 0 173824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1667941163
transform 1 0 177744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _030_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 16464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _031_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 25536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _032_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 27328 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _033_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 9520 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _034_
timestamp 1667941163
transform 1 0 11200 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _035_
timestamp 1667941163
transform 1 0 26656 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _036_
timestamp 1667941163
transform 1 0 33264 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _037_
timestamp 1667941163
transform 1 0 48944 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _038_
timestamp 1667941163
transform 1 0 60704 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _039_
timestamp 1667941163
transform -1 0 80640 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _040_
timestamp 1667941163
transform 1 0 91840 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _242_
timestamp 1667941163
transform 1 0 94304 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _243_
timestamp 1667941163
transform 1 0 95424 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout11 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 21504 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout12
timestamp 1667941163
transform 1 0 21728 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  fanout13 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 21728 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout14 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 17920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1680 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1667941163
transform 1 0 6160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1667941163
transform 1 0 10304 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1667941163
transform 1 0 15568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1667941163
transform 1 0 21280 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1667941163
transform 1 0 25200 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1667941163
transform 1 0 31248 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1667941163
transform 1 0 36960 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1667941163
transform 1 0 39088 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1667941163
transform 1 0 44800 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[0\].pdn_15 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 61824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[0\].pdn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 61712 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[0\].pdp_16
timestamp 1667941163
transform -1 0 41888 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[0\].pdp
timestamp 1667941163
transform -1 0 40320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[1\].pdn_17
timestamp 1667941163
transform -1 0 62048 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[1\].pdn
timestamp 1667941163
transform -1 0 60480 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[1\].pdp
timestamp 1667941163
transform -1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[1\].pdp_18
timestamp 1667941163
transform -1 0 41888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[2\].pdn
timestamp 1667941163
transform 1 0 62944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[2\].pdn_19
timestamp 1667941163
transform 1 0 62048 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[2\].pdp
timestamp 1667941163
transform -1 0 39648 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[2\].pdp_20
timestamp 1667941163
transform -1 0 40992 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[3\].pdn_21
timestamp 1667941163
transform -1 0 62384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[3\].pdn
timestamp 1667941163
transform -1 0 62160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[3\].pdp
timestamp 1667941163
transform 1 0 40656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[3\].pdp_22
timestamp 1667941163
transform 1 0 39984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[4\].pdn_23
timestamp 1667941163
transform -1 0 62720 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[4\].pdn
timestamp 1667941163
transform -1 0 60816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[4\].pdp_24
timestamp 1667941163
transform -1 0 40208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[4\].pdp
timestamp 1667941163
transform -1 0 39536 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[5\].pdn
timestamp 1667941163
transform 1 0 61488 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[5\].pdn_25
timestamp 1667941163
transform 1 0 60704 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[5\].pdp_26
timestamp 1667941163
transform -1 0 43008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[5\].pdp
timestamp 1667941163
transform -1 0 40768 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[6\].pdn_27
timestamp 1667941163
transform -1 0 63504 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[6\].pdn
timestamp 1667941163
transform -1 0 63280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[6\].pdp_28
timestamp 1667941163
transform -1 0 40880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[6\].pdp
timestamp 1667941163
transform -1 0 40768 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[7\].pdn_29
timestamp 1667941163
transform -1 0 64176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[7\].pdn
timestamp 1667941163
transform -1 0 63952 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[7\].pdp
timestamp 1667941163
transform 1 0 41888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[7\].pdp_30
timestamp 1667941163
transform 1 0 41216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[0\].pun pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 21616 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[0\].pup
timestamp 1667941163
transform 1 0 22400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[1\].pun
timestamp 1667941163
transform 1 0 19936 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[1\].pup
timestamp 1667941163
transform 1 0 18032 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[2\].pun
timestamp 1667941163
transform 1 0 20720 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[2\].pup
timestamp 1667941163
transform 1 0 21504 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[3\].pun
timestamp 1667941163
transform 1 0 23408 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[3\].pup
timestamp 1667941163
transform 1 0 20384 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[4\].pun
timestamp 1667941163
transform 1 0 21616 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[4\].pup
timestamp 1667941163
transform 1 0 20720 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[5\].pun
timestamp 1667941163
transform 1 0 24640 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[5\].pup
timestamp 1667941163
transform -1 0 22400 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[6\].pun
timestamp 1667941163
transform 1 0 22512 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[6\].pup
timestamp 1667941163
transform 1 0 16464 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[7\].pun
timestamp 1667941163
transform 1 0 22512 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[7\].pup
timestamp 1667941163
transform 1 0 24304 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[8\].pun
timestamp 1667941163
transform 1 0 20832 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[8\].pup
timestamp 1667941163
transform 1 0 19488 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[9\].pun
timestamp 1667941163
transform 1 0 22512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[9\].pup
timestamp 1667941163
transform -1 0 20496 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[10\].pun
timestamp 1667941163
transform 1 0 21616 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[10\].pup
timestamp 1667941163
transform 1 0 20720 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[11\].pun
timestamp 1667941163
transform 1 0 18592 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[11\].pup
timestamp 1667941163
transform -1 0 19600 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[12\].pun
timestamp 1667941163
transform 1 0 19824 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[12\].pup
timestamp 1667941163
transform -1 0 21504 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[13\].pun
timestamp 1667941163
transform 1 0 23072 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[13\].pup
timestamp 1667941163
transform 1 0 19040 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[14\].pun
timestamp 1667941163
transform 1 0 19488 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[14\].pup
timestamp 1667941163
transform 1 0 20384 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[15\].pun
timestamp 1667941163
transform 1 0 22512 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[15\].pup
timestamp 1667941163
transform 1 0 18592 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[16\].pun
timestamp 1667941163
transform 1 0 23408 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[16\].pup
timestamp 1667941163
transform 1 0 20384 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[17\].pun
timestamp 1667941163
transform 1 0 20384 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[17\].pup
timestamp 1667941163
transform 1 0 18928 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[18\].pun
timestamp 1667941163
transform 1 0 21616 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[18\].pup
timestamp 1667941163
transform 1 0 17696 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ntrimn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 52640 0 1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[0\].ntrimn_31
timestamp 1667941163
transform 1 0 53424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[0\].ntrimp_32
timestamp 1667941163
transform -1 0 54320 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ntrimp
timestamp 1667941163
transform 1 0 51744 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ptrimn
timestamp 1667941163
transform 1 0 17136 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ptrimp
timestamp 1667941163
transform 1 0 17584 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[1\].ntrimn_33
timestamp 1667941163
transform -1 0 64960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ntrimn
timestamp 1667941163
transform 1 0 62832 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[1\].ntrimp_34
timestamp 1667941163
transform -1 0 65744 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ntrimp
timestamp 1667941163
transform 1 0 62832 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ptrimn
timestamp 1667941163
transform 1 0 15008 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ptrimp
timestamp 1667941163
transform 1 0 16240 0 1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[2\].ntrimn_35
timestamp 1667941163
transform 1 0 73472 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ntrimn
timestamp 1667941163
transform 1 0 72352 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[2\].ntrimp_36
timestamp 1667941163
transform 1 0 74144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ntrimp
timestamp 1667941163
transform 1 0 73248 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ptrimn
timestamp 1667941163
transform -1 0 31024 0 1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ptrimp
timestamp 1667941163
transform 1 0 30128 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[3\].ntrimn_37
timestamp 1667941163
transform 1 0 89824 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ntrimn
timestamp 1667941163
transform 1 0 89152 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[3\].ntrimp_38
timestamp 1667941163
transform -1 0 90944 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ntrimp
timestamp 1667941163
transform 1 0 88032 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ptrimn
timestamp 1667941163
transform -1 0 36064 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ptrimp
timestamp 1667941163
transform -1 0 36064 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.nsijn
timestamp 1667941163
transform -1 0 26768 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_inj.nsijp_214 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 52752 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.nsijp
timestamp 1667941163
transform -1 0 52640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_inj.psijn_215
timestamp 1667941163
transform -1 0 53760 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.psijn
timestamp 1667941163
transform -1 0 52080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.psijp
timestamp 1667941163
transform -1 0 26656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.siginv_39
timestamp 1667941163
transform -1 0 28000 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  u_inj.siginv pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 26096 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_40
timestamp 1667941163
transform -1 0 66416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_41
timestamp 1667941163
transform -1 0 68768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_42
timestamp 1667941163
transform -1 0 69776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_43
timestamp 1667941163
transform -1 0 71456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_44
timestamp 1667941163
transform -1 0 73136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_45
timestamp 1667941163
transform -1 0 74816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_46
timestamp 1667941163
transform -1 0 76608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_47
timestamp 1667941163
transform -1 0 78176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_48
timestamp 1667941163
transform -1 0 80528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_49
timestamp 1667941163
transform -1 0 81536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_50
timestamp 1667941163
transform -1 0 83216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_51
timestamp 1667941163
transform -1 0 84896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_52
timestamp 1667941163
transform -1 0 86576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_53
timestamp 1667941163
transform -1 0 88368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_54
timestamp 1667941163
transform -1 0 89936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_55
timestamp 1667941163
transform -1 0 92288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_56
timestamp 1667941163
transform -1 0 93296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_57
timestamp 1667941163
transform -1 0 94976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_58
timestamp 1667941163
transform -1 0 96656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_59
timestamp 1667941163
transform -1 0 98336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_60
timestamp 1667941163
transform -1 0 100128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_61
timestamp 1667941163
transform -1 0 101696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_62
timestamp 1667941163
transform -1 0 104048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_63
timestamp 1667941163
transform -1 0 105056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_64
timestamp 1667941163
transform -1 0 106736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_65
timestamp 1667941163
transform -1 0 108416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_66
timestamp 1667941163
transform -1 0 110096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_67
timestamp 1667941163
transform -1 0 111888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_68
timestamp 1667941163
transform -1 0 113456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_69
timestamp 1667941163
transform -1 0 115808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_70
timestamp 1667941163
transform -1 0 116816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_71
timestamp 1667941163
transform -1 0 118496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_72
timestamp 1667941163
transform -1 0 123648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_73
timestamp 1667941163
transform -1 0 125216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_74
timestamp 1667941163
transform -1 0 127568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_75
timestamp 1667941163
transform -1 0 128576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_76
timestamp 1667941163
transform -1 0 130256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_77
timestamp 1667941163
transform -1 0 131936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_78
timestamp 1667941163
transform -1 0 133616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_79
timestamp 1667941163
transform -1 0 135408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_80
timestamp 1667941163
transform -1 0 136976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_81
timestamp 1667941163
transform -1 0 139328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_82
timestamp 1667941163
transform -1 0 140336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_83
timestamp 1667941163
transform -1 0 142016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_84
timestamp 1667941163
transform -1 0 143696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_85
timestamp 1667941163
transform -1 0 145376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_86
timestamp 1667941163
transform -1 0 147168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_87
timestamp 1667941163
transform -1 0 148736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_88
timestamp 1667941163
transform -1 0 151088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_89
timestamp 1667941163
transform -1 0 152096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_90
timestamp 1667941163
transform -1 0 153776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_91
timestamp 1667941163
transform -1 0 155456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_92
timestamp 1667941163
transform -1 0 157136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_93
timestamp 1667941163
transform -1 0 158928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_94
timestamp 1667941163
transform -1 0 160496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_95
timestamp 1667941163
transform -1 0 162848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_96
timestamp 1667941163
transform -1 0 163856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_97
timestamp 1667941163
transform -1 0 165536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_98
timestamp 1667941163
transform -1 0 167216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_99
timestamp 1667941163
transform -1 0 168896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_100
timestamp 1667941163
transform -1 0 170688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_101
timestamp 1667941163
transform -1 0 172256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_102
timestamp 1667941163
transform -1 0 173376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_103
timestamp 1667941163
transform -1 0 174608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_104
timestamp 1667941163
transform -1 0 175280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_105
timestamp 1667941163
transform -1 0 5040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_106
timestamp 1667941163
transform 1 0 8624 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_107
timestamp 1667941163
transform -1 0 14448 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_108
timestamp 1667941163
transform -1 0 19488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_109
timestamp 1667941163
transform -1 0 23856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_110
timestamp 1667941163
transform -1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_111
timestamp 1667941163
transform 1 0 32144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_112
timestamp 1667941163
transform -1 0 38304 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_113
timestamp 1667941163
transform -1 0 42672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_114
timestamp 1667941163
transform -1 0 47376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_115
timestamp 1667941163
transform 1 0 51072 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_116
timestamp 1667941163
transform -1 0 57008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_117
timestamp 1667941163
transform -1 0 61488 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_118
timestamp 1667941163
transform -1 0 66192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_119
timestamp 1667941163
transform -1 0 70896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_120
timestamp 1667941163
transform -1 0 75600 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_121
timestamp 1667941163
transform -1 0 80528 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_122
timestamp 1667941163
transform -1 0 85008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_123
timestamp 1667941163
transform -1 0 89600 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_124
timestamp 1667941163
transform -1 0 94416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_125
timestamp 1667941163
transform -1 0 99120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_126
timestamp 1667941163
transform -1 0 104048 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_127
timestamp 1667941163
transform -1 0 108528 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_128
timestamp 1667941163
transform -1 0 113232 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_129
timestamp 1667941163
transform -1 0 117936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_130
timestamp 1667941163
transform -1 0 122640 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_131
timestamp 1667941163
transform -1 0 127568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_132
timestamp 1667941163
transform -1 0 132048 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_133
timestamp 1667941163
transform -1 0 136752 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_134
timestamp 1667941163
transform -1 0 141456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_135
timestamp 1667941163
transform -1 0 146160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_136
timestamp 1667941163
transform -1 0 151088 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_137
timestamp 1667941163
transform -1 0 155568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_138
timestamp 1667941163
transform -1 0 160272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_139
timestamp 1667941163
transform -1 0 164976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_140
timestamp 1667941163
transform -1 0 169680 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_141
timestamp 1667941163
transform -1 0 174608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_142
timestamp 1667941163
transform 1 0 177856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_143
timestamp 1667941163
transform -1 0 3472 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_144
timestamp 1667941163
transform -1 0 8176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_145
timestamp 1667941163
transform -1 0 12880 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_146
timestamp 1667941163
transform 1 0 16464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_147
timestamp 1667941163
transform -1 0 22624 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_148
timestamp 1667941163
transform -1 0 26992 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_149
timestamp 1667941163
transform -1 0 32704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_150
timestamp 1667941163
transform -1 0 36736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_151
timestamp 1667941163
transform -1 0 41328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_152
timestamp 1667941163
transform -1 0 46144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_153
timestamp 1667941163
transform -1 0 50512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_154
timestamp 1667941163
transform -1 0 55216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_155
timestamp 1667941163
transform -1 0 59920 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_156
timestamp 1667941163
transform -1 0 66864 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_157
timestamp 1667941163
transform -1 0 69328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_158
timestamp 1667941163
transform 1 0 72800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_159
timestamp 1667941163
transform -1 0 78736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_160
timestamp 1667941163
transform -1 0 83440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_161
timestamp 1667941163
transform -1 0 88368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_162
timestamp 1667941163
transform -1 0 92848 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_163
timestamp 1667941163
transform -1 0 97552 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_164
timestamp 1667941163
transform -1 0 102256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_165
timestamp 1667941163
transform -1 0 106960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_166
timestamp 1667941163
transform -1 0 111888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_167
timestamp 1667941163
transform -1 0 116368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_168
timestamp 1667941163
transform -1 0 121072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_169
timestamp 1667941163
transform -1 0 125776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_170
timestamp 1667941163
transform -1 0 130480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_171
timestamp 1667941163
transform -1 0 135408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_172
timestamp 1667941163
transform -1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_173
timestamp 1667941163
transform -1 0 144592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_174
timestamp 1667941163
transform -1 0 149296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_175
timestamp 1667941163
transform -1 0 154000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_176
timestamp 1667941163
transform -1 0 158928 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_177
timestamp 1667941163
transform -1 0 163408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_178
timestamp 1667941163
transform -1 0 168112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_179
timestamp 1667941163
transform -1 0 172816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_180
timestamp 1667941163
transform -1 0 177520 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_181
timestamp 1667941163
transform -1 0 7616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_182
timestamp 1667941163
transform -1 0 10976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_183
timestamp 1667941163
transform -1 0 13888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_184
timestamp 1667941163
transform -1 0 15456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_185
timestamp 1667941163
transform -1 0 17808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_186
timestamp 1667941163
transform -1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_187
timestamp 1667941163
transform -1 0 21728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_188
timestamp 1667941163
transform -1 0 23296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_189
timestamp 1667941163
transform -1 0 25648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_190
timestamp 1667941163
transform -1 0 26656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_191
timestamp 1667941163
transform -1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_192
timestamp 1667941163
transform -1 0 30016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_193
timestamp 1667941163
transform -1 0 31696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_194
timestamp 1667941163
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_195
timestamp 1667941163
transform -1 0 35056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_196
timestamp 1667941163
transform -1 0 37408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_197
timestamp 1667941163
transform -1 0 38416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_198
timestamp 1667941163
transform -1 0 40096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_199
timestamp 1667941163
transform -1 0 41776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_200
timestamp 1667941163
transform -1 0 43456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_201
timestamp 1667941163
transform -1 0 45248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_202
timestamp 1667941163
transform -1 0 46816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_203
timestamp 1667941163
transform -1 0 49168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_204
timestamp 1667941163
transform -1 0 50176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_205
timestamp 1667941163
transform -1 0 51856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_206
timestamp 1667941163
transform -1 0 53536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_207
timestamp 1667941163
transform -1 0 55216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_208
timestamp 1667941163
transform -1 0 57008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_209
timestamp 1667941163
transform -1 0 58576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_210
timestamp 1667941163
transform -1 0 60928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_211
timestamp 1667941163
transform -1 0 61936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_212
timestamp 1667941163
transform -1 0 63616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_213
timestamp 1667941163
transform -1 0 65296 0 1 3136
box -86 -86 534 870
<< labels >>
flabel metal2 s 1344 19200 1456 20000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 48384 19200 48496 20000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 53088 19200 53200 20000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 57792 19200 57904 20000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 62496 19200 62608 20000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 67200 19200 67312 20000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 71904 19200 72016 20000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 76608 19200 76720 20000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 81312 19200 81424 20000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 86016 19200 86128 20000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 90720 19200 90832 20000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 6048 19200 6160 20000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 95424 19200 95536 20000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 100128 19200 100240 20000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 104832 19200 104944 20000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 109536 19200 109648 20000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 114240 19200 114352 20000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 118944 19200 119056 20000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 123648 19200 123760 20000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 128352 19200 128464 20000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 133056 19200 133168 20000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 137760 19200 137872 20000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 10752 19200 10864 20000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 142464 19200 142576 20000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 147168 19200 147280 20000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 151872 19200 151984 20000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 156576 19200 156688 20000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 161280 19200 161392 20000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 165984 19200 166096 20000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 170688 19200 170800 20000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 175392 19200 175504 20000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 15456 19200 15568 20000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 20160 19200 20272 20000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 24864 19200 24976 20000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 29568 19200 29680 20000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 34272 19200 34384 20000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 38976 19200 39088 20000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 43680 19200 43792 20000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 2912 19200 3024 20000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 49952 19200 50064 20000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 54656 19200 54768 20000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 59360 19200 59472 20000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 64064 19200 64176 20000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 68768 19200 68880 20000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 73472 19200 73584 20000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 78176 19200 78288 20000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 82880 19200 82992 20000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 87584 19200 87696 20000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 92288 19200 92400 20000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 7616 19200 7728 20000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 96992 19200 97104 20000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 101696 19200 101808 20000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 106400 19200 106512 20000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 111104 19200 111216 20000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 115808 19200 115920 20000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 120512 19200 120624 20000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 125216 19200 125328 20000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 129920 19200 130032 20000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 134624 19200 134736 20000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 139328 19200 139440 20000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 12320 19200 12432 20000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 144032 19200 144144 20000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 148736 19200 148848 20000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 153440 19200 153552 20000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 158144 19200 158256 20000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 162848 19200 162960 20000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 167552 19200 167664 20000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 172256 19200 172368 20000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 176960 19200 177072 20000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 17024 19200 17136 20000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 21728 19200 21840 20000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 26432 19200 26544 20000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 31136 19200 31248 20000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 35840 19200 35952 20000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 40544 19200 40656 20000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 45248 19200 45360 20000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4480 19200 4592 20000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 51520 19200 51632 20000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 56224 19200 56336 20000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 60928 19200 61040 20000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 65632 19200 65744 20000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 70336 19200 70448 20000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 75040 19200 75152 20000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 79744 19200 79856 20000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 84448 19200 84560 20000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 89152 19200 89264 20000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 93856 19200 93968 20000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 9184 19200 9296 20000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 98560 19200 98672 20000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 103264 19200 103376 20000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 107968 19200 108080 20000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 112672 19200 112784 20000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 117376 19200 117488 20000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 122080 19200 122192 20000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 126784 19200 126896 20000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 131488 19200 131600 20000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 136192 19200 136304 20000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 140896 19200 141008 20000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 13888 19200 14000 20000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 145600 19200 145712 20000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 150304 19200 150416 20000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 155008 19200 155120 20000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 159712 19200 159824 20000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 164416 19200 164528 20000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 169120 19200 169232 20000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 173824 19200 173936 20000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 178528 19200 178640 20000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 18592 19200 18704 20000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 23296 19200 23408 20000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 28000 19200 28112 20000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 32704 19200 32816 20000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 37408 19200 37520 20000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 42112 19200 42224 20000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 46816 19200 46928 20000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 172816 0 172928 800 0 FreeSans 448 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 173376 0 173488 800 0 FreeSans 448 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 173936 0 174048 800 0 FreeSans 448 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 65296 0 65408 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 82096 0 82208 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 118 nsew signal input
flabel metal2 s 83776 0 83888 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 119 nsew signal input
flabel metal2 s 85456 0 85568 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 120 nsew signal input
flabel metal2 s 87136 0 87248 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 121 nsew signal input
flabel metal2 s 88816 0 88928 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 122 nsew signal input
flabel metal2 s 90496 0 90608 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 123 nsew signal input
flabel metal2 s 92176 0 92288 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 124 nsew signal input
flabel metal2 s 93856 0 93968 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 125 nsew signal input
flabel metal2 s 95536 0 95648 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 126 nsew signal input
flabel metal2 s 97216 0 97328 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 127 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 128 nsew signal input
flabel metal2 s 98896 0 99008 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 129 nsew signal input
flabel metal2 s 100576 0 100688 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 130 nsew signal input
flabel metal2 s 102256 0 102368 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 131 nsew signal input
flabel metal2 s 103936 0 104048 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 132 nsew signal input
flabel metal2 s 105616 0 105728 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 133 nsew signal input
flabel metal2 s 107296 0 107408 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 134 nsew signal input
flabel metal2 s 108976 0 109088 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 135 nsew signal input
flabel metal2 s 110656 0 110768 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 136 nsew signal input
flabel metal2 s 112336 0 112448 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 137 nsew signal input
flabel metal2 s 114016 0 114128 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 138 nsew signal input
flabel metal2 s 68656 0 68768 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 139 nsew signal input
flabel metal2 s 115696 0 115808 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 140 nsew signal input
flabel metal2 s 117376 0 117488 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 141 nsew signal input
flabel metal2 s 119056 0 119168 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 142 nsew signal input
flabel metal2 s 120736 0 120848 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 143 nsew signal input
flabel metal2 s 122416 0 122528 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 144 nsew signal input
flabel metal2 s 124096 0 124208 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 145 nsew signal input
flabel metal2 s 125776 0 125888 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 146 nsew signal input
flabel metal2 s 127456 0 127568 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 147 nsew signal input
flabel metal2 s 129136 0 129248 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 148 nsew signal input
flabel metal2 s 130816 0 130928 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 149 nsew signal input
flabel metal2 s 70336 0 70448 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 150 nsew signal input
flabel metal2 s 132496 0 132608 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 151 nsew signal input
flabel metal2 s 134176 0 134288 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 152 nsew signal input
flabel metal2 s 135856 0 135968 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 153 nsew signal input
flabel metal2 s 137536 0 137648 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 154 nsew signal input
flabel metal2 s 139216 0 139328 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 155 nsew signal input
flabel metal2 s 140896 0 141008 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 156 nsew signal input
flabel metal2 s 142576 0 142688 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 157 nsew signal input
flabel metal2 s 144256 0 144368 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 158 nsew signal input
flabel metal2 s 145936 0 146048 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 159 nsew signal input
flabel metal2 s 147616 0 147728 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 160 nsew signal input
flabel metal2 s 72016 0 72128 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 161 nsew signal input
flabel metal2 s 149296 0 149408 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 162 nsew signal input
flabel metal2 s 150976 0 151088 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 163 nsew signal input
flabel metal2 s 152656 0 152768 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 164 nsew signal input
flabel metal2 s 154336 0 154448 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 165 nsew signal input
flabel metal2 s 156016 0 156128 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 166 nsew signal input
flabel metal2 s 157696 0 157808 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 167 nsew signal input
flabel metal2 s 159376 0 159488 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 168 nsew signal input
flabel metal2 s 161056 0 161168 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 169 nsew signal input
flabel metal2 s 162736 0 162848 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 170 nsew signal input
flabel metal2 s 164416 0 164528 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 171 nsew signal input
flabel metal2 s 73696 0 73808 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 172 nsew signal input
flabel metal2 s 166096 0 166208 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 173 nsew signal input
flabel metal2 s 167776 0 167888 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 174 nsew signal input
flabel metal2 s 169456 0 169568 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 175 nsew signal input
flabel metal2 s 171136 0 171248 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 176 nsew signal input
flabel metal2 s 75376 0 75488 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 177 nsew signal input
flabel metal2 s 77056 0 77168 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 178 nsew signal input
flabel metal2 s 78736 0 78848 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 179 nsew signal input
flabel metal2 s 80416 0 80528 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 180 nsew signal input
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_out[0]
port 181 nsew signal tristate
flabel metal2 s 82656 0 82768 800 0 FreeSans 448 90 0 0 la_data_out[10]
port 182 nsew signal tristate
flabel metal2 s 84336 0 84448 800 0 FreeSans 448 90 0 0 la_data_out[11]
port 183 nsew signal tristate
flabel metal2 s 86016 0 86128 800 0 FreeSans 448 90 0 0 la_data_out[12]
port 184 nsew signal tristate
flabel metal2 s 87696 0 87808 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 185 nsew signal tristate
flabel metal2 s 89376 0 89488 800 0 FreeSans 448 90 0 0 la_data_out[14]
port 186 nsew signal tristate
flabel metal2 s 91056 0 91168 800 0 FreeSans 448 90 0 0 la_data_out[15]
port 187 nsew signal tristate
flabel metal2 s 92736 0 92848 800 0 FreeSans 448 90 0 0 la_data_out[16]
port 188 nsew signal tristate
flabel metal2 s 94416 0 94528 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 189 nsew signal tristate
flabel metal2 s 96096 0 96208 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 190 nsew signal tristate
flabel metal2 s 97776 0 97888 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 191 nsew signal tristate
flabel metal2 s 67536 0 67648 800 0 FreeSans 448 90 0 0 la_data_out[1]
port 192 nsew signal tristate
flabel metal2 s 99456 0 99568 800 0 FreeSans 448 90 0 0 la_data_out[20]
port 193 nsew signal tristate
flabel metal2 s 101136 0 101248 800 0 FreeSans 448 90 0 0 la_data_out[21]
port 194 nsew signal tristate
flabel metal2 s 102816 0 102928 800 0 FreeSans 448 90 0 0 la_data_out[22]
port 195 nsew signal tristate
flabel metal2 s 104496 0 104608 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 196 nsew signal tristate
flabel metal2 s 106176 0 106288 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 197 nsew signal tristate
flabel metal2 s 107856 0 107968 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 198 nsew signal tristate
flabel metal2 s 109536 0 109648 800 0 FreeSans 448 90 0 0 la_data_out[26]
port 199 nsew signal tristate
flabel metal2 s 111216 0 111328 800 0 FreeSans 448 90 0 0 la_data_out[27]
port 200 nsew signal tristate
flabel metal2 s 112896 0 113008 800 0 FreeSans 448 90 0 0 la_data_out[28]
port 201 nsew signal tristate
flabel metal2 s 114576 0 114688 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 202 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_out[2]
port 203 nsew signal tristate
flabel metal2 s 116256 0 116368 800 0 FreeSans 448 90 0 0 la_data_out[30]
port 204 nsew signal tristate
flabel metal2 s 117936 0 118048 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 205 nsew signal tristate
flabel metal2 s 119616 0 119728 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 206 nsew signal tristate
flabel metal2 s 121296 0 121408 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 207 nsew signal tristate
flabel metal2 s 122976 0 123088 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 208 nsew signal tristate
flabel metal2 s 124656 0 124768 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 209 nsew signal tristate
flabel metal2 s 126336 0 126448 800 0 FreeSans 448 90 0 0 la_data_out[36]
port 210 nsew signal tristate
flabel metal2 s 128016 0 128128 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 211 nsew signal tristate
flabel metal2 s 129696 0 129808 800 0 FreeSans 448 90 0 0 la_data_out[38]
port 212 nsew signal tristate
flabel metal2 s 131376 0 131488 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 213 nsew signal tristate
flabel metal2 s 70896 0 71008 800 0 FreeSans 448 90 0 0 la_data_out[3]
port 214 nsew signal tristate
flabel metal2 s 133056 0 133168 800 0 FreeSans 448 90 0 0 la_data_out[40]
port 215 nsew signal tristate
flabel metal2 s 134736 0 134848 800 0 FreeSans 448 90 0 0 la_data_out[41]
port 216 nsew signal tristate
flabel metal2 s 136416 0 136528 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 217 nsew signal tristate
flabel metal2 s 138096 0 138208 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 218 nsew signal tristate
flabel metal2 s 139776 0 139888 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 219 nsew signal tristate
flabel metal2 s 141456 0 141568 800 0 FreeSans 448 90 0 0 la_data_out[45]
port 220 nsew signal tristate
flabel metal2 s 143136 0 143248 800 0 FreeSans 448 90 0 0 la_data_out[46]
port 221 nsew signal tristate
flabel metal2 s 144816 0 144928 800 0 FreeSans 448 90 0 0 la_data_out[47]
port 222 nsew signal tristate
flabel metal2 s 146496 0 146608 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 223 nsew signal tristate
flabel metal2 s 148176 0 148288 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 224 nsew signal tristate
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_out[4]
port 225 nsew signal tristate
flabel metal2 s 149856 0 149968 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 226 nsew signal tristate
flabel metal2 s 151536 0 151648 800 0 FreeSans 448 90 0 0 la_data_out[51]
port 227 nsew signal tristate
flabel metal2 s 153216 0 153328 800 0 FreeSans 448 90 0 0 la_data_out[52]
port 228 nsew signal tristate
flabel metal2 s 154896 0 155008 800 0 FreeSans 448 90 0 0 la_data_out[53]
port 229 nsew signal tristate
flabel metal2 s 156576 0 156688 800 0 FreeSans 448 90 0 0 la_data_out[54]
port 230 nsew signal tristate
flabel metal2 s 158256 0 158368 800 0 FreeSans 448 90 0 0 la_data_out[55]
port 231 nsew signal tristate
flabel metal2 s 159936 0 160048 800 0 FreeSans 448 90 0 0 la_data_out[56]
port 232 nsew signal tristate
flabel metal2 s 161616 0 161728 800 0 FreeSans 448 90 0 0 la_data_out[57]
port 233 nsew signal tristate
flabel metal2 s 163296 0 163408 800 0 FreeSans 448 90 0 0 la_data_out[58]
port 234 nsew signal tristate
flabel metal2 s 164976 0 165088 800 0 FreeSans 448 90 0 0 la_data_out[59]
port 235 nsew signal tristate
flabel metal2 s 74256 0 74368 800 0 FreeSans 448 90 0 0 la_data_out[5]
port 236 nsew signal tristate
flabel metal2 s 166656 0 166768 800 0 FreeSans 448 90 0 0 la_data_out[60]
port 237 nsew signal tristate
flabel metal2 s 168336 0 168448 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 238 nsew signal tristate
flabel metal2 s 170016 0 170128 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 239 nsew signal tristate
flabel metal2 s 171696 0 171808 800 0 FreeSans 448 90 0 0 la_data_out[63]
port 240 nsew signal tristate
flabel metal2 s 75936 0 76048 800 0 FreeSans 448 90 0 0 la_data_out[6]
port 241 nsew signal tristate
flabel metal2 s 77616 0 77728 800 0 FreeSans 448 90 0 0 la_data_out[7]
port 242 nsew signal tristate
flabel metal2 s 79296 0 79408 800 0 FreeSans 448 90 0 0 la_data_out[8]
port 243 nsew signal tristate
flabel metal2 s 80976 0 81088 800 0 FreeSans 448 90 0 0 la_data_out[9]
port 244 nsew signal tristate
flabel metal2 s 66416 0 66528 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 245 nsew signal input
flabel metal2 s 83216 0 83328 800 0 FreeSans 448 90 0 0 la_oenb[10]
port 246 nsew signal input
flabel metal2 s 84896 0 85008 800 0 FreeSans 448 90 0 0 la_oenb[11]
port 247 nsew signal input
flabel metal2 s 86576 0 86688 800 0 FreeSans 448 90 0 0 la_oenb[12]
port 248 nsew signal input
flabel metal2 s 88256 0 88368 800 0 FreeSans 448 90 0 0 la_oenb[13]
port 249 nsew signal input
flabel metal2 s 89936 0 90048 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 250 nsew signal input
flabel metal2 s 91616 0 91728 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 251 nsew signal input
flabel metal2 s 93296 0 93408 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 252 nsew signal input
flabel metal2 s 94976 0 95088 800 0 FreeSans 448 90 0 0 la_oenb[17]
port 253 nsew signal input
flabel metal2 s 96656 0 96768 800 0 FreeSans 448 90 0 0 la_oenb[18]
port 254 nsew signal input
flabel metal2 s 98336 0 98448 800 0 FreeSans 448 90 0 0 la_oenb[19]
port 255 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 256 nsew signal input
flabel metal2 s 100016 0 100128 800 0 FreeSans 448 90 0 0 la_oenb[20]
port 257 nsew signal input
flabel metal2 s 101696 0 101808 800 0 FreeSans 448 90 0 0 la_oenb[21]
port 258 nsew signal input
flabel metal2 s 103376 0 103488 800 0 FreeSans 448 90 0 0 la_oenb[22]
port 259 nsew signal input
flabel metal2 s 105056 0 105168 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 260 nsew signal input
flabel metal2 s 106736 0 106848 800 0 FreeSans 448 90 0 0 la_oenb[24]
port 261 nsew signal input
flabel metal2 s 108416 0 108528 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 262 nsew signal input
flabel metal2 s 110096 0 110208 800 0 FreeSans 448 90 0 0 la_oenb[26]
port 263 nsew signal input
flabel metal2 s 111776 0 111888 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 264 nsew signal input
flabel metal2 s 113456 0 113568 800 0 FreeSans 448 90 0 0 la_oenb[28]
port 265 nsew signal input
flabel metal2 s 115136 0 115248 800 0 FreeSans 448 90 0 0 la_oenb[29]
port 266 nsew signal input
flabel metal2 s 69776 0 69888 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 267 nsew signal input
flabel metal2 s 116816 0 116928 800 0 FreeSans 448 90 0 0 la_oenb[30]
port 268 nsew signal input
flabel metal2 s 118496 0 118608 800 0 FreeSans 448 90 0 0 la_oenb[31]
port 269 nsew signal input
flabel metal2 s 120176 0 120288 800 0 FreeSans 448 90 0 0 la_oenb[32]
port 270 nsew signal input
flabel metal2 s 121856 0 121968 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 271 nsew signal input
flabel metal2 s 123536 0 123648 800 0 FreeSans 448 90 0 0 la_oenb[34]
port 272 nsew signal input
flabel metal2 s 125216 0 125328 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 273 nsew signal input
flabel metal2 s 126896 0 127008 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 274 nsew signal input
flabel metal2 s 128576 0 128688 800 0 FreeSans 448 90 0 0 la_oenb[37]
port 275 nsew signal input
flabel metal2 s 130256 0 130368 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 276 nsew signal input
flabel metal2 s 131936 0 132048 800 0 FreeSans 448 90 0 0 la_oenb[39]
port 277 nsew signal input
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 278 nsew signal input
flabel metal2 s 133616 0 133728 800 0 FreeSans 448 90 0 0 la_oenb[40]
port 279 nsew signal input
flabel metal2 s 135296 0 135408 800 0 FreeSans 448 90 0 0 la_oenb[41]
port 280 nsew signal input
flabel metal2 s 136976 0 137088 800 0 FreeSans 448 90 0 0 la_oenb[42]
port 281 nsew signal input
flabel metal2 s 138656 0 138768 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 282 nsew signal input
flabel metal2 s 140336 0 140448 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 283 nsew signal input
flabel metal2 s 142016 0 142128 800 0 FreeSans 448 90 0 0 la_oenb[45]
port 284 nsew signal input
flabel metal2 s 143696 0 143808 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 285 nsew signal input
flabel metal2 s 145376 0 145488 800 0 FreeSans 448 90 0 0 la_oenb[47]
port 286 nsew signal input
flabel metal2 s 147056 0 147168 800 0 FreeSans 448 90 0 0 la_oenb[48]
port 287 nsew signal input
flabel metal2 s 148736 0 148848 800 0 FreeSans 448 90 0 0 la_oenb[49]
port 288 nsew signal input
flabel metal2 s 73136 0 73248 800 0 FreeSans 448 90 0 0 la_oenb[4]
port 289 nsew signal input
flabel metal2 s 150416 0 150528 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 290 nsew signal input
flabel metal2 s 152096 0 152208 800 0 FreeSans 448 90 0 0 la_oenb[51]
port 291 nsew signal input
flabel metal2 s 153776 0 153888 800 0 FreeSans 448 90 0 0 la_oenb[52]
port 292 nsew signal input
flabel metal2 s 155456 0 155568 800 0 FreeSans 448 90 0 0 la_oenb[53]
port 293 nsew signal input
flabel metal2 s 157136 0 157248 800 0 FreeSans 448 90 0 0 la_oenb[54]
port 294 nsew signal input
flabel metal2 s 158816 0 158928 800 0 FreeSans 448 90 0 0 la_oenb[55]
port 295 nsew signal input
flabel metal2 s 160496 0 160608 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 296 nsew signal input
flabel metal2 s 162176 0 162288 800 0 FreeSans 448 90 0 0 la_oenb[57]
port 297 nsew signal input
flabel metal2 s 163856 0 163968 800 0 FreeSans 448 90 0 0 la_oenb[58]
port 298 nsew signal input
flabel metal2 s 165536 0 165648 800 0 FreeSans 448 90 0 0 la_oenb[59]
port 299 nsew signal input
flabel metal2 s 74816 0 74928 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 300 nsew signal input
flabel metal2 s 167216 0 167328 800 0 FreeSans 448 90 0 0 la_oenb[60]
port 301 nsew signal input
flabel metal2 s 168896 0 169008 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 302 nsew signal input
flabel metal2 s 170576 0 170688 800 0 FreeSans 448 90 0 0 la_oenb[62]
port 303 nsew signal input
flabel metal2 s 172256 0 172368 800 0 FreeSans 448 90 0 0 la_oenb[63]
port 304 nsew signal input
flabel metal2 s 76496 0 76608 800 0 FreeSans 448 90 0 0 la_oenb[6]
port 305 nsew signal input
flabel metal2 s 78176 0 78288 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 306 nsew signal input
flabel metal2 s 79856 0 79968 800 0 FreeSans 448 90 0 0 la_oenb[8]
port 307 nsew signal input
flabel metal2 s 81536 0 81648 800 0 FreeSans 448 90 0 0 la_oenb[9]
port 308 nsew signal input
flabel metal4 s 23346 3076 23666 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 67670 3076 67990 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 111994 3076 112314 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 156318 3076 156638 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 45508 3076 45828 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 89832 3076 90152 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 134156 3076 134476 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 178480 3076 178800 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 wb_clk_i
port 311 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 wb_rst_i
port 312 nsew signal input
flabel metal2 s 7056 0 7168 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 313 nsew signal tristate
flabel metal2 s 9296 0 9408 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 314 nsew signal input
flabel metal2 s 28336 0 28448 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 315 nsew signal input
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 316 nsew signal input
flabel metal2 s 31696 0 31808 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 317 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 318 nsew signal input
flabel metal2 s 35056 0 35168 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 319 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 320 nsew signal input
flabel metal2 s 38416 0 38528 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 321 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 322 nsew signal input
flabel metal2 s 41776 0 41888 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 323 nsew signal input
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 324 nsew signal input
flabel metal2 s 11536 0 11648 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 325 nsew signal input
flabel metal2 s 45136 0 45248 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 326 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 327 nsew signal input
flabel metal2 s 48496 0 48608 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 328 nsew signal input
flabel metal2 s 50176 0 50288 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 329 nsew signal input
flabel metal2 s 51856 0 51968 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 330 nsew signal input
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 331 nsew signal input
flabel metal2 s 55216 0 55328 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 332 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 333 nsew signal input
flabel metal2 s 58576 0 58688 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 334 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 335 nsew signal input
flabel metal2 s 13776 0 13888 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 336 nsew signal input
flabel metal2 s 61936 0 62048 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 337 nsew signal input
flabel metal2 s 63616 0 63728 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 338 nsew signal input
flabel metal2 s 16016 0 16128 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 339 nsew signal input
flabel metal2 s 18256 0 18368 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 340 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 341 nsew signal input
flabel metal2 s 21616 0 21728 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 342 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 343 nsew signal input
flabel metal2 s 24976 0 25088 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 344 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 345 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 346 nsew signal input
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 347 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 348 nsew signal input
flabel metal2 s 30576 0 30688 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 349 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 350 nsew signal input
flabel metal2 s 33936 0 34048 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 351 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 352 nsew signal input
flabel metal2 s 37296 0 37408 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 353 nsew signal input
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 354 nsew signal input
flabel metal2 s 40656 0 40768 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 355 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 356 nsew signal input
flabel metal2 s 44016 0 44128 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 357 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 358 nsew signal input
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 359 nsew signal input
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 360 nsew signal input
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 361 nsew signal input
flabel metal2 s 50736 0 50848 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 362 nsew signal input
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 363 nsew signal input
flabel metal2 s 54096 0 54208 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 364 nsew signal input
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 365 nsew signal input
flabel metal2 s 57456 0 57568 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 366 nsew signal input
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 367 nsew signal input
flabel metal2 s 60816 0 60928 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 368 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 369 nsew signal input
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 370 nsew signal input
flabel metal2 s 64176 0 64288 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 371 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 372 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 373 nsew signal input
flabel metal2 s 20496 0 20608 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 374 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 375 nsew signal input
flabel metal2 s 23856 0 23968 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 376 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 377 nsew signal input
flabel metal2 s 27216 0 27328 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 378 nsew signal input
flabel metal2 s 10416 0 10528 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 379 nsew signal tristate
flabel metal2 s 29456 0 29568 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 380 nsew signal tristate
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 381 nsew signal tristate
flabel metal2 s 32816 0 32928 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 382 nsew signal tristate
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 383 nsew signal tristate
flabel metal2 s 36176 0 36288 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 384 nsew signal tristate
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 385 nsew signal tristate
flabel metal2 s 39536 0 39648 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 386 nsew signal tristate
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 387 nsew signal tristate
flabel metal2 s 42896 0 43008 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 388 nsew signal tristate
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 389 nsew signal tristate
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 390 nsew signal tristate
flabel metal2 s 46256 0 46368 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 391 nsew signal tristate
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 392 nsew signal tristate
flabel metal2 s 49616 0 49728 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 393 nsew signal tristate
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 394 nsew signal tristate
flabel metal2 s 52976 0 53088 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 395 nsew signal tristate
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 396 nsew signal tristate
flabel metal2 s 56336 0 56448 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 397 nsew signal tristate
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 398 nsew signal tristate
flabel metal2 s 59696 0 59808 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 399 nsew signal tristate
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 400 nsew signal tristate
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 401 nsew signal tristate
flabel metal2 s 63056 0 63168 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 402 nsew signal tristate
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 403 nsew signal tristate
flabel metal2 s 17136 0 17248 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 404 nsew signal tristate
flabel metal2 s 19376 0 19488 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 405 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 406 nsew signal tristate
flabel metal2 s 22736 0 22848 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 407 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 408 nsew signal tristate
flabel metal2 s 26096 0 26208 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 409 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 410 nsew signal tristate
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 411 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 412 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 413 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 414 nsew signal input
flabel metal2 s 8176 0 8288 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 415 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_we_i
port 416 nsew signal input
rlabel metal1 89992 16464 89992 16464 0 vdd
rlabel via1 90072 15680 90072 15680 0 vss
rlabel metal3 17416 15512 17416 15512 0 _000_
rlabel metal2 26824 12600 26824 12600 0 _001_
rlabel metal3 26712 12376 26712 12376 0 _002_
rlabel metal2 1848 16296 1848 16296 0 io_in[0]
rlabel metal2 5992 16184 5992 16184 0 io_in[1]
rlabel metal2 10584 15792 10584 15792 0 io_in[2]
rlabel metal2 15400 16184 15400 16184 0 io_in[3]
rlabel metal2 20216 17738 20216 17738 0 io_in[4]
rlabel metal2 24808 16184 24808 16184 0 io_in[5]
rlabel metal2 31416 16352 31416 16352 0 io_in[6]
rlabel via1 37128 15512 37128 15512 0 io_in[7]
rlabel metal2 38920 16184 38920 16184 0 io_in[8]
rlabel via1 44184 16632 44184 16632 0 io_in[9]
rlabel metal2 119672 2534 119672 2534 0 la_data_out[32]
rlabel metal2 121352 2478 121352 2478 0 la_data_out[33]
rlabel metal2 16016 15512 16016 15512 0 net1
rlabel metal2 26936 15456 26936 15456 0 net10
rlabel metal2 170072 2030 170072 2030 0 net100
rlabel metal2 171752 2030 171752 2030 0 net101
rlabel metal2 172872 2030 172872 2030 0 net102
rlabel metal2 173432 1246 173432 1246 0 net103
rlabel metal2 173992 2030 173992 2030 0 net104
rlabel metal2 4648 15960 4648 15960 0 net105
rlabel metal2 9072 15960 9072 15960 0 net106
rlabel metal2 14056 15960 14056 15960 0 net107
rlabel metal2 19208 16296 19208 16296 0 net108
rlabel metal2 23408 15960 23408 15960 0 net109
rlabel metal2 21896 8008 21896 8008 0 net11
rlabel metal2 28168 15960 28168 15960 0 net110
rlabel metal2 32592 15960 32592 15960 0 net111
rlabel metal2 38024 16296 38024 16296 0 net112
rlabel metal2 42280 15960 42280 15960 0 net113
rlabel metal2 46984 15960 46984 15960 0 net114
rlabel metal2 51464 15512 51464 15512 0 net115
rlabel metal2 56728 16800 56728 16800 0 net116
rlabel metal2 61096 15512 61096 15512 0 net117
rlabel metal2 65800 15960 65800 15960 0 net118
rlabel metal2 70504 15960 70504 15960 0 net119
rlabel metal2 21896 10248 21896 10248 0 net12
rlabel metal2 75208 15960 75208 15960 0 net120
rlabel metal2 80248 16800 80248 16800 0 net121
rlabel metal2 84616 15960 84616 15960 0 net122
rlabel metal2 89264 15960 89264 15960 0 net123
rlabel metal2 94024 15512 94024 15512 0 net124
rlabel metal2 98728 15960 98728 15960 0 net125
rlabel metal2 103768 16800 103768 16800 0 net126
rlabel metal2 108136 15960 108136 15960 0 net127
rlabel metal2 112840 15960 112840 15960 0 net128
rlabel metal2 117544 15960 117544 15960 0 net129
rlabel metal2 20552 10976 20552 10976 0 net13
rlabel metal2 122248 15960 122248 15960 0 net130
rlabel metal2 127288 16800 127288 16800 0 net131
rlabel metal2 131656 15960 131656 15960 0 net132
rlabel metal2 136360 15960 136360 15960 0 net133
rlabel metal2 141064 15960 141064 15960 0 net134
rlabel metal2 145768 15960 145768 15960 0 net135
rlabel metal2 150808 16800 150808 16800 0 net136
rlabel metal2 155176 15960 155176 15960 0 net137
rlabel metal2 159880 15960 159880 15960 0 net138
rlabel metal2 164584 15960 164584 15960 0 net139
rlabel metal2 25592 13664 25592 13664 0 net14
rlabel metal2 169288 15960 169288 15960 0 net140
rlabel metal2 174328 16800 174328 16800 0 net141
rlabel metal2 178136 16464 178136 16464 0 net142
rlabel metal2 3080 15960 3080 15960 0 net143
rlabel metal2 7784 15960 7784 15960 0 net144
rlabel metal2 12488 14392 12488 14392 0 net145
rlabel metal2 16744 16296 16744 16296 0 net146
rlabel metal2 22344 16016 22344 16016 0 net147
rlabel metal2 26600 15960 26600 15960 0 net148
rlabel metal2 31192 17402 31192 17402 0 net149
rlabel metal2 61544 11816 61544 11816 0 net15
rlabel metal2 36456 16072 36456 16072 0 net150
rlabel metal2 41048 16800 41048 16800 0 net151
rlabel metal2 45864 16016 45864 16016 0 net152
rlabel metal2 50120 15512 50120 15512 0 net153
rlabel metal2 54824 15960 54824 15960 0 net154
rlabel metal2 59528 15960 59528 15960 0 net155
rlabel metal2 66584 16016 66584 16016 0 net156
rlabel metal2 69048 16296 69048 16296 0 net157
rlabel metal2 73080 16800 73080 16800 0 net158
rlabel metal2 78344 15960 78344 15960 0 net159
rlabel metal2 40152 11816 40152 11816 0 net16
rlabel metal2 83048 15960 83048 15960 0 net160
rlabel metal2 88088 16800 88088 16800 0 net161
rlabel metal2 92568 16072 92568 16072 0 net162
rlabel metal2 97160 15960 97160 15960 0 net163
rlabel metal2 101864 15960 101864 15960 0 net164
rlabel metal2 106568 15960 106568 15960 0 net165
rlabel metal2 111608 16800 111608 16800 0 net166
rlabel metal2 116088 16296 116088 16296 0 net167
rlabel metal2 120680 15960 120680 15960 0 net168
rlabel metal2 125384 15960 125384 15960 0 net169
rlabel metal3 61040 12264 61040 12264 0 net17
rlabel metal2 130088 15960 130088 15960 0 net170
rlabel metal2 135128 16800 135128 16800 0 net171
rlabel metal2 139608 16296 139608 16296 0 net172
rlabel metal2 144200 15960 144200 15960 0 net173
rlabel metal2 148904 15960 148904 15960 0 net174
rlabel metal2 153608 15960 153608 15960 0 net175
rlabel metal2 158648 16800 158648 16800 0 net176
rlabel metal2 163128 16296 163128 16296 0 net177
rlabel metal2 167720 15960 167720 15960 0 net178
rlabel metal2 172424 15960 172424 15960 0 net179
rlabel metal3 40768 10696 40768 10696 0 net18
rlabel metal2 177128 15960 177128 15960 0 net180
rlabel metal2 7112 2030 7112 2030 0 net181
rlabel metal2 10472 2030 10472 2030 0 net182
rlabel metal2 12712 2030 12712 2030 0 net183
rlabel metal2 14952 2030 14952 2030 0 net184
rlabel metal2 17192 2030 17192 2030 0 net185
rlabel metal2 19432 2030 19432 2030 0 net186
rlabel metal2 21112 2030 21112 2030 0 net187
rlabel metal2 22792 2030 22792 2030 0 net188
rlabel metal2 24472 2030 24472 2030 0 net189
rlabel metal2 62440 12376 62440 12376 0 net19
rlabel metal2 26152 2030 26152 2030 0 net190
rlabel metal2 27832 2030 27832 2030 0 net191
rlabel metal2 29512 2030 29512 2030 0 net192
rlabel metal2 31192 2030 31192 2030 0 net193
rlabel metal2 32872 2030 32872 2030 0 net194
rlabel metal2 34552 2030 34552 2030 0 net195
rlabel metal2 36232 2030 36232 2030 0 net196
rlabel metal2 37912 2030 37912 2030 0 net197
rlabel metal2 39592 2030 39592 2030 0 net198
rlabel metal2 41272 2030 41272 2030 0 net199
rlabel metal3 8568 15960 8568 15960 0 net2
rlabel metal3 40096 11256 40096 11256 0 net20
rlabel metal2 42952 2030 42952 2030 0 net200
rlabel metal2 44632 2030 44632 2030 0 net201
rlabel metal2 46312 2030 46312 2030 0 net202
rlabel metal2 47992 2030 47992 2030 0 net203
rlabel metal2 49672 2030 49672 2030 0 net204
rlabel metal2 51352 2030 51352 2030 0 net205
rlabel metal2 53032 2030 53032 2030 0 net206
rlabel metal2 54712 2030 54712 2030 0 net207
rlabel metal2 56392 2030 56392 2030 0 net208
rlabel metal2 58072 2030 58072 2030 0 net209
rlabel metal2 62048 10696 62048 10696 0 net21
rlabel metal2 59752 2030 59752 2030 0 net210
rlabel metal2 61432 2030 61432 2030 0 net211
rlabel metal2 63112 2030 63112 2030 0 net212
rlabel metal2 64792 2030 64792 2030 0 net213
rlabel metal2 52472 11088 52472 11088 0 net214
rlabel metal3 52696 11368 52696 11368 0 net215
rlabel metal3 40544 12824 40544 12824 0 net22
rlabel metal2 60648 12040 60648 12040 0 net23
rlabel metal2 39648 12264 39648 12264 0 net24
rlabel metal2 60984 13048 60984 13048 0 net25
rlabel metal2 40600 10080 40600 10080 0 net26
rlabel metal2 63168 11368 63168 11368 0 net27
rlabel metal2 40600 11480 40600 11480 0 net28
rlabel metal2 63784 11816 63784 11816 0 net29
rlabel metal3 11480 15400 11480 15400 0 net3
rlabel metal3 41776 11256 41776 11256 0 net30
rlabel metal2 53704 14784 53704 14784 0 net31
rlabel metal2 53816 15288 53816 15288 0 net32
rlabel metal2 64568 15176 64568 15176 0 net33
rlabel metal2 65072 15288 65072 15288 0 net34
rlabel metal2 73864 15848 73864 15848 0 net35
rlabel metal2 74424 15568 74424 15568 0 net36
rlabel metal2 90776 15568 90776 15568 0 net37
rlabel metal2 90272 14504 90272 14504 0 net38
rlabel metal3 26824 11368 26824 11368 0 net39
rlabel metal2 26264 15624 26264 15624 0 net4
rlabel metal2 65912 2030 65912 2030 0 net40
rlabel metal2 67592 1246 67592 1246 0 net41
rlabel metal2 69272 2030 69272 2030 0 net42
rlabel metal2 70952 2030 70952 2030 0 net43
rlabel metal2 72632 2030 72632 2030 0 net44
rlabel metal2 74312 2030 74312 2030 0 net45
rlabel metal2 75992 2030 75992 2030 0 net46
rlabel metal2 77672 2030 77672 2030 0 net47
rlabel metal2 79352 1246 79352 1246 0 net48
rlabel metal2 81032 2030 81032 2030 0 net49
rlabel metal2 21672 15176 21672 15176 0 net5
rlabel metal2 82712 2030 82712 2030 0 net50
rlabel metal2 84392 2030 84392 2030 0 net51
rlabel metal2 86072 2030 86072 2030 0 net52
rlabel metal2 87752 2030 87752 2030 0 net53
rlabel metal2 89432 2030 89432 2030 0 net54
rlabel metal2 91112 1246 91112 1246 0 net55
rlabel metal2 92792 2030 92792 2030 0 net56
rlabel metal2 94472 2030 94472 2030 0 net57
rlabel metal2 96152 2030 96152 2030 0 net58
rlabel metal2 97832 2030 97832 2030 0 net59
rlabel metal2 25704 16072 25704 16072 0 net6
rlabel metal2 99512 2030 99512 2030 0 net60
rlabel metal2 101192 2030 101192 2030 0 net61
rlabel metal2 102872 1246 102872 1246 0 net62
rlabel metal2 104552 2030 104552 2030 0 net63
rlabel metal2 106232 2030 106232 2030 0 net64
rlabel metal2 107912 2030 107912 2030 0 net65
rlabel metal2 109592 2030 109592 2030 0 net66
rlabel metal2 111272 2030 111272 2030 0 net67
rlabel metal2 112952 2030 112952 2030 0 net68
rlabel metal2 114632 1246 114632 1246 0 net69
rlabel metal2 31752 16184 31752 16184 0 net7
rlabel metal2 116312 2030 116312 2030 0 net70
rlabel metal2 117992 2030 117992 2030 0 net71
rlabel metal2 123032 2030 123032 2030 0 net72
rlabel metal2 124712 2030 124712 2030 0 net73
rlabel metal2 126392 1246 126392 1246 0 net74
rlabel metal2 128072 2030 128072 2030 0 net75
rlabel metal2 129752 2030 129752 2030 0 net76
rlabel metal2 131432 2030 131432 2030 0 net77
rlabel metal2 133112 2030 133112 2030 0 net78
rlabel metal2 134792 2030 134792 2030 0 net79
rlabel metal2 77000 15736 77000 15736 0 net8
rlabel metal2 136472 2030 136472 2030 0 net80
rlabel metal2 138152 1246 138152 1246 0 net81
rlabel metal2 139832 2030 139832 2030 0 net82
rlabel metal2 141512 2030 141512 2030 0 net83
rlabel metal2 143192 2030 143192 2030 0 net84
rlabel metal2 144872 2030 144872 2030 0 net85
rlabel metal2 146552 2030 146552 2030 0 net86
rlabel metal2 148232 2030 148232 2030 0 net87
rlabel metal2 149912 1246 149912 1246 0 net88
rlabel metal2 151592 2030 151592 2030 0 net89
rlabel metal2 91784 15736 91784 15736 0 net9
rlabel metal2 153272 2030 153272 2030 0 net90
rlabel metal2 154952 2030 154952 2030 0 net91
rlabel metal2 156632 2030 156632 2030 0 net92
rlabel metal2 158312 2030 158312 2030 0 net93
rlabel metal2 159992 2030 159992 2030 0 net94
rlabel metal2 161672 1246 161672 1246 0 net95
rlabel metal2 163352 2030 163352 2030 0 net96
rlabel metal2 165032 2030 165032 2030 0 net97
rlabel metal2 166712 2030 166712 2030 0 net98
rlabel metal2 168392 2030 168392 2030 0 net99
rlabel metal2 30128 15960 30128 15960 0 u_inj.outn
rlabel metal2 21000 10976 21000 10976 0 u_inj.outp
rlabel metal2 25872 11592 25872 11592 0 u_inj.signal_n
rlabel metal2 52024 16128 52024 16128 0 u_inj.trim_n_r\[0\]
rlabel metal2 63224 15736 63224 15736 0 u_inj.trim_n_r\[1\]
rlabel metal3 75600 15288 75600 15288 0 u_inj.trim_n_r\[2\]
rlabel metal2 94920 15736 94920 15736 0 u_inj.trim_n_r\[3\]
rlabel metal2 17752 15736 17752 15736 0 u_inj.trim_p_r\[0\]
rlabel metal2 15400 13720 15400 13720 0 u_inj.trim_p_r\[1\]
rlabel metal2 30576 15288 30576 15288 0 u_inj.trim_p_r\[2\]
rlabel metal2 36120 15288 36120 15288 0 u_inj.trim_p_r\[3\]
<< properties >>
string FIXED_BBOX 0 0 180000 20000
<< end >>
