* NGSPICE file created from caparray_s1.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

.subckt caparray_s1 cap_series_gygyn cap_series_gygyp cap_series_gyn cap_series_gyp
+ cap_shunt_gyn cap_shunt_gyp cap_shunt_n cap_shunt_p tune_series_gy[0] tune_series_gy[1]
+ tune_series_gy[2] tune_series_gy[3] tune_series_gy[4] tune_series_gy[5] tune_series_gygy[0]
+ tune_series_gygy[1] tune_series_gygy[2] tune_series_gygy[3] tune_series_gygy[4]
+ tune_series_gygy[5] tune_shunt[0] tune_shunt[1] tune_shunt[2] tune_shunt[3] tune_shunt[4]
+ tune_shunt[5] tune_shunt[6] tune_shunt[7] tune_shunt_gy[0] tune_shunt_gy[1] tune_shunt_gy[2]
+ tune_shunt_gy[3] tune_shunt_gy[4] tune_shunt_gy[5] tune_shunt_gy[6] vdd vss
XFILLER_54_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[12\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[12\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[72\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[72\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[7\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[7\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g8\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[0] gen_shunt_g8\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g1\[3\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[3\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g2\[3\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[3\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[88\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[88\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[37\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[37\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[71\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[71\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_series_gy_g1\[12\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[12\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[0\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[0\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[39\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[39\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[5\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[5\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[87\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[87\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[3\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[3\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[36\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[36\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[70\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[70\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g1\[5\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[5\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[89\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[89\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[38\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[38\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[86\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[86\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[35\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[35\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[3\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[3\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[88\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[88\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g4\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[37\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[37\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[85\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[85\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g3\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[0\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[0\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[34\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[34\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[87\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[87\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[36\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[36\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[5\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[5\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g2\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[84\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[84\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g3\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[33\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[33\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[86\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[86\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[35\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[35\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[83\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[83\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[32\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[32\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[13\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[13\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gygy_g3\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[3]
+ gen_shunt_gygy_g3\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[85\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[85\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[34\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[34\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[82\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[82\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_43_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[84\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[84\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g3\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[13\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[13\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g2\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g2\[39\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[39\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[33\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[33\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[6\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[6\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[81\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[81\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[49\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[49\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[83\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[83\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[32\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[32\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[38\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[38\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[6\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[6\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[13\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[13\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g3\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[3]
+ gen_shunt_gygy_g3\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[80\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[80\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g7\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[1] gen_shunt_g7\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[48\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[48\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[82\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[82\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[37\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[37\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[6\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[6\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[13\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[13\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[1\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[1\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g2\[39\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[39\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g7\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[1] gen_shunt_g7\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[47\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[47\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g2\[2\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[2\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[6\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[6\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[81\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[81\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[36\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[36\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[49\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[49\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g2\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[38\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[38\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[6\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[6\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[46\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[46\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g3\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[80\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[80\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[2\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[2\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g7\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[1] gen_shunt_g7\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[35\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[35\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[48\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[48\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[37\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[37\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[45\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[45\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[6\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[6\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[1\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[1\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g7\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[1] gen_shunt_g7\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[34\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[34\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[2\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[2\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[47\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[47\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g3\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[2] gen_shunt_gy_g3\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[2\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[2\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[2]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[95\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[95\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g3\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[36\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[36\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[44\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[44\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g4\[0\].u_shunt_n cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[0] gen_shunt_gy_g4\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[33\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[33\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[46\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[46\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[2\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[2\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_gy_g3\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[1] gen_shunt_gy_g3\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[94\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[94\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[35\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[35\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp2 cap_series_gygyp cap_series_gygyp tune_series_gygy[1]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gygy_g1\[4\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[4\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[43\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[43\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[32\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[32\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[45\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[45\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[14\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[14\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[93\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[93\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g2\[34\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[34\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[2\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[2\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gy_g3\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[2] gen_shunt_gy_g3\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[42\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[42\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[2]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp3 cap_series_gygyp cap_series_gygyp tune_series_gygy[0]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp3/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[95\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[95\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g3\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g3\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[44\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[44\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g4\[0\].u_shunt_p cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[0] gen_shunt_gy_g4\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[14\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[14\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[92\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[92\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[33\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[33\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[41\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[41\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g1\[7\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[7\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g3\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[1] gen_shunt_gy_g3\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[94\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[94\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn2 cap_series_gygyn cap_series_gygyn tune_series_gygy[1]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[3\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[3\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g1\[4\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[4\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[43\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[43\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gygy_g1\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[91\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[91\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[32\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[32\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[14\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[14\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[40\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[40\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[59\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[59\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[93\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[93\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g1\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[42\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[42\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn3 cap_series_gygyn cap_series_gygyn tune_series_gygy[0]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn3/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g2\[3\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[3\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[90\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[90\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[58\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[58\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[92\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[92\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[14\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[14\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[2\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[2\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[41\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[41\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[47\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[47\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[7\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[7\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[3\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[3\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[57\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[57\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[91\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[91\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_51_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g5\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[0]
+ gen_series_gy_g5\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[40\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[40\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[46\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[46\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[59\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[59\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g6\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[56\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[56\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[3\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[3\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[90\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[90\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[5\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[5\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[45\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[45\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[58\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[58\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[2\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[2\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[47\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[47\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[55\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[55\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[44\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[44\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[57\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[57\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g1\[5\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[5\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g5\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[0]
+ gen_series_gy_g5\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[46\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[46\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[54\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[54\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g6\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[43\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[43\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[56\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[56\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[5\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[5\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[45\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[45\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_series_gy_g1\[15\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[15\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[7\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[7\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[53\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[53\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g6\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[8\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[8\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[42\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[42\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[55\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[55\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[44\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[44\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[5\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[5\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[52\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[52\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[15\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[15\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g3\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[2] gen_shunt_gy_g3\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[41\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[41\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[54\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[54\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[8\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[8\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[43\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[43\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[51\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[51\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[10\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[10\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[40\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[40\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[15\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[15\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[7\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[7\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[53\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[53\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gy_g3\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[1] gen_shunt_gy_g3\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g4\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[1]
+ gen_series_gy_g4\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[3\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[3\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[8\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[8\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[42\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[42\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[50\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[50\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[69\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[69\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[10\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[10\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[52\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[52\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[15\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[15\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[3\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[3\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g3\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[2] gen_shunt_gy_g3\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[41\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[41\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[8\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[8\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[68\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[68\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[51\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[51\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[10\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[10\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g2\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[40\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[40\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g3\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[1] gen_shunt_gy_g3\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g4\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[1]
+ gen_series_gy_g4\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[67\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[67\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[2\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[2\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[3\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[3\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[50\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[50\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[69\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[69\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[10\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[10\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[66\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[66\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[3\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[3\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_51_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[2\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[2\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g5\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[68\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[68\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[65\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[65\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[67\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[67\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[2\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[2\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[64\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[64\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[66\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[66\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[9\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[9\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_gy_g2\[2\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[2\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g3\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g5\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[63\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[63\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[4\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g5\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[65\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[65\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g5\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[9\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[9\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[62\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[62\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[4\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[4\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[64\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[64\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_51_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[11\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[11\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[61\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[61\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g4\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[1]
+ gen_series_gy_g4\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[9\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[9\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g3\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[63\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[63\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[4\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[11\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[11\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[6\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[6\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[60\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[60\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[79\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[79\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[4\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[4\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[9\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[9\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[62\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[62\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[4\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[11\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[11\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g2\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[78\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[78\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g2\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[61\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[61\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g4\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[1]
+ gen_series_gy_g4\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[77\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[77\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[6\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[6\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[11\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[11\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[60\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[60\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[2\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[2\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[79\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[79\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[4\].u_series_gyn2 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g1\[4\].u_series_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[76\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[76\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_series_gy_g2\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g4\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g2\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[78\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[78\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g3\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[3]
+ gen_shunt_gygy_g3\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[75\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[75\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[77\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[77\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g1\[2\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[2\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_58_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[74\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[74\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_43_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[76\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[76\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g4\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[73\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[73\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[7\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[7\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gy_g2\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g3\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[3]
+ gen_shunt_gygy_g3\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[75\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[75\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[12\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[12\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[72\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[72\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[7\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[7\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g8\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[0] gen_shunt_g8\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[74\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[74\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g2\[3\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[3\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[71\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[71\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[12\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[12\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[39\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[39\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[73\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[73\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[7\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[7\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[5\].u_series_gyp2 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g1\[5\].u_series_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[3\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[3\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[70\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[70\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[89\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[89\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_43_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[38\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[38\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

