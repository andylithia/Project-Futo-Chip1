magic
tech gf180mcuC
magscale 1 5
timestamp 1670230239
<< metal1 >>
rect 672 18437 39312 18454
rect 672 18411 2074 18437
rect 2100 18411 2136 18437
rect 2162 18411 2198 18437
rect 2224 18411 2260 18437
rect 2286 18411 2322 18437
rect 2348 18411 2384 18437
rect 2410 18411 2446 18437
rect 2472 18411 2508 18437
rect 2534 18411 7074 18437
rect 7100 18411 7136 18437
rect 7162 18411 7198 18437
rect 7224 18411 7260 18437
rect 7286 18411 7322 18437
rect 7348 18411 7384 18437
rect 7410 18411 7446 18437
rect 7472 18411 7508 18437
rect 7534 18411 12074 18437
rect 12100 18411 12136 18437
rect 12162 18411 12198 18437
rect 12224 18411 12260 18437
rect 12286 18411 12322 18437
rect 12348 18411 12384 18437
rect 12410 18411 12446 18437
rect 12472 18411 12508 18437
rect 12534 18411 17074 18437
rect 17100 18411 17136 18437
rect 17162 18411 17198 18437
rect 17224 18411 17260 18437
rect 17286 18411 17322 18437
rect 17348 18411 17384 18437
rect 17410 18411 17446 18437
rect 17472 18411 17508 18437
rect 17534 18411 22074 18437
rect 22100 18411 22136 18437
rect 22162 18411 22198 18437
rect 22224 18411 22260 18437
rect 22286 18411 22322 18437
rect 22348 18411 22384 18437
rect 22410 18411 22446 18437
rect 22472 18411 22508 18437
rect 22534 18411 27074 18437
rect 27100 18411 27136 18437
rect 27162 18411 27198 18437
rect 27224 18411 27260 18437
rect 27286 18411 27322 18437
rect 27348 18411 27384 18437
rect 27410 18411 27446 18437
rect 27472 18411 27508 18437
rect 27534 18411 32074 18437
rect 32100 18411 32136 18437
rect 32162 18411 32198 18437
rect 32224 18411 32260 18437
rect 32286 18411 32322 18437
rect 32348 18411 32384 18437
rect 32410 18411 32446 18437
rect 32472 18411 32508 18437
rect 32534 18411 37074 18437
rect 37100 18411 37136 18437
rect 37162 18411 37198 18437
rect 37224 18411 37260 18437
rect 37286 18411 37322 18437
rect 37348 18411 37384 18437
rect 37410 18411 37446 18437
rect 37472 18411 37508 18437
rect 37534 18411 39312 18437
rect 672 18394 39312 18411
rect 672 18045 39312 18062
rect 672 18019 4574 18045
rect 4600 18019 4636 18045
rect 4662 18019 4698 18045
rect 4724 18019 4760 18045
rect 4786 18019 4822 18045
rect 4848 18019 4884 18045
rect 4910 18019 4946 18045
rect 4972 18019 5008 18045
rect 5034 18019 9574 18045
rect 9600 18019 9636 18045
rect 9662 18019 9698 18045
rect 9724 18019 9760 18045
rect 9786 18019 9822 18045
rect 9848 18019 9884 18045
rect 9910 18019 9946 18045
rect 9972 18019 10008 18045
rect 10034 18019 14574 18045
rect 14600 18019 14636 18045
rect 14662 18019 14698 18045
rect 14724 18019 14760 18045
rect 14786 18019 14822 18045
rect 14848 18019 14884 18045
rect 14910 18019 14946 18045
rect 14972 18019 15008 18045
rect 15034 18019 19574 18045
rect 19600 18019 19636 18045
rect 19662 18019 19698 18045
rect 19724 18019 19760 18045
rect 19786 18019 19822 18045
rect 19848 18019 19884 18045
rect 19910 18019 19946 18045
rect 19972 18019 20008 18045
rect 20034 18019 24574 18045
rect 24600 18019 24636 18045
rect 24662 18019 24698 18045
rect 24724 18019 24760 18045
rect 24786 18019 24822 18045
rect 24848 18019 24884 18045
rect 24910 18019 24946 18045
rect 24972 18019 25008 18045
rect 25034 18019 29574 18045
rect 29600 18019 29636 18045
rect 29662 18019 29698 18045
rect 29724 18019 29760 18045
rect 29786 18019 29822 18045
rect 29848 18019 29884 18045
rect 29910 18019 29946 18045
rect 29972 18019 30008 18045
rect 30034 18019 34574 18045
rect 34600 18019 34636 18045
rect 34662 18019 34698 18045
rect 34724 18019 34760 18045
rect 34786 18019 34822 18045
rect 34848 18019 34884 18045
rect 34910 18019 34946 18045
rect 34972 18019 35008 18045
rect 35034 18019 39312 18045
rect 672 18002 39312 18019
rect 672 17653 39312 17670
rect 672 17627 2074 17653
rect 2100 17627 2136 17653
rect 2162 17627 2198 17653
rect 2224 17627 2260 17653
rect 2286 17627 2322 17653
rect 2348 17627 2384 17653
rect 2410 17627 2446 17653
rect 2472 17627 2508 17653
rect 2534 17627 7074 17653
rect 7100 17627 7136 17653
rect 7162 17627 7198 17653
rect 7224 17627 7260 17653
rect 7286 17627 7322 17653
rect 7348 17627 7384 17653
rect 7410 17627 7446 17653
rect 7472 17627 7508 17653
rect 7534 17627 12074 17653
rect 12100 17627 12136 17653
rect 12162 17627 12198 17653
rect 12224 17627 12260 17653
rect 12286 17627 12322 17653
rect 12348 17627 12384 17653
rect 12410 17627 12446 17653
rect 12472 17627 12508 17653
rect 12534 17627 17074 17653
rect 17100 17627 17136 17653
rect 17162 17627 17198 17653
rect 17224 17627 17260 17653
rect 17286 17627 17322 17653
rect 17348 17627 17384 17653
rect 17410 17627 17446 17653
rect 17472 17627 17508 17653
rect 17534 17627 22074 17653
rect 22100 17627 22136 17653
rect 22162 17627 22198 17653
rect 22224 17627 22260 17653
rect 22286 17627 22322 17653
rect 22348 17627 22384 17653
rect 22410 17627 22446 17653
rect 22472 17627 22508 17653
rect 22534 17627 27074 17653
rect 27100 17627 27136 17653
rect 27162 17627 27198 17653
rect 27224 17627 27260 17653
rect 27286 17627 27322 17653
rect 27348 17627 27384 17653
rect 27410 17627 27446 17653
rect 27472 17627 27508 17653
rect 27534 17627 32074 17653
rect 32100 17627 32136 17653
rect 32162 17627 32198 17653
rect 32224 17627 32260 17653
rect 32286 17627 32322 17653
rect 32348 17627 32384 17653
rect 32410 17627 32446 17653
rect 32472 17627 32508 17653
rect 32534 17627 37074 17653
rect 37100 17627 37136 17653
rect 37162 17627 37198 17653
rect 37224 17627 37260 17653
rect 37286 17627 37322 17653
rect 37348 17627 37384 17653
rect 37410 17627 37446 17653
rect 37472 17627 37508 17653
rect 37534 17627 39312 17653
rect 672 17610 39312 17627
rect 12497 17431 12503 17457
rect 12529 17431 12535 17457
rect 13281 17431 13287 17457
rect 13313 17431 13319 17457
rect 13281 17375 13287 17401
rect 13313 17375 13319 17401
rect 672 17261 39312 17278
rect 672 17235 4574 17261
rect 4600 17235 4636 17261
rect 4662 17235 4698 17261
rect 4724 17235 4760 17261
rect 4786 17235 4822 17261
rect 4848 17235 4884 17261
rect 4910 17235 4946 17261
rect 4972 17235 5008 17261
rect 5034 17235 9574 17261
rect 9600 17235 9636 17261
rect 9662 17235 9698 17261
rect 9724 17235 9760 17261
rect 9786 17235 9822 17261
rect 9848 17235 9884 17261
rect 9910 17235 9946 17261
rect 9972 17235 10008 17261
rect 10034 17235 14574 17261
rect 14600 17235 14636 17261
rect 14662 17235 14698 17261
rect 14724 17235 14760 17261
rect 14786 17235 14822 17261
rect 14848 17235 14884 17261
rect 14910 17235 14946 17261
rect 14972 17235 15008 17261
rect 15034 17235 19574 17261
rect 19600 17235 19636 17261
rect 19662 17235 19698 17261
rect 19724 17235 19760 17261
rect 19786 17235 19822 17261
rect 19848 17235 19884 17261
rect 19910 17235 19946 17261
rect 19972 17235 20008 17261
rect 20034 17235 24574 17261
rect 24600 17235 24636 17261
rect 24662 17235 24698 17261
rect 24724 17235 24760 17261
rect 24786 17235 24822 17261
rect 24848 17235 24884 17261
rect 24910 17235 24946 17261
rect 24972 17235 25008 17261
rect 25034 17235 29574 17261
rect 29600 17235 29636 17261
rect 29662 17235 29698 17261
rect 29724 17235 29760 17261
rect 29786 17235 29822 17261
rect 29848 17235 29884 17261
rect 29910 17235 29946 17261
rect 29972 17235 30008 17261
rect 30034 17235 34574 17261
rect 34600 17235 34636 17261
rect 34662 17235 34698 17261
rect 34724 17235 34760 17261
rect 34786 17235 34822 17261
rect 34848 17235 34884 17261
rect 34910 17235 34946 17261
rect 34972 17235 35008 17261
rect 35034 17235 39312 17261
rect 672 17218 39312 17235
rect 10593 17095 10599 17121
rect 10625 17095 10631 17121
rect 12049 17095 12055 17121
rect 12081 17095 12087 17121
rect 9641 17039 9647 17065
rect 9673 17039 9679 17065
rect 10425 17039 10431 17065
rect 10457 17039 10463 17065
rect 11097 17039 11103 17065
rect 11129 17039 11135 17065
rect 11993 17039 11999 17065
rect 12025 17039 12031 17065
rect 12833 17039 12839 17065
rect 12865 17039 12871 17065
rect 13281 17039 13287 17065
rect 13313 17039 13319 17065
rect 13505 17039 13511 17065
rect 13537 17039 13543 17065
rect 672 16869 39312 16886
rect 672 16843 2074 16869
rect 2100 16843 2136 16869
rect 2162 16843 2198 16869
rect 2224 16843 2260 16869
rect 2286 16843 2322 16869
rect 2348 16843 2384 16869
rect 2410 16843 2446 16869
rect 2472 16843 2508 16869
rect 2534 16843 7074 16869
rect 7100 16843 7136 16869
rect 7162 16843 7198 16869
rect 7224 16843 7260 16869
rect 7286 16843 7322 16869
rect 7348 16843 7384 16869
rect 7410 16843 7446 16869
rect 7472 16843 7508 16869
rect 7534 16843 12074 16869
rect 12100 16843 12136 16869
rect 12162 16843 12198 16869
rect 12224 16843 12260 16869
rect 12286 16843 12322 16869
rect 12348 16843 12384 16869
rect 12410 16843 12446 16869
rect 12472 16843 12508 16869
rect 12534 16843 17074 16869
rect 17100 16843 17136 16869
rect 17162 16843 17198 16869
rect 17224 16843 17260 16869
rect 17286 16843 17322 16869
rect 17348 16843 17384 16869
rect 17410 16843 17446 16869
rect 17472 16843 17508 16869
rect 17534 16843 22074 16869
rect 22100 16843 22136 16869
rect 22162 16843 22198 16869
rect 22224 16843 22260 16869
rect 22286 16843 22322 16869
rect 22348 16843 22384 16869
rect 22410 16843 22446 16869
rect 22472 16843 22508 16869
rect 22534 16843 27074 16869
rect 27100 16843 27136 16869
rect 27162 16843 27198 16869
rect 27224 16843 27260 16869
rect 27286 16843 27322 16869
rect 27348 16843 27384 16869
rect 27410 16843 27446 16869
rect 27472 16843 27508 16869
rect 27534 16843 32074 16869
rect 32100 16843 32136 16869
rect 32162 16843 32198 16869
rect 32224 16843 32260 16869
rect 32286 16843 32322 16869
rect 32348 16843 32384 16869
rect 32410 16843 32446 16869
rect 32472 16843 32508 16869
rect 32534 16843 37074 16869
rect 37100 16843 37136 16869
rect 37162 16843 37198 16869
rect 37224 16843 37260 16869
rect 37286 16843 37322 16869
rect 37348 16843 37384 16869
rect 37410 16843 37446 16869
rect 37472 16843 37508 16869
rect 37534 16843 39312 16869
rect 672 16826 39312 16843
rect 9529 16647 9535 16673
rect 9561 16647 9567 16673
rect 10425 16647 10431 16673
rect 10457 16647 10463 16673
rect 10929 16647 10935 16673
rect 10961 16647 10967 16673
rect 11377 16647 11383 16673
rect 11409 16647 11415 16673
rect 11489 16647 11495 16673
rect 11521 16647 11527 16673
rect 12553 16647 12559 16673
rect 12585 16647 12591 16673
rect 13449 16647 13455 16673
rect 13481 16647 13487 16673
rect 10425 16591 10431 16617
rect 10457 16591 10463 16617
rect 13449 16591 13455 16617
rect 13481 16591 13487 16617
rect 672 16477 39312 16494
rect 672 16451 4574 16477
rect 4600 16451 4636 16477
rect 4662 16451 4698 16477
rect 4724 16451 4760 16477
rect 4786 16451 4822 16477
rect 4848 16451 4884 16477
rect 4910 16451 4946 16477
rect 4972 16451 5008 16477
rect 5034 16451 9574 16477
rect 9600 16451 9636 16477
rect 9662 16451 9698 16477
rect 9724 16451 9760 16477
rect 9786 16451 9822 16477
rect 9848 16451 9884 16477
rect 9910 16451 9946 16477
rect 9972 16451 10008 16477
rect 10034 16451 14574 16477
rect 14600 16451 14636 16477
rect 14662 16451 14698 16477
rect 14724 16451 14760 16477
rect 14786 16451 14822 16477
rect 14848 16451 14884 16477
rect 14910 16451 14946 16477
rect 14972 16451 15008 16477
rect 15034 16451 19574 16477
rect 19600 16451 19636 16477
rect 19662 16451 19698 16477
rect 19724 16451 19760 16477
rect 19786 16451 19822 16477
rect 19848 16451 19884 16477
rect 19910 16451 19946 16477
rect 19972 16451 20008 16477
rect 20034 16451 24574 16477
rect 24600 16451 24636 16477
rect 24662 16451 24698 16477
rect 24724 16451 24760 16477
rect 24786 16451 24822 16477
rect 24848 16451 24884 16477
rect 24910 16451 24946 16477
rect 24972 16451 25008 16477
rect 25034 16451 29574 16477
rect 29600 16451 29636 16477
rect 29662 16451 29698 16477
rect 29724 16451 29760 16477
rect 29786 16451 29822 16477
rect 29848 16451 29884 16477
rect 29910 16451 29946 16477
rect 29972 16451 30008 16477
rect 30034 16451 34574 16477
rect 34600 16451 34636 16477
rect 34662 16451 34698 16477
rect 34724 16451 34760 16477
rect 34786 16451 34822 16477
rect 34848 16451 34884 16477
rect 34910 16451 34946 16477
rect 34972 16451 35008 16477
rect 35034 16451 39312 16477
rect 672 16434 39312 16451
rect 7009 16311 7015 16337
rect 7041 16311 7047 16337
rect 8353 16311 8359 16337
rect 8385 16311 8391 16337
rect 10817 16311 10823 16337
rect 10849 16311 10855 16337
rect 12329 16311 12335 16337
rect 12361 16311 12367 16337
rect 13785 16311 13791 16337
rect 13817 16311 13823 16337
rect 15465 16311 15471 16337
rect 15497 16311 15503 16337
rect 6113 16255 6119 16281
rect 6145 16255 6151 16281
rect 7009 16255 7015 16281
rect 7041 16255 7047 16281
rect 7513 16255 7519 16281
rect 7545 16255 7551 16281
rect 8353 16255 8359 16281
rect 8385 16255 8391 16281
rect 9977 16255 9983 16281
rect 10009 16255 10015 16281
rect 10817 16255 10823 16281
rect 10849 16255 10855 16281
rect 11153 16255 11159 16281
rect 11185 16255 11191 16281
rect 12329 16255 12335 16281
rect 12361 16255 12367 16281
rect 12833 16255 12839 16281
rect 12865 16255 12871 16281
rect 13785 16255 13791 16281
rect 13817 16255 13823 16281
rect 14289 16255 14295 16281
rect 14321 16255 14327 16281
rect 15465 16255 15471 16281
rect 15497 16255 15503 16281
rect 672 16085 39312 16102
rect 672 16059 2074 16085
rect 2100 16059 2136 16085
rect 2162 16059 2198 16085
rect 2224 16059 2260 16085
rect 2286 16059 2322 16085
rect 2348 16059 2384 16085
rect 2410 16059 2446 16085
rect 2472 16059 2508 16085
rect 2534 16059 7074 16085
rect 7100 16059 7136 16085
rect 7162 16059 7198 16085
rect 7224 16059 7260 16085
rect 7286 16059 7322 16085
rect 7348 16059 7384 16085
rect 7410 16059 7446 16085
rect 7472 16059 7508 16085
rect 7534 16059 12074 16085
rect 12100 16059 12136 16085
rect 12162 16059 12198 16085
rect 12224 16059 12260 16085
rect 12286 16059 12322 16085
rect 12348 16059 12384 16085
rect 12410 16059 12446 16085
rect 12472 16059 12508 16085
rect 12534 16059 17074 16085
rect 17100 16059 17136 16085
rect 17162 16059 17198 16085
rect 17224 16059 17260 16085
rect 17286 16059 17322 16085
rect 17348 16059 17384 16085
rect 17410 16059 17446 16085
rect 17472 16059 17508 16085
rect 17534 16059 22074 16085
rect 22100 16059 22136 16085
rect 22162 16059 22198 16085
rect 22224 16059 22260 16085
rect 22286 16059 22322 16085
rect 22348 16059 22384 16085
rect 22410 16059 22446 16085
rect 22472 16059 22508 16085
rect 22534 16059 27074 16085
rect 27100 16059 27136 16085
rect 27162 16059 27198 16085
rect 27224 16059 27260 16085
rect 27286 16059 27322 16085
rect 27348 16059 27384 16085
rect 27410 16059 27446 16085
rect 27472 16059 27508 16085
rect 27534 16059 32074 16085
rect 32100 16059 32136 16085
rect 32162 16059 32198 16085
rect 32224 16059 32260 16085
rect 32286 16059 32322 16085
rect 32348 16059 32384 16085
rect 32410 16059 32446 16085
rect 32472 16059 32508 16085
rect 32534 16059 37074 16085
rect 37100 16059 37136 16085
rect 37162 16059 37198 16085
rect 37224 16059 37260 16085
rect 37286 16059 37322 16085
rect 37348 16059 37384 16085
rect 37410 16059 37446 16085
rect 37472 16059 37508 16085
rect 37534 16059 39312 16085
rect 672 16042 39312 16059
rect 5273 15863 5279 15889
rect 5305 15863 5311 15889
rect 6449 15863 6455 15889
rect 6481 15863 6487 15889
rect 7793 15863 7799 15889
rect 7825 15863 7831 15889
rect 8353 15863 8359 15889
rect 8385 15863 8391 15889
rect 8465 15863 8471 15889
rect 8497 15863 8503 15889
rect 9249 15863 9255 15889
rect 9281 15863 9287 15889
rect 10145 15863 10151 15889
rect 10177 15863 10183 15889
rect 11657 15863 11663 15889
rect 11689 15863 11695 15889
rect 12833 15863 12839 15889
rect 12865 15863 12871 15889
rect 13113 15863 13119 15889
rect 13145 15863 13151 15889
rect 14009 15863 14015 15889
rect 14041 15863 14047 15889
rect 15073 15863 15079 15889
rect 15105 15863 15111 15889
rect 15521 15863 15527 15889
rect 15553 15863 15559 15889
rect 16473 15863 16479 15889
rect 16505 15863 16511 15889
rect 16809 15863 16815 15889
rect 16841 15863 16847 15889
rect 16921 15863 16927 15889
rect 16953 15863 16959 15889
rect 6449 15807 6455 15833
rect 6481 15807 6487 15833
rect 10201 15807 10207 15833
rect 10233 15807 10239 15833
rect 12833 15807 12839 15833
rect 12865 15807 12871 15833
rect 14065 15807 14071 15833
rect 14097 15807 14103 15833
rect 15745 15807 15751 15833
rect 15777 15807 15783 15833
rect 672 15693 39312 15710
rect 672 15667 4574 15693
rect 4600 15667 4636 15693
rect 4662 15667 4698 15693
rect 4724 15667 4760 15693
rect 4786 15667 4822 15693
rect 4848 15667 4884 15693
rect 4910 15667 4946 15693
rect 4972 15667 5008 15693
rect 5034 15667 9574 15693
rect 9600 15667 9636 15693
rect 9662 15667 9698 15693
rect 9724 15667 9760 15693
rect 9786 15667 9822 15693
rect 9848 15667 9884 15693
rect 9910 15667 9946 15693
rect 9972 15667 10008 15693
rect 10034 15667 14574 15693
rect 14600 15667 14636 15693
rect 14662 15667 14698 15693
rect 14724 15667 14760 15693
rect 14786 15667 14822 15693
rect 14848 15667 14884 15693
rect 14910 15667 14946 15693
rect 14972 15667 15008 15693
rect 15034 15667 19574 15693
rect 19600 15667 19636 15693
rect 19662 15667 19698 15693
rect 19724 15667 19760 15693
rect 19786 15667 19822 15693
rect 19848 15667 19884 15693
rect 19910 15667 19946 15693
rect 19972 15667 20008 15693
rect 20034 15667 24574 15693
rect 24600 15667 24636 15693
rect 24662 15667 24698 15693
rect 24724 15667 24760 15693
rect 24786 15667 24822 15693
rect 24848 15667 24884 15693
rect 24910 15667 24946 15693
rect 24972 15667 25008 15693
rect 25034 15667 29574 15693
rect 29600 15667 29636 15693
rect 29662 15667 29698 15693
rect 29724 15667 29760 15693
rect 29786 15667 29822 15693
rect 29848 15667 29884 15693
rect 29910 15667 29946 15693
rect 29972 15667 30008 15693
rect 30034 15667 34574 15693
rect 34600 15667 34636 15693
rect 34662 15667 34698 15693
rect 34724 15667 34760 15693
rect 34786 15667 34822 15693
rect 34848 15667 34884 15693
rect 34910 15667 34946 15693
rect 34972 15667 35008 15693
rect 35034 15667 39312 15693
rect 672 15650 39312 15667
rect 6897 15527 6903 15553
rect 6929 15527 6935 15553
rect 8353 15527 8359 15553
rect 8385 15527 8391 15553
rect 10873 15527 10879 15553
rect 10905 15527 10911 15553
rect 12441 15527 12447 15553
rect 12473 15527 12479 15553
rect 14009 15527 14015 15553
rect 14041 15527 14047 15553
rect 15353 15527 15359 15553
rect 15385 15527 15391 15553
rect 5833 15471 5839 15497
rect 5865 15471 5871 15497
rect 6897 15471 6903 15497
rect 6929 15471 6935 15497
rect 7289 15471 7295 15497
rect 7321 15471 7327 15497
rect 8353 15471 8359 15497
rect 8385 15471 8391 15497
rect 9809 15471 9815 15497
rect 9841 15471 9847 15497
rect 10873 15471 10879 15497
rect 10905 15471 10911 15497
rect 11545 15471 11551 15497
rect 11577 15471 11583 15497
rect 12441 15471 12447 15497
rect 12473 15471 12479 15497
rect 13113 15471 13119 15497
rect 13145 15471 13151 15497
rect 14009 15471 14015 15497
rect 14041 15471 14047 15497
rect 14289 15471 14295 15497
rect 14321 15471 14327 15497
rect 15353 15471 15359 15497
rect 15385 15471 15391 15497
rect 672 15301 39312 15318
rect 672 15275 2074 15301
rect 2100 15275 2136 15301
rect 2162 15275 2198 15301
rect 2224 15275 2260 15301
rect 2286 15275 2322 15301
rect 2348 15275 2384 15301
rect 2410 15275 2446 15301
rect 2472 15275 2508 15301
rect 2534 15275 7074 15301
rect 7100 15275 7136 15301
rect 7162 15275 7198 15301
rect 7224 15275 7260 15301
rect 7286 15275 7322 15301
rect 7348 15275 7384 15301
rect 7410 15275 7446 15301
rect 7472 15275 7508 15301
rect 7534 15275 12074 15301
rect 12100 15275 12136 15301
rect 12162 15275 12198 15301
rect 12224 15275 12260 15301
rect 12286 15275 12322 15301
rect 12348 15275 12384 15301
rect 12410 15275 12446 15301
rect 12472 15275 12508 15301
rect 12534 15275 17074 15301
rect 17100 15275 17136 15301
rect 17162 15275 17198 15301
rect 17224 15275 17260 15301
rect 17286 15275 17322 15301
rect 17348 15275 17384 15301
rect 17410 15275 17446 15301
rect 17472 15275 17508 15301
rect 17534 15275 22074 15301
rect 22100 15275 22136 15301
rect 22162 15275 22198 15301
rect 22224 15275 22260 15301
rect 22286 15275 22322 15301
rect 22348 15275 22384 15301
rect 22410 15275 22446 15301
rect 22472 15275 22508 15301
rect 22534 15275 27074 15301
rect 27100 15275 27136 15301
rect 27162 15275 27198 15301
rect 27224 15275 27260 15301
rect 27286 15275 27322 15301
rect 27348 15275 27384 15301
rect 27410 15275 27446 15301
rect 27472 15275 27508 15301
rect 27534 15275 32074 15301
rect 32100 15275 32136 15301
rect 32162 15275 32198 15301
rect 32224 15275 32260 15301
rect 32286 15275 32322 15301
rect 32348 15275 32384 15301
rect 32410 15275 32446 15301
rect 32472 15275 32508 15301
rect 32534 15275 37074 15301
rect 37100 15275 37136 15301
rect 37162 15275 37198 15301
rect 37224 15275 37260 15301
rect 37286 15275 37322 15301
rect 37348 15275 37384 15301
rect 37410 15275 37446 15301
rect 37472 15275 37508 15301
rect 37534 15275 39312 15301
rect 672 15258 39312 15275
rect 1801 15079 1807 15105
rect 1833 15079 1839 15105
rect 1913 15079 1919 15105
rect 1945 15079 1951 15105
rect 2417 15079 2423 15105
rect 2449 15079 2455 15105
rect 3817 15079 3823 15105
rect 3849 15079 3855 15105
rect 4377 15079 4383 15105
rect 4409 15079 4415 15105
rect 4489 15079 4495 15105
rect 4521 15079 4527 15105
rect 5273 15079 5279 15105
rect 5305 15079 5311 15105
rect 6393 15079 6399 15105
rect 6425 15079 6431 15105
rect 7793 15079 7799 15105
rect 7825 15079 7831 15105
rect 8969 15079 8975 15105
rect 9001 15079 9007 15105
rect 9249 15079 9255 15105
rect 9281 15079 9287 15105
rect 10425 15079 10431 15105
rect 10457 15079 10463 15105
rect 11937 15079 11943 15105
rect 11969 15079 11975 15105
rect 12833 15079 12839 15105
rect 12865 15079 12871 15105
rect 13113 15079 13119 15105
rect 13145 15079 13151 15105
rect 14009 15079 14015 15105
rect 14041 15079 14047 15105
rect 14793 15079 14799 15105
rect 14825 15079 14831 15105
rect 15353 15079 15359 15105
rect 15385 15079 15391 15105
rect 15521 15079 15527 15105
rect 15553 15079 15559 15105
rect 16473 15079 16479 15105
rect 16505 15079 16511 15105
rect 17425 15079 17431 15105
rect 17457 15079 17463 15105
rect 18769 15079 18775 15105
rect 18801 15079 18807 15105
rect 19329 15079 19335 15105
rect 19361 15079 19367 15105
rect 19441 15079 19447 15105
rect 19473 15079 19479 15105
rect 6393 15023 6399 15049
rect 6425 15023 6431 15049
rect 8969 15023 8975 15049
rect 9001 15023 9007 15049
rect 10425 15023 10431 15049
rect 10457 15023 10463 15049
rect 12833 15023 12839 15049
rect 12865 15023 12871 15049
rect 14065 15023 14071 15049
rect 14097 15023 14103 15049
rect 17425 15023 17431 15049
rect 17457 15023 17463 15049
rect 672 14909 39312 14926
rect 672 14883 4574 14909
rect 4600 14883 4636 14909
rect 4662 14883 4698 14909
rect 4724 14883 4760 14909
rect 4786 14883 4822 14909
rect 4848 14883 4884 14909
rect 4910 14883 4946 14909
rect 4972 14883 5008 14909
rect 5034 14883 9574 14909
rect 9600 14883 9636 14909
rect 9662 14883 9698 14909
rect 9724 14883 9760 14909
rect 9786 14883 9822 14909
rect 9848 14883 9884 14909
rect 9910 14883 9946 14909
rect 9972 14883 10008 14909
rect 10034 14883 14574 14909
rect 14600 14883 14636 14909
rect 14662 14883 14698 14909
rect 14724 14883 14760 14909
rect 14786 14883 14822 14909
rect 14848 14883 14884 14909
rect 14910 14883 14946 14909
rect 14972 14883 15008 14909
rect 15034 14883 19574 14909
rect 19600 14883 19636 14909
rect 19662 14883 19698 14909
rect 19724 14883 19760 14909
rect 19786 14883 19822 14909
rect 19848 14883 19884 14909
rect 19910 14883 19946 14909
rect 19972 14883 20008 14909
rect 20034 14883 24574 14909
rect 24600 14883 24636 14909
rect 24662 14883 24698 14909
rect 24724 14883 24760 14909
rect 24786 14883 24822 14909
rect 24848 14883 24884 14909
rect 24910 14883 24946 14909
rect 24972 14883 25008 14909
rect 25034 14883 29574 14909
rect 29600 14883 29636 14909
rect 29662 14883 29698 14909
rect 29724 14883 29760 14909
rect 29786 14883 29822 14909
rect 29848 14883 29884 14909
rect 29910 14883 29946 14909
rect 29972 14883 30008 14909
rect 30034 14883 34574 14909
rect 34600 14883 34636 14909
rect 34662 14883 34698 14909
rect 34724 14883 34760 14909
rect 34786 14883 34822 14909
rect 34848 14883 34884 14909
rect 34910 14883 34946 14909
rect 34972 14883 35008 14909
rect 35034 14883 39312 14909
rect 672 14866 39312 14883
rect 1857 14743 1863 14769
rect 1889 14743 1895 14769
rect 4489 14743 4495 14769
rect 4521 14743 4527 14769
rect 6897 14743 6903 14769
rect 6929 14743 6935 14769
rect 8353 14743 8359 14769
rect 8385 14743 8391 14769
rect 10873 14743 10879 14769
rect 10905 14743 10911 14769
rect 12441 14743 12447 14769
rect 12473 14743 12479 14769
rect 14009 14743 14015 14769
rect 14041 14743 14047 14769
rect 15297 14743 15303 14769
rect 15329 14743 15335 14769
rect 17761 14743 17767 14769
rect 17793 14743 17799 14769
rect 1857 14687 1863 14713
rect 1889 14687 1895 14713
rect 3033 14687 3039 14713
rect 3065 14687 3071 14713
rect 3593 14687 3599 14713
rect 3625 14687 3631 14713
rect 4489 14687 4495 14713
rect 4521 14687 4527 14713
rect 5833 14687 5839 14713
rect 5865 14687 5871 14713
rect 6897 14687 6903 14713
rect 6929 14687 6935 14713
rect 7289 14687 7295 14713
rect 7321 14687 7327 14713
rect 8353 14687 8359 14713
rect 8385 14687 8391 14713
rect 9809 14687 9815 14713
rect 9841 14687 9847 14713
rect 10873 14687 10879 14713
rect 10905 14687 10911 14713
rect 11545 14687 11551 14713
rect 11577 14687 11583 14713
rect 12441 14687 12447 14713
rect 12473 14687 12479 14713
rect 13113 14687 13119 14713
rect 13145 14687 13151 14713
rect 14009 14687 14015 14713
rect 14041 14687 14047 14713
rect 14345 14687 14351 14713
rect 14377 14687 14383 14713
rect 15297 14687 15303 14713
rect 15329 14687 15335 14713
rect 17089 14687 17095 14713
rect 17121 14687 17127 14713
rect 17761 14687 17767 14713
rect 17793 14687 17799 14713
rect 18265 14687 18271 14713
rect 18297 14687 18303 14713
rect 18713 14687 18719 14713
rect 18745 14687 18751 14713
rect 18937 14687 18943 14713
rect 18969 14687 18975 14713
rect 672 14517 39312 14534
rect 672 14491 2074 14517
rect 2100 14491 2136 14517
rect 2162 14491 2198 14517
rect 2224 14491 2260 14517
rect 2286 14491 2322 14517
rect 2348 14491 2384 14517
rect 2410 14491 2446 14517
rect 2472 14491 2508 14517
rect 2534 14491 7074 14517
rect 7100 14491 7136 14517
rect 7162 14491 7198 14517
rect 7224 14491 7260 14517
rect 7286 14491 7322 14517
rect 7348 14491 7384 14517
rect 7410 14491 7446 14517
rect 7472 14491 7508 14517
rect 7534 14491 12074 14517
rect 12100 14491 12136 14517
rect 12162 14491 12198 14517
rect 12224 14491 12260 14517
rect 12286 14491 12322 14517
rect 12348 14491 12384 14517
rect 12410 14491 12446 14517
rect 12472 14491 12508 14517
rect 12534 14491 17074 14517
rect 17100 14491 17136 14517
rect 17162 14491 17198 14517
rect 17224 14491 17260 14517
rect 17286 14491 17322 14517
rect 17348 14491 17384 14517
rect 17410 14491 17446 14517
rect 17472 14491 17508 14517
rect 17534 14491 22074 14517
rect 22100 14491 22136 14517
rect 22162 14491 22198 14517
rect 22224 14491 22260 14517
rect 22286 14491 22322 14517
rect 22348 14491 22384 14517
rect 22410 14491 22446 14517
rect 22472 14491 22508 14517
rect 22534 14491 27074 14517
rect 27100 14491 27136 14517
rect 27162 14491 27198 14517
rect 27224 14491 27260 14517
rect 27286 14491 27322 14517
rect 27348 14491 27384 14517
rect 27410 14491 27446 14517
rect 27472 14491 27508 14517
rect 27534 14491 32074 14517
rect 32100 14491 32136 14517
rect 32162 14491 32198 14517
rect 32224 14491 32260 14517
rect 32286 14491 32322 14517
rect 32348 14491 32384 14517
rect 32410 14491 32446 14517
rect 32472 14491 32508 14517
rect 32534 14491 37074 14517
rect 37100 14491 37136 14517
rect 37162 14491 37198 14517
rect 37224 14491 37260 14517
rect 37286 14491 37322 14517
rect 37348 14491 37384 14517
rect 37410 14491 37446 14517
rect 37472 14491 37508 14517
rect 37534 14491 39312 14517
rect 672 14474 39312 14491
rect 1801 14295 1807 14321
rect 1833 14295 1839 14321
rect 1913 14295 1919 14321
rect 1945 14295 1951 14321
rect 2417 14295 2423 14321
rect 2449 14295 2455 14321
rect 3817 14295 3823 14321
rect 3849 14295 3855 14321
rect 4993 14295 4999 14321
rect 5025 14295 5031 14321
rect 5273 14295 5279 14321
rect 5305 14295 5311 14321
rect 6393 14295 6399 14321
rect 6425 14295 6431 14321
rect 7793 14295 7799 14321
rect 7825 14295 7831 14321
rect 8969 14295 8975 14321
rect 9001 14295 9007 14321
rect 9249 14295 9255 14321
rect 9281 14295 9287 14321
rect 10425 14295 10431 14321
rect 10457 14295 10463 14321
rect 11993 14295 11999 14321
rect 12025 14295 12031 14321
rect 12889 14295 12895 14321
rect 12921 14295 12927 14321
rect 13225 14295 13231 14321
rect 13257 14295 13263 14321
rect 14009 14295 14015 14321
rect 14041 14295 14047 14321
rect 14793 14295 14799 14321
rect 14825 14295 14831 14321
rect 15297 14295 15303 14321
rect 15329 14295 15335 14321
rect 15465 14295 15471 14321
rect 15497 14295 15503 14321
rect 16529 14295 16535 14321
rect 16561 14295 16567 14321
rect 17425 14295 17431 14321
rect 17457 14295 17463 14321
rect 18769 14295 18775 14321
rect 18801 14295 18807 14321
rect 19329 14295 19335 14321
rect 19361 14295 19367 14321
rect 19441 14295 19447 14321
rect 19473 14295 19479 14321
rect 20225 14295 20231 14321
rect 20257 14295 20263 14321
rect 21009 14295 21015 14321
rect 21041 14295 21047 14321
rect 23025 14295 23031 14321
rect 23057 14295 23063 14321
rect 23865 14295 23871 14321
rect 23897 14295 23903 14321
rect 24425 14295 24431 14321
rect 24457 14295 24463 14321
rect 25153 14295 25159 14321
rect 25185 14295 25191 14321
rect 4993 14239 4999 14265
rect 5025 14239 5031 14265
rect 6393 14239 6399 14265
rect 6425 14239 6431 14265
rect 8969 14239 8975 14265
rect 9001 14239 9007 14265
rect 10425 14239 10431 14265
rect 10457 14239 10463 14265
rect 12889 14239 12895 14265
rect 12921 14239 12927 14265
rect 14177 14239 14183 14265
rect 14209 14239 14215 14265
rect 17425 14239 17431 14265
rect 17457 14239 17463 14265
rect 21177 14239 21183 14265
rect 21209 14239 21215 14265
rect 23865 14239 23871 14265
rect 23897 14239 23903 14265
rect 25209 14239 25215 14265
rect 25241 14239 25247 14265
rect 672 14125 39312 14142
rect 672 14099 4574 14125
rect 4600 14099 4636 14125
rect 4662 14099 4698 14125
rect 4724 14099 4760 14125
rect 4786 14099 4822 14125
rect 4848 14099 4884 14125
rect 4910 14099 4946 14125
rect 4972 14099 5008 14125
rect 5034 14099 9574 14125
rect 9600 14099 9636 14125
rect 9662 14099 9698 14125
rect 9724 14099 9760 14125
rect 9786 14099 9822 14125
rect 9848 14099 9884 14125
rect 9910 14099 9946 14125
rect 9972 14099 10008 14125
rect 10034 14099 14574 14125
rect 14600 14099 14636 14125
rect 14662 14099 14698 14125
rect 14724 14099 14760 14125
rect 14786 14099 14822 14125
rect 14848 14099 14884 14125
rect 14910 14099 14946 14125
rect 14972 14099 15008 14125
rect 15034 14099 19574 14125
rect 19600 14099 19636 14125
rect 19662 14099 19698 14125
rect 19724 14099 19760 14125
rect 19786 14099 19822 14125
rect 19848 14099 19884 14125
rect 19910 14099 19946 14125
rect 19972 14099 20008 14125
rect 20034 14099 24574 14125
rect 24600 14099 24636 14125
rect 24662 14099 24698 14125
rect 24724 14099 24760 14125
rect 24786 14099 24822 14125
rect 24848 14099 24884 14125
rect 24910 14099 24946 14125
rect 24972 14099 25008 14125
rect 25034 14099 29574 14125
rect 29600 14099 29636 14125
rect 29662 14099 29698 14125
rect 29724 14099 29760 14125
rect 29786 14099 29822 14125
rect 29848 14099 29884 14125
rect 29910 14099 29946 14125
rect 29972 14099 30008 14125
rect 30034 14099 34574 14125
rect 34600 14099 34636 14125
rect 34662 14099 34698 14125
rect 34724 14099 34760 14125
rect 34786 14099 34822 14125
rect 34848 14099 34884 14125
rect 34910 14099 34946 14125
rect 34972 14099 35008 14125
rect 35034 14099 39312 14125
rect 672 14082 39312 14099
rect 4489 13959 4495 13985
rect 4521 13959 4527 13985
rect 6897 13959 6903 13985
rect 6929 13959 6935 13985
rect 8465 13959 8471 13985
rect 8497 13959 8503 13985
rect 10873 13959 10879 13985
rect 10905 13959 10911 13985
rect 12441 13959 12447 13985
rect 12473 13959 12479 13985
rect 14009 13959 14015 13985
rect 14041 13959 14047 13985
rect 15465 13959 15471 13985
rect 15497 13959 15503 13985
rect 17761 13959 17767 13985
rect 17793 13959 17799 13985
rect 19441 13959 19447 13985
rect 19473 13959 19479 13985
rect 21737 13959 21743 13985
rect 21769 13959 21775 13985
rect 23417 13959 23423 13985
rect 23449 13959 23455 13985
rect 2361 13903 2367 13929
rect 2393 13903 2399 13929
rect 2473 13903 2479 13929
rect 2505 13903 2511 13929
rect 3033 13903 3039 13929
rect 3065 13903 3071 13929
rect 3369 13903 3375 13929
rect 3401 13903 3407 13929
rect 4489 13903 4495 13929
rect 4521 13903 4527 13929
rect 5833 13903 5839 13929
rect 5865 13903 5871 13929
rect 6897 13903 6903 13929
rect 6929 13903 6935 13929
rect 7569 13903 7575 13929
rect 7601 13903 7607 13929
rect 8465 13903 8471 13929
rect 8497 13903 8503 13929
rect 9809 13903 9815 13929
rect 9841 13903 9847 13929
rect 10873 13903 10879 13929
rect 10905 13903 10911 13929
rect 11545 13903 11551 13929
rect 11577 13903 11583 13929
rect 12441 13903 12447 13929
rect 12473 13903 12479 13929
rect 13113 13903 13119 13929
rect 13145 13903 13151 13929
rect 14009 13903 14015 13929
rect 14041 13903 14047 13929
rect 14569 13903 14575 13929
rect 14601 13903 14607 13929
rect 15465 13903 15471 13929
rect 15497 13903 15503 13929
rect 16977 13903 16983 13929
rect 17009 13903 17015 13929
rect 17761 13903 17767 13929
rect 17793 13903 17799 13929
rect 18545 13903 18551 13929
rect 18577 13903 18583 13929
rect 19441 13903 19447 13929
rect 19473 13903 19479 13929
rect 20785 13903 20791 13929
rect 20817 13903 20823 13929
rect 21737 13903 21743 13929
rect 21769 13903 21775 13929
rect 22521 13903 22527 13929
rect 22553 13903 22559 13929
rect 23417 13903 23423 13929
rect 23449 13903 23455 13929
rect 25041 13903 25047 13929
rect 25073 13903 25079 13929
rect 25209 13903 25215 13929
rect 25241 13903 25247 13929
rect 25433 13903 25439 13929
rect 25465 13903 25471 13929
rect 672 13733 39312 13750
rect 672 13707 2074 13733
rect 2100 13707 2136 13733
rect 2162 13707 2198 13733
rect 2224 13707 2260 13733
rect 2286 13707 2322 13733
rect 2348 13707 2384 13733
rect 2410 13707 2446 13733
rect 2472 13707 2508 13733
rect 2534 13707 7074 13733
rect 7100 13707 7136 13733
rect 7162 13707 7198 13733
rect 7224 13707 7260 13733
rect 7286 13707 7322 13733
rect 7348 13707 7384 13733
rect 7410 13707 7446 13733
rect 7472 13707 7508 13733
rect 7534 13707 12074 13733
rect 12100 13707 12136 13733
rect 12162 13707 12198 13733
rect 12224 13707 12260 13733
rect 12286 13707 12322 13733
rect 12348 13707 12384 13733
rect 12410 13707 12446 13733
rect 12472 13707 12508 13733
rect 12534 13707 17074 13733
rect 17100 13707 17136 13733
rect 17162 13707 17198 13733
rect 17224 13707 17260 13733
rect 17286 13707 17322 13733
rect 17348 13707 17384 13733
rect 17410 13707 17446 13733
rect 17472 13707 17508 13733
rect 17534 13707 22074 13733
rect 22100 13707 22136 13733
rect 22162 13707 22198 13733
rect 22224 13707 22260 13733
rect 22286 13707 22322 13733
rect 22348 13707 22384 13733
rect 22410 13707 22446 13733
rect 22472 13707 22508 13733
rect 22534 13707 27074 13733
rect 27100 13707 27136 13733
rect 27162 13707 27198 13733
rect 27224 13707 27260 13733
rect 27286 13707 27322 13733
rect 27348 13707 27384 13733
rect 27410 13707 27446 13733
rect 27472 13707 27508 13733
rect 27534 13707 32074 13733
rect 32100 13707 32136 13733
rect 32162 13707 32198 13733
rect 32224 13707 32260 13733
rect 32286 13707 32322 13733
rect 32348 13707 32384 13733
rect 32410 13707 32446 13733
rect 32472 13707 32508 13733
rect 32534 13707 37074 13733
rect 37100 13707 37136 13733
rect 37162 13707 37198 13733
rect 37224 13707 37260 13733
rect 37286 13707 37322 13733
rect 37348 13707 37384 13733
rect 37410 13707 37446 13733
rect 37472 13707 37508 13733
rect 37534 13707 39312 13733
rect 672 13690 39312 13707
rect 1801 13511 1807 13537
rect 1833 13511 1839 13537
rect 1913 13511 1919 13537
rect 1945 13511 1951 13537
rect 2473 13511 2479 13537
rect 2505 13511 2511 13537
rect 3817 13511 3823 13537
rect 3849 13511 3855 13537
rect 4377 13511 4383 13537
rect 4409 13511 4415 13537
rect 4489 13511 4495 13537
rect 4521 13511 4527 13537
rect 5273 13511 5279 13537
rect 5305 13511 5311 13537
rect 6393 13511 6399 13537
rect 6425 13511 6431 13537
rect 7793 13511 7799 13537
rect 7825 13511 7831 13537
rect 8353 13511 8359 13537
rect 8385 13511 8391 13537
rect 8465 13511 8471 13537
rect 8497 13511 8503 13537
rect 9249 13511 9255 13537
rect 9281 13511 9287 13537
rect 10425 13511 10431 13537
rect 10457 13511 10463 13537
rect 11209 13511 11215 13537
rect 11241 13511 11247 13537
rect 12105 13511 12111 13537
rect 12137 13511 12143 13537
rect 12665 13511 12671 13537
rect 12697 13511 12703 13537
rect 13393 13511 13399 13537
rect 13425 13511 13431 13537
rect 14793 13511 14799 13537
rect 14825 13511 14831 13537
rect 15857 13511 15863 13537
rect 15889 13511 15895 13537
rect 16529 13511 16535 13537
rect 16561 13511 16567 13537
rect 17425 13511 17431 13537
rect 17457 13511 17463 13537
rect 19049 13511 19055 13537
rect 19081 13511 19087 13537
rect 19329 13511 19335 13537
rect 19361 13511 19367 13537
rect 19441 13511 19447 13537
rect 19473 13511 19479 13537
rect 20225 13511 20231 13537
rect 20257 13511 20263 13537
rect 21009 13511 21015 13537
rect 21041 13511 21047 13537
rect 23025 13511 23031 13537
rect 23057 13511 23063 13537
rect 23865 13511 23871 13537
rect 23897 13511 23903 13537
rect 24425 13511 24431 13537
rect 24457 13511 24463 13537
rect 25209 13511 25215 13537
rect 25241 13511 25247 13537
rect 6393 13455 6399 13481
rect 6425 13455 6431 13481
rect 10425 13455 10431 13481
rect 10457 13455 10463 13481
rect 12105 13455 12111 13481
rect 12137 13455 12143 13481
rect 13393 13455 13399 13481
rect 13425 13455 13431 13481
rect 15857 13455 15863 13481
rect 15889 13455 15895 13481
rect 17425 13455 17431 13481
rect 17457 13455 17463 13481
rect 21177 13455 21183 13481
rect 21209 13455 21215 13481
rect 23865 13455 23871 13481
rect 23897 13455 23903 13481
rect 25209 13455 25215 13481
rect 25241 13455 25247 13481
rect 672 13341 39312 13358
rect 672 13315 4574 13341
rect 4600 13315 4636 13341
rect 4662 13315 4698 13341
rect 4724 13315 4760 13341
rect 4786 13315 4822 13341
rect 4848 13315 4884 13341
rect 4910 13315 4946 13341
rect 4972 13315 5008 13341
rect 5034 13315 9574 13341
rect 9600 13315 9636 13341
rect 9662 13315 9698 13341
rect 9724 13315 9760 13341
rect 9786 13315 9822 13341
rect 9848 13315 9884 13341
rect 9910 13315 9946 13341
rect 9972 13315 10008 13341
rect 10034 13315 14574 13341
rect 14600 13315 14636 13341
rect 14662 13315 14698 13341
rect 14724 13315 14760 13341
rect 14786 13315 14822 13341
rect 14848 13315 14884 13341
rect 14910 13315 14946 13341
rect 14972 13315 15008 13341
rect 15034 13315 19574 13341
rect 19600 13315 19636 13341
rect 19662 13315 19698 13341
rect 19724 13315 19760 13341
rect 19786 13315 19822 13341
rect 19848 13315 19884 13341
rect 19910 13315 19946 13341
rect 19972 13315 20008 13341
rect 20034 13315 24574 13341
rect 24600 13315 24636 13341
rect 24662 13315 24698 13341
rect 24724 13315 24760 13341
rect 24786 13315 24822 13341
rect 24848 13315 24884 13341
rect 24910 13315 24946 13341
rect 24972 13315 25008 13341
rect 25034 13315 29574 13341
rect 29600 13315 29636 13341
rect 29662 13315 29698 13341
rect 29724 13315 29760 13341
rect 29786 13315 29822 13341
rect 29848 13315 29884 13341
rect 29910 13315 29946 13341
rect 29972 13315 30008 13341
rect 30034 13315 34574 13341
rect 34600 13315 34636 13341
rect 34662 13315 34698 13341
rect 34724 13315 34760 13341
rect 34786 13315 34822 13341
rect 34848 13315 34884 13341
rect 34910 13315 34946 13341
rect 34972 13315 35008 13341
rect 35034 13315 39312 13341
rect 672 13298 39312 13315
rect 4489 13175 4495 13201
rect 4521 13175 4527 13201
rect 6953 13175 6959 13201
rect 6985 13175 6991 13201
rect 8353 13175 8359 13201
rect 8385 13175 8391 13201
rect 10873 13175 10879 13201
rect 10905 13175 10911 13201
rect 12441 13175 12447 13201
rect 12473 13175 12479 13201
rect 14009 13175 14015 13201
rect 14041 13175 14047 13201
rect 15297 13175 15303 13201
rect 15329 13175 15335 13201
rect 17761 13175 17767 13201
rect 17793 13175 17799 13201
rect 19441 13175 19447 13201
rect 19473 13175 19479 13201
rect 23417 13175 23423 13201
rect 23449 13175 23455 13201
rect 25937 13175 25943 13201
rect 25969 13175 25975 13201
rect 2361 13119 2367 13145
rect 2393 13119 2399 13145
rect 2585 13119 2591 13145
rect 2617 13119 2623 13145
rect 2753 13119 2759 13145
rect 2785 13119 2791 13145
rect 3313 13119 3319 13145
rect 3345 13119 3351 13145
rect 4489 13119 4495 13145
rect 4521 13119 4527 13145
rect 5833 13119 5839 13145
rect 5865 13119 5871 13145
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 7569 13119 7575 13145
rect 7601 13119 7607 13145
rect 8353 13119 8359 13145
rect 8385 13119 8391 13145
rect 9809 13119 9815 13145
rect 9841 13119 9847 13145
rect 10873 13119 10879 13145
rect 10905 13119 10911 13145
rect 11545 13119 11551 13145
rect 11577 13119 11583 13145
rect 12441 13119 12447 13145
rect 12473 13119 12479 13145
rect 13113 13119 13119 13145
rect 13145 13119 13151 13145
rect 14009 13119 14015 13145
rect 14041 13119 14047 13145
rect 14457 13119 14463 13145
rect 14489 13119 14495 13145
rect 15297 13119 15303 13145
rect 15329 13119 15335 13145
rect 17089 13119 17095 13145
rect 17121 13119 17127 13145
rect 17593 13119 17599 13145
rect 17625 13119 17631 13145
rect 18545 13119 18551 13145
rect 18577 13119 18583 13145
rect 19441 13119 19447 13145
rect 19473 13119 19479 13145
rect 20953 13119 20959 13145
rect 20985 13119 20991 13145
rect 21289 13119 21295 13145
rect 21321 13119 21327 13145
rect 21457 13119 21463 13145
rect 21489 13119 21495 13145
rect 22521 13119 22527 13145
rect 22553 13119 22559 13145
rect 23417 13119 23423 13145
rect 23449 13119 23455 13145
rect 25041 13119 25047 13145
rect 25073 13119 25079 13145
rect 25937 13119 25943 13145
rect 25969 13119 25975 13145
rect 672 12949 39312 12966
rect 672 12923 2074 12949
rect 2100 12923 2136 12949
rect 2162 12923 2198 12949
rect 2224 12923 2260 12949
rect 2286 12923 2322 12949
rect 2348 12923 2384 12949
rect 2410 12923 2446 12949
rect 2472 12923 2508 12949
rect 2534 12923 7074 12949
rect 7100 12923 7136 12949
rect 7162 12923 7198 12949
rect 7224 12923 7260 12949
rect 7286 12923 7322 12949
rect 7348 12923 7384 12949
rect 7410 12923 7446 12949
rect 7472 12923 7508 12949
rect 7534 12923 12074 12949
rect 12100 12923 12136 12949
rect 12162 12923 12198 12949
rect 12224 12923 12260 12949
rect 12286 12923 12322 12949
rect 12348 12923 12384 12949
rect 12410 12923 12446 12949
rect 12472 12923 12508 12949
rect 12534 12923 17074 12949
rect 17100 12923 17136 12949
rect 17162 12923 17198 12949
rect 17224 12923 17260 12949
rect 17286 12923 17322 12949
rect 17348 12923 17384 12949
rect 17410 12923 17446 12949
rect 17472 12923 17508 12949
rect 17534 12923 22074 12949
rect 22100 12923 22136 12949
rect 22162 12923 22198 12949
rect 22224 12923 22260 12949
rect 22286 12923 22322 12949
rect 22348 12923 22384 12949
rect 22410 12923 22446 12949
rect 22472 12923 22508 12949
rect 22534 12923 27074 12949
rect 27100 12923 27136 12949
rect 27162 12923 27198 12949
rect 27224 12923 27260 12949
rect 27286 12923 27322 12949
rect 27348 12923 27384 12949
rect 27410 12923 27446 12949
rect 27472 12923 27508 12949
rect 27534 12923 32074 12949
rect 32100 12923 32136 12949
rect 32162 12923 32198 12949
rect 32224 12923 32260 12949
rect 32286 12923 32322 12949
rect 32348 12923 32384 12949
rect 32410 12923 32446 12949
rect 32472 12923 32508 12949
rect 32534 12923 37074 12949
rect 37100 12923 37136 12949
rect 37162 12923 37198 12949
rect 37224 12923 37260 12949
rect 37286 12923 37322 12949
rect 37348 12923 37384 12949
rect 37410 12923 37446 12949
rect 37472 12923 37508 12949
rect 37534 12923 39312 12949
rect 672 12906 39312 12923
rect 1801 12727 1807 12753
rect 1833 12727 1839 12753
rect 1969 12727 1975 12753
rect 2001 12727 2007 12753
rect 2193 12727 2199 12753
rect 2225 12727 2231 12753
rect 4097 12727 4103 12753
rect 4129 12727 4135 12753
rect 4377 12727 4383 12753
rect 4409 12727 4415 12753
rect 4489 12727 4495 12753
rect 4521 12727 4527 12753
rect 5273 12727 5279 12753
rect 5305 12727 5311 12753
rect 6449 12727 6455 12753
rect 6481 12727 6487 12753
rect 7793 12727 7799 12753
rect 7825 12727 7831 12753
rect 8353 12727 8359 12753
rect 8385 12727 8391 12753
rect 8465 12727 8471 12753
rect 8497 12727 8503 12753
rect 9249 12727 9255 12753
rect 9281 12727 9287 12753
rect 10425 12727 10431 12753
rect 10457 12727 10463 12753
rect 11993 12727 11999 12753
rect 12025 12727 12031 12753
rect 12889 12727 12895 12753
rect 12921 12727 12927 12753
rect 13337 12727 13343 12753
rect 13369 12727 13375 12753
rect 14233 12727 14239 12753
rect 14265 12727 14271 12753
rect 14793 12727 14799 12753
rect 14825 12727 14831 12753
rect 15297 12727 15303 12753
rect 15329 12727 15335 12753
rect 15465 12727 15471 12753
rect 15497 12727 15503 12753
rect 16529 12727 16535 12753
rect 16561 12727 16567 12753
rect 17425 12727 17431 12753
rect 17457 12727 17463 12753
rect 19049 12727 19055 12753
rect 19081 12727 19087 12753
rect 19329 12727 19335 12753
rect 19361 12727 19367 12753
rect 19441 12727 19447 12753
rect 19473 12727 19479 12753
rect 20505 12727 20511 12753
rect 20537 12727 20543 12753
rect 21289 12727 21295 12753
rect 21321 12727 21327 12753
rect 22969 12727 22975 12753
rect 23001 12727 23007 12753
rect 23865 12727 23871 12753
rect 23897 12727 23903 12753
rect 24481 12727 24487 12753
rect 24513 12727 24519 12753
rect 25153 12727 25159 12753
rect 25185 12727 25191 12753
rect 29633 12727 29639 12753
rect 29665 12727 29671 12753
rect 29745 12727 29751 12753
rect 29777 12727 29783 12753
rect 30193 12727 30199 12753
rect 30225 12727 30231 12753
rect 6449 12671 6455 12697
rect 6481 12671 6487 12697
rect 10425 12671 10431 12697
rect 10457 12671 10463 12697
rect 12889 12671 12895 12697
rect 12921 12671 12927 12697
rect 14233 12671 14239 12697
rect 14265 12671 14271 12697
rect 17425 12671 17431 12697
rect 17457 12671 17463 12697
rect 21289 12671 21295 12697
rect 21321 12671 21327 12697
rect 23865 12671 23871 12697
rect 23897 12671 23903 12697
rect 25153 12671 25159 12697
rect 25185 12671 25191 12697
rect 672 12557 39312 12574
rect 672 12531 4574 12557
rect 4600 12531 4636 12557
rect 4662 12531 4698 12557
rect 4724 12531 4760 12557
rect 4786 12531 4822 12557
rect 4848 12531 4884 12557
rect 4910 12531 4946 12557
rect 4972 12531 5008 12557
rect 5034 12531 9574 12557
rect 9600 12531 9636 12557
rect 9662 12531 9698 12557
rect 9724 12531 9760 12557
rect 9786 12531 9822 12557
rect 9848 12531 9884 12557
rect 9910 12531 9946 12557
rect 9972 12531 10008 12557
rect 10034 12531 14574 12557
rect 14600 12531 14636 12557
rect 14662 12531 14698 12557
rect 14724 12531 14760 12557
rect 14786 12531 14822 12557
rect 14848 12531 14884 12557
rect 14910 12531 14946 12557
rect 14972 12531 15008 12557
rect 15034 12531 19574 12557
rect 19600 12531 19636 12557
rect 19662 12531 19698 12557
rect 19724 12531 19760 12557
rect 19786 12531 19822 12557
rect 19848 12531 19884 12557
rect 19910 12531 19946 12557
rect 19972 12531 20008 12557
rect 20034 12531 24574 12557
rect 24600 12531 24636 12557
rect 24662 12531 24698 12557
rect 24724 12531 24760 12557
rect 24786 12531 24822 12557
rect 24848 12531 24884 12557
rect 24910 12531 24946 12557
rect 24972 12531 25008 12557
rect 25034 12531 29574 12557
rect 29600 12531 29636 12557
rect 29662 12531 29698 12557
rect 29724 12531 29760 12557
rect 29786 12531 29822 12557
rect 29848 12531 29884 12557
rect 29910 12531 29946 12557
rect 29972 12531 30008 12557
rect 30034 12531 34574 12557
rect 34600 12531 34636 12557
rect 34662 12531 34698 12557
rect 34724 12531 34760 12557
rect 34786 12531 34822 12557
rect 34848 12531 34884 12557
rect 34910 12531 34946 12557
rect 34972 12531 35008 12557
rect 35034 12531 39312 12557
rect 672 12514 39312 12531
rect 1857 12391 1863 12417
rect 1889 12391 1895 12417
rect 4489 12391 4495 12417
rect 4521 12391 4527 12417
rect 7009 12391 7015 12417
rect 7041 12391 7047 12417
rect 8353 12391 8359 12417
rect 8385 12391 8391 12417
rect 10873 12391 10879 12417
rect 10905 12391 10911 12417
rect 12441 12391 12447 12417
rect 12473 12391 12479 12417
rect 14401 12391 14407 12417
rect 14433 12391 14439 12417
rect 17985 12391 17991 12417
rect 18017 12391 18023 12417
rect 19441 12391 19447 12417
rect 19473 12391 19479 12417
rect 21793 12391 21799 12417
rect 21825 12391 21831 12417
rect 23417 12391 23423 12417
rect 23449 12391 23455 12417
rect 25937 12391 25943 12417
rect 25969 12391 25975 12417
rect 27393 12391 27399 12417
rect 27425 12391 27431 12417
rect 31593 12391 31599 12417
rect 31625 12391 31631 12417
rect 1857 12335 1863 12361
rect 1889 12335 1895 12361
rect 2753 12335 2759 12361
rect 2785 12335 2791 12361
rect 3593 12335 3599 12361
rect 3625 12335 3631 12361
rect 4489 12335 4495 12361
rect 4521 12335 4527 12361
rect 5833 12335 5839 12361
rect 5865 12335 5871 12361
rect 7009 12335 7015 12361
rect 7041 12335 7047 12361
rect 7569 12335 7575 12361
rect 7601 12335 7607 12361
rect 8353 12335 8359 12361
rect 8385 12335 8391 12361
rect 9809 12335 9815 12361
rect 9841 12335 9847 12361
rect 10873 12335 10879 12361
rect 10905 12335 10911 12361
rect 11545 12335 11551 12361
rect 11577 12335 11583 12361
rect 12441 12335 12447 12361
rect 12473 12335 12479 12361
rect 13337 12335 13343 12361
rect 13369 12335 13375 12361
rect 14401 12335 14407 12361
rect 14433 12335 14439 12361
rect 14737 12335 14743 12361
rect 14769 12335 14775 12361
rect 15297 12335 15303 12361
rect 15329 12335 15335 12361
rect 15409 12335 15415 12361
rect 15441 12335 15447 12361
rect 16809 12335 16815 12361
rect 16841 12335 16847 12361
rect 17985 12335 17991 12361
rect 18017 12335 18023 12361
rect 18545 12335 18551 12361
rect 18577 12335 18583 12361
rect 19441 12335 19447 12361
rect 19473 12335 19479 12361
rect 20897 12335 20903 12361
rect 20929 12335 20935 12361
rect 21793 12335 21799 12361
rect 21825 12335 21831 12361
rect 22521 12335 22527 12361
rect 22553 12335 22559 12361
rect 23417 12335 23423 12361
rect 23449 12335 23455 12361
rect 24761 12335 24767 12361
rect 24793 12335 24799 12361
rect 25937 12335 25943 12361
rect 25969 12335 25975 12361
rect 26497 12335 26503 12361
rect 26529 12335 26535 12361
rect 27393 12335 27399 12361
rect 27425 12335 27431 12361
rect 29689 12335 29695 12361
rect 29721 12335 29727 12361
rect 29913 12335 29919 12361
rect 29945 12335 29951 12361
rect 30361 12335 30367 12361
rect 30393 12335 30399 12361
rect 30697 12335 30703 12361
rect 30729 12335 30735 12361
rect 31593 12335 31599 12361
rect 31625 12335 31631 12361
rect 672 12165 39312 12182
rect 672 12139 2074 12165
rect 2100 12139 2136 12165
rect 2162 12139 2198 12165
rect 2224 12139 2260 12165
rect 2286 12139 2322 12165
rect 2348 12139 2384 12165
rect 2410 12139 2446 12165
rect 2472 12139 2508 12165
rect 2534 12139 7074 12165
rect 7100 12139 7136 12165
rect 7162 12139 7198 12165
rect 7224 12139 7260 12165
rect 7286 12139 7322 12165
rect 7348 12139 7384 12165
rect 7410 12139 7446 12165
rect 7472 12139 7508 12165
rect 7534 12139 12074 12165
rect 12100 12139 12136 12165
rect 12162 12139 12198 12165
rect 12224 12139 12260 12165
rect 12286 12139 12322 12165
rect 12348 12139 12384 12165
rect 12410 12139 12446 12165
rect 12472 12139 12508 12165
rect 12534 12139 17074 12165
rect 17100 12139 17136 12165
rect 17162 12139 17198 12165
rect 17224 12139 17260 12165
rect 17286 12139 17322 12165
rect 17348 12139 17384 12165
rect 17410 12139 17446 12165
rect 17472 12139 17508 12165
rect 17534 12139 22074 12165
rect 22100 12139 22136 12165
rect 22162 12139 22198 12165
rect 22224 12139 22260 12165
rect 22286 12139 22322 12165
rect 22348 12139 22384 12165
rect 22410 12139 22446 12165
rect 22472 12139 22508 12165
rect 22534 12139 27074 12165
rect 27100 12139 27136 12165
rect 27162 12139 27198 12165
rect 27224 12139 27260 12165
rect 27286 12139 27322 12165
rect 27348 12139 27384 12165
rect 27410 12139 27446 12165
rect 27472 12139 27508 12165
rect 27534 12139 32074 12165
rect 32100 12139 32136 12165
rect 32162 12139 32198 12165
rect 32224 12139 32260 12165
rect 32286 12139 32322 12165
rect 32348 12139 32384 12165
rect 32410 12139 32446 12165
rect 32472 12139 32508 12165
rect 32534 12139 37074 12165
rect 37100 12139 37136 12165
rect 37162 12139 37198 12165
rect 37224 12139 37260 12165
rect 37286 12139 37322 12165
rect 37348 12139 37384 12165
rect 37410 12139 37446 12165
rect 37472 12139 37508 12165
rect 37534 12139 39312 12165
rect 672 12122 39312 12139
rect 1801 11943 1807 11969
rect 1833 11943 1839 11969
rect 1913 11943 1919 11969
rect 1945 11943 1951 11969
rect 2193 11943 2199 11969
rect 2225 11943 2231 11969
rect 4097 11943 4103 11969
rect 4129 11943 4135 11969
rect 4321 11943 4327 11969
rect 4353 11943 4359 11969
rect 4489 11943 4495 11969
rect 4521 11943 4527 11969
rect 5273 11943 5279 11969
rect 5305 11943 5311 11969
rect 6393 11943 6399 11969
rect 6425 11943 6431 11969
rect 7793 11943 7799 11969
rect 7825 11943 7831 11969
rect 8353 11943 8359 11969
rect 8385 11943 8391 11969
rect 8465 11943 8471 11969
rect 8497 11943 8503 11969
rect 9249 11943 9255 11969
rect 9281 11943 9287 11969
rect 10425 11943 10431 11969
rect 10457 11943 10463 11969
rect 11993 11943 11999 11969
rect 12025 11943 12031 11969
rect 12945 11943 12951 11969
rect 12977 11943 12983 11969
rect 13337 11943 13343 11969
rect 13369 11943 13375 11969
rect 14401 11943 14407 11969
rect 14433 11943 14439 11969
rect 14793 11943 14799 11969
rect 14825 11943 14831 11969
rect 15857 11943 15863 11969
rect 15889 11943 15895 11969
rect 16529 11943 16535 11969
rect 16561 11943 16567 11969
rect 17425 11943 17431 11969
rect 17457 11943 17463 11969
rect 19049 11943 19055 11969
rect 19081 11943 19087 11969
rect 19945 11943 19951 11969
rect 19977 11943 19983 11969
rect 20505 11943 20511 11969
rect 20537 11943 20543 11969
rect 21401 11943 21407 11969
rect 21433 11943 21439 11969
rect 23025 11943 23031 11969
rect 23057 11943 23063 11969
rect 23305 11943 23311 11969
rect 23337 11943 23343 11969
rect 23417 11943 23423 11969
rect 23449 11943 23455 11969
rect 24481 11943 24487 11969
rect 24513 11943 24519 11969
rect 25153 11943 25159 11969
rect 25185 11943 25191 11969
rect 26721 11943 26727 11969
rect 26753 11943 26759 11969
rect 27673 11943 27679 11969
rect 27705 11943 27711 11969
rect 28233 11943 28239 11969
rect 28265 11943 28271 11969
rect 29353 11943 29359 11969
rect 29385 11943 29391 11969
rect 30697 11943 30703 11969
rect 30729 11943 30735 11969
rect 31593 11943 31599 11969
rect 31625 11943 31631 11969
rect 32433 11943 32439 11969
rect 32465 11943 32471 11969
rect 32825 11943 32831 11969
rect 32857 11943 32863 11969
rect 6393 11887 6399 11913
rect 6425 11887 6431 11913
rect 10425 11887 10431 11913
rect 10457 11887 10463 11913
rect 12945 11887 12951 11913
rect 12977 11887 12983 11913
rect 14401 11887 14407 11913
rect 14433 11887 14439 11913
rect 15857 11887 15863 11913
rect 15889 11887 15895 11913
rect 17425 11887 17431 11913
rect 17457 11887 17463 11913
rect 19945 11887 19951 11913
rect 19977 11887 19983 11913
rect 21401 11887 21407 11913
rect 21433 11887 21439 11913
rect 25153 11887 25159 11913
rect 25185 11887 25191 11913
rect 27673 11887 27679 11913
rect 27705 11887 27711 11913
rect 29353 11887 29359 11913
rect 29385 11887 29391 11913
rect 31649 11887 31655 11913
rect 31681 11887 31687 11913
rect 33105 11887 33111 11913
rect 33137 11887 33143 11913
rect 672 11773 39312 11790
rect 672 11747 4574 11773
rect 4600 11747 4636 11773
rect 4662 11747 4698 11773
rect 4724 11747 4760 11773
rect 4786 11747 4822 11773
rect 4848 11747 4884 11773
rect 4910 11747 4946 11773
rect 4972 11747 5008 11773
rect 5034 11747 9574 11773
rect 9600 11747 9636 11773
rect 9662 11747 9698 11773
rect 9724 11747 9760 11773
rect 9786 11747 9822 11773
rect 9848 11747 9884 11773
rect 9910 11747 9946 11773
rect 9972 11747 10008 11773
rect 10034 11747 14574 11773
rect 14600 11747 14636 11773
rect 14662 11747 14698 11773
rect 14724 11747 14760 11773
rect 14786 11747 14822 11773
rect 14848 11747 14884 11773
rect 14910 11747 14946 11773
rect 14972 11747 15008 11773
rect 15034 11747 19574 11773
rect 19600 11747 19636 11773
rect 19662 11747 19698 11773
rect 19724 11747 19760 11773
rect 19786 11747 19822 11773
rect 19848 11747 19884 11773
rect 19910 11747 19946 11773
rect 19972 11747 20008 11773
rect 20034 11747 24574 11773
rect 24600 11747 24636 11773
rect 24662 11747 24698 11773
rect 24724 11747 24760 11773
rect 24786 11747 24822 11773
rect 24848 11747 24884 11773
rect 24910 11747 24946 11773
rect 24972 11747 25008 11773
rect 25034 11747 29574 11773
rect 29600 11747 29636 11773
rect 29662 11747 29698 11773
rect 29724 11747 29760 11773
rect 29786 11747 29822 11773
rect 29848 11747 29884 11773
rect 29910 11747 29946 11773
rect 29972 11747 30008 11773
rect 30034 11747 34574 11773
rect 34600 11747 34636 11773
rect 34662 11747 34698 11773
rect 34724 11747 34760 11773
rect 34786 11747 34822 11773
rect 34848 11747 34884 11773
rect 34910 11747 34946 11773
rect 34972 11747 35008 11773
rect 35034 11747 39312 11773
rect 672 11730 39312 11747
rect 1857 11607 1863 11633
rect 1889 11607 1895 11633
rect 4433 11607 4439 11633
rect 4465 11607 4471 11633
rect 7009 11607 7015 11633
rect 7041 11607 7047 11633
rect 8353 11607 8359 11633
rect 8385 11607 8391 11633
rect 10761 11607 10767 11633
rect 10793 11607 10799 11633
rect 12441 11607 12447 11633
rect 12473 11607 12479 11633
rect 14457 11607 14463 11633
rect 14489 11607 14495 11633
rect 15857 11607 15863 11633
rect 15889 11607 15895 11633
rect 17985 11607 17991 11633
rect 18017 11607 18023 11633
rect 23305 11607 23311 11633
rect 23337 11607 23343 11633
rect 28345 11607 28351 11633
rect 28377 11607 28383 11633
rect 31481 11607 31487 11633
rect 31513 11607 31519 11633
rect 1857 11551 1863 11577
rect 1889 11551 1895 11577
rect 3033 11551 3039 11577
rect 3065 11551 3071 11577
rect 3593 11551 3599 11577
rect 3625 11551 3631 11577
rect 4433 11551 4439 11577
rect 4465 11551 4471 11577
rect 5833 11551 5839 11577
rect 5865 11551 5871 11577
rect 7009 11551 7015 11577
rect 7041 11551 7047 11577
rect 7569 11551 7575 11577
rect 7601 11551 7607 11577
rect 8353 11551 8359 11577
rect 8385 11551 8391 11577
rect 10033 11551 10039 11577
rect 10065 11551 10071 11577
rect 10761 11551 10767 11577
rect 10793 11551 10799 11577
rect 11545 11551 11551 11577
rect 11577 11551 11583 11577
rect 12441 11551 12447 11577
rect 12473 11551 12479 11577
rect 13449 11551 13455 11577
rect 13481 11551 13487 11577
rect 14457 11551 14463 11577
rect 14489 11551 14495 11577
rect 15073 11551 15079 11577
rect 15105 11551 15111 11577
rect 15857 11551 15863 11577
rect 15889 11551 15895 11577
rect 16809 11551 16815 11577
rect 16841 11551 16847 11577
rect 17985 11551 17991 11577
rect 18017 11551 18023 11577
rect 18545 11551 18551 11577
rect 18577 11551 18583 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 18937 11551 18943 11577
rect 18969 11551 18975 11577
rect 20785 11551 20791 11577
rect 20817 11551 20823 11577
rect 21345 11551 21351 11577
rect 21377 11551 21383 11577
rect 21457 11551 21463 11577
rect 21489 11551 21495 11577
rect 22521 11551 22527 11577
rect 22553 11551 22559 11577
rect 23305 11551 23311 11577
rect 23337 11551 23343 11577
rect 24761 11551 24767 11577
rect 24793 11551 24799 11577
rect 25209 11551 25215 11577
rect 25241 11551 25247 11577
rect 25433 11551 25439 11577
rect 25465 11551 25471 11577
rect 27449 11551 27455 11577
rect 27481 11551 27487 11577
rect 28345 11551 28351 11577
rect 28377 11551 28383 11577
rect 28849 11551 28855 11577
rect 28881 11551 28887 11577
rect 29409 11551 29415 11577
rect 29441 11551 29447 11577
rect 29521 11551 29527 11577
rect 29553 11551 29559 11577
rect 30585 11551 30591 11577
rect 30617 11551 30623 11577
rect 31481 11551 31487 11577
rect 31513 11551 31519 11577
rect 32769 11551 32775 11577
rect 32801 11551 32807 11577
rect 33161 11551 33167 11577
rect 33193 11551 33199 11577
rect 33609 11551 33615 11577
rect 33641 11551 33647 11577
rect 672 11381 39312 11398
rect 672 11355 2074 11381
rect 2100 11355 2136 11381
rect 2162 11355 2198 11381
rect 2224 11355 2260 11381
rect 2286 11355 2322 11381
rect 2348 11355 2384 11381
rect 2410 11355 2446 11381
rect 2472 11355 2508 11381
rect 2534 11355 7074 11381
rect 7100 11355 7136 11381
rect 7162 11355 7198 11381
rect 7224 11355 7260 11381
rect 7286 11355 7322 11381
rect 7348 11355 7384 11381
rect 7410 11355 7446 11381
rect 7472 11355 7508 11381
rect 7534 11355 12074 11381
rect 12100 11355 12136 11381
rect 12162 11355 12198 11381
rect 12224 11355 12260 11381
rect 12286 11355 12322 11381
rect 12348 11355 12384 11381
rect 12410 11355 12446 11381
rect 12472 11355 12508 11381
rect 12534 11355 17074 11381
rect 17100 11355 17136 11381
rect 17162 11355 17198 11381
rect 17224 11355 17260 11381
rect 17286 11355 17322 11381
rect 17348 11355 17384 11381
rect 17410 11355 17446 11381
rect 17472 11355 17508 11381
rect 17534 11355 22074 11381
rect 22100 11355 22136 11381
rect 22162 11355 22198 11381
rect 22224 11355 22260 11381
rect 22286 11355 22322 11381
rect 22348 11355 22384 11381
rect 22410 11355 22446 11381
rect 22472 11355 22508 11381
rect 22534 11355 27074 11381
rect 27100 11355 27136 11381
rect 27162 11355 27198 11381
rect 27224 11355 27260 11381
rect 27286 11355 27322 11381
rect 27348 11355 27384 11381
rect 27410 11355 27446 11381
rect 27472 11355 27508 11381
rect 27534 11355 32074 11381
rect 32100 11355 32136 11381
rect 32162 11355 32198 11381
rect 32224 11355 32260 11381
rect 32286 11355 32322 11381
rect 32348 11355 32384 11381
rect 32410 11355 32446 11381
rect 32472 11355 32508 11381
rect 32534 11355 37074 11381
rect 37100 11355 37136 11381
rect 37162 11355 37198 11381
rect 37224 11355 37260 11381
rect 37286 11355 37322 11381
rect 37348 11355 37384 11381
rect 37410 11355 37446 11381
rect 37472 11355 37508 11381
rect 37534 11355 39312 11381
rect 672 11338 39312 11355
rect 1801 11159 1807 11185
rect 1833 11159 1839 11185
rect 1913 11159 1919 11185
rect 1945 11159 1951 11185
rect 2473 11159 2479 11185
rect 2505 11159 2511 11185
rect 3817 11159 3823 11185
rect 3849 11159 3855 11185
rect 4377 11159 4383 11185
rect 4409 11159 4415 11185
rect 4489 11159 4495 11185
rect 4521 11159 4527 11185
rect 5273 11159 5279 11185
rect 5305 11159 5311 11185
rect 6449 11159 6455 11185
rect 6481 11159 6487 11185
rect 7793 11159 7799 11185
rect 7825 11159 7831 11185
rect 8353 11159 8359 11185
rect 8385 11159 8391 11185
rect 8465 11159 8471 11185
rect 8497 11159 8503 11185
rect 9249 11159 9255 11185
rect 9281 11159 9287 11185
rect 10425 11159 10431 11185
rect 10457 11159 10463 11185
rect 11993 11159 11999 11185
rect 12025 11159 12031 11185
rect 12945 11159 12951 11185
rect 12977 11159 12983 11185
rect 13337 11159 13343 11185
rect 13369 11159 13375 11185
rect 14401 11159 14407 11185
rect 14433 11159 14439 11185
rect 15073 11159 15079 11185
rect 15105 11159 15111 11185
rect 15297 11159 15303 11185
rect 15329 11159 15335 11185
rect 15465 11159 15471 11185
rect 15497 11159 15503 11185
rect 16529 11159 16535 11185
rect 16561 11159 16567 11185
rect 17257 11159 17263 11185
rect 17289 11159 17295 11185
rect 18769 11159 18775 11185
rect 18801 11159 18807 11185
rect 19217 11159 19223 11185
rect 19249 11159 19255 11185
rect 19945 11159 19951 11185
rect 19977 11159 19983 11185
rect 20225 11159 20231 11185
rect 20257 11159 20263 11185
rect 21345 11159 21351 11185
rect 21377 11159 21383 11185
rect 23025 11159 23031 11185
rect 23057 11159 23063 11185
rect 23305 11159 23311 11185
rect 23337 11159 23343 11185
rect 23417 11159 23423 11185
rect 23449 11159 23455 11185
rect 24369 11159 24375 11185
rect 24401 11159 24407 11185
rect 25153 11159 25159 11185
rect 25185 11159 25191 11185
rect 27561 11159 27567 11185
rect 27593 11159 27599 11185
rect 28513 11159 28519 11185
rect 28545 11159 28551 11185
rect 28793 11159 28799 11185
rect 28825 11159 28831 11185
rect 29969 11159 29975 11185
rect 30001 11159 30007 11185
rect 30753 11159 30759 11185
rect 30785 11159 30791 11185
rect 31481 11159 31487 11185
rect 31513 11159 31519 11185
rect 32433 11159 32439 11185
rect 32465 11159 32471 11185
rect 33105 11159 33111 11185
rect 33137 11159 33143 11185
rect 34953 11159 34959 11185
rect 34985 11159 34991 11185
rect 35121 11159 35127 11185
rect 35153 11159 35159 11185
rect 35345 11159 35351 11185
rect 35377 11159 35383 11185
rect 36129 11159 36135 11185
rect 36161 11159 36167 11185
rect 37305 11159 37311 11185
rect 37337 11159 37343 11185
rect 6449 11103 6455 11129
rect 6481 11103 6487 11129
rect 10425 11103 10431 11129
rect 10457 11103 10463 11129
rect 12945 11103 12951 11129
rect 12977 11103 12983 11129
rect 14401 11103 14407 11129
rect 14433 11103 14439 11129
rect 17257 11103 17263 11129
rect 17289 11103 17295 11129
rect 21345 11103 21351 11129
rect 21377 11103 21383 11129
rect 25153 11103 25159 11129
rect 25185 11103 25191 11129
rect 28513 11103 28519 11129
rect 28545 11103 28551 11129
rect 29969 11103 29975 11129
rect 30001 11103 30007 11129
rect 31649 11103 31655 11129
rect 31681 11103 31687 11129
rect 33105 11103 33111 11129
rect 33137 11103 33143 11129
rect 37305 11103 37311 11129
rect 37337 11103 37343 11129
rect 672 10989 39312 11006
rect 672 10963 4574 10989
rect 4600 10963 4636 10989
rect 4662 10963 4698 10989
rect 4724 10963 4760 10989
rect 4786 10963 4822 10989
rect 4848 10963 4884 10989
rect 4910 10963 4946 10989
rect 4972 10963 5008 10989
rect 5034 10963 9574 10989
rect 9600 10963 9636 10989
rect 9662 10963 9698 10989
rect 9724 10963 9760 10989
rect 9786 10963 9822 10989
rect 9848 10963 9884 10989
rect 9910 10963 9946 10989
rect 9972 10963 10008 10989
rect 10034 10963 14574 10989
rect 14600 10963 14636 10989
rect 14662 10963 14698 10989
rect 14724 10963 14760 10989
rect 14786 10963 14822 10989
rect 14848 10963 14884 10989
rect 14910 10963 14946 10989
rect 14972 10963 15008 10989
rect 15034 10963 19574 10989
rect 19600 10963 19636 10989
rect 19662 10963 19698 10989
rect 19724 10963 19760 10989
rect 19786 10963 19822 10989
rect 19848 10963 19884 10989
rect 19910 10963 19946 10989
rect 19972 10963 20008 10989
rect 20034 10963 24574 10989
rect 24600 10963 24636 10989
rect 24662 10963 24698 10989
rect 24724 10963 24760 10989
rect 24786 10963 24822 10989
rect 24848 10963 24884 10989
rect 24910 10963 24946 10989
rect 24972 10963 25008 10989
rect 25034 10963 29574 10989
rect 29600 10963 29636 10989
rect 29662 10963 29698 10989
rect 29724 10963 29760 10989
rect 29786 10963 29822 10989
rect 29848 10963 29884 10989
rect 29910 10963 29946 10989
rect 29972 10963 30008 10989
rect 30034 10963 34574 10989
rect 34600 10963 34636 10989
rect 34662 10963 34698 10989
rect 34724 10963 34760 10989
rect 34786 10963 34822 10989
rect 34848 10963 34884 10989
rect 34910 10963 34946 10989
rect 34972 10963 35008 10989
rect 35034 10963 39312 10989
rect 672 10946 39312 10963
rect 2081 10823 2087 10849
rect 2113 10823 2119 10849
rect 4433 10823 4439 10849
rect 4465 10823 4471 10849
rect 7009 10823 7015 10849
rect 7041 10823 7047 10849
rect 8465 10823 8471 10849
rect 8497 10823 8503 10849
rect 10761 10823 10767 10849
rect 10793 10823 10799 10849
rect 12217 10823 12223 10849
rect 12249 10823 12255 10849
rect 14457 10823 14463 10849
rect 14489 10823 14495 10849
rect 19273 10823 19279 10849
rect 19305 10823 19311 10849
rect 23417 10823 23423 10849
rect 23449 10823 23455 10849
rect 28289 10823 28295 10849
rect 28321 10823 28327 10849
rect 29969 10823 29975 10849
rect 30001 10823 30007 10849
rect 31425 10823 31431 10849
rect 31457 10823 31463 10849
rect 37641 10823 37647 10849
rect 37673 10823 37679 10849
rect 2081 10767 2087 10793
rect 2113 10767 2119 10793
rect 3033 10767 3039 10793
rect 3065 10767 3071 10793
rect 3593 10767 3599 10793
rect 3625 10767 3631 10793
rect 4433 10767 4439 10793
rect 4465 10767 4471 10793
rect 5833 10767 5839 10793
rect 5865 10767 5871 10793
rect 7009 10767 7015 10793
rect 7041 10767 7047 10793
rect 7289 10767 7295 10793
rect 7321 10767 7327 10793
rect 8465 10767 8471 10793
rect 8497 10767 8503 10793
rect 10033 10767 10039 10793
rect 10065 10767 10071 10793
rect 10761 10767 10767 10793
rect 10793 10767 10799 10793
rect 11545 10767 11551 10793
rect 11577 10767 11583 10793
rect 12217 10767 12223 10793
rect 12249 10767 12255 10793
rect 13449 10767 13455 10793
rect 13481 10767 13487 10793
rect 14457 10767 14463 10793
rect 14489 10767 14495 10793
rect 15073 10767 15079 10793
rect 15105 10767 15111 10793
rect 15353 10767 15359 10793
rect 15385 10767 15391 10793
rect 15577 10767 15583 10793
rect 15609 10767 15615 10793
rect 16809 10767 16815 10793
rect 16841 10767 16847 10793
rect 17257 10767 17263 10793
rect 17289 10767 17295 10793
rect 17481 10767 17487 10793
rect 17513 10767 17519 10793
rect 18545 10767 18551 10793
rect 18577 10767 18583 10793
rect 19273 10767 19279 10793
rect 19305 10767 19311 10793
rect 20785 10767 20791 10793
rect 20817 10767 20823 10793
rect 21345 10767 21351 10793
rect 21377 10767 21383 10793
rect 21457 10767 21463 10793
rect 21489 10767 21495 10793
rect 22521 10767 22527 10793
rect 22553 10767 22559 10793
rect 23417 10767 23423 10793
rect 23449 10767 23455 10793
rect 25041 10767 25047 10793
rect 25073 10767 25079 10793
rect 25321 10767 25327 10793
rect 25353 10767 25359 10793
rect 25433 10767 25439 10793
rect 25465 10767 25471 10793
rect 27449 10767 27455 10793
rect 27481 10767 27487 10793
rect 28289 10767 28295 10793
rect 28321 10767 28327 10793
rect 28793 10767 28799 10793
rect 28825 10767 28831 10793
rect 29969 10767 29975 10793
rect 30001 10767 30007 10793
rect 30305 10767 30311 10793
rect 30337 10767 30343 10793
rect 31425 10767 31431 10793
rect 31457 10767 31463 10793
rect 32769 10767 32775 10793
rect 32801 10767 32807 10793
rect 33161 10767 33167 10793
rect 33193 10767 33199 10793
rect 33385 10767 33391 10793
rect 33417 10767 33423 10793
rect 34449 10767 34455 10793
rect 34481 10767 34487 10793
rect 34617 10767 34623 10793
rect 34649 10767 34655 10793
rect 34841 10767 34847 10793
rect 34873 10767 34879 10793
rect 36689 10767 36695 10793
rect 36721 10767 36727 10793
rect 37641 10767 37647 10793
rect 37673 10767 37679 10793
rect 672 10597 39312 10614
rect 672 10571 2074 10597
rect 2100 10571 2136 10597
rect 2162 10571 2198 10597
rect 2224 10571 2260 10597
rect 2286 10571 2322 10597
rect 2348 10571 2384 10597
rect 2410 10571 2446 10597
rect 2472 10571 2508 10597
rect 2534 10571 7074 10597
rect 7100 10571 7136 10597
rect 7162 10571 7198 10597
rect 7224 10571 7260 10597
rect 7286 10571 7322 10597
rect 7348 10571 7384 10597
rect 7410 10571 7446 10597
rect 7472 10571 7508 10597
rect 7534 10571 12074 10597
rect 12100 10571 12136 10597
rect 12162 10571 12198 10597
rect 12224 10571 12260 10597
rect 12286 10571 12322 10597
rect 12348 10571 12384 10597
rect 12410 10571 12446 10597
rect 12472 10571 12508 10597
rect 12534 10571 17074 10597
rect 17100 10571 17136 10597
rect 17162 10571 17198 10597
rect 17224 10571 17260 10597
rect 17286 10571 17322 10597
rect 17348 10571 17384 10597
rect 17410 10571 17446 10597
rect 17472 10571 17508 10597
rect 17534 10571 22074 10597
rect 22100 10571 22136 10597
rect 22162 10571 22198 10597
rect 22224 10571 22260 10597
rect 22286 10571 22322 10597
rect 22348 10571 22384 10597
rect 22410 10571 22446 10597
rect 22472 10571 22508 10597
rect 22534 10571 27074 10597
rect 27100 10571 27136 10597
rect 27162 10571 27198 10597
rect 27224 10571 27260 10597
rect 27286 10571 27322 10597
rect 27348 10571 27384 10597
rect 27410 10571 27446 10597
rect 27472 10571 27508 10597
rect 27534 10571 32074 10597
rect 32100 10571 32136 10597
rect 32162 10571 32198 10597
rect 32224 10571 32260 10597
rect 32286 10571 32322 10597
rect 32348 10571 32384 10597
rect 32410 10571 32446 10597
rect 32472 10571 32508 10597
rect 32534 10571 37074 10597
rect 37100 10571 37136 10597
rect 37162 10571 37198 10597
rect 37224 10571 37260 10597
rect 37286 10571 37322 10597
rect 37348 10571 37384 10597
rect 37410 10571 37446 10597
rect 37472 10571 37508 10597
rect 37534 10571 39312 10597
rect 672 10554 39312 10571
rect 1633 10375 1639 10401
rect 1665 10375 1671 10401
rect 2473 10375 2479 10401
rect 2505 10375 2511 10401
rect 3817 10375 3823 10401
rect 3849 10375 3855 10401
rect 4377 10375 4383 10401
rect 4409 10375 4415 10401
rect 4489 10375 4495 10401
rect 4521 10375 4527 10401
rect 5273 10375 5279 10401
rect 5305 10375 5311 10401
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 7793 10375 7799 10401
rect 7825 10375 7831 10401
rect 8745 10375 8751 10401
rect 8777 10375 8783 10401
rect 9249 10375 9255 10401
rect 9281 10375 9287 10401
rect 10425 10375 10431 10401
rect 10457 10375 10463 10401
rect 11937 10375 11943 10401
rect 11969 10375 11975 10401
rect 12665 10375 12671 10401
rect 12697 10375 12703 10401
rect 13337 10375 13343 10401
rect 13369 10375 13375 10401
rect 14289 10375 14295 10401
rect 14321 10375 14327 10401
rect 15073 10375 15079 10401
rect 15105 10375 15111 10401
rect 15353 10375 15359 10401
rect 15385 10375 15391 10401
rect 15465 10375 15471 10401
rect 15497 10375 15503 10401
rect 16529 10375 16535 10401
rect 16561 10375 16567 10401
rect 16809 10375 16815 10401
rect 16841 10375 16847 10401
rect 16921 10375 16927 10401
rect 16953 10375 16959 10401
rect 18769 10375 18775 10401
rect 18801 10375 18807 10401
rect 19273 10375 19279 10401
rect 19305 10375 19311 10401
rect 19497 10375 19503 10401
rect 19529 10375 19535 10401
rect 20225 10375 20231 10401
rect 20257 10375 20263 10401
rect 21345 10375 21351 10401
rect 21377 10375 21383 10401
rect 23025 10375 23031 10401
rect 23057 10375 23063 10401
rect 23865 10375 23871 10401
rect 23897 10375 23903 10401
rect 24369 10375 24375 10401
rect 24401 10375 24407 10401
rect 24649 10375 24655 10401
rect 24681 10375 24687 10401
rect 24873 10375 24879 10401
rect 24905 10375 24911 10401
rect 27673 10375 27679 10401
rect 27705 10375 27711 10401
rect 28065 10375 28071 10401
rect 28097 10375 28103 10401
rect 28513 10375 28519 10401
rect 28545 10375 28551 10401
rect 28793 10375 28799 10401
rect 28825 10375 28831 10401
rect 29969 10375 29975 10401
rect 30001 10375 30007 10401
rect 30697 10375 30703 10401
rect 30729 10375 30735 10401
rect 31257 10375 31263 10401
rect 31289 10375 31295 10401
rect 31425 10375 31431 10401
rect 31457 10375 31463 10401
rect 32153 10375 32159 10401
rect 32185 10375 32191 10401
rect 33105 10375 33111 10401
rect 33137 10375 33143 10401
rect 34953 10375 34959 10401
rect 34985 10375 34991 10401
rect 35233 10375 35239 10401
rect 35265 10375 35271 10401
rect 35345 10375 35351 10401
rect 35377 10375 35383 10401
rect 36129 10375 36135 10401
rect 36161 10375 36167 10401
rect 37305 10375 37311 10401
rect 37337 10375 37343 10401
rect 1521 10319 1527 10345
rect 1553 10319 1559 10345
rect 6449 10319 6455 10345
rect 6481 10319 6487 10345
rect 8745 10319 8751 10345
rect 8777 10319 8783 10345
rect 10425 10319 10431 10345
rect 10457 10319 10463 10345
rect 12665 10319 12671 10345
rect 12697 10319 12703 10345
rect 14289 10319 14295 10345
rect 14321 10319 14327 10345
rect 21345 10319 21351 10345
rect 21377 10319 21383 10345
rect 23865 10319 23871 10345
rect 23897 10319 23903 10345
rect 29969 10319 29975 10345
rect 30001 10319 30007 10345
rect 33105 10319 33111 10345
rect 33137 10319 33143 10345
rect 37305 10319 37311 10345
rect 37337 10319 37343 10345
rect 672 10205 39312 10222
rect 672 10179 4574 10205
rect 4600 10179 4636 10205
rect 4662 10179 4698 10205
rect 4724 10179 4760 10205
rect 4786 10179 4822 10205
rect 4848 10179 4884 10205
rect 4910 10179 4946 10205
rect 4972 10179 5008 10205
rect 5034 10179 9574 10205
rect 9600 10179 9636 10205
rect 9662 10179 9698 10205
rect 9724 10179 9760 10205
rect 9786 10179 9822 10205
rect 9848 10179 9884 10205
rect 9910 10179 9946 10205
rect 9972 10179 10008 10205
rect 10034 10179 14574 10205
rect 14600 10179 14636 10205
rect 14662 10179 14698 10205
rect 14724 10179 14760 10205
rect 14786 10179 14822 10205
rect 14848 10179 14884 10205
rect 14910 10179 14946 10205
rect 14972 10179 15008 10205
rect 15034 10179 19574 10205
rect 19600 10179 19636 10205
rect 19662 10179 19698 10205
rect 19724 10179 19760 10205
rect 19786 10179 19822 10205
rect 19848 10179 19884 10205
rect 19910 10179 19946 10205
rect 19972 10179 20008 10205
rect 20034 10179 24574 10205
rect 24600 10179 24636 10205
rect 24662 10179 24698 10205
rect 24724 10179 24760 10205
rect 24786 10179 24822 10205
rect 24848 10179 24884 10205
rect 24910 10179 24946 10205
rect 24972 10179 25008 10205
rect 25034 10179 29574 10205
rect 29600 10179 29636 10205
rect 29662 10179 29698 10205
rect 29724 10179 29760 10205
rect 29786 10179 29822 10205
rect 29848 10179 29884 10205
rect 29910 10179 29946 10205
rect 29972 10179 30008 10205
rect 30034 10179 34574 10205
rect 34600 10179 34636 10205
rect 34662 10179 34698 10205
rect 34724 10179 34760 10205
rect 34786 10179 34822 10205
rect 34848 10179 34884 10205
rect 34910 10179 34946 10205
rect 34972 10179 35008 10205
rect 35034 10179 39312 10205
rect 672 10162 39312 10179
rect 1857 10039 1863 10065
rect 1889 10039 1895 10065
rect 7009 10039 7015 10065
rect 7041 10039 7047 10065
rect 8465 10039 8471 10065
rect 8497 10039 8503 10065
rect 17985 10039 17991 10065
rect 18017 10039 18023 10065
rect 19441 10039 19447 10065
rect 19473 10039 19479 10065
rect 23417 10039 23423 10065
rect 23449 10039 23455 10065
rect 25937 10039 25943 10065
rect 25969 10039 25975 10065
rect 37641 10039 37647 10065
rect 37673 10039 37679 10065
rect 1857 9983 1863 10009
rect 1889 9983 1895 10009
rect 2753 9983 2759 10009
rect 2785 9983 2791 10009
rect 3593 9983 3599 10009
rect 3625 9983 3631 10009
rect 3817 9983 3823 10009
rect 3849 9983 3855 10009
rect 3985 9983 3991 10009
rect 4017 9983 4023 10009
rect 5889 9983 5895 10009
rect 5921 9983 5927 10009
rect 7009 9983 7015 10009
rect 7041 9983 7047 10009
rect 7569 9983 7575 10009
rect 7601 9983 7607 10009
rect 8465 9983 8471 10009
rect 8497 9983 8503 10009
rect 10033 9983 10039 10009
rect 10065 9983 10071 10009
rect 10369 9983 10375 10009
rect 10401 9983 10407 10009
rect 10537 9983 10543 10009
rect 10569 9983 10575 10009
rect 11545 9983 11551 10009
rect 11577 9983 11583 10009
rect 11769 9983 11775 10009
rect 11801 9983 11807 10009
rect 11937 9983 11943 10009
rect 11969 9983 11975 10009
rect 13617 9983 13623 10009
rect 13649 9983 13655 10009
rect 14065 9983 14071 10009
rect 14097 9983 14103 10009
rect 14289 9983 14295 10009
rect 14321 9983 14327 10009
rect 15073 9983 15079 10009
rect 15105 9983 15111 10009
rect 15521 9983 15527 10009
rect 15553 9983 15559 10009
rect 15745 9983 15751 10009
rect 15777 9983 15783 10009
rect 16809 9983 16815 10009
rect 16841 9983 16847 10009
rect 17985 9983 17991 10009
rect 18017 9983 18023 10009
rect 18265 9983 18271 10009
rect 18297 9983 18303 10009
rect 19441 9983 19447 10009
rect 19473 9983 19479 10009
rect 20785 9983 20791 10009
rect 20817 9983 20823 10009
rect 21345 9983 21351 10009
rect 21377 9983 21383 10009
rect 21457 9983 21463 10009
rect 21489 9983 21495 10009
rect 22241 9983 22247 10009
rect 22273 9983 22279 10009
rect 23417 9983 23423 10009
rect 23449 9983 23455 10009
rect 25937 9983 25943 10009
rect 25969 9983 25975 10009
rect 26833 9983 26839 10009
rect 26865 9983 26871 10009
rect 27673 9983 27679 10009
rect 27705 9983 27711 10009
rect 27897 9983 27903 10009
rect 27929 9983 27935 10009
rect 28345 9983 28351 10009
rect 28377 9983 28383 10009
rect 29409 9983 29415 10009
rect 29441 9983 29447 10009
rect 29801 9983 29807 10009
rect 29833 9983 29839 10009
rect 30025 9983 30031 10009
rect 30057 9983 30063 10009
rect 30809 9983 30815 10009
rect 30841 9983 30847 10009
rect 31369 9983 31375 10009
rect 31401 9983 31407 10009
rect 31481 9983 31487 10009
rect 31513 9983 31519 10009
rect 32825 9983 32831 10009
rect 32857 9983 32863 10009
rect 33161 9983 33167 10009
rect 33193 9983 33199 10009
rect 33609 9983 33615 10009
rect 33641 9983 33647 10009
rect 34449 9983 34455 10009
rect 34481 9983 34487 10009
rect 34617 9983 34623 10009
rect 34649 9983 34655 10009
rect 34841 9983 34847 10009
rect 34873 9983 34879 10009
rect 36689 9983 36695 10009
rect 36721 9983 36727 10009
rect 37641 9983 37647 10009
rect 37673 9983 37679 10009
rect 672 9813 39312 9830
rect 672 9787 2074 9813
rect 2100 9787 2136 9813
rect 2162 9787 2198 9813
rect 2224 9787 2260 9813
rect 2286 9787 2322 9813
rect 2348 9787 2384 9813
rect 2410 9787 2446 9813
rect 2472 9787 2508 9813
rect 2534 9787 7074 9813
rect 7100 9787 7136 9813
rect 7162 9787 7198 9813
rect 7224 9787 7260 9813
rect 7286 9787 7322 9813
rect 7348 9787 7384 9813
rect 7410 9787 7446 9813
rect 7472 9787 7508 9813
rect 7534 9787 12074 9813
rect 12100 9787 12136 9813
rect 12162 9787 12198 9813
rect 12224 9787 12260 9813
rect 12286 9787 12322 9813
rect 12348 9787 12384 9813
rect 12410 9787 12446 9813
rect 12472 9787 12508 9813
rect 12534 9787 17074 9813
rect 17100 9787 17136 9813
rect 17162 9787 17198 9813
rect 17224 9787 17260 9813
rect 17286 9787 17322 9813
rect 17348 9787 17384 9813
rect 17410 9787 17446 9813
rect 17472 9787 17508 9813
rect 17534 9787 22074 9813
rect 22100 9787 22136 9813
rect 22162 9787 22198 9813
rect 22224 9787 22260 9813
rect 22286 9787 22322 9813
rect 22348 9787 22384 9813
rect 22410 9787 22446 9813
rect 22472 9787 22508 9813
rect 22534 9787 27074 9813
rect 27100 9787 27136 9813
rect 27162 9787 27198 9813
rect 27224 9787 27260 9813
rect 27286 9787 27322 9813
rect 27348 9787 27384 9813
rect 27410 9787 27446 9813
rect 27472 9787 27508 9813
rect 27534 9787 32074 9813
rect 32100 9787 32136 9813
rect 32162 9787 32198 9813
rect 32224 9787 32260 9813
rect 32286 9787 32322 9813
rect 32348 9787 32384 9813
rect 32410 9787 32446 9813
rect 32472 9787 32508 9813
rect 32534 9787 37074 9813
rect 37100 9787 37136 9813
rect 37162 9787 37198 9813
rect 37224 9787 37260 9813
rect 37286 9787 37322 9813
rect 37348 9787 37384 9813
rect 37410 9787 37446 9813
rect 37472 9787 37508 9813
rect 37534 9787 39312 9813
rect 672 9770 39312 9787
rect 1801 9591 1807 9617
rect 1833 9591 1839 9617
rect 2025 9591 2031 9617
rect 2057 9591 2063 9617
rect 2473 9591 2479 9617
rect 2505 9591 2511 9617
rect 3817 9591 3823 9617
rect 3849 9591 3855 9617
rect 4993 9591 4999 9617
rect 5025 9591 5031 9617
rect 5273 9591 5279 9617
rect 5305 9591 5311 9617
rect 5945 9591 5951 9617
rect 5977 9591 5983 9617
rect 7793 9591 7799 9617
rect 7825 9591 7831 9617
rect 8745 9591 8751 9617
rect 8777 9591 8783 9617
rect 9249 9591 9255 9617
rect 9281 9591 9287 9617
rect 10425 9591 10431 9617
rect 10457 9591 10463 9617
rect 11601 9591 11607 9617
rect 11633 9591 11639 9617
rect 12049 9591 12055 9617
rect 12081 9591 12087 9617
rect 12273 9591 12279 9617
rect 12305 9591 12311 9617
rect 13337 9591 13343 9617
rect 13369 9591 13375 9617
rect 14009 9591 14015 9617
rect 14041 9591 14047 9617
rect 14793 9591 14799 9617
rect 14825 9591 14831 9617
rect 15241 9591 15247 9617
rect 15273 9591 15279 9617
rect 15465 9591 15471 9617
rect 15497 9591 15503 9617
rect 16249 9591 16255 9617
rect 16281 9591 16287 9617
rect 16809 9591 16815 9617
rect 16841 9591 16847 9617
rect 16921 9591 16927 9617
rect 16953 9591 16959 9617
rect 18769 9591 18775 9617
rect 18801 9591 18807 9617
rect 19329 9591 19335 9617
rect 19361 9591 19367 9617
rect 19441 9591 19447 9617
rect 19473 9591 19479 9617
rect 20225 9591 20231 9617
rect 20257 9591 20263 9617
rect 21345 9591 21351 9617
rect 21377 9591 21383 9617
rect 22745 9591 22751 9617
rect 22777 9591 22783 9617
rect 23865 9591 23871 9617
rect 23897 9591 23903 9617
rect 24425 9591 24431 9617
rect 24457 9591 24463 9617
rect 25377 9591 25383 9617
rect 25409 9591 25415 9617
rect 28177 9591 28183 9617
rect 28209 9591 28215 9617
rect 28401 9591 28407 9617
rect 28433 9591 28439 9617
rect 28793 9591 28799 9617
rect 28825 9591 28831 9617
rect 29409 9591 29415 9617
rect 29441 9591 29447 9617
rect 29689 9591 29695 9617
rect 29721 9591 29727 9617
rect 29801 9591 29807 9617
rect 29833 9591 29839 9617
rect 30977 9591 30983 9617
rect 31009 9591 31015 9617
rect 31145 9591 31151 9617
rect 31177 9591 31183 9617
rect 31369 9591 31375 9617
rect 31401 9591 31407 9617
rect 32153 9591 32159 9617
rect 32185 9591 32191 9617
rect 32825 9591 32831 9617
rect 32857 9591 32863 9617
rect 34953 9591 34959 9617
rect 34985 9591 34991 9617
rect 35121 9591 35127 9617
rect 35153 9591 35159 9617
rect 35345 9591 35351 9617
rect 35377 9591 35383 9617
rect 36409 9591 36415 9617
rect 36441 9591 36447 9617
rect 37305 9591 37311 9617
rect 37337 9591 37343 9617
rect 3817 9535 3823 9561
rect 3849 9535 3855 9561
rect 6225 9535 6231 9561
rect 6257 9535 6263 9561
rect 8745 9535 8751 9561
rect 8777 9535 8783 9561
rect 10425 9535 10431 9561
rect 10457 9535 10463 9561
rect 14009 9535 14015 9561
rect 14041 9535 14047 9561
rect 21345 9535 21351 9561
rect 21377 9535 21383 9561
rect 23865 9535 23871 9561
rect 23897 9535 23903 9561
rect 25377 9535 25383 9561
rect 25409 9535 25415 9561
rect 33105 9535 33111 9561
rect 33137 9535 33143 9561
rect 37305 9535 37311 9561
rect 37337 9535 37343 9561
rect 672 9421 39312 9438
rect 672 9395 4574 9421
rect 4600 9395 4636 9421
rect 4662 9395 4698 9421
rect 4724 9395 4760 9421
rect 4786 9395 4822 9421
rect 4848 9395 4884 9421
rect 4910 9395 4946 9421
rect 4972 9395 5008 9421
rect 5034 9395 9574 9421
rect 9600 9395 9636 9421
rect 9662 9395 9698 9421
rect 9724 9395 9760 9421
rect 9786 9395 9822 9421
rect 9848 9395 9884 9421
rect 9910 9395 9946 9421
rect 9972 9395 10008 9421
rect 10034 9395 14574 9421
rect 14600 9395 14636 9421
rect 14662 9395 14698 9421
rect 14724 9395 14760 9421
rect 14786 9395 14822 9421
rect 14848 9395 14884 9421
rect 14910 9395 14946 9421
rect 14972 9395 15008 9421
rect 15034 9395 19574 9421
rect 19600 9395 19636 9421
rect 19662 9395 19698 9421
rect 19724 9395 19760 9421
rect 19786 9395 19822 9421
rect 19848 9395 19884 9421
rect 19910 9395 19946 9421
rect 19972 9395 20008 9421
rect 20034 9395 24574 9421
rect 24600 9395 24636 9421
rect 24662 9395 24698 9421
rect 24724 9395 24760 9421
rect 24786 9395 24822 9421
rect 24848 9395 24884 9421
rect 24910 9395 24946 9421
rect 24972 9395 25008 9421
rect 25034 9395 29574 9421
rect 29600 9395 29636 9421
rect 29662 9395 29698 9421
rect 29724 9395 29760 9421
rect 29786 9395 29822 9421
rect 29848 9395 29884 9421
rect 29910 9395 29946 9421
rect 29972 9395 30008 9421
rect 30034 9395 34574 9421
rect 34600 9395 34636 9421
rect 34662 9395 34698 9421
rect 34724 9395 34760 9421
rect 34786 9395 34822 9421
rect 34848 9395 34884 9421
rect 34910 9395 34946 9421
rect 34972 9395 35008 9421
rect 35034 9395 39312 9421
rect 672 9378 39312 9395
rect 1857 9255 1863 9281
rect 1889 9255 1895 9281
rect 3369 9255 3375 9281
rect 3401 9255 3407 9281
rect 8409 9255 8415 9281
rect 8441 9255 8447 9281
rect 15745 9255 15751 9281
rect 15777 9255 15783 9281
rect 17985 9255 17991 9281
rect 18017 9255 18023 9281
rect 19329 9255 19335 9281
rect 19361 9255 19367 9281
rect 23417 9255 23423 9281
rect 23449 9255 23455 9281
rect 25937 9255 25943 9281
rect 25969 9255 25975 9281
rect 27729 9255 27735 9281
rect 27761 9255 27767 9281
rect 30193 9255 30199 9281
rect 30225 9255 30231 9281
rect 35233 9255 35239 9281
rect 35265 9255 35271 9281
rect 37641 9255 37647 9281
rect 37673 9255 37679 9281
rect 1857 9199 1863 9225
rect 1889 9199 1895 9225
rect 3033 9199 3039 9225
rect 3065 9199 3071 9225
rect 3369 9199 3375 9225
rect 3401 9199 3407 9225
rect 4489 9199 4495 9225
rect 4521 9199 4527 9225
rect 6113 9199 6119 9225
rect 6145 9199 6151 9225
rect 6281 9199 6287 9225
rect 6313 9199 6319 9225
rect 6505 9199 6511 9225
rect 6537 9199 6543 9225
rect 7569 9199 7575 9225
rect 7601 9199 7607 9225
rect 8409 9199 8415 9225
rect 8441 9199 8447 9225
rect 10033 9199 10039 9225
rect 10065 9199 10071 9225
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 10481 9199 10487 9225
rect 10513 9199 10519 9225
rect 11433 9199 11439 9225
rect 11465 9199 11471 9225
rect 11769 9199 11775 9225
rect 11801 9199 11807 9225
rect 11937 9199 11943 9225
rect 11969 9199 11975 9225
rect 13337 9199 13343 9225
rect 13369 9199 13375 9225
rect 13785 9199 13791 9225
rect 13817 9199 13823 9225
rect 14009 9199 14015 9225
rect 14041 9199 14047 9225
rect 14793 9199 14799 9225
rect 14825 9199 14831 9225
rect 15745 9199 15751 9225
rect 15777 9199 15783 9225
rect 16809 9199 16815 9225
rect 16841 9199 16847 9225
rect 17985 9199 17991 9225
rect 18017 9199 18023 9225
rect 18265 9199 18271 9225
rect 18297 9199 18303 9225
rect 19273 9199 19279 9225
rect 19305 9199 19311 9225
rect 20785 9199 20791 9225
rect 20817 9199 20823 9225
rect 21345 9199 21351 9225
rect 21377 9199 21383 9225
rect 21457 9199 21463 9225
rect 21489 9199 21495 9225
rect 22521 9199 22527 9225
rect 22553 9199 22559 9225
rect 23417 9199 23423 9225
rect 23449 9199 23455 9225
rect 25041 9199 25047 9225
rect 25073 9199 25079 9225
rect 25937 9199 25943 9225
rect 25969 9199 25975 9225
rect 26945 9199 26951 9225
rect 26977 9199 26983 9225
rect 27617 9199 27623 9225
rect 27649 9199 27655 9225
rect 29521 9199 29527 9225
rect 29553 9199 29559 9225
rect 30193 9199 30199 9225
rect 30225 9199 30231 9225
rect 30977 9199 30983 9225
rect 31009 9199 31015 9225
rect 31145 9199 31151 9225
rect 31177 9199 31183 9225
rect 31369 9199 31375 9225
rect 31401 9199 31407 9225
rect 32825 9199 32831 9225
rect 32857 9199 32863 9225
rect 33161 9199 33167 9225
rect 33193 9199 33199 9225
rect 33609 9199 33615 9225
rect 33641 9199 33647 9225
rect 34169 9199 34175 9225
rect 34201 9199 34207 9225
rect 35233 9199 35239 9225
rect 35265 9199 35271 9225
rect 36689 9199 36695 9225
rect 36721 9199 36727 9225
rect 37641 9199 37647 9225
rect 37673 9199 37679 9225
rect 672 9029 39312 9046
rect 672 9003 2074 9029
rect 2100 9003 2136 9029
rect 2162 9003 2198 9029
rect 2224 9003 2260 9029
rect 2286 9003 2322 9029
rect 2348 9003 2384 9029
rect 2410 9003 2446 9029
rect 2472 9003 2508 9029
rect 2534 9003 7074 9029
rect 7100 9003 7136 9029
rect 7162 9003 7198 9029
rect 7224 9003 7260 9029
rect 7286 9003 7322 9029
rect 7348 9003 7384 9029
rect 7410 9003 7446 9029
rect 7472 9003 7508 9029
rect 7534 9003 12074 9029
rect 12100 9003 12136 9029
rect 12162 9003 12198 9029
rect 12224 9003 12260 9029
rect 12286 9003 12322 9029
rect 12348 9003 12384 9029
rect 12410 9003 12446 9029
rect 12472 9003 12508 9029
rect 12534 9003 17074 9029
rect 17100 9003 17136 9029
rect 17162 9003 17198 9029
rect 17224 9003 17260 9029
rect 17286 9003 17322 9029
rect 17348 9003 17384 9029
rect 17410 9003 17446 9029
rect 17472 9003 17508 9029
rect 17534 9003 22074 9029
rect 22100 9003 22136 9029
rect 22162 9003 22198 9029
rect 22224 9003 22260 9029
rect 22286 9003 22322 9029
rect 22348 9003 22384 9029
rect 22410 9003 22446 9029
rect 22472 9003 22508 9029
rect 22534 9003 27074 9029
rect 27100 9003 27136 9029
rect 27162 9003 27198 9029
rect 27224 9003 27260 9029
rect 27286 9003 27322 9029
rect 27348 9003 27384 9029
rect 27410 9003 27446 9029
rect 27472 9003 27508 9029
rect 27534 9003 32074 9029
rect 32100 9003 32136 9029
rect 32162 9003 32198 9029
rect 32224 9003 32260 9029
rect 32286 9003 32322 9029
rect 32348 9003 32384 9029
rect 32410 9003 32446 9029
rect 32472 9003 32508 9029
rect 32534 9003 37074 9029
rect 37100 9003 37136 9029
rect 37162 9003 37198 9029
rect 37224 9003 37260 9029
rect 37286 9003 37322 9029
rect 37348 9003 37384 9029
rect 37410 9003 37446 9029
rect 37472 9003 37508 9029
rect 37534 9003 39312 9029
rect 672 8986 39312 9003
rect 1409 8807 1415 8833
rect 1441 8807 1447 8833
rect 2473 8807 2479 8833
rect 2505 8807 2511 8833
rect 3817 8807 3823 8833
rect 3849 8807 3855 8833
rect 4993 8807 4999 8833
rect 5025 8807 5031 8833
rect 5553 8807 5559 8833
rect 5585 8807 5591 8833
rect 6449 8807 6455 8833
rect 6481 8807 6487 8833
rect 7793 8807 7799 8833
rect 7825 8807 7831 8833
rect 8745 8807 8751 8833
rect 8777 8807 8783 8833
rect 9249 8807 9255 8833
rect 9281 8807 9287 8833
rect 10313 8807 10319 8833
rect 10345 8807 10351 8833
rect 11601 8807 11607 8833
rect 11633 8807 11639 8833
rect 12049 8807 12055 8833
rect 12081 8807 12087 8833
rect 12273 8807 12279 8833
rect 12305 8807 12311 8833
rect 13057 8807 13063 8833
rect 13089 8807 13095 8833
rect 13505 8807 13511 8833
rect 13537 8807 13543 8833
rect 13729 8807 13735 8833
rect 13761 8807 13767 8833
rect 14793 8807 14799 8833
rect 14825 8807 14831 8833
rect 15241 8807 15247 8833
rect 15273 8807 15279 8833
rect 15465 8807 15471 8833
rect 15497 8807 15503 8833
rect 16249 8807 16255 8833
rect 16281 8807 16287 8833
rect 16809 8807 16815 8833
rect 16841 8807 16847 8833
rect 16921 8807 16927 8833
rect 16953 8807 16959 8833
rect 18769 8807 18775 8833
rect 18801 8807 18807 8833
rect 19329 8807 19335 8833
rect 19361 8807 19367 8833
rect 19441 8807 19447 8833
rect 19473 8807 19479 8833
rect 20225 8807 20231 8833
rect 20257 8807 20263 8833
rect 21401 8807 21407 8833
rect 21433 8807 21439 8833
rect 22745 8807 22751 8833
rect 22777 8807 22783 8833
rect 23865 8807 23871 8833
rect 23897 8807 23903 8833
rect 24481 8807 24487 8833
rect 24513 8807 24519 8833
rect 25377 8807 25383 8833
rect 25409 8807 25415 8833
rect 27729 8807 27735 8833
rect 27761 8807 27767 8833
rect 28849 8807 28855 8833
rect 28881 8807 28887 8833
rect 29409 8807 29415 8833
rect 29441 8807 29447 8833
rect 30193 8807 30199 8833
rect 30225 8807 30231 8833
rect 30977 8807 30983 8833
rect 31009 8807 31015 8833
rect 31145 8807 31151 8833
rect 31177 8807 31183 8833
rect 31369 8807 31375 8833
rect 31401 8807 31407 8833
rect 32153 8807 32159 8833
rect 32185 8807 32191 8833
rect 32825 8807 32831 8833
rect 32857 8807 32863 8833
rect 34673 8807 34679 8833
rect 34705 8807 34711 8833
rect 35849 8807 35855 8833
rect 35881 8807 35887 8833
rect 36409 8807 36415 8833
rect 36441 8807 36447 8833
rect 37305 8807 37311 8833
rect 37337 8807 37343 8833
rect 1409 8751 1415 8777
rect 1441 8751 1447 8777
rect 3817 8751 3823 8777
rect 3849 8751 3855 8777
rect 6449 8751 6455 8777
rect 6481 8751 6487 8777
rect 8745 8751 8751 8777
rect 8777 8751 8783 8777
rect 10313 8751 10319 8777
rect 10345 8751 10351 8777
rect 21401 8751 21407 8777
rect 21433 8751 21439 8777
rect 23865 8751 23871 8777
rect 23897 8751 23903 8777
rect 25377 8751 25383 8777
rect 25409 8751 25415 8777
rect 27729 8751 27735 8777
rect 27761 8751 27767 8777
rect 30193 8751 30199 8777
rect 30225 8751 30231 8777
rect 33105 8751 33111 8777
rect 33137 8751 33143 8777
rect 35849 8751 35855 8777
rect 35881 8751 35887 8777
rect 37305 8751 37311 8777
rect 37337 8751 37343 8777
rect 672 8637 39312 8654
rect 672 8611 4574 8637
rect 4600 8611 4636 8637
rect 4662 8611 4698 8637
rect 4724 8611 4760 8637
rect 4786 8611 4822 8637
rect 4848 8611 4884 8637
rect 4910 8611 4946 8637
rect 4972 8611 5008 8637
rect 5034 8611 9574 8637
rect 9600 8611 9636 8637
rect 9662 8611 9698 8637
rect 9724 8611 9760 8637
rect 9786 8611 9822 8637
rect 9848 8611 9884 8637
rect 9910 8611 9946 8637
rect 9972 8611 10008 8637
rect 10034 8611 14574 8637
rect 14600 8611 14636 8637
rect 14662 8611 14698 8637
rect 14724 8611 14760 8637
rect 14786 8611 14822 8637
rect 14848 8611 14884 8637
rect 14910 8611 14946 8637
rect 14972 8611 15008 8637
rect 15034 8611 19574 8637
rect 19600 8611 19636 8637
rect 19662 8611 19698 8637
rect 19724 8611 19760 8637
rect 19786 8611 19822 8637
rect 19848 8611 19884 8637
rect 19910 8611 19946 8637
rect 19972 8611 20008 8637
rect 20034 8611 24574 8637
rect 24600 8611 24636 8637
rect 24662 8611 24698 8637
rect 24724 8611 24760 8637
rect 24786 8611 24822 8637
rect 24848 8611 24884 8637
rect 24910 8611 24946 8637
rect 24972 8611 25008 8637
rect 25034 8611 29574 8637
rect 29600 8611 29636 8637
rect 29662 8611 29698 8637
rect 29724 8611 29760 8637
rect 29786 8611 29822 8637
rect 29848 8611 29884 8637
rect 29910 8611 29946 8637
rect 29972 8611 30008 8637
rect 30034 8611 34574 8637
rect 34600 8611 34636 8637
rect 34662 8611 34698 8637
rect 34724 8611 34760 8637
rect 34786 8611 34822 8637
rect 34848 8611 34884 8637
rect 34910 8611 34946 8637
rect 34972 8611 35008 8637
rect 35034 8611 39312 8637
rect 672 8594 39312 8611
rect 1857 8471 1863 8497
rect 1889 8471 1895 8497
rect 4489 8471 4495 8497
rect 4521 8471 4527 8497
rect 8409 8471 8415 8497
rect 8441 8471 8447 8497
rect 17985 8471 17991 8497
rect 18017 8471 18023 8497
rect 19441 8471 19447 8497
rect 19473 8471 19479 8497
rect 21793 8471 21799 8497
rect 21825 8471 21831 8497
rect 23417 8471 23423 8497
rect 23449 8471 23455 8497
rect 25937 8471 25943 8497
rect 25969 8471 25975 8497
rect 27393 8471 27399 8497
rect 27425 8471 27431 8497
rect 35345 8471 35351 8497
rect 35377 8471 35383 8497
rect 37641 8471 37647 8497
rect 37673 8471 37679 8497
rect 1857 8415 1863 8441
rect 1889 8415 1895 8441
rect 3033 8415 3039 8441
rect 3065 8415 3071 8441
rect 3593 8415 3599 8441
rect 3625 8415 3631 8441
rect 4489 8415 4495 8441
rect 4521 8415 4527 8441
rect 6113 8415 6119 8441
rect 6145 8415 6151 8441
rect 6393 8415 6399 8441
rect 6425 8415 6431 8441
rect 6505 8415 6511 8441
rect 6537 8415 6543 8441
rect 7569 8415 7575 8441
rect 7601 8415 7607 8441
rect 8409 8415 8415 8441
rect 8441 8415 8447 8441
rect 9809 8415 9815 8441
rect 9841 8415 9847 8441
rect 10313 8415 10319 8441
rect 10345 8415 10351 8441
rect 10481 8415 10487 8441
rect 10513 8415 10519 8441
rect 11433 8415 11439 8441
rect 11465 8415 11471 8441
rect 11769 8415 11775 8441
rect 11801 8415 11807 8441
rect 11937 8415 11943 8441
rect 11969 8415 11975 8441
rect 13001 8415 13007 8441
rect 13033 8415 13039 8441
rect 13449 8415 13455 8441
rect 13481 8415 13487 8441
rect 13673 8415 13679 8441
rect 13705 8415 13711 8441
rect 14457 8415 14463 8441
rect 14489 8415 14495 8441
rect 15017 8415 15023 8441
rect 15049 8415 15055 8441
rect 15129 8415 15135 8441
rect 15161 8415 15167 8441
rect 16809 8415 16815 8441
rect 16841 8415 16847 8441
rect 17985 8415 17991 8441
rect 18017 8415 18023 8441
rect 18265 8415 18271 8441
rect 18297 8415 18303 8441
rect 19441 8415 19447 8441
rect 19473 8415 19479 8441
rect 20785 8415 20791 8441
rect 20817 8415 20823 8441
rect 21793 8415 21799 8441
rect 21825 8415 21831 8441
rect 22521 8415 22527 8441
rect 22553 8415 22559 8441
rect 23417 8415 23423 8441
rect 23449 8415 23455 8441
rect 24761 8415 24767 8441
rect 24793 8415 24799 8441
rect 25937 8415 25943 8441
rect 25969 8415 25975 8441
rect 26217 8415 26223 8441
rect 26249 8415 26255 8441
rect 27393 8415 27399 8441
rect 27425 8415 27431 8441
rect 29409 8415 29415 8441
rect 29441 8415 29447 8441
rect 29857 8415 29863 8441
rect 29889 8415 29895 8441
rect 30081 8415 30087 8441
rect 30113 8415 30119 8441
rect 31033 8415 31039 8441
rect 31065 8415 31071 8441
rect 31313 8415 31319 8441
rect 31345 8415 31351 8441
rect 31425 8415 31431 8441
rect 31457 8415 31463 8441
rect 32713 8415 32719 8441
rect 32745 8415 32751 8441
rect 33161 8415 33167 8441
rect 33193 8415 33199 8441
rect 33609 8415 33615 8441
rect 33641 8415 33647 8441
rect 34169 8415 34175 8441
rect 34201 8415 34207 8441
rect 35345 8415 35351 8441
rect 35377 8415 35383 8441
rect 36689 8415 36695 8441
rect 36721 8415 36727 8441
rect 37641 8415 37647 8441
rect 37673 8415 37679 8441
rect 672 8245 39312 8262
rect 672 8219 2074 8245
rect 2100 8219 2136 8245
rect 2162 8219 2198 8245
rect 2224 8219 2260 8245
rect 2286 8219 2322 8245
rect 2348 8219 2384 8245
rect 2410 8219 2446 8245
rect 2472 8219 2508 8245
rect 2534 8219 7074 8245
rect 7100 8219 7136 8245
rect 7162 8219 7198 8245
rect 7224 8219 7260 8245
rect 7286 8219 7322 8245
rect 7348 8219 7384 8245
rect 7410 8219 7446 8245
rect 7472 8219 7508 8245
rect 7534 8219 12074 8245
rect 12100 8219 12136 8245
rect 12162 8219 12198 8245
rect 12224 8219 12260 8245
rect 12286 8219 12322 8245
rect 12348 8219 12384 8245
rect 12410 8219 12446 8245
rect 12472 8219 12508 8245
rect 12534 8219 17074 8245
rect 17100 8219 17136 8245
rect 17162 8219 17198 8245
rect 17224 8219 17260 8245
rect 17286 8219 17322 8245
rect 17348 8219 17384 8245
rect 17410 8219 17446 8245
rect 17472 8219 17508 8245
rect 17534 8219 22074 8245
rect 22100 8219 22136 8245
rect 22162 8219 22198 8245
rect 22224 8219 22260 8245
rect 22286 8219 22322 8245
rect 22348 8219 22384 8245
rect 22410 8219 22446 8245
rect 22472 8219 22508 8245
rect 22534 8219 27074 8245
rect 27100 8219 27136 8245
rect 27162 8219 27198 8245
rect 27224 8219 27260 8245
rect 27286 8219 27322 8245
rect 27348 8219 27384 8245
rect 27410 8219 27446 8245
rect 27472 8219 27508 8245
rect 27534 8219 32074 8245
rect 32100 8219 32136 8245
rect 32162 8219 32198 8245
rect 32224 8219 32260 8245
rect 32286 8219 32322 8245
rect 32348 8219 32384 8245
rect 32410 8219 32446 8245
rect 32472 8219 32508 8245
rect 32534 8219 37074 8245
rect 37100 8219 37136 8245
rect 37162 8219 37198 8245
rect 37224 8219 37260 8245
rect 37286 8219 37322 8245
rect 37348 8219 37384 8245
rect 37410 8219 37446 8245
rect 37472 8219 37508 8245
rect 37534 8219 39312 8245
rect 672 8202 39312 8219
rect 33615 8049 33641 8055
rect 1801 8023 1807 8049
rect 1833 8023 1839 8049
rect 2473 8023 2479 8049
rect 2505 8023 2511 8049
rect 4097 8023 4103 8049
rect 4129 8023 4135 8049
rect 4377 8023 4383 8049
rect 4409 8023 4415 8049
rect 4489 8023 4495 8049
rect 4521 8023 4527 8049
rect 5553 8023 5559 8049
rect 5585 8023 5591 8049
rect 6449 8023 6455 8049
rect 6481 8023 6487 8049
rect 7793 8023 7799 8049
rect 7825 8023 7831 8049
rect 8745 8023 8751 8049
rect 8777 8023 8783 8049
rect 9249 8023 9255 8049
rect 9281 8023 9287 8049
rect 10425 8023 10431 8049
rect 10457 8023 10463 8049
rect 11433 8023 11439 8049
rect 11465 8023 11471 8049
rect 11769 8023 11775 8049
rect 11801 8023 11807 8049
rect 11881 8023 11887 8049
rect 11913 8023 11919 8049
rect 12889 8023 12895 8049
rect 12921 8023 12927 8049
rect 13449 8023 13455 8049
rect 13481 8023 13487 8049
rect 13561 8023 13567 8049
rect 13593 8023 13599 8049
rect 14961 8023 14967 8049
rect 14993 8023 14999 8049
rect 15745 8023 15751 8049
rect 15777 8023 15783 8049
rect 16249 8023 16255 8049
rect 16281 8023 16287 8049
rect 16809 8023 16815 8049
rect 16841 8023 16847 8049
rect 16921 8023 16927 8049
rect 16953 8023 16959 8049
rect 18769 8023 18775 8049
rect 18801 8023 18807 8049
rect 19945 8023 19951 8049
rect 19977 8023 19983 8049
rect 20225 8023 20231 8049
rect 20257 8023 20263 8049
rect 21401 8023 21407 8049
rect 21433 8023 21439 8049
rect 22745 8023 22751 8049
rect 22777 8023 22783 8049
rect 23865 8023 23871 8049
rect 23897 8023 23903 8049
rect 24481 8023 24487 8049
rect 24513 8023 24519 8049
rect 25153 8023 25159 8049
rect 25185 8023 25191 8049
rect 26721 8023 26727 8049
rect 26753 8023 26759 8049
rect 27673 8023 27679 8049
rect 27705 8023 27711 8049
rect 29353 8023 29359 8049
rect 29385 8023 29391 8049
rect 29857 8023 29863 8049
rect 29889 8023 29895 8049
rect 30753 8023 30759 8049
rect 30785 8023 30791 8049
rect 31145 8023 31151 8049
rect 31177 8023 31183 8049
rect 31369 8023 31375 8049
rect 31401 8023 31407 8049
rect 32433 8023 32439 8049
rect 32465 8023 32471 8049
rect 33161 8023 33167 8049
rect 33193 8023 33199 8049
rect 33615 8017 33641 8023
rect 33727 8049 33753 8055
rect 34673 8023 34679 8049
rect 34705 8023 34711 8049
rect 35849 8023 35855 8049
rect 35881 8023 35887 8049
rect 36129 8023 36135 8049
rect 36161 8023 36167 8049
rect 36969 8023 36975 8049
rect 37001 8023 37007 8049
rect 33727 8017 33753 8023
rect 33895 7993 33921 7999
rect 1521 7967 1527 7993
rect 1553 7967 1559 7993
rect 6449 7967 6455 7993
rect 6481 7967 6487 7993
rect 8745 7967 8751 7993
rect 8777 7967 8783 7993
rect 10425 7967 10431 7993
rect 10457 7967 10463 7993
rect 15745 7967 15751 7993
rect 15777 7967 15783 7993
rect 19945 7967 19951 7993
rect 19977 7967 19983 7993
rect 21401 7967 21407 7993
rect 21433 7967 21439 7993
rect 23865 7967 23871 7993
rect 23897 7967 23903 7993
rect 25153 7967 25159 7993
rect 25185 7967 25191 7993
rect 27673 7967 27679 7993
rect 27705 7967 27711 7993
rect 30081 7967 30087 7993
rect 30113 7967 30119 7993
rect 33161 7967 33167 7993
rect 33193 7967 33199 7993
rect 35849 7967 35855 7993
rect 35881 7967 35887 7993
rect 37081 7967 37087 7993
rect 37113 7967 37119 7993
rect 33895 7961 33921 7967
rect 672 7853 39312 7870
rect 672 7827 4574 7853
rect 4600 7827 4636 7853
rect 4662 7827 4698 7853
rect 4724 7827 4760 7853
rect 4786 7827 4822 7853
rect 4848 7827 4884 7853
rect 4910 7827 4946 7853
rect 4972 7827 5008 7853
rect 5034 7827 9574 7853
rect 9600 7827 9636 7853
rect 9662 7827 9698 7853
rect 9724 7827 9760 7853
rect 9786 7827 9822 7853
rect 9848 7827 9884 7853
rect 9910 7827 9946 7853
rect 9972 7827 10008 7853
rect 10034 7827 14574 7853
rect 14600 7827 14636 7853
rect 14662 7827 14698 7853
rect 14724 7827 14760 7853
rect 14786 7827 14822 7853
rect 14848 7827 14884 7853
rect 14910 7827 14946 7853
rect 14972 7827 15008 7853
rect 15034 7827 19574 7853
rect 19600 7827 19636 7853
rect 19662 7827 19698 7853
rect 19724 7827 19760 7853
rect 19786 7827 19822 7853
rect 19848 7827 19884 7853
rect 19910 7827 19946 7853
rect 19972 7827 20008 7853
rect 20034 7827 24574 7853
rect 24600 7827 24636 7853
rect 24662 7827 24698 7853
rect 24724 7827 24760 7853
rect 24786 7827 24822 7853
rect 24848 7827 24884 7853
rect 24910 7827 24946 7853
rect 24972 7827 25008 7853
rect 25034 7827 29574 7853
rect 29600 7827 29636 7853
rect 29662 7827 29698 7853
rect 29724 7827 29760 7853
rect 29786 7827 29822 7853
rect 29848 7827 29884 7853
rect 29910 7827 29946 7853
rect 29972 7827 30008 7853
rect 30034 7827 34574 7853
rect 34600 7827 34636 7853
rect 34662 7827 34698 7853
rect 34724 7827 34760 7853
rect 34786 7827 34822 7853
rect 34848 7827 34884 7853
rect 34910 7827 34946 7853
rect 34972 7827 35008 7853
rect 35034 7827 39312 7853
rect 672 7810 39312 7827
rect 1857 7687 1863 7713
rect 1889 7687 1895 7713
rect 4489 7687 4495 7713
rect 4521 7687 4527 7713
rect 15241 7687 15247 7713
rect 15273 7687 15279 7713
rect 18377 7687 18383 7713
rect 18409 7687 18415 7713
rect 20001 7687 20007 7713
rect 20033 7687 20039 7713
rect 21793 7687 21799 7713
rect 21825 7687 21831 7713
rect 23417 7687 23423 7713
rect 23449 7687 23455 7713
rect 25937 7687 25943 7713
rect 25969 7687 25975 7713
rect 27393 7687 27399 7713
rect 27425 7687 27431 7713
rect 30193 7687 30199 7713
rect 30225 7687 30231 7713
rect 35233 7687 35239 7713
rect 35265 7687 35271 7713
rect 1857 7631 1863 7657
rect 1889 7631 1895 7657
rect 3033 7631 3039 7657
rect 3065 7631 3071 7657
rect 3593 7631 3599 7657
rect 3625 7631 3631 7657
rect 4489 7631 4495 7657
rect 4521 7631 4527 7657
rect 6113 7631 6119 7657
rect 6145 7631 6151 7657
rect 6393 7631 6399 7657
rect 6425 7631 6431 7657
rect 6505 7631 6511 7657
rect 6537 7631 6543 7657
rect 7289 7631 7295 7657
rect 7321 7631 7327 7657
rect 7737 7631 7743 7657
rect 7769 7631 7775 7657
rect 7961 7631 7967 7657
rect 7993 7631 7999 7657
rect 10033 7631 10039 7657
rect 10065 7631 10071 7657
rect 10201 7631 10207 7657
rect 10233 7631 10239 7657
rect 10425 7631 10431 7657
rect 10457 7631 10463 7657
rect 11433 7631 11439 7657
rect 11465 7631 11471 7657
rect 11769 7631 11775 7657
rect 11801 7631 11807 7657
rect 11881 7631 11887 7657
rect 11913 7631 11919 7657
rect 12833 7631 12839 7657
rect 12865 7631 12871 7657
rect 13393 7631 13399 7657
rect 13425 7631 13431 7657
rect 13505 7631 13511 7657
rect 13537 7631 13543 7657
rect 14401 7631 14407 7657
rect 14433 7631 14439 7657
rect 15241 7631 15247 7657
rect 15273 7631 15279 7657
rect 17593 7631 17599 7657
rect 17625 7631 17631 7657
rect 18377 7631 18383 7657
rect 18409 7631 18415 7657
rect 19105 7631 19111 7657
rect 19137 7631 19143 7657
rect 20001 7631 20007 7657
rect 20033 7631 20039 7657
rect 20953 7631 20959 7657
rect 20985 7631 20991 7657
rect 21793 7631 21799 7657
rect 21825 7631 21831 7657
rect 22521 7631 22527 7657
rect 22553 7631 22559 7657
rect 23417 7631 23423 7657
rect 23449 7631 23455 7657
rect 24817 7631 24823 7657
rect 24849 7631 24855 7657
rect 25937 7631 25943 7657
rect 25969 7631 25975 7657
rect 26217 7631 26223 7657
rect 26249 7631 26255 7657
rect 27393 7631 27399 7657
rect 27425 7631 27431 7657
rect 29353 7631 29359 7657
rect 29385 7631 29391 7657
rect 30193 7631 30199 7657
rect 30225 7631 30231 7657
rect 30753 7631 30759 7657
rect 30785 7631 30791 7657
rect 31201 7631 31207 7657
rect 31233 7631 31239 7657
rect 31369 7631 31375 7657
rect 31401 7631 31407 7657
rect 32993 7631 32999 7657
rect 33025 7631 33031 7657
rect 33161 7631 33167 7657
rect 33193 7631 33199 7657
rect 33385 7631 33391 7657
rect 33417 7631 33423 7657
rect 34393 7631 34399 7657
rect 34425 7631 34431 7657
rect 35233 7631 35239 7657
rect 35265 7631 35271 7657
rect 36689 7631 36695 7657
rect 36721 7631 36727 7657
rect 37137 7631 37143 7657
rect 37169 7631 37175 7657
rect 37361 7631 37367 7657
rect 37393 7631 37399 7657
rect 672 7461 39312 7478
rect 672 7435 2074 7461
rect 2100 7435 2136 7461
rect 2162 7435 2198 7461
rect 2224 7435 2260 7461
rect 2286 7435 2322 7461
rect 2348 7435 2384 7461
rect 2410 7435 2446 7461
rect 2472 7435 2508 7461
rect 2534 7435 7074 7461
rect 7100 7435 7136 7461
rect 7162 7435 7198 7461
rect 7224 7435 7260 7461
rect 7286 7435 7322 7461
rect 7348 7435 7384 7461
rect 7410 7435 7446 7461
rect 7472 7435 7508 7461
rect 7534 7435 12074 7461
rect 12100 7435 12136 7461
rect 12162 7435 12198 7461
rect 12224 7435 12260 7461
rect 12286 7435 12322 7461
rect 12348 7435 12384 7461
rect 12410 7435 12446 7461
rect 12472 7435 12508 7461
rect 12534 7435 17074 7461
rect 17100 7435 17136 7461
rect 17162 7435 17198 7461
rect 17224 7435 17260 7461
rect 17286 7435 17322 7461
rect 17348 7435 17384 7461
rect 17410 7435 17446 7461
rect 17472 7435 17508 7461
rect 17534 7435 22074 7461
rect 22100 7435 22136 7461
rect 22162 7435 22198 7461
rect 22224 7435 22260 7461
rect 22286 7435 22322 7461
rect 22348 7435 22384 7461
rect 22410 7435 22446 7461
rect 22472 7435 22508 7461
rect 22534 7435 27074 7461
rect 27100 7435 27136 7461
rect 27162 7435 27198 7461
rect 27224 7435 27260 7461
rect 27286 7435 27322 7461
rect 27348 7435 27384 7461
rect 27410 7435 27446 7461
rect 27472 7435 27508 7461
rect 27534 7435 32074 7461
rect 32100 7435 32136 7461
rect 32162 7435 32198 7461
rect 32224 7435 32260 7461
rect 32286 7435 32322 7461
rect 32348 7435 32384 7461
rect 32410 7435 32446 7461
rect 32472 7435 32508 7461
rect 32534 7435 37074 7461
rect 37100 7435 37136 7461
rect 37162 7435 37198 7461
rect 37224 7435 37260 7461
rect 37286 7435 37322 7461
rect 37348 7435 37384 7461
rect 37410 7435 37446 7461
rect 37472 7435 37508 7461
rect 37534 7435 39312 7461
rect 672 7418 39312 7435
rect 33783 7265 33809 7271
rect 1801 7239 1807 7265
rect 1833 7239 1839 7265
rect 2473 7239 2479 7265
rect 2505 7239 2511 7265
rect 4097 7239 4103 7265
rect 4129 7239 4135 7265
rect 4993 7239 4999 7265
rect 5025 7239 5031 7265
rect 5553 7239 5559 7265
rect 5585 7239 5591 7265
rect 6449 7239 6455 7265
rect 6481 7239 6487 7265
rect 7793 7239 7799 7265
rect 7825 7239 7831 7265
rect 8241 7239 8247 7265
rect 8273 7239 8279 7265
rect 8465 7239 8471 7265
rect 8497 7239 8503 7265
rect 9473 7239 9479 7265
rect 9505 7239 9511 7265
rect 10145 7239 10151 7265
rect 10177 7239 10183 7265
rect 11433 7239 11439 7265
rect 11465 7239 11471 7265
rect 11769 7239 11775 7265
rect 11801 7239 11807 7265
rect 11881 7239 11887 7265
rect 11913 7239 11919 7265
rect 12777 7239 12783 7265
rect 12809 7239 12815 7265
rect 13113 7239 13119 7265
rect 13145 7239 13151 7265
rect 13449 7239 13455 7265
rect 13481 7239 13487 7265
rect 15073 7239 15079 7265
rect 15105 7239 15111 7265
rect 15241 7239 15247 7265
rect 15273 7239 15279 7265
rect 15465 7239 15471 7265
rect 15497 7239 15503 7265
rect 17481 7239 17487 7265
rect 17513 7239 17519 7265
rect 18377 7239 18383 7265
rect 18409 7239 18415 7265
rect 19049 7239 19055 7265
rect 19081 7239 19087 7265
rect 19945 7239 19951 7265
rect 19977 7239 19983 7265
rect 20505 7239 20511 7265
rect 20537 7239 20543 7265
rect 21345 7239 21351 7265
rect 21377 7239 21383 7265
rect 22745 7239 22751 7265
rect 22777 7239 22783 7265
rect 23529 7239 23535 7265
rect 23561 7239 23567 7265
rect 24369 7239 24375 7265
rect 24401 7239 24407 7265
rect 24649 7239 24655 7265
rect 24681 7239 24687 7265
rect 24873 7239 24879 7265
rect 24905 7239 24911 7265
rect 27673 7239 27679 7265
rect 27705 7239 27711 7265
rect 28849 7239 28855 7265
rect 28881 7239 28887 7265
rect 29353 7239 29359 7265
rect 29385 7239 29391 7265
rect 30193 7239 30199 7265
rect 30225 7239 30231 7265
rect 30921 7239 30927 7265
rect 30953 7239 30959 7265
rect 31593 7239 31599 7265
rect 31625 7239 31631 7265
rect 32433 7239 32439 7265
rect 32465 7239 32471 7265
rect 33329 7239 33335 7265
rect 33361 7239 33367 7265
rect 34953 7239 34959 7265
rect 34985 7239 34991 7265
rect 35793 7239 35799 7265
rect 35825 7239 35831 7265
rect 36129 7239 36135 7265
rect 36161 7239 36167 7265
rect 37305 7239 37311 7265
rect 37337 7239 37343 7265
rect 33783 7233 33809 7239
rect 33615 7209 33641 7215
rect 1521 7183 1527 7209
rect 1553 7183 1559 7209
rect 4993 7183 4999 7209
rect 5025 7183 5031 7209
rect 6449 7183 6455 7209
rect 6481 7183 6487 7209
rect 10201 7183 10207 7209
rect 10233 7183 10239 7209
rect 18377 7183 18383 7209
rect 18409 7183 18415 7209
rect 19945 7183 19951 7209
rect 19977 7183 19983 7209
rect 21345 7183 21351 7209
rect 21377 7183 21383 7209
rect 23697 7183 23703 7209
rect 23729 7183 23735 7209
rect 27673 7183 27679 7209
rect 27705 7183 27711 7209
rect 30193 7183 30199 7209
rect 30225 7183 30231 7209
rect 31649 7183 31655 7209
rect 31681 7183 31687 7209
rect 33329 7183 33335 7209
rect 33361 7183 33367 7209
rect 33615 7177 33641 7183
rect 33895 7209 33921 7215
rect 35793 7183 35799 7209
rect 35825 7183 35831 7209
rect 37305 7183 37311 7209
rect 37337 7183 37343 7209
rect 33895 7177 33921 7183
rect 672 7069 39312 7086
rect 672 7043 4574 7069
rect 4600 7043 4636 7069
rect 4662 7043 4698 7069
rect 4724 7043 4760 7069
rect 4786 7043 4822 7069
rect 4848 7043 4884 7069
rect 4910 7043 4946 7069
rect 4972 7043 5008 7069
rect 5034 7043 9574 7069
rect 9600 7043 9636 7069
rect 9662 7043 9698 7069
rect 9724 7043 9760 7069
rect 9786 7043 9822 7069
rect 9848 7043 9884 7069
rect 9910 7043 9946 7069
rect 9972 7043 10008 7069
rect 10034 7043 14574 7069
rect 14600 7043 14636 7069
rect 14662 7043 14698 7069
rect 14724 7043 14760 7069
rect 14786 7043 14822 7069
rect 14848 7043 14884 7069
rect 14910 7043 14946 7069
rect 14972 7043 15008 7069
rect 15034 7043 19574 7069
rect 19600 7043 19636 7069
rect 19662 7043 19698 7069
rect 19724 7043 19760 7069
rect 19786 7043 19822 7069
rect 19848 7043 19884 7069
rect 19910 7043 19946 7069
rect 19972 7043 20008 7069
rect 20034 7043 24574 7069
rect 24600 7043 24636 7069
rect 24662 7043 24698 7069
rect 24724 7043 24760 7069
rect 24786 7043 24822 7069
rect 24848 7043 24884 7069
rect 24910 7043 24946 7069
rect 24972 7043 25008 7069
rect 25034 7043 29574 7069
rect 29600 7043 29636 7069
rect 29662 7043 29698 7069
rect 29724 7043 29760 7069
rect 29786 7043 29822 7069
rect 29848 7043 29884 7069
rect 29910 7043 29946 7069
rect 29972 7043 30008 7069
rect 30034 7043 34574 7069
rect 34600 7043 34636 7069
rect 34662 7043 34698 7069
rect 34724 7043 34760 7069
rect 34786 7043 34822 7069
rect 34848 7043 34884 7069
rect 34910 7043 34946 7069
rect 34972 7043 35008 7069
rect 35034 7043 39312 7069
rect 672 7026 39312 7043
rect 1857 6903 1863 6929
rect 1889 6903 1895 6929
rect 6953 6903 6959 6929
rect 6985 6903 6991 6929
rect 8241 6903 8247 6929
rect 8273 6903 8279 6929
rect 15241 6903 15247 6929
rect 15273 6903 15279 6929
rect 18433 6903 18439 6929
rect 18465 6903 18471 6929
rect 20001 6903 20007 6929
rect 20033 6903 20039 6929
rect 21737 6903 21743 6929
rect 21769 6903 21775 6929
rect 23193 6903 23199 6929
rect 23225 6903 23231 6929
rect 30193 6903 30199 6929
rect 30225 6903 30231 6929
rect 31593 6903 31599 6929
rect 31625 6903 31631 6929
rect 33889 6903 33895 6929
rect 33921 6903 33927 6929
rect 35289 6903 35295 6929
rect 35321 6903 35327 6929
rect 37641 6903 37647 6929
rect 37673 6903 37679 6929
rect 35687 6873 35713 6879
rect 1857 6847 1863 6873
rect 1889 6847 1895 6873
rect 3033 6847 3039 6873
rect 3065 6847 3071 6873
rect 3593 6847 3599 6873
rect 3625 6847 3631 6873
rect 3817 6847 3823 6873
rect 3849 6847 3855 6873
rect 3985 6847 3991 6873
rect 4017 6847 4023 6873
rect 6001 6847 6007 6873
rect 6033 6847 6039 6873
rect 6953 6847 6959 6873
rect 6985 6847 6991 6873
rect 7513 6847 7519 6873
rect 7545 6847 7551 6873
rect 8241 6847 8247 6873
rect 8273 6847 8279 6873
rect 9697 6847 9703 6873
rect 9729 6847 9735 6873
rect 10201 6847 10207 6873
rect 10233 6847 10239 6873
rect 10369 6847 10375 6873
rect 10401 6847 10407 6873
rect 11433 6847 11439 6873
rect 11465 6847 11471 6873
rect 11713 6847 11719 6873
rect 11745 6847 11751 6873
rect 11825 6847 11831 6873
rect 11857 6847 11863 6873
rect 13113 6847 13119 6873
rect 13145 6847 13151 6873
rect 13393 6847 13399 6873
rect 13425 6847 13431 6873
rect 13505 6847 13511 6873
rect 13537 6847 13543 6873
rect 14401 6847 14407 6873
rect 14433 6847 14439 6873
rect 15129 6847 15135 6873
rect 15161 6847 15167 6873
rect 17593 6847 17599 6873
rect 17625 6847 17631 6873
rect 18433 6847 18439 6873
rect 18465 6847 18471 6873
rect 19105 6847 19111 6873
rect 19137 6847 19143 6873
rect 20001 6847 20007 6873
rect 20033 6847 20039 6873
rect 20953 6847 20959 6873
rect 20985 6847 20991 6873
rect 21737 6847 21743 6873
rect 21769 6847 21775 6873
rect 22521 6847 22527 6873
rect 22553 6847 22559 6873
rect 23193 6847 23199 6873
rect 23225 6847 23231 6873
rect 24761 6847 24767 6873
rect 24793 6847 24799 6873
rect 25209 6847 25215 6873
rect 25241 6847 25247 6873
rect 25433 6847 25439 6873
rect 25465 6847 25471 6873
rect 27561 6847 27567 6873
rect 27593 6847 27599 6873
rect 27785 6847 27791 6873
rect 27817 6847 27823 6873
rect 28345 6847 28351 6873
rect 28377 6847 28383 6873
rect 29353 6847 29359 6873
rect 29385 6847 29391 6873
rect 30193 6847 30199 6873
rect 30225 6847 30231 6873
rect 30921 6847 30927 6873
rect 30953 6847 30959 6873
rect 31593 6847 31599 6873
rect 31625 6847 31631 6873
rect 32993 6847 32999 6873
rect 33025 6847 33031 6873
rect 33889 6847 33895 6873
rect 33921 6847 33927 6873
rect 34393 6847 34399 6873
rect 34425 6847 34431 6873
rect 35289 6847 35295 6873
rect 35321 6847 35327 6873
rect 35687 6841 35713 6847
rect 35799 6873 35825 6879
rect 35799 6841 35825 6847
rect 35911 6873 35937 6879
rect 36689 6847 36695 6873
rect 36721 6847 36727 6873
rect 37641 6847 37647 6873
rect 37673 6847 37679 6873
rect 35911 6841 35937 6847
rect 672 6677 39312 6694
rect 672 6651 2074 6677
rect 2100 6651 2136 6677
rect 2162 6651 2198 6677
rect 2224 6651 2260 6677
rect 2286 6651 2322 6677
rect 2348 6651 2384 6677
rect 2410 6651 2446 6677
rect 2472 6651 2508 6677
rect 2534 6651 7074 6677
rect 7100 6651 7136 6677
rect 7162 6651 7198 6677
rect 7224 6651 7260 6677
rect 7286 6651 7322 6677
rect 7348 6651 7384 6677
rect 7410 6651 7446 6677
rect 7472 6651 7508 6677
rect 7534 6651 12074 6677
rect 12100 6651 12136 6677
rect 12162 6651 12198 6677
rect 12224 6651 12260 6677
rect 12286 6651 12322 6677
rect 12348 6651 12384 6677
rect 12410 6651 12446 6677
rect 12472 6651 12508 6677
rect 12534 6651 17074 6677
rect 17100 6651 17136 6677
rect 17162 6651 17198 6677
rect 17224 6651 17260 6677
rect 17286 6651 17322 6677
rect 17348 6651 17384 6677
rect 17410 6651 17446 6677
rect 17472 6651 17508 6677
rect 17534 6651 22074 6677
rect 22100 6651 22136 6677
rect 22162 6651 22198 6677
rect 22224 6651 22260 6677
rect 22286 6651 22322 6677
rect 22348 6651 22384 6677
rect 22410 6651 22446 6677
rect 22472 6651 22508 6677
rect 22534 6651 27074 6677
rect 27100 6651 27136 6677
rect 27162 6651 27198 6677
rect 27224 6651 27260 6677
rect 27286 6651 27322 6677
rect 27348 6651 27384 6677
rect 27410 6651 27446 6677
rect 27472 6651 27508 6677
rect 27534 6651 32074 6677
rect 32100 6651 32136 6677
rect 32162 6651 32198 6677
rect 32224 6651 32260 6677
rect 32286 6651 32322 6677
rect 32348 6651 32384 6677
rect 32410 6651 32446 6677
rect 32472 6651 32508 6677
rect 32534 6651 37074 6677
rect 37100 6651 37136 6677
rect 37162 6651 37198 6677
rect 37224 6651 37260 6677
rect 37286 6651 37322 6677
rect 37348 6651 37384 6677
rect 37410 6651 37446 6677
rect 37472 6651 37508 6677
rect 37534 6651 39312 6677
rect 672 6634 39312 6651
rect 33671 6481 33697 6487
rect 1801 6455 1807 6481
rect 1833 6455 1839 6481
rect 2193 6455 2199 6481
rect 2225 6455 2231 6481
rect 4097 6455 4103 6481
rect 4129 6455 4135 6481
rect 4265 6455 4271 6481
rect 4297 6455 4303 6481
rect 4489 6455 4495 6481
rect 4521 6455 4527 6481
rect 5553 6455 5559 6481
rect 5585 6455 5591 6481
rect 6449 6455 6455 6481
rect 6481 6455 6487 6481
rect 8073 6455 8079 6481
rect 8105 6455 8111 6481
rect 8241 6455 8247 6481
rect 8273 6455 8279 6481
rect 8465 6455 8471 6481
rect 8497 6455 8503 6481
rect 9473 6455 9479 6481
rect 9505 6455 9511 6481
rect 10369 6455 10375 6481
rect 10401 6455 10407 6481
rect 11489 6455 11495 6481
rect 11521 6455 11527 6481
rect 11993 6455 11999 6481
rect 12025 6455 12031 6481
rect 12161 6455 12167 6481
rect 12193 6455 12199 6481
rect 13113 6455 13119 6481
rect 13145 6455 13151 6481
rect 13449 6455 13455 6481
rect 13481 6455 13487 6481
rect 13617 6455 13623 6481
rect 13649 6455 13655 6481
rect 15745 6455 15751 6481
rect 15777 6455 15783 6481
rect 16753 6455 16759 6481
rect 16785 6455 16791 6481
rect 17481 6455 17487 6481
rect 17513 6455 17519 6481
rect 18377 6455 18383 6481
rect 18409 6455 18415 6481
rect 19049 6455 19055 6481
rect 19081 6455 19087 6481
rect 19945 6455 19951 6481
rect 19977 6455 19983 6481
rect 20505 6455 20511 6481
rect 20537 6455 20543 6481
rect 21401 6455 21407 6481
rect 21433 6455 21439 6481
rect 23025 6455 23031 6481
rect 23057 6455 23063 6481
rect 23193 6455 23199 6481
rect 23225 6455 23231 6481
rect 23529 6455 23535 6481
rect 23561 6455 23567 6481
rect 24481 6455 24487 6481
rect 24513 6455 24519 6481
rect 25153 6455 25159 6481
rect 25185 6455 25191 6481
rect 27841 6455 27847 6481
rect 27873 6455 27879 6481
rect 28849 6455 28855 6481
rect 28881 6455 28887 6481
rect 29353 6455 29359 6481
rect 29385 6455 29391 6481
rect 30193 6455 30199 6481
rect 30225 6455 30231 6481
rect 30977 6455 30983 6481
rect 31009 6455 31015 6481
rect 31817 6455 31823 6481
rect 31849 6455 31855 6481
rect 32433 6455 32439 6481
rect 32465 6455 32471 6481
rect 33329 6455 33335 6481
rect 33361 6455 33367 6481
rect 33671 6449 33697 6455
rect 33727 6481 33753 6487
rect 33727 6449 33753 6455
rect 33895 6481 33921 6487
rect 34673 6455 34679 6481
rect 34705 6455 34711 6481
rect 35625 6455 35631 6481
rect 35657 6455 35663 6481
rect 36409 6455 36415 6481
rect 36441 6455 36447 6481
rect 37249 6455 37255 6481
rect 37281 6455 37287 6481
rect 33895 6449 33921 6455
rect 1521 6399 1527 6425
rect 1553 6399 1559 6425
rect 6449 6399 6455 6425
rect 6481 6399 6487 6425
rect 10369 6399 10375 6425
rect 10401 6399 10407 6425
rect 16753 6399 16759 6425
rect 16785 6399 16791 6425
rect 18377 6399 18383 6425
rect 18409 6399 18415 6425
rect 19945 6399 19951 6425
rect 19977 6399 19983 6425
rect 21401 6399 21407 6425
rect 21433 6399 21439 6425
rect 25153 6399 25159 6425
rect 25185 6399 25191 6425
rect 27841 6399 27847 6425
rect 27873 6399 27879 6425
rect 30193 6399 30199 6425
rect 30225 6399 30231 6425
rect 31817 6399 31823 6425
rect 31849 6399 31855 6425
rect 33329 6399 33335 6425
rect 33361 6399 33367 6425
rect 35625 6399 35631 6425
rect 35657 6399 35663 6425
rect 37249 6399 37255 6425
rect 37281 6399 37287 6425
rect 672 6285 39312 6302
rect 672 6259 4574 6285
rect 4600 6259 4636 6285
rect 4662 6259 4698 6285
rect 4724 6259 4760 6285
rect 4786 6259 4822 6285
rect 4848 6259 4884 6285
rect 4910 6259 4946 6285
rect 4972 6259 5008 6285
rect 5034 6259 9574 6285
rect 9600 6259 9636 6285
rect 9662 6259 9698 6285
rect 9724 6259 9760 6285
rect 9786 6259 9822 6285
rect 9848 6259 9884 6285
rect 9910 6259 9946 6285
rect 9972 6259 10008 6285
rect 10034 6259 14574 6285
rect 14600 6259 14636 6285
rect 14662 6259 14698 6285
rect 14724 6259 14760 6285
rect 14786 6259 14822 6285
rect 14848 6259 14884 6285
rect 14910 6259 14946 6285
rect 14972 6259 15008 6285
rect 15034 6259 19574 6285
rect 19600 6259 19636 6285
rect 19662 6259 19698 6285
rect 19724 6259 19760 6285
rect 19786 6259 19822 6285
rect 19848 6259 19884 6285
rect 19910 6259 19946 6285
rect 19972 6259 20008 6285
rect 20034 6259 24574 6285
rect 24600 6259 24636 6285
rect 24662 6259 24698 6285
rect 24724 6259 24760 6285
rect 24786 6259 24822 6285
rect 24848 6259 24884 6285
rect 24910 6259 24946 6285
rect 24972 6259 25008 6285
rect 25034 6259 29574 6285
rect 29600 6259 29636 6285
rect 29662 6259 29698 6285
rect 29724 6259 29760 6285
rect 29786 6259 29822 6285
rect 29848 6259 29884 6285
rect 29910 6259 29946 6285
rect 29972 6259 30008 6285
rect 30034 6259 34574 6285
rect 34600 6259 34636 6285
rect 34662 6259 34698 6285
rect 34724 6259 34760 6285
rect 34786 6259 34822 6285
rect 34848 6259 34884 6285
rect 34910 6259 34946 6285
rect 34972 6259 35008 6285
rect 35034 6259 39312 6285
rect 672 6242 39312 6259
rect 1857 6119 1863 6145
rect 1889 6119 1895 6145
rect 8241 6119 8247 6145
rect 8273 6119 8279 6145
rect 16417 6119 16423 6145
rect 16449 6119 16455 6145
rect 18433 6119 18439 6145
rect 18465 6119 18471 6145
rect 20001 6119 20007 6145
rect 20033 6119 20039 6145
rect 21793 6119 21799 6145
rect 21825 6119 21831 6145
rect 23417 6119 23423 6145
rect 23449 6119 23455 6145
rect 27393 6119 27399 6145
rect 27425 6119 27431 6145
rect 30193 6119 30199 6145
rect 30225 6119 30231 6145
rect 31817 6119 31823 6145
rect 31849 6119 31855 6145
rect 35345 6119 35351 6145
rect 35377 6119 35383 6145
rect 35631 6089 35657 6095
rect 1857 6063 1863 6089
rect 1889 6063 1895 6089
rect 2753 6063 2759 6089
rect 2785 6063 2791 6089
rect 3593 6063 3599 6089
rect 3625 6063 3631 6089
rect 3873 6063 3879 6089
rect 3905 6063 3911 6089
rect 3985 6063 3991 6089
rect 4017 6063 4023 6089
rect 6001 6063 6007 6089
rect 6033 6063 6039 6089
rect 6393 6063 6399 6089
rect 6425 6063 6431 6089
rect 6505 6063 6511 6089
rect 6537 6063 6543 6089
rect 7569 6063 7575 6089
rect 7601 6063 7607 6089
rect 8241 6063 8247 6089
rect 8273 6063 8279 6089
rect 10033 6063 10039 6089
rect 10065 6063 10071 6089
rect 10369 6063 10375 6089
rect 10401 6063 10407 6089
rect 10481 6063 10487 6089
rect 10513 6063 10519 6089
rect 11545 6063 11551 6089
rect 11577 6063 11583 6089
rect 11825 6063 11831 6089
rect 11857 6063 11863 6089
rect 11937 6063 11943 6089
rect 11969 6063 11975 6089
rect 13113 6063 13119 6089
rect 13145 6063 13151 6089
rect 13281 6063 13287 6089
rect 13313 6063 13319 6089
rect 13505 6063 13511 6089
rect 13537 6063 13543 6089
rect 15521 6063 15527 6089
rect 15553 6063 15559 6089
rect 16417 6063 16423 6089
rect 16449 6063 16455 6089
rect 17593 6063 17599 6089
rect 17625 6063 17631 6089
rect 18433 6063 18439 6089
rect 18465 6063 18471 6089
rect 19105 6063 19111 6089
rect 19137 6063 19143 6089
rect 20001 6063 20007 6089
rect 20033 6063 20039 6089
rect 20785 6063 20791 6089
rect 20817 6063 20823 6089
rect 21793 6063 21799 6089
rect 21825 6063 21831 6089
rect 22521 6063 22527 6089
rect 22553 6063 22559 6089
rect 23417 6063 23423 6089
rect 23449 6063 23455 6089
rect 25041 6063 25047 6089
rect 25073 6063 25079 6089
rect 25209 6063 25215 6089
rect 25241 6063 25247 6089
rect 25433 6063 25439 6089
rect 25465 6063 25471 6089
rect 26217 6063 26223 6089
rect 26249 6063 26255 6089
rect 27393 6063 27399 6089
rect 27425 6063 27431 6089
rect 29353 6063 29359 6089
rect 29385 6063 29391 6089
rect 30193 6063 30199 6089
rect 30225 6063 30231 6089
rect 30921 6063 30927 6089
rect 30953 6063 30959 6089
rect 31817 6063 31823 6089
rect 31849 6063 31855 6089
rect 32713 6063 32719 6089
rect 32745 6063 32751 6089
rect 33273 6063 33279 6089
rect 33305 6063 33311 6089
rect 33385 6063 33391 6089
rect 33417 6063 33423 6089
rect 34449 6063 34455 6089
rect 34481 6063 34487 6089
rect 35345 6063 35351 6089
rect 35377 6063 35383 6089
rect 35631 6057 35657 6063
rect 35743 6089 35769 6095
rect 35743 6057 35769 6063
rect 35911 6089 35937 6095
rect 36689 6063 36695 6089
rect 36721 6063 36727 6089
rect 37249 6063 37255 6089
rect 37281 6063 37287 6089
rect 37361 6063 37367 6089
rect 37393 6063 37399 6089
rect 35911 6057 35937 6063
rect 672 5893 39312 5910
rect 672 5867 2074 5893
rect 2100 5867 2136 5893
rect 2162 5867 2198 5893
rect 2224 5867 2260 5893
rect 2286 5867 2322 5893
rect 2348 5867 2384 5893
rect 2410 5867 2446 5893
rect 2472 5867 2508 5893
rect 2534 5867 7074 5893
rect 7100 5867 7136 5893
rect 7162 5867 7198 5893
rect 7224 5867 7260 5893
rect 7286 5867 7322 5893
rect 7348 5867 7384 5893
rect 7410 5867 7446 5893
rect 7472 5867 7508 5893
rect 7534 5867 12074 5893
rect 12100 5867 12136 5893
rect 12162 5867 12198 5893
rect 12224 5867 12260 5893
rect 12286 5867 12322 5893
rect 12348 5867 12384 5893
rect 12410 5867 12446 5893
rect 12472 5867 12508 5893
rect 12534 5867 17074 5893
rect 17100 5867 17136 5893
rect 17162 5867 17198 5893
rect 17224 5867 17260 5893
rect 17286 5867 17322 5893
rect 17348 5867 17384 5893
rect 17410 5867 17446 5893
rect 17472 5867 17508 5893
rect 17534 5867 22074 5893
rect 22100 5867 22136 5893
rect 22162 5867 22198 5893
rect 22224 5867 22260 5893
rect 22286 5867 22322 5893
rect 22348 5867 22384 5893
rect 22410 5867 22446 5893
rect 22472 5867 22508 5893
rect 22534 5867 27074 5893
rect 27100 5867 27136 5893
rect 27162 5867 27198 5893
rect 27224 5867 27260 5893
rect 27286 5867 27322 5893
rect 27348 5867 27384 5893
rect 27410 5867 27446 5893
rect 27472 5867 27508 5893
rect 27534 5867 32074 5893
rect 32100 5867 32136 5893
rect 32162 5867 32198 5893
rect 32224 5867 32260 5893
rect 32286 5867 32322 5893
rect 32348 5867 32384 5893
rect 32410 5867 32446 5893
rect 32472 5867 32508 5893
rect 32534 5867 37074 5893
rect 37100 5867 37136 5893
rect 37162 5867 37198 5893
rect 37224 5867 37260 5893
rect 37286 5867 37322 5893
rect 37348 5867 37384 5893
rect 37410 5867 37446 5893
rect 37472 5867 37508 5893
rect 37534 5867 39312 5893
rect 672 5850 39312 5867
rect 33671 5697 33697 5703
rect 1801 5671 1807 5697
rect 1833 5671 1839 5697
rect 1913 5671 1919 5697
rect 1945 5671 1951 5697
rect 2473 5671 2479 5697
rect 2505 5671 2511 5697
rect 4097 5671 4103 5697
rect 4129 5671 4135 5697
rect 4377 5671 4383 5697
rect 4409 5671 4415 5697
rect 4489 5671 4495 5697
rect 4521 5671 4527 5697
rect 5553 5671 5559 5697
rect 5585 5671 5591 5697
rect 6449 5671 6455 5697
rect 6481 5671 6487 5697
rect 8073 5671 8079 5697
rect 8105 5671 8111 5697
rect 8969 5671 8975 5697
rect 9001 5671 9007 5697
rect 9529 5671 9535 5697
rect 9561 5671 9567 5697
rect 10425 5671 10431 5697
rect 10457 5671 10463 5697
rect 12329 5671 12335 5697
rect 12361 5671 12367 5697
rect 12497 5671 12503 5697
rect 12529 5671 12535 5697
rect 12721 5671 12727 5697
rect 12753 5671 12759 5697
rect 15745 5671 15751 5697
rect 15777 5671 15783 5697
rect 16753 5671 16759 5697
rect 16785 5671 16791 5697
rect 17481 5671 17487 5697
rect 17513 5671 17519 5697
rect 18377 5671 18383 5697
rect 18409 5671 18415 5697
rect 19049 5671 19055 5697
rect 19081 5671 19087 5697
rect 19945 5671 19951 5697
rect 19977 5671 19983 5697
rect 20505 5671 20511 5697
rect 20537 5671 20543 5697
rect 21345 5671 21351 5697
rect 21377 5671 21383 5697
rect 23025 5671 23031 5697
rect 23057 5671 23063 5697
rect 23865 5671 23871 5697
rect 23897 5671 23903 5697
rect 24425 5671 24431 5697
rect 24457 5671 24463 5697
rect 25153 5671 25159 5697
rect 25185 5671 25191 5697
rect 26889 5671 26895 5697
rect 26921 5671 26927 5697
rect 27617 5671 27623 5697
rect 27649 5671 27655 5697
rect 29353 5671 29359 5697
rect 29385 5671 29391 5697
rect 30193 5671 30199 5697
rect 30225 5671 30231 5697
rect 30977 5671 30983 5697
rect 31009 5671 31015 5697
rect 31873 5671 31879 5697
rect 31905 5671 31911 5697
rect 32433 5671 32439 5697
rect 32465 5671 32471 5697
rect 33329 5671 33335 5697
rect 33361 5671 33367 5697
rect 33671 5665 33697 5671
rect 33895 5697 33921 5703
rect 34673 5671 34679 5697
rect 34705 5671 34711 5697
rect 35233 5671 35239 5697
rect 35265 5671 35271 5697
rect 35345 5671 35351 5697
rect 35377 5671 35383 5697
rect 36129 5671 36135 5697
rect 36161 5671 36167 5697
rect 37305 5671 37311 5697
rect 37337 5671 37343 5697
rect 33895 5665 33921 5671
rect 33727 5641 33753 5647
rect 37591 5641 37617 5647
rect 6449 5615 6455 5641
rect 6481 5615 6487 5641
rect 8969 5615 8975 5641
rect 9001 5615 9007 5641
rect 10425 5615 10431 5641
rect 10457 5615 10463 5641
rect 16753 5615 16759 5641
rect 16785 5615 16791 5641
rect 18377 5615 18383 5641
rect 18409 5615 18415 5641
rect 19945 5615 19951 5641
rect 19977 5615 19983 5641
rect 21345 5615 21351 5641
rect 21377 5615 21383 5641
rect 23865 5615 23871 5641
rect 23897 5615 23903 5641
rect 25153 5615 25159 5641
rect 25185 5615 25191 5641
rect 27673 5615 27679 5641
rect 27705 5615 27711 5641
rect 30193 5615 30199 5641
rect 30225 5615 30231 5641
rect 31873 5615 31879 5641
rect 31905 5615 31911 5641
rect 33329 5615 33335 5641
rect 33361 5615 33367 5641
rect 37305 5615 37311 5641
rect 37337 5615 37343 5641
rect 33727 5609 33753 5615
rect 37591 5609 37617 5615
rect 37703 5641 37729 5647
rect 37703 5609 37729 5615
rect 37871 5641 37897 5647
rect 37871 5609 37897 5615
rect 672 5501 39312 5518
rect 672 5475 4574 5501
rect 4600 5475 4636 5501
rect 4662 5475 4698 5501
rect 4724 5475 4760 5501
rect 4786 5475 4822 5501
rect 4848 5475 4884 5501
rect 4910 5475 4946 5501
rect 4972 5475 5008 5501
rect 5034 5475 9574 5501
rect 9600 5475 9636 5501
rect 9662 5475 9698 5501
rect 9724 5475 9760 5501
rect 9786 5475 9822 5501
rect 9848 5475 9884 5501
rect 9910 5475 9946 5501
rect 9972 5475 10008 5501
rect 10034 5475 14574 5501
rect 14600 5475 14636 5501
rect 14662 5475 14698 5501
rect 14724 5475 14760 5501
rect 14786 5475 14822 5501
rect 14848 5475 14884 5501
rect 14910 5475 14946 5501
rect 14972 5475 15008 5501
rect 15034 5475 19574 5501
rect 19600 5475 19636 5501
rect 19662 5475 19698 5501
rect 19724 5475 19760 5501
rect 19786 5475 19822 5501
rect 19848 5475 19884 5501
rect 19910 5475 19946 5501
rect 19972 5475 20008 5501
rect 20034 5475 24574 5501
rect 24600 5475 24636 5501
rect 24662 5475 24698 5501
rect 24724 5475 24760 5501
rect 24786 5475 24822 5501
rect 24848 5475 24884 5501
rect 24910 5475 24946 5501
rect 24972 5475 25008 5501
rect 25034 5475 29574 5501
rect 29600 5475 29636 5501
rect 29662 5475 29698 5501
rect 29724 5475 29760 5501
rect 29786 5475 29822 5501
rect 29848 5475 29884 5501
rect 29910 5475 29946 5501
rect 29972 5475 30008 5501
rect 30034 5475 34574 5501
rect 34600 5475 34636 5501
rect 34662 5475 34698 5501
rect 34724 5475 34760 5501
rect 34786 5475 34822 5501
rect 34848 5475 34884 5501
rect 34910 5475 34946 5501
rect 34972 5475 35008 5501
rect 35034 5475 39312 5501
rect 672 5458 39312 5475
rect 35911 5361 35937 5367
rect 1857 5335 1863 5361
rect 1889 5335 1895 5361
rect 4433 5335 4439 5361
rect 4465 5335 4471 5361
rect 16417 5335 16423 5361
rect 16449 5335 16455 5361
rect 18433 5335 18439 5361
rect 18465 5335 18471 5361
rect 20001 5335 20007 5361
rect 20033 5335 20039 5361
rect 23417 5335 23423 5361
rect 23449 5335 23455 5361
rect 30193 5335 30199 5361
rect 30225 5335 30231 5361
rect 31817 5335 31823 5361
rect 31849 5335 31855 5361
rect 37641 5335 37647 5361
rect 37673 5335 37679 5361
rect 35911 5329 35937 5335
rect 35631 5305 35657 5311
rect 1857 5279 1863 5305
rect 1889 5279 1895 5305
rect 2753 5279 2759 5305
rect 2785 5279 2791 5305
rect 3593 5279 3599 5305
rect 3625 5279 3631 5305
rect 4433 5279 4439 5305
rect 4465 5279 4471 5305
rect 6001 5279 6007 5305
rect 6033 5279 6039 5305
rect 6393 5279 6399 5305
rect 6425 5279 6431 5305
rect 6505 5279 6511 5305
rect 6537 5279 6543 5305
rect 7513 5279 7519 5305
rect 7545 5279 7551 5305
rect 7737 5279 7743 5305
rect 7769 5279 7775 5305
rect 7961 5279 7967 5305
rect 7993 5279 7999 5305
rect 9809 5279 9815 5305
rect 9841 5279 9847 5305
rect 10257 5279 10263 5305
rect 10289 5279 10295 5305
rect 10481 5279 10487 5305
rect 10513 5279 10519 5305
rect 11545 5279 11551 5305
rect 11577 5279 11583 5305
rect 11825 5279 11831 5305
rect 11857 5279 11863 5305
rect 11937 5279 11943 5305
rect 11969 5279 11975 5305
rect 13113 5279 13119 5305
rect 13145 5279 13151 5305
rect 13281 5279 13287 5305
rect 13313 5279 13319 5305
rect 13505 5279 13511 5305
rect 13537 5279 13543 5305
rect 15353 5279 15359 5305
rect 15385 5279 15391 5305
rect 16417 5279 16423 5305
rect 16449 5279 16455 5305
rect 17593 5279 17599 5305
rect 17625 5279 17631 5305
rect 18433 5279 18439 5305
rect 18465 5279 18471 5305
rect 19049 5279 19055 5305
rect 19081 5279 19087 5305
rect 20001 5279 20007 5305
rect 20033 5279 20039 5305
rect 20841 5279 20847 5305
rect 20873 5279 20879 5305
rect 21345 5279 21351 5305
rect 21377 5279 21383 5305
rect 21457 5279 21463 5305
rect 21489 5279 21495 5305
rect 22521 5279 22527 5305
rect 22553 5279 22559 5305
rect 23417 5279 23423 5305
rect 23449 5279 23455 5305
rect 25041 5279 25047 5305
rect 25073 5279 25079 5305
rect 25209 5279 25215 5305
rect 25241 5279 25247 5305
rect 25433 5279 25439 5305
rect 25465 5279 25471 5305
rect 26497 5279 26503 5305
rect 26529 5279 26535 5305
rect 26777 5279 26783 5305
rect 26809 5279 26815 5305
rect 26889 5279 26895 5305
rect 26921 5279 26927 5305
rect 29353 5279 29359 5305
rect 29385 5279 29391 5305
rect 30193 5279 30199 5305
rect 30225 5279 30231 5305
rect 30921 5279 30927 5305
rect 30953 5279 30959 5305
rect 31817 5279 31823 5305
rect 31849 5279 31855 5305
rect 32713 5279 32719 5305
rect 32745 5279 32751 5305
rect 33273 5279 33279 5305
rect 33305 5279 33311 5305
rect 33385 5279 33391 5305
rect 33417 5279 33423 5305
rect 34169 5279 34175 5305
rect 34201 5279 34207 5305
rect 34617 5279 34623 5305
rect 34649 5279 34655 5305
rect 34841 5279 34847 5305
rect 34873 5279 34879 5305
rect 35631 5273 35657 5279
rect 35743 5305 35769 5311
rect 36689 5279 36695 5305
rect 36721 5279 36727 5305
rect 37641 5279 37647 5305
rect 37673 5279 37679 5305
rect 35743 5273 35769 5279
rect 672 5109 39312 5126
rect 672 5083 2074 5109
rect 2100 5083 2136 5109
rect 2162 5083 2198 5109
rect 2224 5083 2260 5109
rect 2286 5083 2322 5109
rect 2348 5083 2384 5109
rect 2410 5083 2446 5109
rect 2472 5083 2508 5109
rect 2534 5083 7074 5109
rect 7100 5083 7136 5109
rect 7162 5083 7198 5109
rect 7224 5083 7260 5109
rect 7286 5083 7322 5109
rect 7348 5083 7384 5109
rect 7410 5083 7446 5109
rect 7472 5083 7508 5109
rect 7534 5083 12074 5109
rect 12100 5083 12136 5109
rect 12162 5083 12198 5109
rect 12224 5083 12260 5109
rect 12286 5083 12322 5109
rect 12348 5083 12384 5109
rect 12410 5083 12446 5109
rect 12472 5083 12508 5109
rect 12534 5083 17074 5109
rect 17100 5083 17136 5109
rect 17162 5083 17198 5109
rect 17224 5083 17260 5109
rect 17286 5083 17322 5109
rect 17348 5083 17384 5109
rect 17410 5083 17446 5109
rect 17472 5083 17508 5109
rect 17534 5083 22074 5109
rect 22100 5083 22136 5109
rect 22162 5083 22198 5109
rect 22224 5083 22260 5109
rect 22286 5083 22322 5109
rect 22348 5083 22384 5109
rect 22410 5083 22446 5109
rect 22472 5083 22508 5109
rect 22534 5083 27074 5109
rect 27100 5083 27136 5109
rect 27162 5083 27198 5109
rect 27224 5083 27260 5109
rect 27286 5083 27322 5109
rect 27348 5083 27384 5109
rect 27410 5083 27446 5109
rect 27472 5083 27508 5109
rect 27534 5083 32074 5109
rect 32100 5083 32136 5109
rect 32162 5083 32198 5109
rect 32224 5083 32260 5109
rect 32286 5083 32322 5109
rect 32348 5083 32384 5109
rect 32410 5083 32446 5109
rect 32472 5083 32508 5109
rect 32534 5083 37074 5109
rect 37100 5083 37136 5109
rect 37162 5083 37198 5109
rect 37224 5083 37260 5109
rect 37286 5083 37322 5109
rect 37348 5083 37384 5109
rect 37410 5083 37446 5109
rect 37472 5083 37508 5109
rect 37534 5083 39312 5109
rect 672 5066 39312 5083
rect 30143 4913 30169 4919
rect 1801 4887 1807 4913
rect 1833 4887 1839 4913
rect 1913 4887 1919 4913
rect 1945 4887 1951 4913
rect 2473 4887 2479 4913
rect 2505 4887 2511 4913
rect 4097 4887 4103 4913
rect 4129 4887 4135 4913
rect 4377 4887 4383 4913
rect 4409 4887 4415 4913
rect 4489 4887 4495 4913
rect 4521 4887 4527 4913
rect 5553 4887 5559 4913
rect 5585 4887 5591 4913
rect 6393 4887 6399 4913
rect 6425 4887 6431 4913
rect 7793 4887 7799 4913
rect 7825 4887 7831 4913
rect 8241 4887 8247 4913
rect 8273 4887 8279 4913
rect 8465 4887 8471 4913
rect 8497 4887 8503 4913
rect 9529 4887 9535 4913
rect 9561 4887 9567 4913
rect 10257 4887 10263 4913
rect 10289 4887 10295 4913
rect 12329 4887 12335 4913
rect 12361 4887 12367 4913
rect 12609 4887 12615 4913
rect 12641 4887 12647 4913
rect 12721 4887 12727 4913
rect 12753 4887 12759 4913
rect 15745 4887 15751 4913
rect 15777 4887 15783 4913
rect 16753 4887 16759 4913
rect 16785 4887 16791 4913
rect 17481 4887 17487 4913
rect 17513 4887 17519 4913
rect 18377 4887 18383 4913
rect 18409 4887 18415 4913
rect 19049 4887 19055 4913
rect 19081 4887 19087 4913
rect 19945 4887 19951 4913
rect 19977 4887 19983 4913
rect 20505 4887 20511 4913
rect 20537 4887 20543 4913
rect 21345 4887 21351 4913
rect 21377 4887 21383 4913
rect 23025 4887 23031 4913
rect 23057 4887 23063 4913
rect 23865 4887 23871 4913
rect 23897 4887 23903 4913
rect 24481 4887 24487 4913
rect 24513 4887 24519 4913
rect 24649 4887 24655 4913
rect 24681 4887 24687 4913
rect 24873 4887 24879 4913
rect 24905 4887 24911 4913
rect 26889 4887 26895 4913
rect 26921 4887 26927 4913
rect 27169 4887 27175 4913
rect 27201 4887 27207 4913
rect 27393 4887 27399 4913
rect 27425 4887 27431 4913
rect 28457 4887 28463 4913
rect 28489 4887 28495 4913
rect 29297 4887 29303 4913
rect 29329 4887 29335 4913
rect 30143 4881 30169 4887
rect 30367 4913 30393 4919
rect 33671 4913 33697 4919
rect 30977 4887 30983 4913
rect 31009 4887 31015 4913
rect 31873 4887 31879 4913
rect 31905 4887 31911 4913
rect 32153 4887 32159 4913
rect 32185 4887 32191 4913
rect 33329 4887 33335 4913
rect 33361 4887 33367 4913
rect 34673 4887 34679 4913
rect 34705 4887 34711 4913
rect 35233 4887 35239 4913
rect 35265 4887 35271 4913
rect 35345 4887 35351 4913
rect 35377 4887 35383 4913
rect 36129 4887 36135 4913
rect 36161 4887 36167 4913
rect 37305 4887 37311 4913
rect 37337 4887 37343 4913
rect 30367 4881 30393 4887
rect 33671 4881 33697 4887
rect 30031 4857 30057 4863
rect 33727 4857 33753 4863
rect 6393 4831 6399 4857
rect 6425 4831 6431 4857
rect 10257 4831 10263 4857
rect 10289 4831 10295 4857
rect 16753 4831 16759 4857
rect 16785 4831 16791 4857
rect 18377 4831 18383 4857
rect 18409 4831 18415 4857
rect 19945 4831 19951 4857
rect 19977 4831 19983 4857
rect 21345 4831 21351 4857
rect 21377 4831 21383 4857
rect 23865 4831 23871 4857
rect 23897 4831 23903 4857
rect 29297 4831 29303 4857
rect 29329 4831 29335 4857
rect 31873 4831 31879 4857
rect 31905 4831 31911 4857
rect 33329 4831 33335 4857
rect 33361 4831 33367 4857
rect 30031 4825 30057 4831
rect 33727 4825 33753 4831
rect 33895 4857 33921 4863
rect 37591 4857 37617 4863
rect 37305 4831 37311 4857
rect 37337 4831 37343 4857
rect 33895 4825 33921 4831
rect 37591 4825 37617 4831
rect 37703 4857 37729 4863
rect 37703 4825 37729 4831
rect 37871 4857 37897 4863
rect 37871 4825 37897 4831
rect 38655 4857 38681 4863
rect 38655 4825 38681 4831
rect 38767 4857 38793 4863
rect 38767 4825 38793 4831
rect 38935 4857 38961 4863
rect 38935 4825 38961 4831
rect 672 4717 39312 4734
rect 672 4691 4574 4717
rect 4600 4691 4636 4717
rect 4662 4691 4698 4717
rect 4724 4691 4760 4717
rect 4786 4691 4822 4717
rect 4848 4691 4884 4717
rect 4910 4691 4946 4717
rect 4972 4691 5008 4717
rect 5034 4691 9574 4717
rect 9600 4691 9636 4717
rect 9662 4691 9698 4717
rect 9724 4691 9760 4717
rect 9786 4691 9822 4717
rect 9848 4691 9884 4717
rect 9910 4691 9946 4717
rect 9972 4691 10008 4717
rect 10034 4691 14574 4717
rect 14600 4691 14636 4717
rect 14662 4691 14698 4717
rect 14724 4691 14760 4717
rect 14786 4691 14822 4717
rect 14848 4691 14884 4717
rect 14910 4691 14946 4717
rect 14972 4691 15008 4717
rect 15034 4691 19574 4717
rect 19600 4691 19636 4717
rect 19662 4691 19698 4717
rect 19724 4691 19760 4717
rect 19786 4691 19822 4717
rect 19848 4691 19884 4717
rect 19910 4691 19946 4717
rect 19972 4691 20008 4717
rect 20034 4691 24574 4717
rect 24600 4691 24636 4717
rect 24662 4691 24698 4717
rect 24724 4691 24760 4717
rect 24786 4691 24822 4717
rect 24848 4691 24884 4717
rect 24910 4691 24946 4717
rect 24972 4691 25008 4717
rect 25034 4691 29574 4717
rect 29600 4691 29636 4717
rect 29662 4691 29698 4717
rect 29724 4691 29760 4717
rect 29786 4691 29822 4717
rect 29848 4691 29884 4717
rect 29910 4691 29946 4717
rect 29972 4691 30008 4717
rect 30034 4691 34574 4717
rect 34600 4691 34636 4717
rect 34662 4691 34698 4717
rect 34724 4691 34760 4717
rect 34786 4691 34822 4717
rect 34848 4691 34884 4717
rect 34910 4691 34946 4717
rect 34972 4691 35008 4717
rect 35034 4691 39312 4717
rect 672 4674 39312 4691
rect 28071 4577 28097 4583
rect 1857 4551 1863 4577
rect 1889 4551 1895 4577
rect 4433 4551 4439 4577
rect 4465 4551 4471 4577
rect 6953 4551 6959 4577
rect 6985 4551 6991 4577
rect 8241 4551 8247 4577
rect 8273 4551 8279 4577
rect 14737 4551 14743 4577
rect 14769 4551 14775 4577
rect 16417 4551 16423 4577
rect 16449 4551 16455 4577
rect 18433 4551 18439 4577
rect 18465 4551 18471 4577
rect 20001 4551 20007 4577
rect 20033 4551 20039 4577
rect 21793 4551 21799 4577
rect 21825 4551 21831 4577
rect 27169 4551 27175 4577
rect 27201 4551 27207 4577
rect 28071 4545 28097 4551
rect 28239 4577 28265 4583
rect 31369 4551 31375 4577
rect 31401 4551 31407 4577
rect 35345 4551 35351 4577
rect 35377 4551 35383 4577
rect 37641 4551 37647 4577
rect 37673 4551 37679 4577
rect 28239 4545 28265 4551
rect 28351 4521 28377 4527
rect 32047 4521 32073 4527
rect 1857 4495 1863 4521
rect 1889 4495 1895 4521
rect 2753 4495 2759 4521
rect 2785 4495 2791 4521
rect 3313 4495 3319 4521
rect 3345 4495 3351 4521
rect 4433 4495 4439 4521
rect 4465 4495 4471 4521
rect 6001 4495 6007 4521
rect 6033 4495 6039 4521
rect 6953 4495 6959 4521
rect 6985 4495 6991 4521
rect 7289 4495 7295 4521
rect 7321 4495 7327 4521
rect 8241 4495 8247 4521
rect 8273 4495 8279 4521
rect 10033 4495 10039 4521
rect 10065 4495 10071 4521
rect 10257 4495 10263 4521
rect 10289 4495 10295 4521
rect 10481 4495 10487 4521
rect 10513 4495 10519 4521
rect 11489 4495 11495 4521
rect 11521 4495 11527 4521
rect 11769 4495 11775 4521
rect 11801 4495 11807 4521
rect 11937 4495 11943 4521
rect 11969 4495 11975 4521
rect 14065 4495 14071 4521
rect 14097 4495 14103 4521
rect 14737 4495 14743 4521
rect 14769 4495 14775 4521
rect 15353 4495 15359 4521
rect 15385 4495 15391 4521
rect 16417 4495 16423 4521
rect 16449 4495 16455 4521
rect 17593 4495 17599 4521
rect 17625 4495 17631 4521
rect 18433 4495 18439 4521
rect 18465 4495 18471 4521
rect 19105 4495 19111 4521
rect 19137 4495 19143 4521
rect 20001 4495 20007 4521
rect 20033 4495 20039 4521
rect 20841 4495 20847 4521
rect 20873 4495 20879 4521
rect 21793 4495 21799 4521
rect 21825 4495 21831 4521
rect 22521 4495 22527 4521
rect 22553 4495 22559 4521
rect 22689 4495 22695 4521
rect 22721 4495 22727 4521
rect 22913 4495 22919 4521
rect 22945 4495 22951 4521
rect 24761 4495 24767 4521
rect 24793 4495 24799 4521
rect 25209 4495 25215 4521
rect 25241 4495 25247 4521
rect 25433 4495 25439 4521
rect 25465 4495 25471 4521
rect 26497 4495 26503 4521
rect 26529 4495 26535 4521
rect 26889 4495 26895 4521
rect 26921 4495 26927 4521
rect 28737 4495 28743 4521
rect 28769 4495 28775 4521
rect 29297 4495 29303 4521
rect 29329 4495 29335 4521
rect 29409 4495 29415 4521
rect 29441 4495 29447 4521
rect 30473 4495 30479 4521
rect 30505 4495 30511 4521
rect 31369 4495 31375 4521
rect 31401 4495 31407 4521
rect 28351 4489 28377 4495
rect 32047 4489 32073 4495
rect 32159 4521 32185 4527
rect 32159 4489 32185 4495
rect 32327 4521 32353 4527
rect 35687 4521 35713 4527
rect 32713 4495 32719 4521
rect 32745 4495 32751 4521
rect 33273 4495 33279 4521
rect 33305 4495 33311 4521
rect 33385 4495 33391 4521
rect 33417 4495 33423 4521
rect 34449 4495 34455 4521
rect 34481 4495 34487 4521
rect 35345 4495 35351 4521
rect 35377 4495 35383 4521
rect 32327 4489 32353 4495
rect 35687 4489 35713 4495
rect 35799 4521 35825 4527
rect 35799 4489 35825 4495
rect 35967 4521 35993 4527
rect 38207 4521 38233 4527
rect 36689 4495 36695 4521
rect 36721 4495 36727 4521
rect 37641 4495 37647 4521
rect 37673 4495 37679 4521
rect 35967 4489 35993 4495
rect 38207 4489 38233 4495
rect 38263 4521 38289 4527
rect 38263 4489 38289 4495
rect 38431 4521 38457 4527
rect 38431 4489 38457 4495
rect 38711 4521 38737 4527
rect 38711 4489 38737 4495
rect 38823 4521 38849 4527
rect 38823 4489 38849 4495
rect 38991 4521 39017 4527
rect 38991 4489 39017 4495
rect 672 4325 39312 4342
rect 672 4299 2074 4325
rect 2100 4299 2136 4325
rect 2162 4299 2198 4325
rect 2224 4299 2260 4325
rect 2286 4299 2322 4325
rect 2348 4299 2384 4325
rect 2410 4299 2446 4325
rect 2472 4299 2508 4325
rect 2534 4299 7074 4325
rect 7100 4299 7136 4325
rect 7162 4299 7198 4325
rect 7224 4299 7260 4325
rect 7286 4299 7322 4325
rect 7348 4299 7384 4325
rect 7410 4299 7446 4325
rect 7472 4299 7508 4325
rect 7534 4299 12074 4325
rect 12100 4299 12136 4325
rect 12162 4299 12198 4325
rect 12224 4299 12260 4325
rect 12286 4299 12322 4325
rect 12348 4299 12384 4325
rect 12410 4299 12446 4325
rect 12472 4299 12508 4325
rect 12534 4299 17074 4325
rect 17100 4299 17136 4325
rect 17162 4299 17198 4325
rect 17224 4299 17260 4325
rect 17286 4299 17322 4325
rect 17348 4299 17384 4325
rect 17410 4299 17446 4325
rect 17472 4299 17508 4325
rect 17534 4299 22074 4325
rect 22100 4299 22136 4325
rect 22162 4299 22198 4325
rect 22224 4299 22260 4325
rect 22286 4299 22322 4325
rect 22348 4299 22384 4325
rect 22410 4299 22446 4325
rect 22472 4299 22508 4325
rect 22534 4299 27074 4325
rect 27100 4299 27136 4325
rect 27162 4299 27198 4325
rect 27224 4299 27260 4325
rect 27286 4299 27322 4325
rect 27348 4299 27384 4325
rect 27410 4299 27446 4325
rect 27472 4299 27508 4325
rect 27534 4299 32074 4325
rect 32100 4299 32136 4325
rect 32162 4299 32198 4325
rect 32224 4299 32260 4325
rect 32286 4299 32322 4325
rect 32348 4299 32384 4325
rect 32410 4299 32446 4325
rect 32472 4299 32508 4325
rect 32534 4299 37074 4325
rect 37100 4299 37136 4325
rect 37162 4299 37198 4325
rect 37224 4299 37260 4325
rect 37286 4299 37322 4325
rect 37348 4299 37384 4325
rect 37410 4299 37446 4325
rect 37472 4299 37508 4325
rect 37534 4299 39312 4325
rect 672 4282 39312 4299
rect 30087 4129 30113 4135
rect 33671 4129 33697 4135
rect 38823 4129 38849 4135
rect 1801 4103 1807 4129
rect 1833 4103 1839 4129
rect 2025 4103 2031 4129
rect 2057 4103 2063 4129
rect 2473 4103 2479 4129
rect 2505 4103 2511 4129
rect 4097 4103 4103 4129
rect 4129 4103 4135 4129
rect 4993 4103 4999 4129
rect 5025 4103 5031 4129
rect 5273 4103 5279 4129
rect 5305 4103 5311 4129
rect 6449 4103 6455 4129
rect 6481 4103 6487 4129
rect 7793 4103 7799 4129
rect 7825 4103 7831 4129
rect 8969 4103 8975 4129
rect 9001 4103 9007 4129
rect 9473 4103 9479 4129
rect 9505 4103 9511 4129
rect 10425 4103 10431 4129
rect 10457 4103 10463 4129
rect 11769 4103 11775 4129
rect 11801 4103 11807 4129
rect 12945 4103 12951 4129
rect 12977 4103 12983 4129
rect 13225 4103 13231 4129
rect 13257 4103 13263 4129
rect 14401 4103 14407 4129
rect 14433 4103 14439 4129
rect 15745 4103 15751 4129
rect 15777 4103 15783 4129
rect 16249 4103 16255 4129
rect 16281 4103 16287 4129
rect 16417 4103 16423 4129
rect 16449 4103 16455 4129
rect 17481 4103 17487 4129
rect 17513 4103 17519 4129
rect 18377 4103 18383 4129
rect 18409 4103 18415 4129
rect 19049 4103 19055 4129
rect 19081 4103 19087 4129
rect 19945 4103 19951 4129
rect 19977 4103 19983 4129
rect 20505 4103 20511 4129
rect 20537 4103 20543 4129
rect 21345 4103 21351 4129
rect 21377 4103 21383 4129
rect 22745 4103 22751 4129
rect 22777 4103 22783 4129
rect 23865 4103 23871 4129
rect 23897 4103 23903 4129
rect 24481 4103 24487 4129
rect 24513 4103 24519 4129
rect 25377 4103 25383 4129
rect 25409 4103 25415 4129
rect 26833 4103 26839 4129
rect 26865 4103 26871 4129
rect 27505 4103 27511 4129
rect 27537 4103 27543 4129
rect 28457 4103 28463 4129
rect 28489 4103 28495 4129
rect 28681 4103 28687 4129
rect 28713 4103 28719 4129
rect 28905 4103 28911 4129
rect 28937 4103 28943 4129
rect 30977 4103 30983 4129
rect 31009 4103 31015 4129
rect 31873 4103 31879 4129
rect 31905 4103 31911 4129
rect 32153 4103 32159 4129
rect 32185 4103 32191 4129
rect 33329 4103 33335 4129
rect 33361 4103 33367 4129
rect 34673 4103 34679 4129
rect 34705 4103 34711 4129
rect 35849 4103 35855 4129
rect 35881 4103 35887 4129
rect 36129 4103 36135 4129
rect 36161 4103 36167 4129
rect 37081 4103 37087 4129
rect 37113 4103 37119 4129
rect 30087 4097 30113 4103
rect 33671 4097 33697 4103
rect 38823 4097 38849 4103
rect 38935 4129 38961 4135
rect 38935 4097 38961 4103
rect 30143 4073 30169 4079
rect 4993 4047 4999 4073
rect 5025 4047 5031 4073
rect 6449 4047 6455 4073
rect 6481 4047 6487 4073
rect 7793 4047 7799 4073
rect 7825 4047 7831 4073
rect 10425 4047 10431 4073
rect 10457 4047 10463 4073
rect 11769 4047 11775 4073
rect 11801 4047 11807 4073
rect 14401 4047 14407 4073
rect 14433 4047 14439 4073
rect 18377 4047 18383 4073
rect 18409 4047 18415 4073
rect 19945 4047 19951 4073
rect 19977 4047 19983 4073
rect 21345 4047 21351 4073
rect 21377 4047 21383 4073
rect 23865 4047 23871 4073
rect 23897 4047 23903 4073
rect 25377 4047 25383 4073
rect 25409 4047 25415 4073
rect 27673 4047 27679 4073
rect 27705 4047 27711 4073
rect 30143 4041 30169 4047
rect 30311 4073 30337 4079
rect 33727 4073 33753 4079
rect 31873 4047 31879 4073
rect 31905 4047 31911 4073
rect 33329 4047 33335 4073
rect 33361 4047 33367 4073
rect 30311 4041 30337 4047
rect 33727 4041 33753 4047
rect 33895 4073 33921 4079
rect 37591 4073 37617 4079
rect 35849 4047 35855 4073
rect 35881 4047 35887 4073
rect 37081 4047 37087 4073
rect 37113 4047 37119 4073
rect 33895 4041 33921 4047
rect 37591 4041 37617 4047
rect 37703 4073 37729 4079
rect 37703 4041 37729 4047
rect 37871 4073 37897 4079
rect 37871 4041 37897 4047
rect 38655 4073 38681 4079
rect 38655 4041 38681 4047
rect 672 3933 39312 3950
rect 672 3907 4574 3933
rect 4600 3907 4636 3933
rect 4662 3907 4698 3933
rect 4724 3907 4760 3933
rect 4786 3907 4822 3933
rect 4848 3907 4884 3933
rect 4910 3907 4946 3933
rect 4972 3907 5008 3933
rect 5034 3907 9574 3933
rect 9600 3907 9636 3933
rect 9662 3907 9698 3933
rect 9724 3907 9760 3933
rect 9786 3907 9822 3933
rect 9848 3907 9884 3933
rect 9910 3907 9946 3933
rect 9972 3907 10008 3933
rect 10034 3907 14574 3933
rect 14600 3907 14636 3933
rect 14662 3907 14698 3933
rect 14724 3907 14760 3933
rect 14786 3907 14822 3933
rect 14848 3907 14884 3933
rect 14910 3907 14946 3933
rect 14972 3907 15008 3933
rect 15034 3907 19574 3933
rect 19600 3907 19636 3933
rect 19662 3907 19698 3933
rect 19724 3907 19760 3933
rect 19786 3907 19822 3933
rect 19848 3907 19884 3933
rect 19910 3907 19946 3933
rect 19972 3907 20008 3933
rect 20034 3907 24574 3933
rect 24600 3907 24636 3933
rect 24662 3907 24698 3933
rect 24724 3907 24760 3933
rect 24786 3907 24822 3933
rect 24848 3907 24884 3933
rect 24910 3907 24946 3933
rect 24972 3907 25008 3933
rect 25034 3907 29574 3933
rect 29600 3907 29636 3933
rect 29662 3907 29698 3933
rect 29724 3907 29760 3933
rect 29786 3907 29822 3933
rect 29848 3907 29884 3933
rect 29910 3907 29946 3933
rect 29972 3907 30008 3933
rect 30034 3907 34574 3933
rect 34600 3907 34636 3933
rect 34662 3907 34698 3933
rect 34724 3907 34760 3933
rect 34786 3907 34822 3933
rect 34848 3907 34884 3933
rect 34910 3907 34946 3933
rect 34972 3907 35008 3933
rect 35034 3907 39312 3933
rect 672 3890 39312 3907
rect 35743 3793 35769 3799
rect 4489 3767 4495 3793
rect 4521 3767 4527 3793
rect 7009 3767 7015 3793
rect 7041 3767 7047 3793
rect 10873 3767 10879 3793
rect 10905 3767 10911 3793
rect 14961 3767 14967 3793
rect 14993 3767 14999 3793
rect 16417 3767 16423 3793
rect 16449 3767 16455 3793
rect 18377 3767 18383 3793
rect 18409 3767 18415 3793
rect 20001 3767 20007 3793
rect 20033 3767 20039 3793
rect 25937 3767 25943 3793
rect 25969 3767 25975 3793
rect 27169 3767 27175 3793
rect 27201 3767 27207 3793
rect 29689 3767 29695 3793
rect 29721 3767 29727 3793
rect 31369 3767 31375 3793
rect 31401 3767 31407 3793
rect 33889 3767 33895 3793
rect 33921 3767 33927 3793
rect 35345 3767 35351 3793
rect 35377 3767 35383 3793
rect 37641 3767 37647 3793
rect 37673 3767 37679 3793
rect 35743 3761 35769 3767
rect 28015 3737 28041 3743
rect 2361 3711 2367 3737
rect 2393 3711 2399 3737
rect 2473 3711 2479 3737
rect 2505 3711 2511 3737
rect 2977 3711 2983 3737
rect 3009 3711 3015 3737
rect 3593 3711 3599 3737
rect 3625 3711 3631 3737
rect 4489 3711 4495 3737
rect 4521 3711 4527 3737
rect 6057 3711 6063 3737
rect 6089 3711 6095 3737
rect 7009 3711 7015 3737
rect 7041 3711 7047 3737
rect 7793 3711 7799 3737
rect 7825 3711 7831 3737
rect 8017 3711 8023 3737
rect 8049 3711 8055 3737
rect 8465 3711 8471 3737
rect 8497 3711 8503 3737
rect 9809 3711 9815 3737
rect 9841 3711 9847 3737
rect 10873 3711 10879 3737
rect 10905 3711 10911 3737
rect 11377 3711 11383 3737
rect 11409 3711 11415 3737
rect 11825 3711 11831 3737
rect 11857 3711 11863 3737
rect 11937 3711 11943 3737
rect 11969 3711 11975 3737
rect 13785 3711 13791 3737
rect 13817 3711 13823 3737
rect 14961 3711 14967 3737
rect 14993 3711 14999 3737
rect 15241 3711 15247 3737
rect 15273 3711 15279 3737
rect 16417 3711 16423 3737
rect 16449 3711 16455 3737
rect 17593 3711 17599 3737
rect 17625 3711 17631 3737
rect 18377 3711 18383 3737
rect 18409 3711 18415 3737
rect 19105 3711 19111 3737
rect 19137 3711 19143 3737
rect 20001 3711 20007 3737
rect 20033 3711 20039 3737
rect 20953 3711 20959 3737
rect 20985 3711 20991 3737
rect 21345 3711 21351 3737
rect 21377 3711 21383 3737
rect 21457 3711 21463 3737
rect 21489 3711 21495 3737
rect 22521 3711 22527 3737
rect 22553 3711 22559 3737
rect 22689 3711 22695 3737
rect 22721 3711 22727 3737
rect 22913 3711 22919 3737
rect 22945 3711 22951 3737
rect 24761 3711 24767 3737
rect 24793 3711 24799 3737
rect 25937 3711 25943 3737
rect 25969 3711 25975 3737
rect 26217 3711 26223 3737
rect 26249 3711 26255 3737
rect 27169 3711 27175 3737
rect 27201 3711 27207 3737
rect 28015 3705 28041 3711
rect 28183 3737 28209 3743
rect 28183 3705 28209 3711
rect 28295 3737 28321 3743
rect 32047 3737 32073 3743
rect 28961 3711 28967 3737
rect 28993 3711 28999 3737
rect 29465 3711 29471 3737
rect 29497 3711 29503 3737
rect 30473 3711 30479 3737
rect 30505 3711 30511 3737
rect 31369 3711 31375 3737
rect 31401 3711 31407 3737
rect 28295 3705 28321 3711
rect 32047 3705 32073 3711
rect 32159 3737 32185 3743
rect 32159 3705 32185 3711
rect 32327 3737 32353 3743
rect 35687 3737 35713 3743
rect 32881 3711 32887 3737
rect 32913 3711 32919 3737
rect 33889 3711 33895 3737
rect 33921 3711 33927 3737
rect 34169 3711 34175 3737
rect 34201 3711 34207 3737
rect 35345 3711 35351 3737
rect 35377 3711 35383 3737
rect 32327 3705 32353 3711
rect 35687 3705 35713 3711
rect 35911 3737 35937 3743
rect 38151 3737 38177 3743
rect 36689 3711 36695 3737
rect 36721 3711 36727 3737
rect 37641 3711 37647 3737
rect 37673 3711 37679 3737
rect 35911 3705 35937 3711
rect 38151 3705 38177 3711
rect 38263 3737 38289 3743
rect 38263 3705 38289 3711
rect 38431 3737 38457 3743
rect 38431 3705 38457 3711
rect 38655 3737 38681 3743
rect 38655 3705 38681 3711
rect 38823 3737 38849 3743
rect 38823 3705 38849 3711
rect 38991 3737 39017 3743
rect 38991 3705 39017 3711
rect 672 3541 39312 3558
rect 672 3515 2074 3541
rect 2100 3515 2136 3541
rect 2162 3515 2198 3541
rect 2224 3515 2260 3541
rect 2286 3515 2322 3541
rect 2348 3515 2384 3541
rect 2410 3515 2446 3541
rect 2472 3515 2508 3541
rect 2534 3515 7074 3541
rect 7100 3515 7136 3541
rect 7162 3515 7198 3541
rect 7224 3515 7260 3541
rect 7286 3515 7322 3541
rect 7348 3515 7384 3541
rect 7410 3515 7446 3541
rect 7472 3515 7508 3541
rect 7534 3515 12074 3541
rect 12100 3515 12136 3541
rect 12162 3515 12198 3541
rect 12224 3515 12260 3541
rect 12286 3515 12322 3541
rect 12348 3515 12384 3541
rect 12410 3515 12446 3541
rect 12472 3515 12508 3541
rect 12534 3515 17074 3541
rect 17100 3515 17136 3541
rect 17162 3515 17198 3541
rect 17224 3515 17260 3541
rect 17286 3515 17322 3541
rect 17348 3515 17384 3541
rect 17410 3515 17446 3541
rect 17472 3515 17508 3541
rect 17534 3515 22074 3541
rect 22100 3515 22136 3541
rect 22162 3515 22198 3541
rect 22224 3515 22260 3541
rect 22286 3515 22322 3541
rect 22348 3515 22384 3541
rect 22410 3515 22446 3541
rect 22472 3515 22508 3541
rect 22534 3515 27074 3541
rect 27100 3515 27136 3541
rect 27162 3515 27198 3541
rect 27224 3515 27260 3541
rect 27286 3515 27322 3541
rect 27348 3515 27384 3541
rect 27410 3515 27446 3541
rect 27472 3515 27508 3541
rect 27534 3515 32074 3541
rect 32100 3515 32136 3541
rect 32162 3515 32198 3541
rect 32224 3515 32260 3541
rect 32286 3515 32322 3541
rect 32348 3515 32384 3541
rect 32410 3515 32446 3541
rect 32472 3515 32508 3541
rect 32534 3515 37074 3541
rect 37100 3515 37136 3541
rect 37162 3515 37198 3541
rect 37224 3515 37260 3541
rect 37286 3515 37322 3541
rect 37348 3515 37384 3541
rect 37410 3515 37446 3541
rect 37472 3515 37508 3541
rect 37534 3515 39312 3541
rect 672 3498 39312 3515
rect 33671 3345 33697 3351
rect 1353 3319 1359 3345
rect 1385 3319 1391 3345
rect 2473 3319 2479 3345
rect 2505 3319 2511 3345
rect 4097 3319 4103 3345
rect 4129 3319 4135 3345
rect 4377 3319 4383 3345
rect 4409 3319 4415 3345
rect 4489 3319 4495 3345
rect 4521 3319 4527 3345
rect 5721 3319 5727 3345
rect 5753 3319 5759 3345
rect 6001 3319 6007 3345
rect 6033 3319 6039 3345
rect 6449 3319 6455 3345
rect 6481 3319 6487 3345
rect 8297 3319 8303 3345
rect 8329 3319 8335 3345
rect 8409 3319 8415 3345
rect 8441 3319 8447 3345
rect 8969 3319 8975 3345
rect 9001 3319 9007 3345
rect 9473 3319 9479 3345
rect 9505 3319 9511 3345
rect 10425 3319 10431 3345
rect 10457 3319 10463 3345
rect 11993 3319 11999 3345
rect 12025 3319 12031 3345
rect 12329 3319 12335 3345
rect 12361 3319 12367 3345
rect 12441 3319 12447 3345
rect 12473 3319 12479 3345
rect 13225 3319 13231 3345
rect 13257 3319 13263 3345
rect 14401 3319 14407 3345
rect 14433 3319 14439 3345
rect 15745 3319 15751 3345
rect 15777 3319 15783 3345
rect 16753 3319 16759 3345
rect 16785 3319 16791 3345
rect 17481 3319 17487 3345
rect 17513 3319 17519 3345
rect 18377 3319 18383 3345
rect 18409 3319 18415 3345
rect 19049 3319 19055 3345
rect 19081 3319 19087 3345
rect 19945 3319 19951 3345
rect 19977 3319 19983 3345
rect 20505 3319 20511 3345
rect 20537 3319 20543 3345
rect 21345 3319 21351 3345
rect 21377 3319 21383 3345
rect 22745 3319 22751 3345
rect 22777 3319 22783 3345
rect 23865 3319 23871 3345
rect 23897 3319 23903 3345
rect 24425 3319 24431 3345
rect 24457 3319 24463 3345
rect 25377 3319 25383 3345
rect 25409 3319 25415 3345
rect 26889 3319 26895 3345
rect 26921 3319 26927 3345
rect 27673 3319 27679 3345
rect 27705 3319 27711 3345
rect 28457 3319 28463 3345
rect 28489 3319 28495 3345
rect 29353 3319 29359 3345
rect 29385 3319 29391 3345
rect 30697 3319 30703 3345
rect 30729 3319 30735 3345
rect 31873 3319 31879 3345
rect 31905 3319 31911 3345
rect 32433 3319 32439 3345
rect 32465 3319 32471 3345
rect 32713 3319 32719 3345
rect 32745 3319 32751 3345
rect 32825 3319 32831 3345
rect 32857 3319 32863 3345
rect 33671 3313 33697 3319
rect 33895 3345 33921 3351
rect 34673 3319 34679 3345
rect 34705 3319 34711 3345
rect 35625 3319 35631 3345
rect 35657 3319 35663 3345
rect 36129 3319 36135 3345
rect 36161 3319 36167 3345
rect 37305 3319 37311 3345
rect 37337 3319 37343 3345
rect 33895 3313 33921 3319
rect 30031 3289 30057 3295
rect 1353 3263 1359 3289
rect 1385 3263 1391 3289
rect 10425 3263 10431 3289
rect 10457 3263 10463 3289
rect 14401 3263 14407 3289
rect 14433 3263 14439 3289
rect 16753 3263 16759 3289
rect 16785 3263 16791 3289
rect 18377 3263 18383 3289
rect 18409 3263 18415 3289
rect 19945 3263 19951 3289
rect 19977 3263 19983 3289
rect 21345 3263 21351 3289
rect 21377 3263 21383 3289
rect 23865 3263 23871 3289
rect 23897 3263 23903 3289
rect 25377 3263 25383 3289
rect 25409 3263 25415 3289
rect 27673 3263 27679 3289
rect 27705 3263 27711 3289
rect 29353 3263 29359 3289
rect 29385 3263 29391 3289
rect 30031 3257 30057 3263
rect 30143 3289 30169 3295
rect 30143 3257 30169 3263
rect 30311 3289 30337 3295
rect 33727 3289 33753 3295
rect 37591 3289 37617 3295
rect 31873 3263 31879 3289
rect 31905 3263 31911 3289
rect 35625 3263 35631 3289
rect 35657 3263 35663 3289
rect 37305 3263 37311 3289
rect 37337 3263 37343 3289
rect 30311 3257 30337 3263
rect 33727 3257 33753 3263
rect 37591 3257 37617 3263
rect 37703 3289 37729 3295
rect 37703 3257 37729 3263
rect 37871 3289 37897 3295
rect 37871 3257 37897 3263
rect 38655 3289 38681 3295
rect 38655 3257 38681 3263
rect 38823 3289 38849 3295
rect 38823 3257 38849 3263
rect 38935 3289 38961 3295
rect 38935 3257 38961 3263
rect 672 3149 39312 3166
rect 672 3123 4574 3149
rect 4600 3123 4636 3149
rect 4662 3123 4698 3149
rect 4724 3123 4760 3149
rect 4786 3123 4822 3149
rect 4848 3123 4884 3149
rect 4910 3123 4946 3149
rect 4972 3123 5008 3149
rect 5034 3123 9574 3149
rect 9600 3123 9636 3149
rect 9662 3123 9698 3149
rect 9724 3123 9760 3149
rect 9786 3123 9822 3149
rect 9848 3123 9884 3149
rect 9910 3123 9946 3149
rect 9972 3123 10008 3149
rect 10034 3123 14574 3149
rect 14600 3123 14636 3149
rect 14662 3123 14698 3149
rect 14724 3123 14760 3149
rect 14786 3123 14822 3149
rect 14848 3123 14884 3149
rect 14910 3123 14946 3149
rect 14972 3123 15008 3149
rect 15034 3123 19574 3149
rect 19600 3123 19636 3149
rect 19662 3123 19698 3149
rect 19724 3123 19760 3149
rect 19786 3123 19822 3149
rect 19848 3123 19884 3149
rect 19910 3123 19946 3149
rect 19972 3123 20008 3149
rect 20034 3123 24574 3149
rect 24600 3123 24636 3149
rect 24662 3123 24698 3149
rect 24724 3123 24760 3149
rect 24786 3123 24822 3149
rect 24848 3123 24884 3149
rect 24910 3123 24946 3149
rect 24972 3123 25008 3149
rect 25034 3123 29574 3149
rect 29600 3123 29636 3149
rect 29662 3123 29698 3149
rect 29724 3123 29760 3149
rect 29786 3123 29822 3149
rect 29848 3123 29884 3149
rect 29910 3123 29946 3149
rect 29972 3123 30008 3149
rect 30034 3123 34574 3149
rect 34600 3123 34636 3149
rect 34662 3123 34698 3149
rect 34724 3123 34760 3149
rect 34786 3123 34822 3149
rect 34848 3123 34884 3149
rect 34910 3123 34946 3149
rect 34972 3123 35008 3149
rect 35034 3123 39312 3149
rect 672 3106 39312 3123
rect 28071 3009 28097 3015
rect 1969 2983 1975 3009
rect 2001 2983 2007 3009
rect 4489 2983 4495 3009
rect 4521 2983 4527 3009
rect 8465 2983 8471 3009
rect 8497 2983 8503 3009
rect 12441 2983 12447 3009
rect 12473 2983 12479 3009
rect 14961 2983 14967 3009
rect 14993 2983 14999 3009
rect 18377 2983 18383 3009
rect 18409 2983 18415 3009
rect 20001 2983 20007 3009
rect 20033 2983 20039 3009
rect 23417 2983 23423 3009
rect 23449 2983 23455 3009
rect 25937 2983 25943 3009
rect 25969 2983 25975 3009
rect 27393 2983 27399 3009
rect 27425 2983 27431 3009
rect 28071 2977 28097 2983
rect 28351 3009 28377 3015
rect 32159 3009 32185 3015
rect 29913 2983 29919 3009
rect 29945 2983 29951 3009
rect 31257 2983 31263 3009
rect 31289 2983 31295 3009
rect 28351 2977 28377 2983
rect 32159 2977 32185 2983
rect 32327 3009 32353 3015
rect 35743 3009 35769 3015
rect 35345 2983 35351 3009
rect 35377 2983 35383 3009
rect 32327 2977 32353 2983
rect 35743 2977 35769 2983
rect 35911 3009 35937 3015
rect 35911 2977 35937 2983
rect 38431 3009 38457 3015
rect 38431 2977 38457 2983
rect 28183 2953 28209 2959
rect 32047 2953 32073 2959
rect 35687 2953 35713 2959
rect 38207 2953 38233 2959
rect 1969 2927 1975 2953
rect 2001 2927 2007 2953
rect 3033 2927 3039 2953
rect 3065 2927 3071 2953
rect 3593 2927 3599 2953
rect 3625 2927 3631 2953
rect 4489 2927 4495 2953
rect 4521 2927 4527 2953
rect 6337 2927 6343 2953
rect 6369 2927 6375 2953
rect 6449 2927 6455 2953
rect 6481 2927 6487 2953
rect 7009 2927 7015 2953
rect 7041 2927 7047 2953
rect 7569 2927 7575 2953
rect 7601 2927 7607 2953
rect 8465 2927 8471 2953
rect 8497 2927 8503 2953
rect 10313 2927 10319 2953
rect 10345 2927 10351 2953
rect 10481 2927 10487 2953
rect 10513 2927 10519 2953
rect 10873 2927 10879 2953
rect 10905 2927 10911 2953
rect 11377 2927 11383 2953
rect 11409 2927 11415 2953
rect 12441 2927 12447 2953
rect 12473 2927 12479 2953
rect 14065 2927 14071 2953
rect 14097 2927 14103 2953
rect 14961 2927 14967 2953
rect 14993 2927 14999 2953
rect 15241 2927 15247 2953
rect 15273 2927 15279 2953
rect 15689 2927 15695 2953
rect 15721 2927 15727 2953
rect 16417 2927 16423 2953
rect 16449 2927 16455 2953
rect 17593 2927 17599 2953
rect 17625 2927 17631 2953
rect 18377 2927 18383 2953
rect 18409 2927 18415 2953
rect 19105 2927 19111 2953
rect 19137 2927 19143 2953
rect 20001 2927 20007 2953
rect 20033 2927 20039 2953
rect 20953 2927 20959 2953
rect 20985 2927 20991 2953
rect 21345 2927 21351 2953
rect 21377 2927 21383 2953
rect 21457 2927 21463 2953
rect 21489 2927 21495 2953
rect 22521 2927 22527 2953
rect 22553 2927 22559 2953
rect 23417 2927 23423 2953
rect 23449 2927 23455 2953
rect 24761 2927 24767 2953
rect 24793 2927 24799 2953
rect 25937 2927 25943 2953
rect 25969 2927 25975 2953
rect 26217 2927 26223 2953
rect 26249 2927 26255 2953
rect 27393 2927 27399 2953
rect 27425 2927 27431 2953
rect 28737 2927 28743 2953
rect 28769 2927 28775 2953
rect 29913 2927 29919 2953
rect 29945 2927 29951 2953
rect 30361 2927 30367 2953
rect 30393 2927 30399 2953
rect 31257 2927 31263 2953
rect 31289 2927 31295 2953
rect 32993 2927 32999 2953
rect 33025 2927 33031 2953
rect 33161 2927 33167 2953
rect 33193 2927 33199 2953
rect 33385 2927 33391 2953
rect 33417 2927 33423 2953
rect 34169 2927 34175 2953
rect 34201 2927 34207 2953
rect 35345 2927 35351 2953
rect 35377 2927 35383 2953
rect 36745 2927 36751 2953
rect 36777 2927 36783 2953
rect 37137 2927 37143 2953
rect 37169 2927 37175 2953
rect 37361 2927 37367 2953
rect 37393 2927 37399 2953
rect 28183 2921 28209 2927
rect 32047 2921 32073 2927
rect 35687 2921 35713 2927
rect 38207 2921 38233 2927
rect 38263 2953 38289 2959
rect 38263 2921 38289 2927
rect 38655 2953 38681 2959
rect 38655 2921 38681 2927
rect 38823 2953 38849 2959
rect 38823 2921 38849 2927
rect 38935 2953 38961 2959
rect 38935 2921 38961 2927
rect 672 2757 39312 2774
rect 672 2731 2074 2757
rect 2100 2731 2136 2757
rect 2162 2731 2198 2757
rect 2224 2731 2260 2757
rect 2286 2731 2322 2757
rect 2348 2731 2384 2757
rect 2410 2731 2446 2757
rect 2472 2731 2508 2757
rect 2534 2731 7074 2757
rect 7100 2731 7136 2757
rect 7162 2731 7198 2757
rect 7224 2731 7260 2757
rect 7286 2731 7322 2757
rect 7348 2731 7384 2757
rect 7410 2731 7446 2757
rect 7472 2731 7508 2757
rect 7534 2731 12074 2757
rect 12100 2731 12136 2757
rect 12162 2731 12198 2757
rect 12224 2731 12260 2757
rect 12286 2731 12322 2757
rect 12348 2731 12384 2757
rect 12410 2731 12446 2757
rect 12472 2731 12508 2757
rect 12534 2731 17074 2757
rect 17100 2731 17136 2757
rect 17162 2731 17198 2757
rect 17224 2731 17260 2757
rect 17286 2731 17322 2757
rect 17348 2731 17384 2757
rect 17410 2731 17446 2757
rect 17472 2731 17508 2757
rect 17534 2731 22074 2757
rect 22100 2731 22136 2757
rect 22162 2731 22198 2757
rect 22224 2731 22260 2757
rect 22286 2731 22322 2757
rect 22348 2731 22384 2757
rect 22410 2731 22446 2757
rect 22472 2731 22508 2757
rect 22534 2731 27074 2757
rect 27100 2731 27136 2757
rect 27162 2731 27198 2757
rect 27224 2731 27260 2757
rect 27286 2731 27322 2757
rect 27348 2731 27384 2757
rect 27410 2731 27446 2757
rect 27472 2731 27508 2757
rect 27534 2731 32074 2757
rect 32100 2731 32136 2757
rect 32162 2731 32198 2757
rect 32224 2731 32260 2757
rect 32286 2731 32322 2757
rect 32348 2731 32384 2757
rect 32410 2731 32446 2757
rect 32472 2731 32508 2757
rect 32534 2731 37074 2757
rect 37100 2731 37136 2757
rect 37162 2731 37198 2757
rect 37224 2731 37260 2757
rect 37286 2731 37322 2757
rect 37348 2731 37384 2757
rect 37410 2731 37446 2757
rect 37472 2731 37508 2757
rect 37534 2731 39312 2757
rect 672 2714 39312 2731
rect 30087 2561 30113 2567
rect 1633 2535 1639 2561
rect 1665 2535 1671 2561
rect 2473 2535 2479 2561
rect 2505 2535 2511 2561
rect 4041 2535 4047 2561
rect 4073 2535 4079 2561
rect 4993 2535 4999 2561
rect 5025 2535 5031 2561
rect 5721 2535 5727 2561
rect 5753 2535 5759 2561
rect 6449 2535 6455 2561
rect 6481 2535 6487 2561
rect 8073 2535 8079 2561
rect 8105 2535 8111 2561
rect 8969 2535 8975 2561
rect 9001 2535 9007 2561
rect 9473 2535 9479 2561
rect 9505 2535 9511 2561
rect 10425 2535 10431 2561
rect 10457 2535 10463 2561
rect 12217 2535 12223 2561
rect 12249 2535 12255 2561
rect 13169 2535 13175 2561
rect 13201 2535 13207 2561
rect 15745 2535 15751 2561
rect 15777 2535 15783 2561
rect 16753 2535 16759 2561
rect 16785 2535 16791 2561
rect 17369 2535 17375 2561
rect 17401 2535 17407 2561
rect 18265 2535 18271 2561
rect 18297 2535 18303 2561
rect 19049 2535 19055 2561
rect 19081 2535 19087 2561
rect 19945 2535 19951 2561
rect 19977 2535 19983 2561
rect 20505 2535 20511 2561
rect 20537 2535 20543 2561
rect 21345 2535 21351 2561
rect 21377 2535 21383 2561
rect 22745 2535 22751 2561
rect 22777 2535 22783 2561
rect 23865 2535 23871 2561
rect 23897 2535 23903 2561
rect 24425 2535 24431 2561
rect 24457 2535 24463 2561
rect 25377 2535 25383 2561
rect 25409 2535 25415 2561
rect 26721 2535 26727 2561
rect 26753 2535 26759 2561
rect 27673 2535 27679 2561
rect 27705 2535 27711 2561
rect 28457 2535 28463 2561
rect 28489 2535 28495 2561
rect 29353 2535 29359 2561
rect 29385 2535 29391 2561
rect 30087 2529 30113 2535
rect 30143 2561 30169 2567
rect 30143 2529 30169 2535
rect 30311 2561 30337 2567
rect 33671 2561 33697 2567
rect 30809 2535 30815 2561
rect 30841 2535 30847 2561
rect 31873 2535 31879 2561
rect 31905 2535 31911 2561
rect 32153 2535 32159 2561
rect 32185 2535 32191 2561
rect 33329 2535 33335 2561
rect 33361 2535 33367 2561
rect 30311 2529 30337 2535
rect 33671 2529 33697 2535
rect 33895 2561 33921 2567
rect 38655 2561 38681 2567
rect 34673 2535 34679 2561
rect 34705 2535 34711 2561
rect 35849 2535 35855 2561
rect 35881 2535 35887 2561
rect 36129 2535 36135 2561
rect 36161 2535 36167 2561
rect 36969 2535 36975 2561
rect 37001 2535 37007 2561
rect 33895 2529 33921 2535
rect 38655 2529 38681 2535
rect 38767 2561 38793 2567
rect 38767 2529 38793 2535
rect 33727 2505 33753 2511
rect 37591 2505 37617 2511
rect 1521 2479 1527 2505
rect 1553 2479 1559 2505
rect 4993 2479 4999 2505
rect 5025 2479 5031 2505
rect 5497 2479 5503 2505
rect 5529 2479 5535 2505
rect 8969 2479 8975 2505
rect 9001 2479 9007 2505
rect 10425 2479 10431 2505
rect 10457 2479 10463 2505
rect 13169 2479 13175 2505
rect 13201 2479 13207 2505
rect 16753 2479 16759 2505
rect 16785 2479 16791 2505
rect 18265 2479 18271 2505
rect 18297 2479 18303 2505
rect 19945 2479 19951 2505
rect 19977 2479 19983 2505
rect 21345 2479 21351 2505
rect 21377 2479 21383 2505
rect 23865 2479 23871 2505
rect 23897 2479 23903 2505
rect 25377 2479 25383 2505
rect 25409 2479 25415 2505
rect 27673 2479 27679 2505
rect 27705 2479 27711 2505
rect 29353 2479 29359 2505
rect 29385 2479 29391 2505
rect 31873 2479 31879 2505
rect 31905 2479 31911 2505
rect 33329 2479 33335 2505
rect 33361 2479 33367 2505
rect 35849 2479 35855 2505
rect 35881 2479 35887 2505
rect 37081 2479 37087 2505
rect 37113 2479 37119 2505
rect 33727 2473 33753 2479
rect 37591 2473 37617 2479
rect 37703 2505 37729 2511
rect 37703 2473 37729 2479
rect 37871 2505 37897 2511
rect 37871 2473 37897 2479
rect 38935 2505 38961 2511
rect 38935 2473 38961 2479
rect 672 2365 39312 2382
rect 672 2339 4574 2365
rect 4600 2339 4636 2365
rect 4662 2339 4698 2365
rect 4724 2339 4760 2365
rect 4786 2339 4822 2365
rect 4848 2339 4884 2365
rect 4910 2339 4946 2365
rect 4972 2339 5008 2365
rect 5034 2339 9574 2365
rect 9600 2339 9636 2365
rect 9662 2339 9698 2365
rect 9724 2339 9760 2365
rect 9786 2339 9822 2365
rect 9848 2339 9884 2365
rect 9910 2339 9946 2365
rect 9972 2339 10008 2365
rect 10034 2339 14574 2365
rect 14600 2339 14636 2365
rect 14662 2339 14698 2365
rect 14724 2339 14760 2365
rect 14786 2339 14822 2365
rect 14848 2339 14884 2365
rect 14910 2339 14946 2365
rect 14972 2339 15008 2365
rect 15034 2339 19574 2365
rect 19600 2339 19636 2365
rect 19662 2339 19698 2365
rect 19724 2339 19760 2365
rect 19786 2339 19822 2365
rect 19848 2339 19884 2365
rect 19910 2339 19946 2365
rect 19972 2339 20008 2365
rect 20034 2339 24574 2365
rect 24600 2339 24636 2365
rect 24662 2339 24698 2365
rect 24724 2339 24760 2365
rect 24786 2339 24822 2365
rect 24848 2339 24884 2365
rect 24910 2339 24946 2365
rect 24972 2339 25008 2365
rect 25034 2339 29574 2365
rect 29600 2339 29636 2365
rect 29662 2339 29698 2365
rect 29724 2339 29760 2365
rect 29786 2339 29822 2365
rect 29848 2339 29884 2365
rect 29910 2339 29946 2365
rect 29972 2339 30008 2365
rect 30034 2339 34574 2365
rect 34600 2339 34636 2365
rect 34662 2339 34698 2365
rect 34724 2339 34760 2365
rect 34786 2339 34822 2365
rect 34848 2339 34884 2365
rect 34910 2339 34946 2365
rect 34972 2339 35008 2365
rect 35034 2339 39312 2365
rect 672 2322 39312 2339
rect 28071 2225 28097 2231
rect 32159 2225 32185 2231
rect 4489 2199 4495 2225
rect 4521 2199 4527 2225
rect 5833 2199 5839 2225
rect 5865 2199 5871 2225
rect 8353 2199 8359 2225
rect 8385 2199 8391 2225
rect 10817 2199 10823 2225
rect 10849 2199 10855 2225
rect 18265 2199 18271 2225
rect 18297 2199 18303 2225
rect 19497 2199 19503 2225
rect 19529 2199 19535 2225
rect 21793 2199 21799 2225
rect 21825 2199 21831 2225
rect 23417 2199 23423 2225
rect 23449 2199 23455 2225
rect 25937 2199 25943 2225
rect 25969 2199 25975 2225
rect 27393 2199 27399 2225
rect 27425 2199 27431 2225
rect 29913 2199 29919 2225
rect 29945 2199 29951 2225
rect 31369 2199 31375 2225
rect 31401 2199 31407 2225
rect 28071 2193 28097 2199
rect 32159 2193 32185 2199
rect 32327 2225 32353 2231
rect 35743 2225 35769 2231
rect 33833 2199 33839 2225
rect 33865 2199 33871 2225
rect 35177 2199 35183 2225
rect 35209 2199 35215 2225
rect 32327 2193 32353 2199
rect 35743 2193 35769 2199
rect 35911 2225 35937 2231
rect 38151 2225 38177 2231
rect 37641 2199 37647 2225
rect 37673 2199 37679 2225
rect 35911 2193 35937 2199
rect 38151 2193 38177 2199
rect 38431 2225 38457 2231
rect 38431 2193 38457 2199
rect 38711 2225 38737 2231
rect 38711 2193 38737 2199
rect 38879 2225 38905 2231
rect 38879 2193 38905 2199
rect 28183 2169 28209 2175
rect 2361 2143 2367 2169
rect 2393 2143 2399 2169
rect 2473 2143 2479 2169
rect 2505 2143 2511 2169
rect 3033 2143 3039 2169
rect 3065 2143 3071 2169
rect 3537 2143 3543 2169
rect 3569 2143 3575 2169
rect 4433 2143 4439 2169
rect 4465 2143 4471 2169
rect 5833 2143 5839 2169
rect 5865 2143 5871 2169
rect 7009 2143 7015 2169
rect 7041 2143 7047 2169
rect 7513 2143 7519 2169
rect 7545 2143 7551 2169
rect 8353 2143 8359 2169
rect 8385 2143 8391 2169
rect 10033 2143 10039 2169
rect 10065 2143 10071 2169
rect 10817 2143 10823 2169
rect 10849 2143 10855 2169
rect 11377 2143 11383 2169
rect 11409 2143 11415 2169
rect 11769 2143 11775 2169
rect 11801 2143 11807 2169
rect 11937 2143 11943 2169
rect 11969 2143 11975 2169
rect 13785 2143 13791 2169
rect 13817 2143 13823 2169
rect 14233 2143 14239 2169
rect 14265 2143 14271 2169
rect 14457 2143 14463 2169
rect 14489 2143 14495 2169
rect 15241 2143 15247 2169
rect 15273 2143 15279 2169
rect 15689 2143 15695 2169
rect 15721 2143 15727 2169
rect 15913 2143 15919 2169
rect 15945 2143 15951 2169
rect 17369 2143 17375 2169
rect 17401 2143 17407 2169
rect 18265 2143 18271 2169
rect 18297 2143 18303 2169
rect 18825 2143 18831 2169
rect 18857 2143 18863 2169
rect 19497 2143 19503 2169
rect 19529 2143 19535 2169
rect 20785 2143 20791 2169
rect 20817 2143 20823 2169
rect 21793 2143 21799 2169
rect 21825 2143 21831 2169
rect 22241 2143 22247 2169
rect 22273 2143 22279 2169
rect 23417 2143 23423 2169
rect 23449 2143 23455 2169
rect 24761 2143 24767 2169
rect 24793 2143 24799 2169
rect 25937 2143 25943 2169
rect 25969 2143 25975 2169
rect 26217 2143 26223 2169
rect 26249 2143 26255 2169
rect 27393 2143 27399 2169
rect 27425 2143 27431 2169
rect 28183 2137 28209 2143
rect 28351 2169 28377 2175
rect 32103 2169 32129 2175
rect 35687 2169 35713 2175
rect 38319 2169 38345 2175
rect 28737 2143 28743 2169
rect 28769 2143 28775 2169
rect 29913 2143 29919 2169
rect 29945 2143 29951 2169
rect 30305 2143 30311 2169
rect 30337 2143 30343 2169
rect 31369 2143 31375 2169
rect 31401 2143 31407 2169
rect 32713 2143 32719 2169
rect 32745 2143 32751 2169
rect 33833 2143 33839 2169
rect 33865 2143 33871 2169
rect 34225 2143 34231 2169
rect 34257 2143 34263 2169
rect 35177 2143 35183 2169
rect 35209 2143 35215 2169
rect 36689 2143 36695 2169
rect 36721 2143 36727 2169
rect 37641 2143 37647 2169
rect 37673 2143 37679 2169
rect 28351 2137 28377 2143
rect 32103 2137 32129 2143
rect 35687 2137 35713 2143
rect 38319 2137 38345 2143
rect 38935 2169 38961 2175
rect 38935 2137 38961 2143
rect 672 1973 39312 1990
rect 672 1947 2074 1973
rect 2100 1947 2136 1973
rect 2162 1947 2198 1973
rect 2224 1947 2260 1973
rect 2286 1947 2322 1973
rect 2348 1947 2384 1973
rect 2410 1947 2446 1973
rect 2472 1947 2508 1973
rect 2534 1947 7074 1973
rect 7100 1947 7136 1973
rect 7162 1947 7198 1973
rect 7224 1947 7260 1973
rect 7286 1947 7322 1973
rect 7348 1947 7384 1973
rect 7410 1947 7446 1973
rect 7472 1947 7508 1973
rect 7534 1947 12074 1973
rect 12100 1947 12136 1973
rect 12162 1947 12198 1973
rect 12224 1947 12260 1973
rect 12286 1947 12322 1973
rect 12348 1947 12384 1973
rect 12410 1947 12446 1973
rect 12472 1947 12508 1973
rect 12534 1947 17074 1973
rect 17100 1947 17136 1973
rect 17162 1947 17198 1973
rect 17224 1947 17260 1973
rect 17286 1947 17322 1973
rect 17348 1947 17384 1973
rect 17410 1947 17446 1973
rect 17472 1947 17508 1973
rect 17534 1947 22074 1973
rect 22100 1947 22136 1973
rect 22162 1947 22198 1973
rect 22224 1947 22260 1973
rect 22286 1947 22322 1973
rect 22348 1947 22384 1973
rect 22410 1947 22446 1973
rect 22472 1947 22508 1973
rect 22534 1947 27074 1973
rect 27100 1947 27136 1973
rect 27162 1947 27198 1973
rect 27224 1947 27260 1973
rect 27286 1947 27322 1973
rect 27348 1947 27384 1973
rect 27410 1947 27446 1973
rect 27472 1947 27508 1973
rect 27534 1947 32074 1973
rect 32100 1947 32136 1973
rect 32162 1947 32198 1973
rect 32224 1947 32260 1973
rect 32286 1947 32322 1973
rect 32348 1947 32384 1973
rect 32410 1947 32446 1973
rect 32472 1947 32508 1973
rect 32534 1947 37074 1973
rect 37100 1947 37136 1973
rect 37162 1947 37198 1973
rect 37224 1947 37260 1973
rect 37286 1947 37322 1973
rect 37348 1947 37384 1973
rect 37410 1947 37446 1973
rect 37472 1947 37508 1973
rect 37534 1947 39312 1973
rect 672 1930 39312 1947
rect 38151 1777 38177 1783
rect 1185 1751 1191 1777
rect 1217 1751 1223 1777
rect 1913 1751 1919 1777
rect 1945 1751 1951 1777
rect 3537 1751 3543 1777
rect 3569 1751 3575 1777
rect 4433 1751 4439 1777
rect 4465 1751 4471 1777
rect 5497 1751 5503 1777
rect 5529 1751 5535 1777
rect 6393 1751 6399 1777
rect 6425 1751 6431 1777
rect 7457 1751 7463 1777
rect 7489 1751 7495 1777
rect 8353 1751 8359 1777
rect 8385 1751 8391 1777
rect 9361 1751 9367 1777
rect 9393 1751 9399 1777
rect 9697 1751 9703 1777
rect 9729 1751 9735 1777
rect 9809 1751 9815 1777
rect 9841 1751 9847 1777
rect 11377 1751 11383 1777
rect 11409 1751 11415 1777
rect 11657 1751 11663 1777
rect 11689 1751 11695 1777
rect 11769 1751 11775 1777
rect 11801 1751 11807 1777
rect 13057 1751 13063 1777
rect 13089 1751 13095 1777
rect 13505 1751 13511 1777
rect 13537 1751 13543 1777
rect 13729 1751 13735 1777
rect 13761 1751 13767 1777
rect 15241 1751 15247 1777
rect 15273 1751 15279 1777
rect 15577 1751 15583 1777
rect 15609 1751 15615 1777
rect 15689 1751 15695 1777
rect 15721 1751 15727 1777
rect 17257 1751 17263 1777
rect 17289 1751 17295 1777
rect 18153 1751 18159 1777
rect 18185 1751 18191 1777
rect 18825 1751 18831 1777
rect 18857 1751 18863 1777
rect 19497 1751 19503 1777
rect 19529 1751 19535 1777
rect 20505 1751 20511 1777
rect 20537 1751 20543 1777
rect 21681 1751 21687 1777
rect 21713 1751 21719 1777
rect 22465 1751 22471 1777
rect 22497 1751 22503 1777
rect 23641 1751 23647 1777
rect 23673 1751 23679 1777
rect 24425 1751 24431 1777
rect 24457 1751 24463 1777
rect 25601 1751 25607 1777
rect 25633 1751 25639 1777
rect 26385 1751 26391 1777
rect 26417 1751 26423 1777
rect 27561 1751 27567 1777
rect 27593 1751 27599 1777
rect 28513 1751 28519 1777
rect 28545 1751 28551 1777
rect 29353 1751 29359 1777
rect 29385 1751 29391 1777
rect 30305 1751 30311 1777
rect 30337 1751 30343 1777
rect 31481 1751 31487 1777
rect 31513 1751 31519 1777
rect 32545 1751 32551 1777
rect 32577 1751 32583 1777
rect 33441 1751 33447 1777
rect 33473 1751 33479 1777
rect 34225 1751 34231 1777
rect 34257 1751 34263 1777
rect 35177 1751 35183 1777
rect 35209 1751 35215 1777
rect 36185 1751 36191 1777
rect 36217 1751 36223 1777
rect 36969 1751 36975 1777
rect 37001 1751 37007 1777
rect 38151 1745 38177 1751
rect 38263 1777 38289 1783
rect 38263 1745 38289 1751
rect 38431 1777 38457 1783
rect 38431 1745 38457 1751
rect 38655 1777 38681 1783
rect 38655 1745 38681 1751
rect 38823 1777 38849 1783
rect 38823 1745 38849 1751
rect 38935 1777 38961 1783
rect 38935 1745 38961 1751
rect 1913 1695 1919 1721
rect 1945 1695 1951 1721
rect 4433 1695 4439 1721
rect 4465 1695 4471 1721
rect 6393 1695 6399 1721
rect 6425 1695 6431 1721
rect 8353 1695 8359 1721
rect 8385 1695 8391 1721
rect 18153 1695 18159 1721
rect 18185 1695 18191 1721
rect 19497 1695 19503 1721
rect 19529 1695 19535 1721
rect 21681 1695 21687 1721
rect 21713 1695 21719 1721
rect 23641 1695 23647 1721
rect 23673 1695 23679 1721
rect 25601 1695 25607 1721
rect 25633 1695 25639 1721
rect 27561 1695 27567 1721
rect 27593 1695 27599 1721
rect 29353 1695 29359 1721
rect 29385 1695 29391 1721
rect 31481 1695 31487 1721
rect 31513 1695 31519 1721
rect 33441 1695 33447 1721
rect 33473 1695 33479 1721
rect 35177 1695 35183 1721
rect 35209 1695 35215 1721
rect 37137 1695 37143 1721
rect 37169 1695 37175 1721
rect 672 1581 39312 1598
rect 672 1555 4574 1581
rect 4600 1555 4636 1581
rect 4662 1555 4698 1581
rect 4724 1555 4760 1581
rect 4786 1555 4822 1581
rect 4848 1555 4884 1581
rect 4910 1555 4946 1581
rect 4972 1555 5008 1581
rect 5034 1555 9574 1581
rect 9600 1555 9636 1581
rect 9662 1555 9698 1581
rect 9724 1555 9760 1581
rect 9786 1555 9822 1581
rect 9848 1555 9884 1581
rect 9910 1555 9946 1581
rect 9972 1555 10008 1581
rect 10034 1555 14574 1581
rect 14600 1555 14636 1581
rect 14662 1555 14698 1581
rect 14724 1555 14760 1581
rect 14786 1555 14822 1581
rect 14848 1555 14884 1581
rect 14910 1555 14946 1581
rect 14972 1555 15008 1581
rect 15034 1555 19574 1581
rect 19600 1555 19636 1581
rect 19662 1555 19698 1581
rect 19724 1555 19760 1581
rect 19786 1555 19822 1581
rect 19848 1555 19884 1581
rect 19910 1555 19946 1581
rect 19972 1555 20008 1581
rect 20034 1555 24574 1581
rect 24600 1555 24636 1581
rect 24662 1555 24698 1581
rect 24724 1555 24760 1581
rect 24786 1555 24822 1581
rect 24848 1555 24884 1581
rect 24910 1555 24946 1581
rect 24972 1555 25008 1581
rect 25034 1555 29574 1581
rect 29600 1555 29636 1581
rect 29662 1555 29698 1581
rect 29724 1555 29760 1581
rect 29786 1555 29822 1581
rect 29848 1555 29884 1581
rect 29910 1555 29946 1581
rect 29972 1555 30008 1581
rect 30034 1555 34574 1581
rect 34600 1555 34636 1581
rect 34662 1555 34698 1581
rect 34724 1555 34760 1581
rect 34786 1555 34822 1581
rect 34848 1555 34884 1581
rect 34910 1555 34946 1581
rect 34972 1555 35008 1581
rect 35034 1555 39312 1581
rect 672 1538 39312 1555
<< via1 >>
rect 2074 18411 2100 18437
rect 2136 18411 2162 18437
rect 2198 18411 2224 18437
rect 2260 18411 2286 18437
rect 2322 18411 2348 18437
rect 2384 18411 2410 18437
rect 2446 18411 2472 18437
rect 2508 18411 2534 18437
rect 7074 18411 7100 18437
rect 7136 18411 7162 18437
rect 7198 18411 7224 18437
rect 7260 18411 7286 18437
rect 7322 18411 7348 18437
rect 7384 18411 7410 18437
rect 7446 18411 7472 18437
rect 7508 18411 7534 18437
rect 12074 18411 12100 18437
rect 12136 18411 12162 18437
rect 12198 18411 12224 18437
rect 12260 18411 12286 18437
rect 12322 18411 12348 18437
rect 12384 18411 12410 18437
rect 12446 18411 12472 18437
rect 12508 18411 12534 18437
rect 17074 18411 17100 18437
rect 17136 18411 17162 18437
rect 17198 18411 17224 18437
rect 17260 18411 17286 18437
rect 17322 18411 17348 18437
rect 17384 18411 17410 18437
rect 17446 18411 17472 18437
rect 17508 18411 17534 18437
rect 22074 18411 22100 18437
rect 22136 18411 22162 18437
rect 22198 18411 22224 18437
rect 22260 18411 22286 18437
rect 22322 18411 22348 18437
rect 22384 18411 22410 18437
rect 22446 18411 22472 18437
rect 22508 18411 22534 18437
rect 27074 18411 27100 18437
rect 27136 18411 27162 18437
rect 27198 18411 27224 18437
rect 27260 18411 27286 18437
rect 27322 18411 27348 18437
rect 27384 18411 27410 18437
rect 27446 18411 27472 18437
rect 27508 18411 27534 18437
rect 32074 18411 32100 18437
rect 32136 18411 32162 18437
rect 32198 18411 32224 18437
rect 32260 18411 32286 18437
rect 32322 18411 32348 18437
rect 32384 18411 32410 18437
rect 32446 18411 32472 18437
rect 32508 18411 32534 18437
rect 37074 18411 37100 18437
rect 37136 18411 37162 18437
rect 37198 18411 37224 18437
rect 37260 18411 37286 18437
rect 37322 18411 37348 18437
rect 37384 18411 37410 18437
rect 37446 18411 37472 18437
rect 37508 18411 37534 18437
rect 4574 18019 4600 18045
rect 4636 18019 4662 18045
rect 4698 18019 4724 18045
rect 4760 18019 4786 18045
rect 4822 18019 4848 18045
rect 4884 18019 4910 18045
rect 4946 18019 4972 18045
rect 5008 18019 5034 18045
rect 9574 18019 9600 18045
rect 9636 18019 9662 18045
rect 9698 18019 9724 18045
rect 9760 18019 9786 18045
rect 9822 18019 9848 18045
rect 9884 18019 9910 18045
rect 9946 18019 9972 18045
rect 10008 18019 10034 18045
rect 14574 18019 14600 18045
rect 14636 18019 14662 18045
rect 14698 18019 14724 18045
rect 14760 18019 14786 18045
rect 14822 18019 14848 18045
rect 14884 18019 14910 18045
rect 14946 18019 14972 18045
rect 15008 18019 15034 18045
rect 19574 18019 19600 18045
rect 19636 18019 19662 18045
rect 19698 18019 19724 18045
rect 19760 18019 19786 18045
rect 19822 18019 19848 18045
rect 19884 18019 19910 18045
rect 19946 18019 19972 18045
rect 20008 18019 20034 18045
rect 24574 18019 24600 18045
rect 24636 18019 24662 18045
rect 24698 18019 24724 18045
rect 24760 18019 24786 18045
rect 24822 18019 24848 18045
rect 24884 18019 24910 18045
rect 24946 18019 24972 18045
rect 25008 18019 25034 18045
rect 29574 18019 29600 18045
rect 29636 18019 29662 18045
rect 29698 18019 29724 18045
rect 29760 18019 29786 18045
rect 29822 18019 29848 18045
rect 29884 18019 29910 18045
rect 29946 18019 29972 18045
rect 30008 18019 30034 18045
rect 34574 18019 34600 18045
rect 34636 18019 34662 18045
rect 34698 18019 34724 18045
rect 34760 18019 34786 18045
rect 34822 18019 34848 18045
rect 34884 18019 34910 18045
rect 34946 18019 34972 18045
rect 35008 18019 35034 18045
rect 2074 17627 2100 17653
rect 2136 17627 2162 17653
rect 2198 17627 2224 17653
rect 2260 17627 2286 17653
rect 2322 17627 2348 17653
rect 2384 17627 2410 17653
rect 2446 17627 2472 17653
rect 2508 17627 2534 17653
rect 7074 17627 7100 17653
rect 7136 17627 7162 17653
rect 7198 17627 7224 17653
rect 7260 17627 7286 17653
rect 7322 17627 7348 17653
rect 7384 17627 7410 17653
rect 7446 17627 7472 17653
rect 7508 17627 7534 17653
rect 12074 17627 12100 17653
rect 12136 17627 12162 17653
rect 12198 17627 12224 17653
rect 12260 17627 12286 17653
rect 12322 17627 12348 17653
rect 12384 17627 12410 17653
rect 12446 17627 12472 17653
rect 12508 17627 12534 17653
rect 17074 17627 17100 17653
rect 17136 17627 17162 17653
rect 17198 17627 17224 17653
rect 17260 17627 17286 17653
rect 17322 17627 17348 17653
rect 17384 17627 17410 17653
rect 17446 17627 17472 17653
rect 17508 17627 17534 17653
rect 22074 17627 22100 17653
rect 22136 17627 22162 17653
rect 22198 17627 22224 17653
rect 22260 17627 22286 17653
rect 22322 17627 22348 17653
rect 22384 17627 22410 17653
rect 22446 17627 22472 17653
rect 22508 17627 22534 17653
rect 27074 17627 27100 17653
rect 27136 17627 27162 17653
rect 27198 17627 27224 17653
rect 27260 17627 27286 17653
rect 27322 17627 27348 17653
rect 27384 17627 27410 17653
rect 27446 17627 27472 17653
rect 27508 17627 27534 17653
rect 32074 17627 32100 17653
rect 32136 17627 32162 17653
rect 32198 17627 32224 17653
rect 32260 17627 32286 17653
rect 32322 17627 32348 17653
rect 32384 17627 32410 17653
rect 32446 17627 32472 17653
rect 32508 17627 32534 17653
rect 37074 17627 37100 17653
rect 37136 17627 37162 17653
rect 37198 17627 37224 17653
rect 37260 17627 37286 17653
rect 37322 17627 37348 17653
rect 37384 17627 37410 17653
rect 37446 17627 37472 17653
rect 37508 17627 37534 17653
rect 12503 17431 12529 17457
rect 13287 17431 13313 17457
rect 13287 17375 13313 17401
rect 4574 17235 4600 17261
rect 4636 17235 4662 17261
rect 4698 17235 4724 17261
rect 4760 17235 4786 17261
rect 4822 17235 4848 17261
rect 4884 17235 4910 17261
rect 4946 17235 4972 17261
rect 5008 17235 5034 17261
rect 9574 17235 9600 17261
rect 9636 17235 9662 17261
rect 9698 17235 9724 17261
rect 9760 17235 9786 17261
rect 9822 17235 9848 17261
rect 9884 17235 9910 17261
rect 9946 17235 9972 17261
rect 10008 17235 10034 17261
rect 14574 17235 14600 17261
rect 14636 17235 14662 17261
rect 14698 17235 14724 17261
rect 14760 17235 14786 17261
rect 14822 17235 14848 17261
rect 14884 17235 14910 17261
rect 14946 17235 14972 17261
rect 15008 17235 15034 17261
rect 19574 17235 19600 17261
rect 19636 17235 19662 17261
rect 19698 17235 19724 17261
rect 19760 17235 19786 17261
rect 19822 17235 19848 17261
rect 19884 17235 19910 17261
rect 19946 17235 19972 17261
rect 20008 17235 20034 17261
rect 24574 17235 24600 17261
rect 24636 17235 24662 17261
rect 24698 17235 24724 17261
rect 24760 17235 24786 17261
rect 24822 17235 24848 17261
rect 24884 17235 24910 17261
rect 24946 17235 24972 17261
rect 25008 17235 25034 17261
rect 29574 17235 29600 17261
rect 29636 17235 29662 17261
rect 29698 17235 29724 17261
rect 29760 17235 29786 17261
rect 29822 17235 29848 17261
rect 29884 17235 29910 17261
rect 29946 17235 29972 17261
rect 30008 17235 30034 17261
rect 34574 17235 34600 17261
rect 34636 17235 34662 17261
rect 34698 17235 34724 17261
rect 34760 17235 34786 17261
rect 34822 17235 34848 17261
rect 34884 17235 34910 17261
rect 34946 17235 34972 17261
rect 35008 17235 35034 17261
rect 10599 17095 10625 17121
rect 12055 17095 12081 17121
rect 9647 17039 9673 17065
rect 10431 17039 10457 17065
rect 11103 17039 11129 17065
rect 11999 17039 12025 17065
rect 12839 17039 12865 17065
rect 13287 17039 13313 17065
rect 13511 17039 13537 17065
rect 2074 16843 2100 16869
rect 2136 16843 2162 16869
rect 2198 16843 2224 16869
rect 2260 16843 2286 16869
rect 2322 16843 2348 16869
rect 2384 16843 2410 16869
rect 2446 16843 2472 16869
rect 2508 16843 2534 16869
rect 7074 16843 7100 16869
rect 7136 16843 7162 16869
rect 7198 16843 7224 16869
rect 7260 16843 7286 16869
rect 7322 16843 7348 16869
rect 7384 16843 7410 16869
rect 7446 16843 7472 16869
rect 7508 16843 7534 16869
rect 12074 16843 12100 16869
rect 12136 16843 12162 16869
rect 12198 16843 12224 16869
rect 12260 16843 12286 16869
rect 12322 16843 12348 16869
rect 12384 16843 12410 16869
rect 12446 16843 12472 16869
rect 12508 16843 12534 16869
rect 17074 16843 17100 16869
rect 17136 16843 17162 16869
rect 17198 16843 17224 16869
rect 17260 16843 17286 16869
rect 17322 16843 17348 16869
rect 17384 16843 17410 16869
rect 17446 16843 17472 16869
rect 17508 16843 17534 16869
rect 22074 16843 22100 16869
rect 22136 16843 22162 16869
rect 22198 16843 22224 16869
rect 22260 16843 22286 16869
rect 22322 16843 22348 16869
rect 22384 16843 22410 16869
rect 22446 16843 22472 16869
rect 22508 16843 22534 16869
rect 27074 16843 27100 16869
rect 27136 16843 27162 16869
rect 27198 16843 27224 16869
rect 27260 16843 27286 16869
rect 27322 16843 27348 16869
rect 27384 16843 27410 16869
rect 27446 16843 27472 16869
rect 27508 16843 27534 16869
rect 32074 16843 32100 16869
rect 32136 16843 32162 16869
rect 32198 16843 32224 16869
rect 32260 16843 32286 16869
rect 32322 16843 32348 16869
rect 32384 16843 32410 16869
rect 32446 16843 32472 16869
rect 32508 16843 32534 16869
rect 37074 16843 37100 16869
rect 37136 16843 37162 16869
rect 37198 16843 37224 16869
rect 37260 16843 37286 16869
rect 37322 16843 37348 16869
rect 37384 16843 37410 16869
rect 37446 16843 37472 16869
rect 37508 16843 37534 16869
rect 9535 16647 9561 16673
rect 10431 16647 10457 16673
rect 10935 16647 10961 16673
rect 11383 16647 11409 16673
rect 11495 16647 11521 16673
rect 12559 16647 12585 16673
rect 13455 16647 13481 16673
rect 10431 16591 10457 16617
rect 13455 16591 13481 16617
rect 4574 16451 4600 16477
rect 4636 16451 4662 16477
rect 4698 16451 4724 16477
rect 4760 16451 4786 16477
rect 4822 16451 4848 16477
rect 4884 16451 4910 16477
rect 4946 16451 4972 16477
rect 5008 16451 5034 16477
rect 9574 16451 9600 16477
rect 9636 16451 9662 16477
rect 9698 16451 9724 16477
rect 9760 16451 9786 16477
rect 9822 16451 9848 16477
rect 9884 16451 9910 16477
rect 9946 16451 9972 16477
rect 10008 16451 10034 16477
rect 14574 16451 14600 16477
rect 14636 16451 14662 16477
rect 14698 16451 14724 16477
rect 14760 16451 14786 16477
rect 14822 16451 14848 16477
rect 14884 16451 14910 16477
rect 14946 16451 14972 16477
rect 15008 16451 15034 16477
rect 19574 16451 19600 16477
rect 19636 16451 19662 16477
rect 19698 16451 19724 16477
rect 19760 16451 19786 16477
rect 19822 16451 19848 16477
rect 19884 16451 19910 16477
rect 19946 16451 19972 16477
rect 20008 16451 20034 16477
rect 24574 16451 24600 16477
rect 24636 16451 24662 16477
rect 24698 16451 24724 16477
rect 24760 16451 24786 16477
rect 24822 16451 24848 16477
rect 24884 16451 24910 16477
rect 24946 16451 24972 16477
rect 25008 16451 25034 16477
rect 29574 16451 29600 16477
rect 29636 16451 29662 16477
rect 29698 16451 29724 16477
rect 29760 16451 29786 16477
rect 29822 16451 29848 16477
rect 29884 16451 29910 16477
rect 29946 16451 29972 16477
rect 30008 16451 30034 16477
rect 34574 16451 34600 16477
rect 34636 16451 34662 16477
rect 34698 16451 34724 16477
rect 34760 16451 34786 16477
rect 34822 16451 34848 16477
rect 34884 16451 34910 16477
rect 34946 16451 34972 16477
rect 35008 16451 35034 16477
rect 7015 16311 7041 16337
rect 8359 16311 8385 16337
rect 10823 16311 10849 16337
rect 12335 16311 12361 16337
rect 13791 16311 13817 16337
rect 15471 16311 15497 16337
rect 6119 16255 6145 16281
rect 7015 16255 7041 16281
rect 7519 16255 7545 16281
rect 8359 16255 8385 16281
rect 9983 16255 10009 16281
rect 10823 16255 10849 16281
rect 11159 16255 11185 16281
rect 12335 16255 12361 16281
rect 12839 16255 12865 16281
rect 13791 16255 13817 16281
rect 14295 16255 14321 16281
rect 15471 16255 15497 16281
rect 2074 16059 2100 16085
rect 2136 16059 2162 16085
rect 2198 16059 2224 16085
rect 2260 16059 2286 16085
rect 2322 16059 2348 16085
rect 2384 16059 2410 16085
rect 2446 16059 2472 16085
rect 2508 16059 2534 16085
rect 7074 16059 7100 16085
rect 7136 16059 7162 16085
rect 7198 16059 7224 16085
rect 7260 16059 7286 16085
rect 7322 16059 7348 16085
rect 7384 16059 7410 16085
rect 7446 16059 7472 16085
rect 7508 16059 7534 16085
rect 12074 16059 12100 16085
rect 12136 16059 12162 16085
rect 12198 16059 12224 16085
rect 12260 16059 12286 16085
rect 12322 16059 12348 16085
rect 12384 16059 12410 16085
rect 12446 16059 12472 16085
rect 12508 16059 12534 16085
rect 17074 16059 17100 16085
rect 17136 16059 17162 16085
rect 17198 16059 17224 16085
rect 17260 16059 17286 16085
rect 17322 16059 17348 16085
rect 17384 16059 17410 16085
rect 17446 16059 17472 16085
rect 17508 16059 17534 16085
rect 22074 16059 22100 16085
rect 22136 16059 22162 16085
rect 22198 16059 22224 16085
rect 22260 16059 22286 16085
rect 22322 16059 22348 16085
rect 22384 16059 22410 16085
rect 22446 16059 22472 16085
rect 22508 16059 22534 16085
rect 27074 16059 27100 16085
rect 27136 16059 27162 16085
rect 27198 16059 27224 16085
rect 27260 16059 27286 16085
rect 27322 16059 27348 16085
rect 27384 16059 27410 16085
rect 27446 16059 27472 16085
rect 27508 16059 27534 16085
rect 32074 16059 32100 16085
rect 32136 16059 32162 16085
rect 32198 16059 32224 16085
rect 32260 16059 32286 16085
rect 32322 16059 32348 16085
rect 32384 16059 32410 16085
rect 32446 16059 32472 16085
rect 32508 16059 32534 16085
rect 37074 16059 37100 16085
rect 37136 16059 37162 16085
rect 37198 16059 37224 16085
rect 37260 16059 37286 16085
rect 37322 16059 37348 16085
rect 37384 16059 37410 16085
rect 37446 16059 37472 16085
rect 37508 16059 37534 16085
rect 5279 15863 5305 15889
rect 6455 15863 6481 15889
rect 7799 15863 7825 15889
rect 8359 15863 8385 15889
rect 8471 15863 8497 15889
rect 9255 15863 9281 15889
rect 10151 15863 10177 15889
rect 11663 15863 11689 15889
rect 12839 15863 12865 15889
rect 13119 15863 13145 15889
rect 14015 15863 14041 15889
rect 15079 15863 15105 15889
rect 15527 15863 15553 15889
rect 16479 15863 16505 15889
rect 16815 15863 16841 15889
rect 16927 15863 16953 15889
rect 6455 15807 6481 15833
rect 10207 15807 10233 15833
rect 12839 15807 12865 15833
rect 14071 15807 14097 15833
rect 15751 15807 15777 15833
rect 4574 15667 4600 15693
rect 4636 15667 4662 15693
rect 4698 15667 4724 15693
rect 4760 15667 4786 15693
rect 4822 15667 4848 15693
rect 4884 15667 4910 15693
rect 4946 15667 4972 15693
rect 5008 15667 5034 15693
rect 9574 15667 9600 15693
rect 9636 15667 9662 15693
rect 9698 15667 9724 15693
rect 9760 15667 9786 15693
rect 9822 15667 9848 15693
rect 9884 15667 9910 15693
rect 9946 15667 9972 15693
rect 10008 15667 10034 15693
rect 14574 15667 14600 15693
rect 14636 15667 14662 15693
rect 14698 15667 14724 15693
rect 14760 15667 14786 15693
rect 14822 15667 14848 15693
rect 14884 15667 14910 15693
rect 14946 15667 14972 15693
rect 15008 15667 15034 15693
rect 19574 15667 19600 15693
rect 19636 15667 19662 15693
rect 19698 15667 19724 15693
rect 19760 15667 19786 15693
rect 19822 15667 19848 15693
rect 19884 15667 19910 15693
rect 19946 15667 19972 15693
rect 20008 15667 20034 15693
rect 24574 15667 24600 15693
rect 24636 15667 24662 15693
rect 24698 15667 24724 15693
rect 24760 15667 24786 15693
rect 24822 15667 24848 15693
rect 24884 15667 24910 15693
rect 24946 15667 24972 15693
rect 25008 15667 25034 15693
rect 29574 15667 29600 15693
rect 29636 15667 29662 15693
rect 29698 15667 29724 15693
rect 29760 15667 29786 15693
rect 29822 15667 29848 15693
rect 29884 15667 29910 15693
rect 29946 15667 29972 15693
rect 30008 15667 30034 15693
rect 34574 15667 34600 15693
rect 34636 15667 34662 15693
rect 34698 15667 34724 15693
rect 34760 15667 34786 15693
rect 34822 15667 34848 15693
rect 34884 15667 34910 15693
rect 34946 15667 34972 15693
rect 35008 15667 35034 15693
rect 6903 15527 6929 15553
rect 8359 15527 8385 15553
rect 10879 15527 10905 15553
rect 12447 15527 12473 15553
rect 14015 15527 14041 15553
rect 15359 15527 15385 15553
rect 5839 15471 5865 15497
rect 6903 15471 6929 15497
rect 7295 15471 7321 15497
rect 8359 15471 8385 15497
rect 9815 15471 9841 15497
rect 10879 15471 10905 15497
rect 11551 15471 11577 15497
rect 12447 15471 12473 15497
rect 13119 15471 13145 15497
rect 14015 15471 14041 15497
rect 14295 15471 14321 15497
rect 15359 15471 15385 15497
rect 2074 15275 2100 15301
rect 2136 15275 2162 15301
rect 2198 15275 2224 15301
rect 2260 15275 2286 15301
rect 2322 15275 2348 15301
rect 2384 15275 2410 15301
rect 2446 15275 2472 15301
rect 2508 15275 2534 15301
rect 7074 15275 7100 15301
rect 7136 15275 7162 15301
rect 7198 15275 7224 15301
rect 7260 15275 7286 15301
rect 7322 15275 7348 15301
rect 7384 15275 7410 15301
rect 7446 15275 7472 15301
rect 7508 15275 7534 15301
rect 12074 15275 12100 15301
rect 12136 15275 12162 15301
rect 12198 15275 12224 15301
rect 12260 15275 12286 15301
rect 12322 15275 12348 15301
rect 12384 15275 12410 15301
rect 12446 15275 12472 15301
rect 12508 15275 12534 15301
rect 17074 15275 17100 15301
rect 17136 15275 17162 15301
rect 17198 15275 17224 15301
rect 17260 15275 17286 15301
rect 17322 15275 17348 15301
rect 17384 15275 17410 15301
rect 17446 15275 17472 15301
rect 17508 15275 17534 15301
rect 22074 15275 22100 15301
rect 22136 15275 22162 15301
rect 22198 15275 22224 15301
rect 22260 15275 22286 15301
rect 22322 15275 22348 15301
rect 22384 15275 22410 15301
rect 22446 15275 22472 15301
rect 22508 15275 22534 15301
rect 27074 15275 27100 15301
rect 27136 15275 27162 15301
rect 27198 15275 27224 15301
rect 27260 15275 27286 15301
rect 27322 15275 27348 15301
rect 27384 15275 27410 15301
rect 27446 15275 27472 15301
rect 27508 15275 27534 15301
rect 32074 15275 32100 15301
rect 32136 15275 32162 15301
rect 32198 15275 32224 15301
rect 32260 15275 32286 15301
rect 32322 15275 32348 15301
rect 32384 15275 32410 15301
rect 32446 15275 32472 15301
rect 32508 15275 32534 15301
rect 37074 15275 37100 15301
rect 37136 15275 37162 15301
rect 37198 15275 37224 15301
rect 37260 15275 37286 15301
rect 37322 15275 37348 15301
rect 37384 15275 37410 15301
rect 37446 15275 37472 15301
rect 37508 15275 37534 15301
rect 1807 15079 1833 15105
rect 1919 15079 1945 15105
rect 2423 15079 2449 15105
rect 3823 15079 3849 15105
rect 4383 15079 4409 15105
rect 4495 15079 4521 15105
rect 5279 15079 5305 15105
rect 6399 15079 6425 15105
rect 7799 15079 7825 15105
rect 8975 15079 9001 15105
rect 9255 15079 9281 15105
rect 10431 15079 10457 15105
rect 11943 15079 11969 15105
rect 12839 15079 12865 15105
rect 13119 15079 13145 15105
rect 14015 15079 14041 15105
rect 14799 15079 14825 15105
rect 15359 15079 15385 15105
rect 15527 15079 15553 15105
rect 16479 15079 16505 15105
rect 17431 15079 17457 15105
rect 18775 15079 18801 15105
rect 19335 15079 19361 15105
rect 19447 15079 19473 15105
rect 6399 15023 6425 15049
rect 8975 15023 9001 15049
rect 10431 15023 10457 15049
rect 12839 15023 12865 15049
rect 14071 15023 14097 15049
rect 17431 15023 17457 15049
rect 4574 14883 4600 14909
rect 4636 14883 4662 14909
rect 4698 14883 4724 14909
rect 4760 14883 4786 14909
rect 4822 14883 4848 14909
rect 4884 14883 4910 14909
rect 4946 14883 4972 14909
rect 5008 14883 5034 14909
rect 9574 14883 9600 14909
rect 9636 14883 9662 14909
rect 9698 14883 9724 14909
rect 9760 14883 9786 14909
rect 9822 14883 9848 14909
rect 9884 14883 9910 14909
rect 9946 14883 9972 14909
rect 10008 14883 10034 14909
rect 14574 14883 14600 14909
rect 14636 14883 14662 14909
rect 14698 14883 14724 14909
rect 14760 14883 14786 14909
rect 14822 14883 14848 14909
rect 14884 14883 14910 14909
rect 14946 14883 14972 14909
rect 15008 14883 15034 14909
rect 19574 14883 19600 14909
rect 19636 14883 19662 14909
rect 19698 14883 19724 14909
rect 19760 14883 19786 14909
rect 19822 14883 19848 14909
rect 19884 14883 19910 14909
rect 19946 14883 19972 14909
rect 20008 14883 20034 14909
rect 24574 14883 24600 14909
rect 24636 14883 24662 14909
rect 24698 14883 24724 14909
rect 24760 14883 24786 14909
rect 24822 14883 24848 14909
rect 24884 14883 24910 14909
rect 24946 14883 24972 14909
rect 25008 14883 25034 14909
rect 29574 14883 29600 14909
rect 29636 14883 29662 14909
rect 29698 14883 29724 14909
rect 29760 14883 29786 14909
rect 29822 14883 29848 14909
rect 29884 14883 29910 14909
rect 29946 14883 29972 14909
rect 30008 14883 30034 14909
rect 34574 14883 34600 14909
rect 34636 14883 34662 14909
rect 34698 14883 34724 14909
rect 34760 14883 34786 14909
rect 34822 14883 34848 14909
rect 34884 14883 34910 14909
rect 34946 14883 34972 14909
rect 35008 14883 35034 14909
rect 1863 14743 1889 14769
rect 4495 14743 4521 14769
rect 6903 14743 6929 14769
rect 8359 14743 8385 14769
rect 10879 14743 10905 14769
rect 12447 14743 12473 14769
rect 14015 14743 14041 14769
rect 15303 14743 15329 14769
rect 17767 14743 17793 14769
rect 1863 14687 1889 14713
rect 3039 14687 3065 14713
rect 3599 14687 3625 14713
rect 4495 14687 4521 14713
rect 5839 14687 5865 14713
rect 6903 14687 6929 14713
rect 7295 14687 7321 14713
rect 8359 14687 8385 14713
rect 9815 14687 9841 14713
rect 10879 14687 10905 14713
rect 11551 14687 11577 14713
rect 12447 14687 12473 14713
rect 13119 14687 13145 14713
rect 14015 14687 14041 14713
rect 14351 14687 14377 14713
rect 15303 14687 15329 14713
rect 17095 14687 17121 14713
rect 17767 14687 17793 14713
rect 18271 14687 18297 14713
rect 18719 14687 18745 14713
rect 18943 14687 18969 14713
rect 2074 14491 2100 14517
rect 2136 14491 2162 14517
rect 2198 14491 2224 14517
rect 2260 14491 2286 14517
rect 2322 14491 2348 14517
rect 2384 14491 2410 14517
rect 2446 14491 2472 14517
rect 2508 14491 2534 14517
rect 7074 14491 7100 14517
rect 7136 14491 7162 14517
rect 7198 14491 7224 14517
rect 7260 14491 7286 14517
rect 7322 14491 7348 14517
rect 7384 14491 7410 14517
rect 7446 14491 7472 14517
rect 7508 14491 7534 14517
rect 12074 14491 12100 14517
rect 12136 14491 12162 14517
rect 12198 14491 12224 14517
rect 12260 14491 12286 14517
rect 12322 14491 12348 14517
rect 12384 14491 12410 14517
rect 12446 14491 12472 14517
rect 12508 14491 12534 14517
rect 17074 14491 17100 14517
rect 17136 14491 17162 14517
rect 17198 14491 17224 14517
rect 17260 14491 17286 14517
rect 17322 14491 17348 14517
rect 17384 14491 17410 14517
rect 17446 14491 17472 14517
rect 17508 14491 17534 14517
rect 22074 14491 22100 14517
rect 22136 14491 22162 14517
rect 22198 14491 22224 14517
rect 22260 14491 22286 14517
rect 22322 14491 22348 14517
rect 22384 14491 22410 14517
rect 22446 14491 22472 14517
rect 22508 14491 22534 14517
rect 27074 14491 27100 14517
rect 27136 14491 27162 14517
rect 27198 14491 27224 14517
rect 27260 14491 27286 14517
rect 27322 14491 27348 14517
rect 27384 14491 27410 14517
rect 27446 14491 27472 14517
rect 27508 14491 27534 14517
rect 32074 14491 32100 14517
rect 32136 14491 32162 14517
rect 32198 14491 32224 14517
rect 32260 14491 32286 14517
rect 32322 14491 32348 14517
rect 32384 14491 32410 14517
rect 32446 14491 32472 14517
rect 32508 14491 32534 14517
rect 37074 14491 37100 14517
rect 37136 14491 37162 14517
rect 37198 14491 37224 14517
rect 37260 14491 37286 14517
rect 37322 14491 37348 14517
rect 37384 14491 37410 14517
rect 37446 14491 37472 14517
rect 37508 14491 37534 14517
rect 1807 14295 1833 14321
rect 1919 14295 1945 14321
rect 2423 14295 2449 14321
rect 3823 14295 3849 14321
rect 4999 14295 5025 14321
rect 5279 14295 5305 14321
rect 6399 14295 6425 14321
rect 7799 14295 7825 14321
rect 8975 14295 9001 14321
rect 9255 14295 9281 14321
rect 10431 14295 10457 14321
rect 11999 14295 12025 14321
rect 12895 14295 12921 14321
rect 13231 14295 13257 14321
rect 14015 14295 14041 14321
rect 14799 14295 14825 14321
rect 15303 14295 15329 14321
rect 15471 14295 15497 14321
rect 16535 14295 16561 14321
rect 17431 14295 17457 14321
rect 18775 14295 18801 14321
rect 19335 14295 19361 14321
rect 19447 14295 19473 14321
rect 20231 14295 20257 14321
rect 21015 14295 21041 14321
rect 23031 14295 23057 14321
rect 23871 14295 23897 14321
rect 24431 14295 24457 14321
rect 25159 14295 25185 14321
rect 4999 14239 5025 14265
rect 6399 14239 6425 14265
rect 8975 14239 9001 14265
rect 10431 14239 10457 14265
rect 12895 14239 12921 14265
rect 14183 14239 14209 14265
rect 17431 14239 17457 14265
rect 21183 14239 21209 14265
rect 23871 14239 23897 14265
rect 25215 14239 25241 14265
rect 4574 14099 4600 14125
rect 4636 14099 4662 14125
rect 4698 14099 4724 14125
rect 4760 14099 4786 14125
rect 4822 14099 4848 14125
rect 4884 14099 4910 14125
rect 4946 14099 4972 14125
rect 5008 14099 5034 14125
rect 9574 14099 9600 14125
rect 9636 14099 9662 14125
rect 9698 14099 9724 14125
rect 9760 14099 9786 14125
rect 9822 14099 9848 14125
rect 9884 14099 9910 14125
rect 9946 14099 9972 14125
rect 10008 14099 10034 14125
rect 14574 14099 14600 14125
rect 14636 14099 14662 14125
rect 14698 14099 14724 14125
rect 14760 14099 14786 14125
rect 14822 14099 14848 14125
rect 14884 14099 14910 14125
rect 14946 14099 14972 14125
rect 15008 14099 15034 14125
rect 19574 14099 19600 14125
rect 19636 14099 19662 14125
rect 19698 14099 19724 14125
rect 19760 14099 19786 14125
rect 19822 14099 19848 14125
rect 19884 14099 19910 14125
rect 19946 14099 19972 14125
rect 20008 14099 20034 14125
rect 24574 14099 24600 14125
rect 24636 14099 24662 14125
rect 24698 14099 24724 14125
rect 24760 14099 24786 14125
rect 24822 14099 24848 14125
rect 24884 14099 24910 14125
rect 24946 14099 24972 14125
rect 25008 14099 25034 14125
rect 29574 14099 29600 14125
rect 29636 14099 29662 14125
rect 29698 14099 29724 14125
rect 29760 14099 29786 14125
rect 29822 14099 29848 14125
rect 29884 14099 29910 14125
rect 29946 14099 29972 14125
rect 30008 14099 30034 14125
rect 34574 14099 34600 14125
rect 34636 14099 34662 14125
rect 34698 14099 34724 14125
rect 34760 14099 34786 14125
rect 34822 14099 34848 14125
rect 34884 14099 34910 14125
rect 34946 14099 34972 14125
rect 35008 14099 35034 14125
rect 4495 13959 4521 13985
rect 6903 13959 6929 13985
rect 8471 13959 8497 13985
rect 10879 13959 10905 13985
rect 12447 13959 12473 13985
rect 14015 13959 14041 13985
rect 15471 13959 15497 13985
rect 17767 13959 17793 13985
rect 19447 13959 19473 13985
rect 21743 13959 21769 13985
rect 23423 13959 23449 13985
rect 2367 13903 2393 13929
rect 2479 13903 2505 13929
rect 3039 13903 3065 13929
rect 3375 13903 3401 13929
rect 4495 13903 4521 13929
rect 5839 13903 5865 13929
rect 6903 13903 6929 13929
rect 7575 13903 7601 13929
rect 8471 13903 8497 13929
rect 9815 13903 9841 13929
rect 10879 13903 10905 13929
rect 11551 13903 11577 13929
rect 12447 13903 12473 13929
rect 13119 13903 13145 13929
rect 14015 13903 14041 13929
rect 14575 13903 14601 13929
rect 15471 13903 15497 13929
rect 16983 13903 17009 13929
rect 17767 13903 17793 13929
rect 18551 13903 18577 13929
rect 19447 13903 19473 13929
rect 20791 13903 20817 13929
rect 21743 13903 21769 13929
rect 22527 13903 22553 13929
rect 23423 13903 23449 13929
rect 25047 13903 25073 13929
rect 25215 13903 25241 13929
rect 25439 13903 25465 13929
rect 2074 13707 2100 13733
rect 2136 13707 2162 13733
rect 2198 13707 2224 13733
rect 2260 13707 2286 13733
rect 2322 13707 2348 13733
rect 2384 13707 2410 13733
rect 2446 13707 2472 13733
rect 2508 13707 2534 13733
rect 7074 13707 7100 13733
rect 7136 13707 7162 13733
rect 7198 13707 7224 13733
rect 7260 13707 7286 13733
rect 7322 13707 7348 13733
rect 7384 13707 7410 13733
rect 7446 13707 7472 13733
rect 7508 13707 7534 13733
rect 12074 13707 12100 13733
rect 12136 13707 12162 13733
rect 12198 13707 12224 13733
rect 12260 13707 12286 13733
rect 12322 13707 12348 13733
rect 12384 13707 12410 13733
rect 12446 13707 12472 13733
rect 12508 13707 12534 13733
rect 17074 13707 17100 13733
rect 17136 13707 17162 13733
rect 17198 13707 17224 13733
rect 17260 13707 17286 13733
rect 17322 13707 17348 13733
rect 17384 13707 17410 13733
rect 17446 13707 17472 13733
rect 17508 13707 17534 13733
rect 22074 13707 22100 13733
rect 22136 13707 22162 13733
rect 22198 13707 22224 13733
rect 22260 13707 22286 13733
rect 22322 13707 22348 13733
rect 22384 13707 22410 13733
rect 22446 13707 22472 13733
rect 22508 13707 22534 13733
rect 27074 13707 27100 13733
rect 27136 13707 27162 13733
rect 27198 13707 27224 13733
rect 27260 13707 27286 13733
rect 27322 13707 27348 13733
rect 27384 13707 27410 13733
rect 27446 13707 27472 13733
rect 27508 13707 27534 13733
rect 32074 13707 32100 13733
rect 32136 13707 32162 13733
rect 32198 13707 32224 13733
rect 32260 13707 32286 13733
rect 32322 13707 32348 13733
rect 32384 13707 32410 13733
rect 32446 13707 32472 13733
rect 32508 13707 32534 13733
rect 37074 13707 37100 13733
rect 37136 13707 37162 13733
rect 37198 13707 37224 13733
rect 37260 13707 37286 13733
rect 37322 13707 37348 13733
rect 37384 13707 37410 13733
rect 37446 13707 37472 13733
rect 37508 13707 37534 13733
rect 1807 13511 1833 13537
rect 1919 13511 1945 13537
rect 2479 13511 2505 13537
rect 3823 13511 3849 13537
rect 4383 13511 4409 13537
rect 4495 13511 4521 13537
rect 5279 13511 5305 13537
rect 6399 13511 6425 13537
rect 7799 13511 7825 13537
rect 8359 13511 8385 13537
rect 8471 13511 8497 13537
rect 9255 13511 9281 13537
rect 10431 13511 10457 13537
rect 11215 13511 11241 13537
rect 12111 13511 12137 13537
rect 12671 13511 12697 13537
rect 13399 13511 13425 13537
rect 14799 13511 14825 13537
rect 15863 13511 15889 13537
rect 16535 13511 16561 13537
rect 17431 13511 17457 13537
rect 19055 13511 19081 13537
rect 19335 13511 19361 13537
rect 19447 13511 19473 13537
rect 20231 13511 20257 13537
rect 21015 13511 21041 13537
rect 23031 13511 23057 13537
rect 23871 13511 23897 13537
rect 24431 13511 24457 13537
rect 25215 13511 25241 13537
rect 6399 13455 6425 13481
rect 10431 13455 10457 13481
rect 12111 13455 12137 13481
rect 13399 13455 13425 13481
rect 15863 13455 15889 13481
rect 17431 13455 17457 13481
rect 21183 13455 21209 13481
rect 23871 13455 23897 13481
rect 25215 13455 25241 13481
rect 4574 13315 4600 13341
rect 4636 13315 4662 13341
rect 4698 13315 4724 13341
rect 4760 13315 4786 13341
rect 4822 13315 4848 13341
rect 4884 13315 4910 13341
rect 4946 13315 4972 13341
rect 5008 13315 5034 13341
rect 9574 13315 9600 13341
rect 9636 13315 9662 13341
rect 9698 13315 9724 13341
rect 9760 13315 9786 13341
rect 9822 13315 9848 13341
rect 9884 13315 9910 13341
rect 9946 13315 9972 13341
rect 10008 13315 10034 13341
rect 14574 13315 14600 13341
rect 14636 13315 14662 13341
rect 14698 13315 14724 13341
rect 14760 13315 14786 13341
rect 14822 13315 14848 13341
rect 14884 13315 14910 13341
rect 14946 13315 14972 13341
rect 15008 13315 15034 13341
rect 19574 13315 19600 13341
rect 19636 13315 19662 13341
rect 19698 13315 19724 13341
rect 19760 13315 19786 13341
rect 19822 13315 19848 13341
rect 19884 13315 19910 13341
rect 19946 13315 19972 13341
rect 20008 13315 20034 13341
rect 24574 13315 24600 13341
rect 24636 13315 24662 13341
rect 24698 13315 24724 13341
rect 24760 13315 24786 13341
rect 24822 13315 24848 13341
rect 24884 13315 24910 13341
rect 24946 13315 24972 13341
rect 25008 13315 25034 13341
rect 29574 13315 29600 13341
rect 29636 13315 29662 13341
rect 29698 13315 29724 13341
rect 29760 13315 29786 13341
rect 29822 13315 29848 13341
rect 29884 13315 29910 13341
rect 29946 13315 29972 13341
rect 30008 13315 30034 13341
rect 34574 13315 34600 13341
rect 34636 13315 34662 13341
rect 34698 13315 34724 13341
rect 34760 13315 34786 13341
rect 34822 13315 34848 13341
rect 34884 13315 34910 13341
rect 34946 13315 34972 13341
rect 35008 13315 35034 13341
rect 4495 13175 4521 13201
rect 6959 13175 6985 13201
rect 8359 13175 8385 13201
rect 10879 13175 10905 13201
rect 12447 13175 12473 13201
rect 14015 13175 14041 13201
rect 15303 13175 15329 13201
rect 17767 13175 17793 13201
rect 19447 13175 19473 13201
rect 23423 13175 23449 13201
rect 25943 13175 25969 13201
rect 2367 13119 2393 13145
rect 2591 13119 2617 13145
rect 2759 13119 2785 13145
rect 3319 13119 3345 13145
rect 4495 13119 4521 13145
rect 5839 13119 5865 13145
rect 6959 13119 6985 13145
rect 7575 13119 7601 13145
rect 8359 13119 8385 13145
rect 9815 13119 9841 13145
rect 10879 13119 10905 13145
rect 11551 13119 11577 13145
rect 12447 13119 12473 13145
rect 13119 13119 13145 13145
rect 14015 13119 14041 13145
rect 14463 13119 14489 13145
rect 15303 13119 15329 13145
rect 17095 13119 17121 13145
rect 17599 13119 17625 13145
rect 18551 13119 18577 13145
rect 19447 13119 19473 13145
rect 20959 13119 20985 13145
rect 21295 13119 21321 13145
rect 21463 13119 21489 13145
rect 22527 13119 22553 13145
rect 23423 13119 23449 13145
rect 25047 13119 25073 13145
rect 25943 13119 25969 13145
rect 2074 12923 2100 12949
rect 2136 12923 2162 12949
rect 2198 12923 2224 12949
rect 2260 12923 2286 12949
rect 2322 12923 2348 12949
rect 2384 12923 2410 12949
rect 2446 12923 2472 12949
rect 2508 12923 2534 12949
rect 7074 12923 7100 12949
rect 7136 12923 7162 12949
rect 7198 12923 7224 12949
rect 7260 12923 7286 12949
rect 7322 12923 7348 12949
rect 7384 12923 7410 12949
rect 7446 12923 7472 12949
rect 7508 12923 7534 12949
rect 12074 12923 12100 12949
rect 12136 12923 12162 12949
rect 12198 12923 12224 12949
rect 12260 12923 12286 12949
rect 12322 12923 12348 12949
rect 12384 12923 12410 12949
rect 12446 12923 12472 12949
rect 12508 12923 12534 12949
rect 17074 12923 17100 12949
rect 17136 12923 17162 12949
rect 17198 12923 17224 12949
rect 17260 12923 17286 12949
rect 17322 12923 17348 12949
rect 17384 12923 17410 12949
rect 17446 12923 17472 12949
rect 17508 12923 17534 12949
rect 22074 12923 22100 12949
rect 22136 12923 22162 12949
rect 22198 12923 22224 12949
rect 22260 12923 22286 12949
rect 22322 12923 22348 12949
rect 22384 12923 22410 12949
rect 22446 12923 22472 12949
rect 22508 12923 22534 12949
rect 27074 12923 27100 12949
rect 27136 12923 27162 12949
rect 27198 12923 27224 12949
rect 27260 12923 27286 12949
rect 27322 12923 27348 12949
rect 27384 12923 27410 12949
rect 27446 12923 27472 12949
rect 27508 12923 27534 12949
rect 32074 12923 32100 12949
rect 32136 12923 32162 12949
rect 32198 12923 32224 12949
rect 32260 12923 32286 12949
rect 32322 12923 32348 12949
rect 32384 12923 32410 12949
rect 32446 12923 32472 12949
rect 32508 12923 32534 12949
rect 37074 12923 37100 12949
rect 37136 12923 37162 12949
rect 37198 12923 37224 12949
rect 37260 12923 37286 12949
rect 37322 12923 37348 12949
rect 37384 12923 37410 12949
rect 37446 12923 37472 12949
rect 37508 12923 37534 12949
rect 1807 12727 1833 12753
rect 1975 12727 2001 12753
rect 2199 12727 2225 12753
rect 4103 12727 4129 12753
rect 4383 12727 4409 12753
rect 4495 12727 4521 12753
rect 5279 12727 5305 12753
rect 6455 12727 6481 12753
rect 7799 12727 7825 12753
rect 8359 12727 8385 12753
rect 8471 12727 8497 12753
rect 9255 12727 9281 12753
rect 10431 12727 10457 12753
rect 11999 12727 12025 12753
rect 12895 12727 12921 12753
rect 13343 12727 13369 12753
rect 14239 12727 14265 12753
rect 14799 12727 14825 12753
rect 15303 12727 15329 12753
rect 15471 12727 15497 12753
rect 16535 12727 16561 12753
rect 17431 12727 17457 12753
rect 19055 12727 19081 12753
rect 19335 12727 19361 12753
rect 19447 12727 19473 12753
rect 20511 12727 20537 12753
rect 21295 12727 21321 12753
rect 22975 12727 23001 12753
rect 23871 12727 23897 12753
rect 24487 12727 24513 12753
rect 25159 12727 25185 12753
rect 29639 12727 29665 12753
rect 29751 12727 29777 12753
rect 30199 12727 30225 12753
rect 6455 12671 6481 12697
rect 10431 12671 10457 12697
rect 12895 12671 12921 12697
rect 14239 12671 14265 12697
rect 17431 12671 17457 12697
rect 21295 12671 21321 12697
rect 23871 12671 23897 12697
rect 25159 12671 25185 12697
rect 4574 12531 4600 12557
rect 4636 12531 4662 12557
rect 4698 12531 4724 12557
rect 4760 12531 4786 12557
rect 4822 12531 4848 12557
rect 4884 12531 4910 12557
rect 4946 12531 4972 12557
rect 5008 12531 5034 12557
rect 9574 12531 9600 12557
rect 9636 12531 9662 12557
rect 9698 12531 9724 12557
rect 9760 12531 9786 12557
rect 9822 12531 9848 12557
rect 9884 12531 9910 12557
rect 9946 12531 9972 12557
rect 10008 12531 10034 12557
rect 14574 12531 14600 12557
rect 14636 12531 14662 12557
rect 14698 12531 14724 12557
rect 14760 12531 14786 12557
rect 14822 12531 14848 12557
rect 14884 12531 14910 12557
rect 14946 12531 14972 12557
rect 15008 12531 15034 12557
rect 19574 12531 19600 12557
rect 19636 12531 19662 12557
rect 19698 12531 19724 12557
rect 19760 12531 19786 12557
rect 19822 12531 19848 12557
rect 19884 12531 19910 12557
rect 19946 12531 19972 12557
rect 20008 12531 20034 12557
rect 24574 12531 24600 12557
rect 24636 12531 24662 12557
rect 24698 12531 24724 12557
rect 24760 12531 24786 12557
rect 24822 12531 24848 12557
rect 24884 12531 24910 12557
rect 24946 12531 24972 12557
rect 25008 12531 25034 12557
rect 29574 12531 29600 12557
rect 29636 12531 29662 12557
rect 29698 12531 29724 12557
rect 29760 12531 29786 12557
rect 29822 12531 29848 12557
rect 29884 12531 29910 12557
rect 29946 12531 29972 12557
rect 30008 12531 30034 12557
rect 34574 12531 34600 12557
rect 34636 12531 34662 12557
rect 34698 12531 34724 12557
rect 34760 12531 34786 12557
rect 34822 12531 34848 12557
rect 34884 12531 34910 12557
rect 34946 12531 34972 12557
rect 35008 12531 35034 12557
rect 1863 12391 1889 12417
rect 4495 12391 4521 12417
rect 7015 12391 7041 12417
rect 8359 12391 8385 12417
rect 10879 12391 10905 12417
rect 12447 12391 12473 12417
rect 14407 12391 14433 12417
rect 17991 12391 18017 12417
rect 19447 12391 19473 12417
rect 21799 12391 21825 12417
rect 23423 12391 23449 12417
rect 25943 12391 25969 12417
rect 27399 12391 27425 12417
rect 31599 12391 31625 12417
rect 1863 12335 1889 12361
rect 2759 12335 2785 12361
rect 3599 12335 3625 12361
rect 4495 12335 4521 12361
rect 5839 12335 5865 12361
rect 7015 12335 7041 12361
rect 7575 12335 7601 12361
rect 8359 12335 8385 12361
rect 9815 12335 9841 12361
rect 10879 12335 10905 12361
rect 11551 12335 11577 12361
rect 12447 12335 12473 12361
rect 13343 12335 13369 12361
rect 14407 12335 14433 12361
rect 14743 12335 14769 12361
rect 15303 12335 15329 12361
rect 15415 12335 15441 12361
rect 16815 12335 16841 12361
rect 17991 12335 18017 12361
rect 18551 12335 18577 12361
rect 19447 12335 19473 12361
rect 20903 12335 20929 12361
rect 21799 12335 21825 12361
rect 22527 12335 22553 12361
rect 23423 12335 23449 12361
rect 24767 12335 24793 12361
rect 25943 12335 25969 12361
rect 26503 12335 26529 12361
rect 27399 12335 27425 12361
rect 29695 12335 29721 12361
rect 29919 12335 29945 12361
rect 30367 12335 30393 12361
rect 30703 12335 30729 12361
rect 31599 12335 31625 12361
rect 2074 12139 2100 12165
rect 2136 12139 2162 12165
rect 2198 12139 2224 12165
rect 2260 12139 2286 12165
rect 2322 12139 2348 12165
rect 2384 12139 2410 12165
rect 2446 12139 2472 12165
rect 2508 12139 2534 12165
rect 7074 12139 7100 12165
rect 7136 12139 7162 12165
rect 7198 12139 7224 12165
rect 7260 12139 7286 12165
rect 7322 12139 7348 12165
rect 7384 12139 7410 12165
rect 7446 12139 7472 12165
rect 7508 12139 7534 12165
rect 12074 12139 12100 12165
rect 12136 12139 12162 12165
rect 12198 12139 12224 12165
rect 12260 12139 12286 12165
rect 12322 12139 12348 12165
rect 12384 12139 12410 12165
rect 12446 12139 12472 12165
rect 12508 12139 12534 12165
rect 17074 12139 17100 12165
rect 17136 12139 17162 12165
rect 17198 12139 17224 12165
rect 17260 12139 17286 12165
rect 17322 12139 17348 12165
rect 17384 12139 17410 12165
rect 17446 12139 17472 12165
rect 17508 12139 17534 12165
rect 22074 12139 22100 12165
rect 22136 12139 22162 12165
rect 22198 12139 22224 12165
rect 22260 12139 22286 12165
rect 22322 12139 22348 12165
rect 22384 12139 22410 12165
rect 22446 12139 22472 12165
rect 22508 12139 22534 12165
rect 27074 12139 27100 12165
rect 27136 12139 27162 12165
rect 27198 12139 27224 12165
rect 27260 12139 27286 12165
rect 27322 12139 27348 12165
rect 27384 12139 27410 12165
rect 27446 12139 27472 12165
rect 27508 12139 27534 12165
rect 32074 12139 32100 12165
rect 32136 12139 32162 12165
rect 32198 12139 32224 12165
rect 32260 12139 32286 12165
rect 32322 12139 32348 12165
rect 32384 12139 32410 12165
rect 32446 12139 32472 12165
rect 32508 12139 32534 12165
rect 37074 12139 37100 12165
rect 37136 12139 37162 12165
rect 37198 12139 37224 12165
rect 37260 12139 37286 12165
rect 37322 12139 37348 12165
rect 37384 12139 37410 12165
rect 37446 12139 37472 12165
rect 37508 12139 37534 12165
rect 1807 11943 1833 11969
rect 1919 11943 1945 11969
rect 2199 11943 2225 11969
rect 4103 11943 4129 11969
rect 4327 11943 4353 11969
rect 4495 11943 4521 11969
rect 5279 11943 5305 11969
rect 6399 11943 6425 11969
rect 7799 11943 7825 11969
rect 8359 11943 8385 11969
rect 8471 11943 8497 11969
rect 9255 11943 9281 11969
rect 10431 11943 10457 11969
rect 11999 11943 12025 11969
rect 12951 11943 12977 11969
rect 13343 11943 13369 11969
rect 14407 11943 14433 11969
rect 14799 11943 14825 11969
rect 15863 11943 15889 11969
rect 16535 11943 16561 11969
rect 17431 11943 17457 11969
rect 19055 11943 19081 11969
rect 19951 11943 19977 11969
rect 20511 11943 20537 11969
rect 21407 11943 21433 11969
rect 23031 11943 23057 11969
rect 23311 11943 23337 11969
rect 23423 11943 23449 11969
rect 24487 11943 24513 11969
rect 25159 11943 25185 11969
rect 26727 11943 26753 11969
rect 27679 11943 27705 11969
rect 28239 11943 28265 11969
rect 29359 11943 29385 11969
rect 30703 11943 30729 11969
rect 31599 11943 31625 11969
rect 32439 11943 32465 11969
rect 32831 11943 32857 11969
rect 6399 11887 6425 11913
rect 10431 11887 10457 11913
rect 12951 11887 12977 11913
rect 14407 11887 14433 11913
rect 15863 11887 15889 11913
rect 17431 11887 17457 11913
rect 19951 11887 19977 11913
rect 21407 11887 21433 11913
rect 25159 11887 25185 11913
rect 27679 11887 27705 11913
rect 29359 11887 29385 11913
rect 31655 11887 31681 11913
rect 33111 11887 33137 11913
rect 4574 11747 4600 11773
rect 4636 11747 4662 11773
rect 4698 11747 4724 11773
rect 4760 11747 4786 11773
rect 4822 11747 4848 11773
rect 4884 11747 4910 11773
rect 4946 11747 4972 11773
rect 5008 11747 5034 11773
rect 9574 11747 9600 11773
rect 9636 11747 9662 11773
rect 9698 11747 9724 11773
rect 9760 11747 9786 11773
rect 9822 11747 9848 11773
rect 9884 11747 9910 11773
rect 9946 11747 9972 11773
rect 10008 11747 10034 11773
rect 14574 11747 14600 11773
rect 14636 11747 14662 11773
rect 14698 11747 14724 11773
rect 14760 11747 14786 11773
rect 14822 11747 14848 11773
rect 14884 11747 14910 11773
rect 14946 11747 14972 11773
rect 15008 11747 15034 11773
rect 19574 11747 19600 11773
rect 19636 11747 19662 11773
rect 19698 11747 19724 11773
rect 19760 11747 19786 11773
rect 19822 11747 19848 11773
rect 19884 11747 19910 11773
rect 19946 11747 19972 11773
rect 20008 11747 20034 11773
rect 24574 11747 24600 11773
rect 24636 11747 24662 11773
rect 24698 11747 24724 11773
rect 24760 11747 24786 11773
rect 24822 11747 24848 11773
rect 24884 11747 24910 11773
rect 24946 11747 24972 11773
rect 25008 11747 25034 11773
rect 29574 11747 29600 11773
rect 29636 11747 29662 11773
rect 29698 11747 29724 11773
rect 29760 11747 29786 11773
rect 29822 11747 29848 11773
rect 29884 11747 29910 11773
rect 29946 11747 29972 11773
rect 30008 11747 30034 11773
rect 34574 11747 34600 11773
rect 34636 11747 34662 11773
rect 34698 11747 34724 11773
rect 34760 11747 34786 11773
rect 34822 11747 34848 11773
rect 34884 11747 34910 11773
rect 34946 11747 34972 11773
rect 35008 11747 35034 11773
rect 1863 11607 1889 11633
rect 4439 11607 4465 11633
rect 7015 11607 7041 11633
rect 8359 11607 8385 11633
rect 10767 11607 10793 11633
rect 12447 11607 12473 11633
rect 14463 11607 14489 11633
rect 15863 11607 15889 11633
rect 17991 11607 18017 11633
rect 23311 11607 23337 11633
rect 28351 11607 28377 11633
rect 31487 11607 31513 11633
rect 1863 11551 1889 11577
rect 3039 11551 3065 11577
rect 3599 11551 3625 11577
rect 4439 11551 4465 11577
rect 5839 11551 5865 11577
rect 7015 11551 7041 11577
rect 7575 11551 7601 11577
rect 8359 11551 8385 11577
rect 10039 11551 10065 11577
rect 10767 11551 10793 11577
rect 11551 11551 11577 11577
rect 12447 11551 12473 11577
rect 13455 11551 13481 11577
rect 14463 11551 14489 11577
rect 15079 11551 15105 11577
rect 15863 11551 15889 11577
rect 16815 11551 16841 11577
rect 17991 11551 18017 11577
rect 18551 11551 18577 11577
rect 18831 11551 18857 11577
rect 18943 11551 18969 11577
rect 20791 11551 20817 11577
rect 21351 11551 21377 11577
rect 21463 11551 21489 11577
rect 22527 11551 22553 11577
rect 23311 11551 23337 11577
rect 24767 11551 24793 11577
rect 25215 11551 25241 11577
rect 25439 11551 25465 11577
rect 27455 11551 27481 11577
rect 28351 11551 28377 11577
rect 28855 11551 28881 11577
rect 29415 11551 29441 11577
rect 29527 11551 29553 11577
rect 30591 11551 30617 11577
rect 31487 11551 31513 11577
rect 32775 11551 32801 11577
rect 33167 11551 33193 11577
rect 33615 11551 33641 11577
rect 2074 11355 2100 11381
rect 2136 11355 2162 11381
rect 2198 11355 2224 11381
rect 2260 11355 2286 11381
rect 2322 11355 2348 11381
rect 2384 11355 2410 11381
rect 2446 11355 2472 11381
rect 2508 11355 2534 11381
rect 7074 11355 7100 11381
rect 7136 11355 7162 11381
rect 7198 11355 7224 11381
rect 7260 11355 7286 11381
rect 7322 11355 7348 11381
rect 7384 11355 7410 11381
rect 7446 11355 7472 11381
rect 7508 11355 7534 11381
rect 12074 11355 12100 11381
rect 12136 11355 12162 11381
rect 12198 11355 12224 11381
rect 12260 11355 12286 11381
rect 12322 11355 12348 11381
rect 12384 11355 12410 11381
rect 12446 11355 12472 11381
rect 12508 11355 12534 11381
rect 17074 11355 17100 11381
rect 17136 11355 17162 11381
rect 17198 11355 17224 11381
rect 17260 11355 17286 11381
rect 17322 11355 17348 11381
rect 17384 11355 17410 11381
rect 17446 11355 17472 11381
rect 17508 11355 17534 11381
rect 22074 11355 22100 11381
rect 22136 11355 22162 11381
rect 22198 11355 22224 11381
rect 22260 11355 22286 11381
rect 22322 11355 22348 11381
rect 22384 11355 22410 11381
rect 22446 11355 22472 11381
rect 22508 11355 22534 11381
rect 27074 11355 27100 11381
rect 27136 11355 27162 11381
rect 27198 11355 27224 11381
rect 27260 11355 27286 11381
rect 27322 11355 27348 11381
rect 27384 11355 27410 11381
rect 27446 11355 27472 11381
rect 27508 11355 27534 11381
rect 32074 11355 32100 11381
rect 32136 11355 32162 11381
rect 32198 11355 32224 11381
rect 32260 11355 32286 11381
rect 32322 11355 32348 11381
rect 32384 11355 32410 11381
rect 32446 11355 32472 11381
rect 32508 11355 32534 11381
rect 37074 11355 37100 11381
rect 37136 11355 37162 11381
rect 37198 11355 37224 11381
rect 37260 11355 37286 11381
rect 37322 11355 37348 11381
rect 37384 11355 37410 11381
rect 37446 11355 37472 11381
rect 37508 11355 37534 11381
rect 1807 11159 1833 11185
rect 1919 11159 1945 11185
rect 2479 11159 2505 11185
rect 3823 11159 3849 11185
rect 4383 11159 4409 11185
rect 4495 11159 4521 11185
rect 5279 11159 5305 11185
rect 6455 11159 6481 11185
rect 7799 11159 7825 11185
rect 8359 11159 8385 11185
rect 8471 11159 8497 11185
rect 9255 11159 9281 11185
rect 10431 11159 10457 11185
rect 11999 11159 12025 11185
rect 12951 11159 12977 11185
rect 13343 11159 13369 11185
rect 14407 11159 14433 11185
rect 15079 11159 15105 11185
rect 15303 11159 15329 11185
rect 15471 11159 15497 11185
rect 16535 11159 16561 11185
rect 17263 11159 17289 11185
rect 18775 11159 18801 11185
rect 19223 11159 19249 11185
rect 19951 11159 19977 11185
rect 20231 11159 20257 11185
rect 21351 11159 21377 11185
rect 23031 11159 23057 11185
rect 23311 11159 23337 11185
rect 23423 11159 23449 11185
rect 24375 11159 24401 11185
rect 25159 11159 25185 11185
rect 27567 11159 27593 11185
rect 28519 11159 28545 11185
rect 28799 11159 28825 11185
rect 29975 11159 30001 11185
rect 30759 11159 30785 11185
rect 31487 11159 31513 11185
rect 32439 11159 32465 11185
rect 33111 11159 33137 11185
rect 34959 11159 34985 11185
rect 35127 11159 35153 11185
rect 35351 11159 35377 11185
rect 36135 11159 36161 11185
rect 37311 11159 37337 11185
rect 6455 11103 6481 11129
rect 10431 11103 10457 11129
rect 12951 11103 12977 11129
rect 14407 11103 14433 11129
rect 17263 11103 17289 11129
rect 21351 11103 21377 11129
rect 25159 11103 25185 11129
rect 28519 11103 28545 11129
rect 29975 11103 30001 11129
rect 31655 11103 31681 11129
rect 33111 11103 33137 11129
rect 37311 11103 37337 11129
rect 4574 10963 4600 10989
rect 4636 10963 4662 10989
rect 4698 10963 4724 10989
rect 4760 10963 4786 10989
rect 4822 10963 4848 10989
rect 4884 10963 4910 10989
rect 4946 10963 4972 10989
rect 5008 10963 5034 10989
rect 9574 10963 9600 10989
rect 9636 10963 9662 10989
rect 9698 10963 9724 10989
rect 9760 10963 9786 10989
rect 9822 10963 9848 10989
rect 9884 10963 9910 10989
rect 9946 10963 9972 10989
rect 10008 10963 10034 10989
rect 14574 10963 14600 10989
rect 14636 10963 14662 10989
rect 14698 10963 14724 10989
rect 14760 10963 14786 10989
rect 14822 10963 14848 10989
rect 14884 10963 14910 10989
rect 14946 10963 14972 10989
rect 15008 10963 15034 10989
rect 19574 10963 19600 10989
rect 19636 10963 19662 10989
rect 19698 10963 19724 10989
rect 19760 10963 19786 10989
rect 19822 10963 19848 10989
rect 19884 10963 19910 10989
rect 19946 10963 19972 10989
rect 20008 10963 20034 10989
rect 24574 10963 24600 10989
rect 24636 10963 24662 10989
rect 24698 10963 24724 10989
rect 24760 10963 24786 10989
rect 24822 10963 24848 10989
rect 24884 10963 24910 10989
rect 24946 10963 24972 10989
rect 25008 10963 25034 10989
rect 29574 10963 29600 10989
rect 29636 10963 29662 10989
rect 29698 10963 29724 10989
rect 29760 10963 29786 10989
rect 29822 10963 29848 10989
rect 29884 10963 29910 10989
rect 29946 10963 29972 10989
rect 30008 10963 30034 10989
rect 34574 10963 34600 10989
rect 34636 10963 34662 10989
rect 34698 10963 34724 10989
rect 34760 10963 34786 10989
rect 34822 10963 34848 10989
rect 34884 10963 34910 10989
rect 34946 10963 34972 10989
rect 35008 10963 35034 10989
rect 2087 10823 2113 10849
rect 4439 10823 4465 10849
rect 7015 10823 7041 10849
rect 8471 10823 8497 10849
rect 10767 10823 10793 10849
rect 12223 10823 12249 10849
rect 14463 10823 14489 10849
rect 19279 10823 19305 10849
rect 23423 10823 23449 10849
rect 28295 10823 28321 10849
rect 29975 10823 30001 10849
rect 31431 10823 31457 10849
rect 37647 10823 37673 10849
rect 2087 10767 2113 10793
rect 3039 10767 3065 10793
rect 3599 10767 3625 10793
rect 4439 10767 4465 10793
rect 5839 10767 5865 10793
rect 7015 10767 7041 10793
rect 7295 10767 7321 10793
rect 8471 10767 8497 10793
rect 10039 10767 10065 10793
rect 10767 10767 10793 10793
rect 11551 10767 11577 10793
rect 12223 10767 12249 10793
rect 13455 10767 13481 10793
rect 14463 10767 14489 10793
rect 15079 10767 15105 10793
rect 15359 10767 15385 10793
rect 15583 10767 15609 10793
rect 16815 10767 16841 10793
rect 17263 10767 17289 10793
rect 17487 10767 17513 10793
rect 18551 10767 18577 10793
rect 19279 10767 19305 10793
rect 20791 10767 20817 10793
rect 21351 10767 21377 10793
rect 21463 10767 21489 10793
rect 22527 10767 22553 10793
rect 23423 10767 23449 10793
rect 25047 10767 25073 10793
rect 25327 10767 25353 10793
rect 25439 10767 25465 10793
rect 27455 10767 27481 10793
rect 28295 10767 28321 10793
rect 28799 10767 28825 10793
rect 29975 10767 30001 10793
rect 30311 10767 30337 10793
rect 31431 10767 31457 10793
rect 32775 10767 32801 10793
rect 33167 10767 33193 10793
rect 33391 10767 33417 10793
rect 34455 10767 34481 10793
rect 34623 10767 34649 10793
rect 34847 10767 34873 10793
rect 36695 10767 36721 10793
rect 37647 10767 37673 10793
rect 2074 10571 2100 10597
rect 2136 10571 2162 10597
rect 2198 10571 2224 10597
rect 2260 10571 2286 10597
rect 2322 10571 2348 10597
rect 2384 10571 2410 10597
rect 2446 10571 2472 10597
rect 2508 10571 2534 10597
rect 7074 10571 7100 10597
rect 7136 10571 7162 10597
rect 7198 10571 7224 10597
rect 7260 10571 7286 10597
rect 7322 10571 7348 10597
rect 7384 10571 7410 10597
rect 7446 10571 7472 10597
rect 7508 10571 7534 10597
rect 12074 10571 12100 10597
rect 12136 10571 12162 10597
rect 12198 10571 12224 10597
rect 12260 10571 12286 10597
rect 12322 10571 12348 10597
rect 12384 10571 12410 10597
rect 12446 10571 12472 10597
rect 12508 10571 12534 10597
rect 17074 10571 17100 10597
rect 17136 10571 17162 10597
rect 17198 10571 17224 10597
rect 17260 10571 17286 10597
rect 17322 10571 17348 10597
rect 17384 10571 17410 10597
rect 17446 10571 17472 10597
rect 17508 10571 17534 10597
rect 22074 10571 22100 10597
rect 22136 10571 22162 10597
rect 22198 10571 22224 10597
rect 22260 10571 22286 10597
rect 22322 10571 22348 10597
rect 22384 10571 22410 10597
rect 22446 10571 22472 10597
rect 22508 10571 22534 10597
rect 27074 10571 27100 10597
rect 27136 10571 27162 10597
rect 27198 10571 27224 10597
rect 27260 10571 27286 10597
rect 27322 10571 27348 10597
rect 27384 10571 27410 10597
rect 27446 10571 27472 10597
rect 27508 10571 27534 10597
rect 32074 10571 32100 10597
rect 32136 10571 32162 10597
rect 32198 10571 32224 10597
rect 32260 10571 32286 10597
rect 32322 10571 32348 10597
rect 32384 10571 32410 10597
rect 32446 10571 32472 10597
rect 32508 10571 32534 10597
rect 37074 10571 37100 10597
rect 37136 10571 37162 10597
rect 37198 10571 37224 10597
rect 37260 10571 37286 10597
rect 37322 10571 37348 10597
rect 37384 10571 37410 10597
rect 37446 10571 37472 10597
rect 37508 10571 37534 10597
rect 1639 10375 1665 10401
rect 2479 10375 2505 10401
rect 3823 10375 3849 10401
rect 4383 10375 4409 10401
rect 4495 10375 4521 10401
rect 5279 10375 5305 10401
rect 6455 10375 6481 10401
rect 7799 10375 7825 10401
rect 8751 10375 8777 10401
rect 9255 10375 9281 10401
rect 10431 10375 10457 10401
rect 11943 10375 11969 10401
rect 12671 10375 12697 10401
rect 13343 10375 13369 10401
rect 14295 10375 14321 10401
rect 15079 10375 15105 10401
rect 15359 10375 15385 10401
rect 15471 10375 15497 10401
rect 16535 10375 16561 10401
rect 16815 10375 16841 10401
rect 16927 10375 16953 10401
rect 18775 10375 18801 10401
rect 19279 10375 19305 10401
rect 19503 10375 19529 10401
rect 20231 10375 20257 10401
rect 21351 10375 21377 10401
rect 23031 10375 23057 10401
rect 23871 10375 23897 10401
rect 24375 10375 24401 10401
rect 24655 10375 24681 10401
rect 24879 10375 24905 10401
rect 27679 10375 27705 10401
rect 28071 10375 28097 10401
rect 28519 10375 28545 10401
rect 28799 10375 28825 10401
rect 29975 10375 30001 10401
rect 30703 10375 30729 10401
rect 31263 10375 31289 10401
rect 31431 10375 31457 10401
rect 32159 10375 32185 10401
rect 33111 10375 33137 10401
rect 34959 10375 34985 10401
rect 35239 10375 35265 10401
rect 35351 10375 35377 10401
rect 36135 10375 36161 10401
rect 37311 10375 37337 10401
rect 1527 10319 1553 10345
rect 6455 10319 6481 10345
rect 8751 10319 8777 10345
rect 10431 10319 10457 10345
rect 12671 10319 12697 10345
rect 14295 10319 14321 10345
rect 21351 10319 21377 10345
rect 23871 10319 23897 10345
rect 29975 10319 30001 10345
rect 33111 10319 33137 10345
rect 37311 10319 37337 10345
rect 4574 10179 4600 10205
rect 4636 10179 4662 10205
rect 4698 10179 4724 10205
rect 4760 10179 4786 10205
rect 4822 10179 4848 10205
rect 4884 10179 4910 10205
rect 4946 10179 4972 10205
rect 5008 10179 5034 10205
rect 9574 10179 9600 10205
rect 9636 10179 9662 10205
rect 9698 10179 9724 10205
rect 9760 10179 9786 10205
rect 9822 10179 9848 10205
rect 9884 10179 9910 10205
rect 9946 10179 9972 10205
rect 10008 10179 10034 10205
rect 14574 10179 14600 10205
rect 14636 10179 14662 10205
rect 14698 10179 14724 10205
rect 14760 10179 14786 10205
rect 14822 10179 14848 10205
rect 14884 10179 14910 10205
rect 14946 10179 14972 10205
rect 15008 10179 15034 10205
rect 19574 10179 19600 10205
rect 19636 10179 19662 10205
rect 19698 10179 19724 10205
rect 19760 10179 19786 10205
rect 19822 10179 19848 10205
rect 19884 10179 19910 10205
rect 19946 10179 19972 10205
rect 20008 10179 20034 10205
rect 24574 10179 24600 10205
rect 24636 10179 24662 10205
rect 24698 10179 24724 10205
rect 24760 10179 24786 10205
rect 24822 10179 24848 10205
rect 24884 10179 24910 10205
rect 24946 10179 24972 10205
rect 25008 10179 25034 10205
rect 29574 10179 29600 10205
rect 29636 10179 29662 10205
rect 29698 10179 29724 10205
rect 29760 10179 29786 10205
rect 29822 10179 29848 10205
rect 29884 10179 29910 10205
rect 29946 10179 29972 10205
rect 30008 10179 30034 10205
rect 34574 10179 34600 10205
rect 34636 10179 34662 10205
rect 34698 10179 34724 10205
rect 34760 10179 34786 10205
rect 34822 10179 34848 10205
rect 34884 10179 34910 10205
rect 34946 10179 34972 10205
rect 35008 10179 35034 10205
rect 1863 10039 1889 10065
rect 7015 10039 7041 10065
rect 8471 10039 8497 10065
rect 17991 10039 18017 10065
rect 19447 10039 19473 10065
rect 23423 10039 23449 10065
rect 25943 10039 25969 10065
rect 37647 10039 37673 10065
rect 1863 9983 1889 10009
rect 2759 9983 2785 10009
rect 3599 9983 3625 10009
rect 3823 9983 3849 10009
rect 3991 9983 4017 10009
rect 5895 9983 5921 10009
rect 7015 9983 7041 10009
rect 7575 9983 7601 10009
rect 8471 9983 8497 10009
rect 10039 9983 10065 10009
rect 10375 9983 10401 10009
rect 10543 9983 10569 10009
rect 11551 9983 11577 10009
rect 11775 9983 11801 10009
rect 11943 9983 11969 10009
rect 13623 9983 13649 10009
rect 14071 9983 14097 10009
rect 14295 9983 14321 10009
rect 15079 9983 15105 10009
rect 15527 9983 15553 10009
rect 15751 9983 15777 10009
rect 16815 9983 16841 10009
rect 17991 9983 18017 10009
rect 18271 9983 18297 10009
rect 19447 9983 19473 10009
rect 20791 9983 20817 10009
rect 21351 9983 21377 10009
rect 21463 9983 21489 10009
rect 22247 9983 22273 10009
rect 23423 9983 23449 10009
rect 25943 9983 25969 10009
rect 26839 9983 26865 10009
rect 27679 9983 27705 10009
rect 27903 9983 27929 10009
rect 28351 9983 28377 10009
rect 29415 9983 29441 10009
rect 29807 9983 29833 10009
rect 30031 9983 30057 10009
rect 30815 9983 30841 10009
rect 31375 9983 31401 10009
rect 31487 9983 31513 10009
rect 32831 9983 32857 10009
rect 33167 9983 33193 10009
rect 33615 9983 33641 10009
rect 34455 9983 34481 10009
rect 34623 9983 34649 10009
rect 34847 9983 34873 10009
rect 36695 9983 36721 10009
rect 37647 9983 37673 10009
rect 2074 9787 2100 9813
rect 2136 9787 2162 9813
rect 2198 9787 2224 9813
rect 2260 9787 2286 9813
rect 2322 9787 2348 9813
rect 2384 9787 2410 9813
rect 2446 9787 2472 9813
rect 2508 9787 2534 9813
rect 7074 9787 7100 9813
rect 7136 9787 7162 9813
rect 7198 9787 7224 9813
rect 7260 9787 7286 9813
rect 7322 9787 7348 9813
rect 7384 9787 7410 9813
rect 7446 9787 7472 9813
rect 7508 9787 7534 9813
rect 12074 9787 12100 9813
rect 12136 9787 12162 9813
rect 12198 9787 12224 9813
rect 12260 9787 12286 9813
rect 12322 9787 12348 9813
rect 12384 9787 12410 9813
rect 12446 9787 12472 9813
rect 12508 9787 12534 9813
rect 17074 9787 17100 9813
rect 17136 9787 17162 9813
rect 17198 9787 17224 9813
rect 17260 9787 17286 9813
rect 17322 9787 17348 9813
rect 17384 9787 17410 9813
rect 17446 9787 17472 9813
rect 17508 9787 17534 9813
rect 22074 9787 22100 9813
rect 22136 9787 22162 9813
rect 22198 9787 22224 9813
rect 22260 9787 22286 9813
rect 22322 9787 22348 9813
rect 22384 9787 22410 9813
rect 22446 9787 22472 9813
rect 22508 9787 22534 9813
rect 27074 9787 27100 9813
rect 27136 9787 27162 9813
rect 27198 9787 27224 9813
rect 27260 9787 27286 9813
rect 27322 9787 27348 9813
rect 27384 9787 27410 9813
rect 27446 9787 27472 9813
rect 27508 9787 27534 9813
rect 32074 9787 32100 9813
rect 32136 9787 32162 9813
rect 32198 9787 32224 9813
rect 32260 9787 32286 9813
rect 32322 9787 32348 9813
rect 32384 9787 32410 9813
rect 32446 9787 32472 9813
rect 32508 9787 32534 9813
rect 37074 9787 37100 9813
rect 37136 9787 37162 9813
rect 37198 9787 37224 9813
rect 37260 9787 37286 9813
rect 37322 9787 37348 9813
rect 37384 9787 37410 9813
rect 37446 9787 37472 9813
rect 37508 9787 37534 9813
rect 1807 9591 1833 9617
rect 2031 9591 2057 9617
rect 2479 9591 2505 9617
rect 3823 9591 3849 9617
rect 4999 9591 5025 9617
rect 5279 9591 5305 9617
rect 5951 9591 5977 9617
rect 7799 9591 7825 9617
rect 8751 9591 8777 9617
rect 9255 9591 9281 9617
rect 10431 9591 10457 9617
rect 11607 9591 11633 9617
rect 12055 9591 12081 9617
rect 12279 9591 12305 9617
rect 13343 9591 13369 9617
rect 14015 9591 14041 9617
rect 14799 9591 14825 9617
rect 15247 9591 15273 9617
rect 15471 9591 15497 9617
rect 16255 9591 16281 9617
rect 16815 9591 16841 9617
rect 16927 9591 16953 9617
rect 18775 9591 18801 9617
rect 19335 9591 19361 9617
rect 19447 9591 19473 9617
rect 20231 9591 20257 9617
rect 21351 9591 21377 9617
rect 22751 9591 22777 9617
rect 23871 9591 23897 9617
rect 24431 9591 24457 9617
rect 25383 9591 25409 9617
rect 28183 9591 28209 9617
rect 28407 9591 28433 9617
rect 28799 9591 28825 9617
rect 29415 9591 29441 9617
rect 29695 9591 29721 9617
rect 29807 9591 29833 9617
rect 30983 9591 31009 9617
rect 31151 9591 31177 9617
rect 31375 9591 31401 9617
rect 32159 9591 32185 9617
rect 32831 9591 32857 9617
rect 34959 9591 34985 9617
rect 35127 9591 35153 9617
rect 35351 9591 35377 9617
rect 36415 9591 36441 9617
rect 37311 9591 37337 9617
rect 3823 9535 3849 9561
rect 6231 9535 6257 9561
rect 8751 9535 8777 9561
rect 10431 9535 10457 9561
rect 14015 9535 14041 9561
rect 21351 9535 21377 9561
rect 23871 9535 23897 9561
rect 25383 9535 25409 9561
rect 33111 9535 33137 9561
rect 37311 9535 37337 9561
rect 4574 9395 4600 9421
rect 4636 9395 4662 9421
rect 4698 9395 4724 9421
rect 4760 9395 4786 9421
rect 4822 9395 4848 9421
rect 4884 9395 4910 9421
rect 4946 9395 4972 9421
rect 5008 9395 5034 9421
rect 9574 9395 9600 9421
rect 9636 9395 9662 9421
rect 9698 9395 9724 9421
rect 9760 9395 9786 9421
rect 9822 9395 9848 9421
rect 9884 9395 9910 9421
rect 9946 9395 9972 9421
rect 10008 9395 10034 9421
rect 14574 9395 14600 9421
rect 14636 9395 14662 9421
rect 14698 9395 14724 9421
rect 14760 9395 14786 9421
rect 14822 9395 14848 9421
rect 14884 9395 14910 9421
rect 14946 9395 14972 9421
rect 15008 9395 15034 9421
rect 19574 9395 19600 9421
rect 19636 9395 19662 9421
rect 19698 9395 19724 9421
rect 19760 9395 19786 9421
rect 19822 9395 19848 9421
rect 19884 9395 19910 9421
rect 19946 9395 19972 9421
rect 20008 9395 20034 9421
rect 24574 9395 24600 9421
rect 24636 9395 24662 9421
rect 24698 9395 24724 9421
rect 24760 9395 24786 9421
rect 24822 9395 24848 9421
rect 24884 9395 24910 9421
rect 24946 9395 24972 9421
rect 25008 9395 25034 9421
rect 29574 9395 29600 9421
rect 29636 9395 29662 9421
rect 29698 9395 29724 9421
rect 29760 9395 29786 9421
rect 29822 9395 29848 9421
rect 29884 9395 29910 9421
rect 29946 9395 29972 9421
rect 30008 9395 30034 9421
rect 34574 9395 34600 9421
rect 34636 9395 34662 9421
rect 34698 9395 34724 9421
rect 34760 9395 34786 9421
rect 34822 9395 34848 9421
rect 34884 9395 34910 9421
rect 34946 9395 34972 9421
rect 35008 9395 35034 9421
rect 1863 9255 1889 9281
rect 3375 9255 3401 9281
rect 8415 9255 8441 9281
rect 15751 9255 15777 9281
rect 17991 9255 18017 9281
rect 19335 9255 19361 9281
rect 23423 9255 23449 9281
rect 25943 9255 25969 9281
rect 27735 9255 27761 9281
rect 30199 9255 30225 9281
rect 35239 9255 35265 9281
rect 37647 9255 37673 9281
rect 1863 9199 1889 9225
rect 3039 9199 3065 9225
rect 3375 9199 3401 9225
rect 4495 9199 4521 9225
rect 6119 9199 6145 9225
rect 6287 9199 6313 9225
rect 6511 9199 6537 9225
rect 7575 9199 7601 9225
rect 8415 9199 8441 9225
rect 10039 9199 10065 9225
rect 10319 9199 10345 9225
rect 10487 9199 10513 9225
rect 11439 9199 11465 9225
rect 11775 9199 11801 9225
rect 11943 9199 11969 9225
rect 13343 9199 13369 9225
rect 13791 9199 13817 9225
rect 14015 9199 14041 9225
rect 14799 9199 14825 9225
rect 15751 9199 15777 9225
rect 16815 9199 16841 9225
rect 17991 9199 18017 9225
rect 18271 9199 18297 9225
rect 19279 9199 19305 9225
rect 20791 9199 20817 9225
rect 21351 9199 21377 9225
rect 21463 9199 21489 9225
rect 22527 9199 22553 9225
rect 23423 9199 23449 9225
rect 25047 9199 25073 9225
rect 25943 9199 25969 9225
rect 26951 9199 26977 9225
rect 27623 9199 27649 9225
rect 29527 9199 29553 9225
rect 30199 9199 30225 9225
rect 30983 9199 31009 9225
rect 31151 9199 31177 9225
rect 31375 9199 31401 9225
rect 32831 9199 32857 9225
rect 33167 9199 33193 9225
rect 33615 9199 33641 9225
rect 34175 9199 34201 9225
rect 35239 9199 35265 9225
rect 36695 9199 36721 9225
rect 37647 9199 37673 9225
rect 2074 9003 2100 9029
rect 2136 9003 2162 9029
rect 2198 9003 2224 9029
rect 2260 9003 2286 9029
rect 2322 9003 2348 9029
rect 2384 9003 2410 9029
rect 2446 9003 2472 9029
rect 2508 9003 2534 9029
rect 7074 9003 7100 9029
rect 7136 9003 7162 9029
rect 7198 9003 7224 9029
rect 7260 9003 7286 9029
rect 7322 9003 7348 9029
rect 7384 9003 7410 9029
rect 7446 9003 7472 9029
rect 7508 9003 7534 9029
rect 12074 9003 12100 9029
rect 12136 9003 12162 9029
rect 12198 9003 12224 9029
rect 12260 9003 12286 9029
rect 12322 9003 12348 9029
rect 12384 9003 12410 9029
rect 12446 9003 12472 9029
rect 12508 9003 12534 9029
rect 17074 9003 17100 9029
rect 17136 9003 17162 9029
rect 17198 9003 17224 9029
rect 17260 9003 17286 9029
rect 17322 9003 17348 9029
rect 17384 9003 17410 9029
rect 17446 9003 17472 9029
rect 17508 9003 17534 9029
rect 22074 9003 22100 9029
rect 22136 9003 22162 9029
rect 22198 9003 22224 9029
rect 22260 9003 22286 9029
rect 22322 9003 22348 9029
rect 22384 9003 22410 9029
rect 22446 9003 22472 9029
rect 22508 9003 22534 9029
rect 27074 9003 27100 9029
rect 27136 9003 27162 9029
rect 27198 9003 27224 9029
rect 27260 9003 27286 9029
rect 27322 9003 27348 9029
rect 27384 9003 27410 9029
rect 27446 9003 27472 9029
rect 27508 9003 27534 9029
rect 32074 9003 32100 9029
rect 32136 9003 32162 9029
rect 32198 9003 32224 9029
rect 32260 9003 32286 9029
rect 32322 9003 32348 9029
rect 32384 9003 32410 9029
rect 32446 9003 32472 9029
rect 32508 9003 32534 9029
rect 37074 9003 37100 9029
rect 37136 9003 37162 9029
rect 37198 9003 37224 9029
rect 37260 9003 37286 9029
rect 37322 9003 37348 9029
rect 37384 9003 37410 9029
rect 37446 9003 37472 9029
rect 37508 9003 37534 9029
rect 1415 8807 1441 8833
rect 2479 8807 2505 8833
rect 3823 8807 3849 8833
rect 4999 8807 5025 8833
rect 5559 8807 5585 8833
rect 6455 8807 6481 8833
rect 7799 8807 7825 8833
rect 8751 8807 8777 8833
rect 9255 8807 9281 8833
rect 10319 8807 10345 8833
rect 11607 8807 11633 8833
rect 12055 8807 12081 8833
rect 12279 8807 12305 8833
rect 13063 8807 13089 8833
rect 13511 8807 13537 8833
rect 13735 8807 13761 8833
rect 14799 8807 14825 8833
rect 15247 8807 15273 8833
rect 15471 8807 15497 8833
rect 16255 8807 16281 8833
rect 16815 8807 16841 8833
rect 16927 8807 16953 8833
rect 18775 8807 18801 8833
rect 19335 8807 19361 8833
rect 19447 8807 19473 8833
rect 20231 8807 20257 8833
rect 21407 8807 21433 8833
rect 22751 8807 22777 8833
rect 23871 8807 23897 8833
rect 24487 8807 24513 8833
rect 25383 8807 25409 8833
rect 27735 8807 27761 8833
rect 28855 8807 28881 8833
rect 29415 8807 29441 8833
rect 30199 8807 30225 8833
rect 30983 8807 31009 8833
rect 31151 8807 31177 8833
rect 31375 8807 31401 8833
rect 32159 8807 32185 8833
rect 32831 8807 32857 8833
rect 34679 8807 34705 8833
rect 35855 8807 35881 8833
rect 36415 8807 36441 8833
rect 37311 8807 37337 8833
rect 1415 8751 1441 8777
rect 3823 8751 3849 8777
rect 6455 8751 6481 8777
rect 8751 8751 8777 8777
rect 10319 8751 10345 8777
rect 21407 8751 21433 8777
rect 23871 8751 23897 8777
rect 25383 8751 25409 8777
rect 27735 8751 27761 8777
rect 30199 8751 30225 8777
rect 33111 8751 33137 8777
rect 35855 8751 35881 8777
rect 37311 8751 37337 8777
rect 4574 8611 4600 8637
rect 4636 8611 4662 8637
rect 4698 8611 4724 8637
rect 4760 8611 4786 8637
rect 4822 8611 4848 8637
rect 4884 8611 4910 8637
rect 4946 8611 4972 8637
rect 5008 8611 5034 8637
rect 9574 8611 9600 8637
rect 9636 8611 9662 8637
rect 9698 8611 9724 8637
rect 9760 8611 9786 8637
rect 9822 8611 9848 8637
rect 9884 8611 9910 8637
rect 9946 8611 9972 8637
rect 10008 8611 10034 8637
rect 14574 8611 14600 8637
rect 14636 8611 14662 8637
rect 14698 8611 14724 8637
rect 14760 8611 14786 8637
rect 14822 8611 14848 8637
rect 14884 8611 14910 8637
rect 14946 8611 14972 8637
rect 15008 8611 15034 8637
rect 19574 8611 19600 8637
rect 19636 8611 19662 8637
rect 19698 8611 19724 8637
rect 19760 8611 19786 8637
rect 19822 8611 19848 8637
rect 19884 8611 19910 8637
rect 19946 8611 19972 8637
rect 20008 8611 20034 8637
rect 24574 8611 24600 8637
rect 24636 8611 24662 8637
rect 24698 8611 24724 8637
rect 24760 8611 24786 8637
rect 24822 8611 24848 8637
rect 24884 8611 24910 8637
rect 24946 8611 24972 8637
rect 25008 8611 25034 8637
rect 29574 8611 29600 8637
rect 29636 8611 29662 8637
rect 29698 8611 29724 8637
rect 29760 8611 29786 8637
rect 29822 8611 29848 8637
rect 29884 8611 29910 8637
rect 29946 8611 29972 8637
rect 30008 8611 30034 8637
rect 34574 8611 34600 8637
rect 34636 8611 34662 8637
rect 34698 8611 34724 8637
rect 34760 8611 34786 8637
rect 34822 8611 34848 8637
rect 34884 8611 34910 8637
rect 34946 8611 34972 8637
rect 35008 8611 35034 8637
rect 1863 8471 1889 8497
rect 4495 8471 4521 8497
rect 8415 8471 8441 8497
rect 17991 8471 18017 8497
rect 19447 8471 19473 8497
rect 21799 8471 21825 8497
rect 23423 8471 23449 8497
rect 25943 8471 25969 8497
rect 27399 8471 27425 8497
rect 35351 8471 35377 8497
rect 37647 8471 37673 8497
rect 1863 8415 1889 8441
rect 3039 8415 3065 8441
rect 3599 8415 3625 8441
rect 4495 8415 4521 8441
rect 6119 8415 6145 8441
rect 6399 8415 6425 8441
rect 6511 8415 6537 8441
rect 7575 8415 7601 8441
rect 8415 8415 8441 8441
rect 9815 8415 9841 8441
rect 10319 8415 10345 8441
rect 10487 8415 10513 8441
rect 11439 8415 11465 8441
rect 11775 8415 11801 8441
rect 11943 8415 11969 8441
rect 13007 8415 13033 8441
rect 13455 8415 13481 8441
rect 13679 8415 13705 8441
rect 14463 8415 14489 8441
rect 15023 8415 15049 8441
rect 15135 8415 15161 8441
rect 16815 8415 16841 8441
rect 17991 8415 18017 8441
rect 18271 8415 18297 8441
rect 19447 8415 19473 8441
rect 20791 8415 20817 8441
rect 21799 8415 21825 8441
rect 22527 8415 22553 8441
rect 23423 8415 23449 8441
rect 24767 8415 24793 8441
rect 25943 8415 25969 8441
rect 26223 8415 26249 8441
rect 27399 8415 27425 8441
rect 29415 8415 29441 8441
rect 29863 8415 29889 8441
rect 30087 8415 30113 8441
rect 31039 8415 31065 8441
rect 31319 8415 31345 8441
rect 31431 8415 31457 8441
rect 32719 8415 32745 8441
rect 33167 8415 33193 8441
rect 33615 8415 33641 8441
rect 34175 8415 34201 8441
rect 35351 8415 35377 8441
rect 36695 8415 36721 8441
rect 37647 8415 37673 8441
rect 2074 8219 2100 8245
rect 2136 8219 2162 8245
rect 2198 8219 2224 8245
rect 2260 8219 2286 8245
rect 2322 8219 2348 8245
rect 2384 8219 2410 8245
rect 2446 8219 2472 8245
rect 2508 8219 2534 8245
rect 7074 8219 7100 8245
rect 7136 8219 7162 8245
rect 7198 8219 7224 8245
rect 7260 8219 7286 8245
rect 7322 8219 7348 8245
rect 7384 8219 7410 8245
rect 7446 8219 7472 8245
rect 7508 8219 7534 8245
rect 12074 8219 12100 8245
rect 12136 8219 12162 8245
rect 12198 8219 12224 8245
rect 12260 8219 12286 8245
rect 12322 8219 12348 8245
rect 12384 8219 12410 8245
rect 12446 8219 12472 8245
rect 12508 8219 12534 8245
rect 17074 8219 17100 8245
rect 17136 8219 17162 8245
rect 17198 8219 17224 8245
rect 17260 8219 17286 8245
rect 17322 8219 17348 8245
rect 17384 8219 17410 8245
rect 17446 8219 17472 8245
rect 17508 8219 17534 8245
rect 22074 8219 22100 8245
rect 22136 8219 22162 8245
rect 22198 8219 22224 8245
rect 22260 8219 22286 8245
rect 22322 8219 22348 8245
rect 22384 8219 22410 8245
rect 22446 8219 22472 8245
rect 22508 8219 22534 8245
rect 27074 8219 27100 8245
rect 27136 8219 27162 8245
rect 27198 8219 27224 8245
rect 27260 8219 27286 8245
rect 27322 8219 27348 8245
rect 27384 8219 27410 8245
rect 27446 8219 27472 8245
rect 27508 8219 27534 8245
rect 32074 8219 32100 8245
rect 32136 8219 32162 8245
rect 32198 8219 32224 8245
rect 32260 8219 32286 8245
rect 32322 8219 32348 8245
rect 32384 8219 32410 8245
rect 32446 8219 32472 8245
rect 32508 8219 32534 8245
rect 37074 8219 37100 8245
rect 37136 8219 37162 8245
rect 37198 8219 37224 8245
rect 37260 8219 37286 8245
rect 37322 8219 37348 8245
rect 37384 8219 37410 8245
rect 37446 8219 37472 8245
rect 37508 8219 37534 8245
rect 1807 8023 1833 8049
rect 2479 8023 2505 8049
rect 4103 8023 4129 8049
rect 4383 8023 4409 8049
rect 4495 8023 4521 8049
rect 5559 8023 5585 8049
rect 6455 8023 6481 8049
rect 7799 8023 7825 8049
rect 8751 8023 8777 8049
rect 9255 8023 9281 8049
rect 10431 8023 10457 8049
rect 11439 8023 11465 8049
rect 11775 8023 11801 8049
rect 11887 8023 11913 8049
rect 12895 8023 12921 8049
rect 13455 8023 13481 8049
rect 13567 8023 13593 8049
rect 14967 8023 14993 8049
rect 15751 8023 15777 8049
rect 16255 8023 16281 8049
rect 16815 8023 16841 8049
rect 16927 8023 16953 8049
rect 18775 8023 18801 8049
rect 19951 8023 19977 8049
rect 20231 8023 20257 8049
rect 21407 8023 21433 8049
rect 22751 8023 22777 8049
rect 23871 8023 23897 8049
rect 24487 8023 24513 8049
rect 25159 8023 25185 8049
rect 26727 8023 26753 8049
rect 27679 8023 27705 8049
rect 29359 8023 29385 8049
rect 29863 8023 29889 8049
rect 30759 8023 30785 8049
rect 31151 8023 31177 8049
rect 31375 8023 31401 8049
rect 32439 8023 32465 8049
rect 33167 8023 33193 8049
rect 33615 8023 33641 8049
rect 33727 8023 33753 8049
rect 34679 8023 34705 8049
rect 35855 8023 35881 8049
rect 36135 8023 36161 8049
rect 36975 8023 37001 8049
rect 1527 7967 1553 7993
rect 6455 7967 6481 7993
rect 8751 7967 8777 7993
rect 10431 7967 10457 7993
rect 15751 7967 15777 7993
rect 19951 7967 19977 7993
rect 21407 7967 21433 7993
rect 23871 7967 23897 7993
rect 25159 7967 25185 7993
rect 27679 7967 27705 7993
rect 30087 7967 30113 7993
rect 33167 7967 33193 7993
rect 33895 7967 33921 7993
rect 35855 7967 35881 7993
rect 37087 7967 37113 7993
rect 4574 7827 4600 7853
rect 4636 7827 4662 7853
rect 4698 7827 4724 7853
rect 4760 7827 4786 7853
rect 4822 7827 4848 7853
rect 4884 7827 4910 7853
rect 4946 7827 4972 7853
rect 5008 7827 5034 7853
rect 9574 7827 9600 7853
rect 9636 7827 9662 7853
rect 9698 7827 9724 7853
rect 9760 7827 9786 7853
rect 9822 7827 9848 7853
rect 9884 7827 9910 7853
rect 9946 7827 9972 7853
rect 10008 7827 10034 7853
rect 14574 7827 14600 7853
rect 14636 7827 14662 7853
rect 14698 7827 14724 7853
rect 14760 7827 14786 7853
rect 14822 7827 14848 7853
rect 14884 7827 14910 7853
rect 14946 7827 14972 7853
rect 15008 7827 15034 7853
rect 19574 7827 19600 7853
rect 19636 7827 19662 7853
rect 19698 7827 19724 7853
rect 19760 7827 19786 7853
rect 19822 7827 19848 7853
rect 19884 7827 19910 7853
rect 19946 7827 19972 7853
rect 20008 7827 20034 7853
rect 24574 7827 24600 7853
rect 24636 7827 24662 7853
rect 24698 7827 24724 7853
rect 24760 7827 24786 7853
rect 24822 7827 24848 7853
rect 24884 7827 24910 7853
rect 24946 7827 24972 7853
rect 25008 7827 25034 7853
rect 29574 7827 29600 7853
rect 29636 7827 29662 7853
rect 29698 7827 29724 7853
rect 29760 7827 29786 7853
rect 29822 7827 29848 7853
rect 29884 7827 29910 7853
rect 29946 7827 29972 7853
rect 30008 7827 30034 7853
rect 34574 7827 34600 7853
rect 34636 7827 34662 7853
rect 34698 7827 34724 7853
rect 34760 7827 34786 7853
rect 34822 7827 34848 7853
rect 34884 7827 34910 7853
rect 34946 7827 34972 7853
rect 35008 7827 35034 7853
rect 1863 7687 1889 7713
rect 4495 7687 4521 7713
rect 15247 7687 15273 7713
rect 18383 7687 18409 7713
rect 20007 7687 20033 7713
rect 21799 7687 21825 7713
rect 23423 7687 23449 7713
rect 25943 7687 25969 7713
rect 27399 7687 27425 7713
rect 30199 7687 30225 7713
rect 35239 7687 35265 7713
rect 1863 7631 1889 7657
rect 3039 7631 3065 7657
rect 3599 7631 3625 7657
rect 4495 7631 4521 7657
rect 6119 7631 6145 7657
rect 6399 7631 6425 7657
rect 6511 7631 6537 7657
rect 7295 7631 7321 7657
rect 7743 7631 7769 7657
rect 7967 7631 7993 7657
rect 10039 7631 10065 7657
rect 10207 7631 10233 7657
rect 10431 7631 10457 7657
rect 11439 7631 11465 7657
rect 11775 7631 11801 7657
rect 11887 7631 11913 7657
rect 12839 7631 12865 7657
rect 13399 7631 13425 7657
rect 13511 7631 13537 7657
rect 14407 7631 14433 7657
rect 15247 7631 15273 7657
rect 17599 7631 17625 7657
rect 18383 7631 18409 7657
rect 19111 7631 19137 7657
rect 20007 7631 20033 7657
rect 20959 7631 20985 7657
rect 21799 7631 21825 7657
rect 22527 7631 22553 7657
rect 23423 7631 23449 7657
rect 24823 7631 24849 7657
rect 25943 7631 25969 7657
rect 26223 7631 26249 7657
rect 27399 7631 27425 7657
rect 29359 7631 29385 7657
rect 30199 7631 30225 7657
rect 30759 7631 30785 7657
rect 31207 7631 31233 7657
rect 31375 7631 31401 7657
rect 32999 7631 33025 7657
rect 33167 7631 33193 7657
rect 33391 7631 33417 7657
rect 34399 7631 34425 7657
rect 35239 7631 35265 7657
rect 36695 7631 36721 7657
rect 37143 7631 37169 7657
rect 37367 7631 37393 7657
rect 2074 7435 2100 7461
rect 2136 7435 2162 7461
rect 2198 7435 2224 7461
rect 2260 7435 2286 7461
rect 2322 7435 2348 7461
rect 2384 7435 2410 7461
rect 2446 7435 2472 7461
rect 2508 7435 2534 7461
rect 7074 7435 7100 7461
rect 7136 7435 7162 7461
rect 7198 7435 7224 7461
rect 7260 7435 7286 7461
rect 7322 7435 7348 7461
rect 7384 7435 7410 7461
rect 7446 7435 7472 7461
rect 7508 7435 7534 7461
rect 12074 7435 12100 7461
rect 12136 7435 12162 7461
rect 12198 7435 12224 7461
rect 12260 7435 12286 7461
rect 12322 7435 12348 7461
rect 12384 7435 12410 7461
rect 12446 7435 12472 7461
rect 12508 7435 12534 7461
rect 17074 7435 17100 7461
rect 17136 7435 17162 7461
rect 17198 7435 17224 7461
rect 17260 7435 17286 7461
rect 17322 7435 17348 7461
rect 17384 7435 17410 7461
rect 17446 7435 17472 7461
rect 17508 7435 17534 7461
rect 22074 7435 22100 7461
rect 22136 7435 22162 7461
rect 22198 7435 22224 7461
rect 22260 7435 22286 7461
rect 22322 7435 22348 7461
rect 22384 7435 22410 7461
rect 22446 7435 22472 7461
rect 22508 7435 22534 7461
rect 27074 7435 27100 7461
rect 27136 7435 27162 7461
rect 27198 7435 27224 7461
rect 27260 7435 27286 7461
rect 27322 7435 27348 7461
rect 27384 7435 27410 7461
rect 27446 7435 27472 7461
rect 27508 7435 27534 7461
rect 32074 7435 32100 7461
rect 32136 7435 32162 7461
rect 32198 7435 32224 7461
rect 32260 7435 32286 7461
rect 32322 7435 32348 7461
rect 32384 7435 32410 7461
rect 32446 7435 32472 7461
rect 32508 7435 32534 7461
rect 37074 7435 37100 7461
rect 37136 7435 37162 7461
rect 37198 7435 37224 7461
rect 37260 7435 37286 7461
rect 37322 7435 37348 7461
rect 37384 7435 37410 7461
rect 37446 7435 37472 7461
rect 37508 7435 37534 7461
rect 1807 7239 1833 7265
rect 2479 7239 2505 7265
rect 4103 7239 4129 7265
rect 4999 7239 5025 7265
rect 5559 7239 5585 7265
rect 6455 7239 6481 7265
rect 7799 7239 7825 7265
rect 8247 7239 8273 7265
rect 8471 7239 8497 7265
rect 9479 7239 9505 7265
rect 10151 7239 10177 7265
rect 11439 7239 11465 7265
rect 11775 7239 11801 7265
rect 11887 7239 11913 7265
rect 12783 7239 12809 7265
rect 13119 7239 13145 7265
rect 13455 7239 13481 7265
rect 15079 7239 15105 7265
rect 15247 7239 15273 7265
rect 15471 7239 15497 7265
rect 17487 7239 17513 7265
rect 18383 7239 18409 7265
rect 19055 7239 19081 7265
rect 19951 7239 19977 7265
rect 20511 7239 20537 7265
rect 21351 7239 21377 7265
rect 22751 7239 22777 7265
rect 23535 7239 23561 7265
rect 24375 7239 24401 7265
rect 24655 7239 24681 7265
rect 24879 7239 24905 7265
rect 27679 7239 27705 7265
rect 28855 7239 28881 7265
rect 29359 7239 29385 7265
rect 30199 7239 30225 7265
rect 30927 7239 30953 7265
rect 31599 7239 31625 7265
rect 32439 7239 32465 7265
rect 33335 7239 33361 7265
rect 33783 7239 33809 7265
rect 34959 7239 34985 7265
rect 35799 7239 35825 7265
rect 36135 7239 36161 7265
rect 37311 7239 37337 7265
rect 1527 7183 1553 7209
rect 4999 7183 5025 7209
rect 6455 7183 6481 7209
rect 10207 7183 10233 7209
rect 18383 7183 18409 7209
rect 19951 7183 19977 7209
rect 21351 7183 21377 7209
rect 23703 7183 23729 7209
rect 27679 7183 27705 7209
rect 30199 7183 30225 7209
rect 31655 7183 31681 7209
rect 33335 7183 33361 7209
rect 33615 7183 33641 7209
rect 33895 7183 33921 7209
rect 35799 7183 35825 7209
rect 37311 7183 37337 7209
rect 4574 7043 4600 7069
rect 4636 7043 4662 7069
rect 4698 7043 4724 7069
rect 4760 7043 4786 7069
rect 4822 7043 4848 7069
rect 4884 7043 4910 7069
rect 4946 7043 4972 7069
rect 5008 7043 5034 7069
rect 9574 7043 9600 7069
rect 9636 7043 9662 7069
rect 9698 7043 9724 7069
rect 9760 7043 9786 7069
rect 9822 7043 9848 7069
rect 9884 7043 9910 7069
rect 9946 7043 9972 7069
rect 10008 7043 10034 7069
rect 14574 7043 14600 7069
rect 14636 7043 14662 7069
rect 14698 7043 14724 7069
rect 14760 7043 14786 7069
rect 14822 7043 14848 7069
rect 14884 7043 14910 7069
rect 14946 7043 14972 7069
rect 15008 7043 15034 7069
rect 19574 7043 19600 7069
rect 19636 7043 19662 7069
rect 19698 7043 19724 7069
rect 19760 7043 19786 7069
rect 19822 7043 19848 7069
rect 19884 7043 19910 7069
rect 19946 7043 19972 7069
rect 20008 7043 20034 7069
rect 24574 7043 24600 7069
rect 24636 7043 24662 7069
rect 24698 7043 24724 7069
rect 24760 7043 24786 7069
rect 24822 7043 24848 7069
rect 24884 7043 24910 7069
rect 24946 7043 24972 7069
rect 25008 7043 25034 7069
rect 29574 7043 29600 7069
rect 29636 7043 29662 7069
rect 29698 7043 29724 7069
rect 29760 7043 29786 7069
rect 29822 7043 29848 7069
rect 29884 7043 29910 7069
rect 29946 7043 29972 7069
rect 30008 7043 30034 7069
rect 34574 7043 34600 7069
rect 34636 7043 34662 7069
rect 34698 7043 34724 7069
rect 34760 7043 34786 7069
rect 34822 7043 34848 7069
rect 34884 7043 34910 7069
rect 34946 7043 34972 7069
rect 35008 7043 35034 7069
rect 1863 6903 1889 6929
rect 6959 6903 6985 6929
rect 8247 6903 8273 6929
rect 15247 6903 15273 6929
rect 18439 6903 18465 6929
rect 20007 6903 20033 6929
rect 21743 6903 21769 6929
rect 23199 6903 23225 6929
rect 30199 6903 30225 6929
rect 31599 6903 31625 6929
rect 33895 6903 33921 6929
rect 35295 6903 35321 6929
rect 37647 6903 37673 6929
rect 1863 6847 1889 6873
rect 3039 6847 3065 6873
rect 3599 6847 3625 6873
rect 3823 6847 3849 6873
rect 3991 6847 4017 6873
rect 6007 6847 6033 6873
rect 6959 6847 6985 6873
rect 7519 6847 7545 6873
rect 8247 6847 8273 6873
rect 9703 6847 9729 6873
rect 10207 6847 10233 6873
rect 10375 6847 10401 6873
rect 11439 6847 11465 6873
rect 11719 6847 11745 6873
rect 11831 6847 11857 6873
rect 13119 6847 13145 6873
rect 13399 6847 13425 6873
rect 13511 6847 13537 6873
rect 14407 6847 14433 6873
rect 15135 6847 15161 6873
rect 17599 6847 17625 6873
rect 18439 6847 18465 6873
rect 19111 6847 19137 6873
rect 20007 6847 20033 6873
rect 20959 6847 20985 6873
rect 21743 6847 21769 6873
rect 22527 6847 22553 6873
rect 23199 6847 23225 6873
rect 24767 6847 24793 6873
rect 25215 6847 25241 6873
rect 25439 6847 25465 6873
rect 27567 6847 27593 6873
rect 27791 6847 27817 6873
rect 28351 6847 28377 6873
rect 29359 6847 29385 6873
rect 30199 6847 30225 6873
rect 30927 6847 30953 6873
rect 31599 6847 31625 6873
rect 32999 6847 33025 6873
rect 33895 6847 33921 6873
rect 34399 6847 34425 6873
rect 35295 6847 35321 6873
rect 35687 6847 35713 6873
rect 35799 6847 35825 6873
rect 35911 6847 35937 6873
rect 36695 6847 36721 6873
rect 37647 6847 37673 6873
rect 2074 6651 2100 6677
rect 2136 6651 2162 6677
rect 2198 6651 2224 6677
rect 2260 6651 2286 6677
rect 2322 6651 2348 6677
rect 2384 6651 2410 6677
rect 2446 6651 2472 6677
rect 2508 6651 2534 6677
rect 7074 6651 7100 6677
rect 7136 6651 7162 6677
rect 7198 6651 7224 6677
rect 7260 6651 7286 6677
rect 7322 6651 7348 6677
rect 7384 6651 7410 6677
rect 7446 6651 7472 6677
rect 7508 6651 7534 6677
rect 12074 6651 12100 6677
rect 12136 6651 12162 6677
rect 12198 6651 12224 6677
rect 12260 6651 12286 6677
rect 12322 6651 12348 6677
rect 12384 6651 12410 6677
rect 12446 6651 12472 6677
rect 12508 6651 12534 6677
rect 17074 6651 17100 6677
rect 17136 6651 17162 6677
rect 17198 6651 17224 6677
rect 17260 6651 17286 6677
rect 17322 6651 17348 6677
rect 17384 6651 17410 6677
rect 17446 6651 17472 6677
rect 17508 6651 17534 6677
rect 22074 6651 22100 6677
rect 22136 6651 22162 6677
rect 22198 6651 22224 6677
rect 22260 6651 22286 6677
rect 22322 6651 22348 6677
rect 22384 6651 22410 6677
rect 22446 6651 22472 6677
rect 22508 6651 22534 6677
rect 27074 6651 27100 6677
rect 27136 6651 27162 6677
rect 27198 6651 27224 6677
rect 27260 6651 27286 6677
rect 27322 6651 27348 6677
rect 27384 6651 27410 6677
rect 27446 6651 27472 6677
rect 27508 6651 27534 6677
rect 32074 6651 32100 6677
rect 32136 6651 32162 6677
rect 32198 6651 32224 6677
rect 32260 6651 32286 6677
rect 32322 6651 32348 6677
rect 32384 6651 32410 6677
rect 32446 6651 32472 6677
rect 32508 6651 32534 6677
rect 37074 6651 37100 6677
rect 37136 6651 37162 6677
rect 37198 6651 37224 6677
rect 37260 6651 37286 6677
rect 37322 6651 37348 6677
rect 37384 6651 37410 6677
rect 37446 6651 37472 6677
rect 37508 6651 37534 6677
rect 1807 6455 1833 6481
rect 2199 6455 2225 6481
rect 4103 6455 4129 6481
rect 4271 6455 4297 6481
rect 4495 6455 4521 6481
rect 5559 6455 5585 6481
rect 6455 6455 6481 6481
rect 8079 6455 8105 6481
rect 8247 6455 8273 6481
rect 8471 6455 8497 6481
rect 9479 6455 9505 6481
rect 10375 6455 10401 6481
rect 11495 6455 11521 6481
rect 11999 6455 12025 6481
rect 12167 6455 12193 6481
rect 13119 6455 13145 6481
rect 13455 6455 13481 6481
rect 13623 6455 13649 6481
rect 15751 6455 15777 6481
rect 16759 6455 16785 6481
rect 17487 6455 17513 6481
rect 18383 6455 18409 6481
rect 19055 6455 19081 6481
rect 19951 6455 19977 6481
rect 20511 6455 20537 6481
rect 21407 6455 21433 6481
rect 23031 6455 23057 6481
rect 23199 6455 23225 6481
rect 23535 6455 23561 6481
rect 24487 6455 24513 6481
rect 25159 6455 25185 6481
rect 27847 6455 27873 6481
rect 28855 6455 28881 6481
rect 29359 6455 29385 6481
rect 30199 6455 30225 6481
rect 30983 6455 31009 6481
rect 31823 6455 31849 6481
rect 32439 6455 32465 6481
rect 33335 6455 33361 6481
rect 33671 6455 33697 6481
rect 33727 6455 33753 6481
rect 33895 6455 33921 6481
rect 34679 6455 34705 6481
rect 35631 6455 35657 6481
rect 36415 6455 36441 6481
rect 37255 6455 37281 6481
rect 1527 6399 1553 6425
rect 6455 6399 6481 6425
rect 10375 6399 10401 6425
rect 16759 6399 16785 6425
rect 18383 6399 18409 6425
rect 19951 6399 19977 6425
rect 21407 6399 21433 6425
rect 25159 6399 25185 6425
rect 27847 6399 27873 6425
rect 30199 6399 30225 6425
rect 31823 6399 31849 6425
rect 33335 6399 33361 6425
rect 35631 6399 35657 6425
rect 37255 6399 37281 6425
rect 4574 6259 4600 6285
rect 4636 6259 4662 6285
rect 4698 6259 4724 6285
rect 4760 6259 4786 6285
rect 4822 6259 4848 6285
rect 4884 6259 4910 6285
rect 4946 6259 4972 6285
rect 5008 6259 5034 6285
rect 9574 6259 9600 6285
rect 9636 6259 9662 6285
rect 9698 6259 9724 6285
rect 9760 6259 9786 6285
rect 9822 6259 9848 6285
rect 9884 6259 9910 6285
rect 9946 6259 9972 6285
rect 10008 6259 10034 6285
rect 14574 6259 14600 6285
rect 14636 6259 14662 6285
rect 14698 6259 14724 6285
rect 14760 6259 14786 6285
rect 14822 6259 14848 6285
rect 14884 6259 14910 6285
rect 14946 6259 14972 6285
rect 15008 6259 15034 6285
rect 19574 6259 19600 6285
rect 19636 6259 19662 6285
rect 19698 6259 19724 6285
rect 19760 6259 19786 6285
rect 19822 6259 19848 6285
rect 19884 6259 19910 6285
rect 19946 6259 19972 6285
rect 20008 6259 20034 6285
rect 24574 6259 24600 6285
rect 24636 6259 24662 6285
rect 24698 6259 24724 6285
rect 24760 6259 24786 6285
rect 24822 6259 24848 6285
rect 24884 6259 24910 6285
rect 24946 6259 24972 6285
rect 25008 6259 25034 6285
rect 29574 6259 29600 6285
rect 29636 6259 29662 6285
rect 29698 6259 29724 6285
rect 29760 6259 29786 6285
rect 29822 6259 29848 6285
rect 29884 6259 29910 6285
rect 29946 6259 29972 6285
rect 30008 6259 30034 6285
rect 34574 6259 34600 6285
rect 34636 6259 34662 6285
rect 34698 6259 34724 6285
rect 34760 6259 34786 6285
rect 34822 6259 34848 6285
rect 34884 6259 34910 6285
rect 34946 6259 34972 6285
rect 35008 6259 35034 6285
rect 1863 6119 1889 6145
rect 8247 6119 8273 6145
rect 16423 6119 16449 6145
rect 18439 6119 18465 6145
rect 20007 6119 20033 6145
rect 21799 6119 21825 6145
rect 23423 6119 23449 6145
rect 27399 6119 27425 6145
rect 30199 6119 30225 6145
rect 31823 6119 31849 6145
rect 35351 6119 35377 6145
rect 1863 6063 1889 6089
rect 2759 6063 2785 6089
rect 3599 6063 3625 6089
rect 3879 6063 3905 6089
rect 3991 6063 4017 6089
rect 6007 6063 6033 6089
rect 6399 6063 6425 6089
rect 6511 6063 6537 6089
rect 7575 6063 7601 6089
rect 8247 6063 8273 6089
rect 10039 6063 10065 6089
rect 10375 6063 10401 6089
rect 10487 6063 10513 6089
rect 11551 6063 11577 6089
rect 11831 6063 11857 6089
rect 11943 6063 11969 6089
rect 13119 6063 13145 6089
rect 13287 6063 13313 6089
rect 13511 6063 13537 6089
rect 15527 6063 15553 6089
rect 16423 6063 16449 6089
rect 17599 6063 17625 6089
rect 18439 6063 18465 6089
rect 19111 6063 19137 6089
rect 20007 6063 20033 6089
rect 20791 6063 20817 6089
rect 21799 6063 21825 6089
rect 22527 6063 22553 6089
rect 23423 6063 23449 6089
rect 25047 6063 25073 6089
rect 25215 6063 25241 6089
rect 25439 6063 25465 6089
rect 26223 6063 26249 6089
rect 27399 6063 27425 6089
rect 29359 6063 29385 6089
rect 30199 6063 30225 6089
rect 30927 6063 30953 6089
rect 31823 6063 31849 6089
rect 32719 6063 32745 6089
rect 33279 6063 33305 6089
rect 33391 6063 33417 6089
rect 34455 6063 34481 6089
rect 35351 6063 35377 6089
rect 35631 6063 35657 6089
rect 35743 6063 35769 6089
rect 35911 6063 35937 6089
rect 36695 6063 36721 6089
rect 37255 6063 37281 6089
rect 37367 6063 37393 6089
rect 2074 5867 2100 5893
rect 2136 5867 2162 5893
rect 2198 5867 2224 5893
rect 2260 5867 2286 5893
rect 2322 5867 2348 5893
rect 2384 5867 2410 5893
rect 2446 5867 2472 5893
rect 2508 5867 2534 5893
rect 7074 5867 7100 5893
rect 7136 5867 7162 5893
rect 7198 5867 7224 5893
rect 7260 5867 7286 5893
rect 7322 5867 7348 5893
rect 7384 5867 7410 5893
rect 7446 5867 7472 5893
rect 7508 5867 7534 5893
rect 12074 5867 12100 5893
rect 12136 5867 12162 5893
rect 12198 5867 12224 5893
rect 12260 5867 12286 5893
rect 12322 5867 12348 5893
rect 12384 5867 12410 5893
rect 12446 5867 12472 5893
rect 12508 5867 12534 5893
rect 17074 5867 17100 5893
rect 17136 5867 17162 5893
rect 17198 5867 17224 5893
rect 17260 5867 17286 5893
rect 17322 5867 17348 5893
rect 17384 5867 17410 5893
rect 17446 5867 17472 5893
rect 17508 5867 17534 5893
rect 22074 5867 22100 5893
rect 22136 5867 22162 5893
rect 22198 5867 22224 5893
rect 22260 5867 22286 5893
rect 22322 5867 22348 5893
rect 22384 5867 22410 5893
rect 22446 5867 22472 5893
rect 22508 5867 22534 5893
rect 27074 5867 27100 5893
rect 27136 5867 27162 5893
rect 27198 5867 27224 5893
rect 27260 5867 27286 5893
rect 27322 5867 27348 5893
rect 27384 5867 27410 5893
rect 27446 5867 27472 5893
rect 27508 5867 27534 5893
rect 32074 5867 32100 5893
rect 32136 5867 32162 5893
rect 32198 5867 32224 5893
rect 32260 5867 32286 5893
rect 32322 5867 32348 5893
rect 32384 5867 32410 5893
rect 32446 5867 32472 5893
rect 32508 5867 32534 5893
rect 37074 5867 37100 5893
rect 37136 5867 37162 5893
rect 37198 5867 37224 5893
rect 37260 5867 37286 5893
rect 37322 5867 37348 5893
rect 37384 5867 37410 5893
rect 37446 5867 37472 5893
rect 37508 5867 37534 5893
rect 1807 5671 1833 5697
rect 1919 5671 1945 5697
rect 2479 5671 2505 5697
rect 4103 5671 4129 5697
rect 4383 5671 4409 5697
rect 4495 5671 4521 5697
rect 5559 5671 5585 5697
rect 6455 5671 6481 5697
rect 8079 5671 8105 5697
rect 8975 5671 9001 5697
rect 9535 5671 9561 5697
rect 10431 5671 10457 5697
rect 12335 5671 12361 5697
rect 12503 5671 12529 5697
rect 12727 5671 12753 5697
rect 15751 5671 15777 5697
rect 16759 5671 16785 5697
rect 17487 5671 17513 5697
rect 18383 5671 18409 5697
rect 19055 5671 19081 5697
rect 19951 5671 19977 5697
rect 20511 5671 20537 5697
rect 21351 5671 21377 5697
rect 23031 5671 23057 5697
rect 23871 5671 23897 5697
rect 24431 5671 24457 5697
rect 25159 5671 25185 5697
rect 26895 5671 26921 5697
rect 27623 5671 27649 5697
rect 29359 5671 29385 5697
rect 30199 5671 30225 5697
rect 30983 5671 31009 5697
rect 31879 5671 31905 5697
rect 32439 5671 32465 5697
rect 33335 5671 33361 5697
rect 33671 5671 33697 5697
rect 33895 5671 33921 5697
rect 34679 5671 34705 5697
rect 35239 5671 35265 5697
rect 35351 5671 35377 5697
rect 36135 5671 36161 5697
rect 37311 5671 37337 5697
rect 6455 5615 6481 5641
rect 8975 5615 9001 5641
rect 10431 5615 10457 5641
rect 16759 5615 16785 5641
rect 18383 5615 18409 5641
rect 19951 5615 19977 5641
rect 21351 5615 21377 5641
rect 23871 5615 23897 5641
rect 25159 5615 25185 5641
rect 27679 5615 27705 5641
rect 30199 5615 30225 5641
rect 31879 5615 31905 5641
rect 33335 5615 33361 5641
rect 33727 5615 33753 5641
rect 37311 5615 37337 5641
rect 37591 5615 37617 5641
rect 37703 5615 37729 5641
rect 37871 5615 37897 5641
rect 4574 5475 4600 5501
rect 4636 5475 4662 5501
rect 4698 5475 4724 5501
rect 4760 5475 4786 5501
rect 4822 5475 4848 5501
rect 4884 5475 4910 5501
rect 4946 5475 4972 5501
rect 5008 5475 5034 5501
rect 9574 5475 9600 5501
rect 9636 5475 9662 5501
rect 9698 5475 9724 5501
rect 9760 5475 9786 5501
rect 9822 5475 9848 5501
rect 9884 5475 9910 5501
rect 9946 5475 9972 5501
rect 10008 5475 10034 5501
rect 14574 5475 14600 5501
rect 14636 5475 14662 5501
rect 14698 5475 14724 5501
rect 14760 5475 14786 5501
rect 14822 5475 14848 5501
rect 14884 5475 14910 5501
rect 14946 5475 14972 5501
rect 15008 5475 15034 5501
rect 19574 5475 19600 5501
rect 19636 5475 19662 5501
rect 19698 5475 19724 5501
rect 19760 5475 19786 5501
rect 19822 5475 19848 5501
rect 19884 5475 19910 5501
rect 19946 5475 19972 5501
rect 20008 5475 20034 5501
rect 24574 5475 24600 5501
rect 24636 5475 24662 5501
rect 24698 5475 24724 5501
rect 24760 5475 24786 5501
rect 24822 5475 24848 5501
rect 24884 5475 24910 5501
rect 24946 5475 24972 5501
rect 25008 5475 25034 5501
rect 29574 5475 29600 5501
rect 29636 5475 29662 5501
rect 29698 5475 29724 5501
rect 29760 5475 29786 5501
rect 29822 5475 29848 5501
rect 29884 5475 29910 5501
rect 29946 5475 29972 5501
rect 30008 5475 30034 5501
rect 34574 5475 34600 5501
rect 34636 5475 34662 5501
rect 34698 5475 34724 5501
rect 34760 5475 34786 5501
rect 34822 5475 34848 5501
rect 34884 5475 34910 5501
rect 34946 5475 34972 5501
rect 35008 5475 35034 5501
rect 1863 5335 1889 5361
rect 4439 5335 4465 5361
rect 16423 5335 16449 5361
rect 18439 5335 18465 5361
rect 20007 5335 20033 5361
rect 23423 5335 23449 5361
rect 30199 5335 30225 5361
rect 31823 5335 31849 5361
rect 35911 5335 35937 5361
rect 37647 5335 37673 5361
rect 1863 5279 1889 5305
rect 2759 5279 2785 5305
rect 3599 5279 3625 5305
rect 4439 5279 4465 5305
rect 6007 5279 6033 5305
rect 6399 5279 6425 5305
rect 6511 5279 6537 5305
rect 7519 5279 7545 5305
rect 7743 5279 7769 5305
rect 7967 5279 7993 5305
rect 9815 5279 9841 5305
rect 10263 5279 10289 5305
rect 10487 5279 10513 5305
rect 11551 5279 11577 5305
rect 11831 5279 11857 5305
rect 11943 5279 11969 5305
rect 13119 5279 13145 5305
rect 13287 5279 13313 5305
rect 13511 5279 13537 5305
rect 15359 5279 15385 5305
rect 16423 5279 16449 5305
rect 17599 5279 17625 5305
rect 18439 5279 18465 5305
rect 19055 5279 19081 5305
rect 20007 5279 20033 5305
rect 20847 5279 20873 5305
rect 21351 5279 21377 5305
rect 21463 5279 21489 5305
rect 22527 5279 22553 5305
rect 23423 5279 23449 5305
rect 25047 5279 25073 5305
rect 25215 5279 25241 5305
rect 25439 5279 25465 5305
rect 26503 5279 26529 5305
rect 26783 5279 26809 5305
rect 26895 5279 26921 5305
rect 29359 5279 29385 5305
rect 30199 5279 30225 5305
rect 30927 5279 30953 5305
rect 31823 5279 31849 5305
rect 32719 5279 32745 5305
rect 33279 5279 33305 5305
rect 33391 5279 33417 5305
rect 34175 5279 34201 5305
rect 34623 5279 34649 5305
rect 34847 5279 34873 5305
rect 35631 5279 35657 5305
rect 35743 5279 35769 5305
rect 36695 5279 36721 5305
rect 37647 5279 37673 5305
rect 2074 5083 2100 5109
rect 2136 5083 2162 5109
rect 2198 5083 2224 5109
rect 2260 5083 2286 5109
rect 2322 5083 2348 5109
rect 2384 5083 2410 5109
rect 2446 5083 2472 5109
rect 2508 5083 2534 5109
rect 7074 5083 7100 5109
rect 7136 5083 7162 5109
rect 7198 5083 7224 5109
rect 7260 5083 7286 5109
rect 7322 5083 7348 5109
rect 7384 5083 7410 5109
rect 7446 5083 7472 5109
rect 7508 5083 7534 5109
rect 12074 5083 12100 5109
rect 12136 5083 12162 5109
rect 12198 5083 12224 5109
rect 12260 5083 12286 5109
rect 12322 5083 12348 5109
rect 12384 5083 12410 5109
rect 12446 5083 12472 5109
rect 12508 5083 12534 5109
rect 17074 5083 17100 5109
rect 17136 5083 17162 5109
rect 17198 5083 17224 5109
rect 17260 5083 17286 5109
rect 17322 5083 17348 5109
rect 17384 5083 17410 5109
rect 17446 5083 17472 5109
rect 17508 5083 17534 5109
rect 22074 5083 22100 5109
rect 22136 5083 22162 5109
rect 22198 5083 22224 5109
rect 22260 5083 22286 5109
rect 22322 5083 22348 5109
rect 22384 5083 22410 5109
rect 22446 5083 22472 5109
rect 22508 5083 22534 5109
rect 27074 5083 27100 5109
rect 27136 5083 27162 5109
rect 27198 5083 27224 5109
rect 27260 5083 27286 5109
rect 27322 5083 27348 5109
rect 27384 5083 27410 5109
rect 27446 5083 27472 5109
rect 27508 5083 27534 5109
rect 32074 5083 32100 5109
rect 32136 5083 32162 5109
rect 32198 5083 32224 5109
rect 32260 5083 32286 5109
rect 32322 5083 32348 5109
rect 32384 5083 32410 5109
rect 32446 5083 32472 5109
rect 32508 5083 32534 5109
rect 37074 5083 37100 5109
rect 37136 5083 37162 5109
rect 37198 5083 37224 5109
rect 37260 5083 37286 5109
rect 37322 5083 37348 5109
rect 37384 5083 37410 5109
rect 37446 5083 37472 5109
rect 37508 5083 37534 5109
rect 1807 4887 1833 4913
rect 1919 4887 1945 4913
rect 2479 4887 2505 4913
rect 4103 4887 4129 4913
rect 4383 4887 4409 4913
rect 4495 4887 4521 4913
rect 5559 4887 5585 4913
rect 6399 4887 6425 4913
rect 7799 4887 7825 4913
rect 8247 4887 8273 4913
rect 8471 4887 8497 4913
rect 9535 4887 9561 4913
rect 10263 4887 10289 4913
rect 12335 4887 12361 4913
rect 12615 4887 12641 4913
rect 12727 4887 12753 4913
rect 15751 4887 15777 4913
rect 16759 4887 16785 4913
rect 17487 4887 17513 4913
rect 18383 4887 18409 4913
rect 19055 4887 19081 4913
rect 19951 4887 19977 4913
rect 20511 4887 20537 4913
rect 21351 4887 21377 4913
rect 23031 4887 23057 4913
rect 23871 4887 23897 4913
rect 24487 4887 24513 4913
rect 24655 4887 24681 4913
rect 24879 4887 24905 4913
rect 26895 4887 26921 4913
rect 27175 4887 27201 4913
rect 27399 4887 27425 4913
rect 28463 4887 28489 4913
rect 29303 4887 29329 4913
rect 30143 4887 30169 4913
rect 30367 4887 30393 4913
rect 30983 4887 31009 4913
rect 31879 4887 31905 4913
rect 32159 4887 32185 4913
rect 33335 4887 33361 4913
rect 33671 4887 33697 4913
rect 34679 4887 34705 4913
rect 35239 4887 35265 4913
rect 35351 4887 35377 4913
rect 36135 4887 36161 4913
rect 37311 4887 37337 4913
rect 6399 4831 6425 4857
rect 10263 4831 10289 4857
rect 16759 4831 16785 4857
rect 18383 4831 18409 4857
rect 19951 4831 19977 4857
rect 21351 4831 21377 4857
rect 23871 4831 23897 4857
rect 29303 4831 29329 4857
rect 30031 4831 30057 4857
rect 31879 4831 31905 4857
rect 33335 4831 33361 4857
rect 33727 4831 33753 4857
rect 33895 4831 33921 4857
rect 37311 4831 37337 4857
rect 37591 4831 37617 4857
rect 37703 4831 37729 4857
rect 37871 4831 37897 4857
rect 38655 4831 38681 4857
rect 38767 4831 38793 4857
rect 38935 4831 38961 4857
rect 4574 4691 4600 4717
rect 4636 4691 4662 4717
rect 4698 4691 4724 4717
rect 4760 4691 4786 4717
rect 4822 4691 4848 4717
rect 4884 4691 4910 4717
rect 4946 4691 4972 4717
rect 5008 4691 5034 4717
rect 9574 4691 9600 4717
rect 9636 4691 9662 4717
rect 9698 4691 9724 4717
rect 9760 4691 9786 4717
rect 9822 4691 9848 4717
rect 9884 4691 9910 4717
rect 9946 4691 9972 4717
rect 10008 4691 10034 4717
rect 14574 4691 14600 4717
rect 14636 4691 14662 4717
rect 14698 4691 14724 4717
rect 14760 4691 14786 4717
rect 14822 4691 14848 4717
rect 14884 4691 14910 4717
rect 14946 4691 14972 4717
rect 15008 4691 15034 4717
rect 19574 4691 19600 4717
rect 19636 4691 19662 4717
rect 19698 4691 19724 4717
rect 19760 4691 19786 4717
rect 19822 4691 19848 4717
rect 19884 4691 19910 4717
rect 19946 4691 19972 4717
rect 20008 4691 20034 4717
rect 24574 4691 24600 4717
rect 24636 4691 24662 4717
rect 24698 4691 24724 4717
rect 24760 4691 24786 4717
rect 24822 4691 24848 4717
rect 24884 4691 24910 4717
rect 24946 4691 24972 4717
rect 25008 4691 25034 4717
rect 29574 4691 29600 4717
rect 29636 4691 29662 4717
rect 29698 4691 29724 4717
rect 29760 4691 29786 4717
rect 29822 4691 29848 4717
rect 29884 4691 29910 4717
rect 29946 4691 29972 4717
rect 30008 4691 30034 4717
rect 34574 4691 34600 4717
rect 34636 4691 34662 4717
rect 34698 4691 34724 4717
rect 34760 4691 34786 4717
rect 34822 4691 34848 4717
rect 34884 4691 34910 4717
rect 34946 4691 34972 4717
rect 35008 4691 35034 4717
rect 1863 4551 1889 4577
rect 4439 4551 4465 4577
rect 6959 4551 6985 4577
rect 8247 4551 8273 4577
rect 14743 4551 14769 4577
rect 16423 4551 16449 4577
rect 18439 4551 18465 4577
rect 20007 4551 20033 4577
rect 21799 4551 21825 4577
rect 27175 4551 27201 4577
rect 28071 4551 28097 4577
rect 28239 4551 28265 4577
rect 31375 4551 31401 4577
rect 35351 4551 35377 4577
rect 37647 4551 37673 4577
rect 1863 4495 1889 4521
rect 2759 4495 2785 4521
rect 3319 4495 3345 4521
rect 4439 4495 4465 4521
rect 6007 4495 6033 4521
rect 6959 4495 6985 4521
rect 7295 4495 7321 4521
rect 8247 4495 8273 4521
rect 10039 4495 10065 4521
rect 10263 4495 10289 4521
rect 10487 4495 10513 4521
rect 11495 4495 11521 4521
rect 11775 4495 11801 4521
rect 11943 4495 11969 4521
rect 14071 4495 14097 4521
rect 14743 4495 14769 4521
rect 15359 4495 15385 4521
rect 16423 4495 16449 4521
rect 17599 4495 17625 4521
rect 18439 4495 18465 4521
rect 19111 4495 19137 4521
rect 20007 4495 20033 4521
rect 20847 4495 20873 4521
rect 21799 4495 21825 4521
rect 22527 4495 22553 4521
rect 22695 4495 22721 4521
rect 22919 4495 22945 4521
rect 24767 4495 24793 4521
rect 25215 4495 25241 4521
rect 25439 4495 25465 4521
rect 26503 4495 26529 4521
rect 26895 4495 26921 4521
rect 28351 4495 28377 4521
rect 28743 4495 28769 4521
rect 29303 4495 29329 4521
rect 29415 4495 29441 4521
rect 30479 4495 30505 4521
rect 31375 4495 31401 4521
rect 32047 4495 32073 4521
rect 32159 4495 32185 4521
rect 32327 4495 32353 4521
rect 32719 4495 32745 4521
rect 33279 4495 33305 4521
rect 33391 4495 33417 4521
rect 34455 4495 34481 4521
rect 35351 4495 35377 4521
rect 35687 4495 35713 4521
rect 35799 4495 35825 4521
rect 35967 4495 35993 4521
rect 36695 4495 36721 4521
rect 37647 4495 37673 4521
rect 38207 4495 38233 4521
rect 38263 4495 38289 4521
rect 38431 4495 38457 4521
rect 38711 4495 38737 4521
rect 38823 4495 38849 4521
rect 38991 4495 39017 4521
rect 2074 4299 2100 4325
rect 2136 4299 2162 4325
rect 2198 4299 2224 4325
rect 2260 4299 2286 4325
rect 2322 4299 2348 4325
rect 2384 4299 2410 4325
rect 2446 4299 2472 4325
rect 2508 4299 2534 4325
rect 7074 4299 7100 4325
rect 7136 4299 7162 4325
rect 7198 4299 7224 4325
rect 7260 4299 7286 4325
rect 7322 4299 7348 4325
rect 7384 4299 7410 4325
rect 7446 4299 7472 4325
rect 7508 4299 7534 4325
rect 12074 4299 12100 4325
rect 12136 4299 12162 4325
rect 12198 4299 12224 4325
rect 12260 4299 12286 4325
rect 12322 4299 12348 4325
rect 12384 4299 12410 4325
rect 12446 4299 12472 4325
rect 12508 4299 12534 4325
rect 17074 4299 17100 4325
rect 17136 4299 17162 4325
rect 17198 4299 17224 4325
rect 17260 4299 17286 4325
rect 17322 4299 17348 4325
rect 17384 4299 17410 4325
rect 17446 4299 17472 4325
rect 17508 4299 17534 4325
rect 22074 4299 22100 4325
rect 22136 4299 22162 4325
rect 22198 4299 22224 4325
rect 22260 4299 22286 4325
rect 22322 4299 22348 4325
rect 22384 4299 22410 4325
rect 22446 4299 22472 4325
rect 22508 4299 22534 4325
rect 27074 4299 27100 4325
rect 27136 4299 27162 4325
rect 27198 4299 27224 4325
rect 27260 4299 27286 4325
rect 27322 4299 27348 4325
rect 27384 4299 27410 4325
rect 27446 4299 27472 4325
rect 27508 4299 27534 4325
rect 32074 4299 32100 4325
rect 32136 4299 32162 4325
rect 32198 4299 32224 4325
rect 32260 4299 32286 4325
rect 32322 4299 32348 4325
rect 32384 4299 32410 4325
rect 32446 4299 32472 4325
rect 32508 4299 32534 4325
rect 37074 4299 37100 4325
rect 37136 4299 37162 4325
rect 37198 4299 37224 4325
rect 37260 4299 37286 4325
rect 37322 4299 37348 4325
rect 37384 4299 37410 4325
rect 37446 4299 37472 4325
rect 37508 4299 37534 4325
rect 1807 4103 1833 4129
rect 2031 4103 2057 4129
rect 2479 4103 2505 4129
rect 4103 4103 4129 4129
rect 4999 4103 5025 4129
rect 5279 4103 5305 4129
rect 6455 4103 6481 4129
rect 7799 4103 7825 4129
rect 8975 4103 9001 4129
rect 9479 4103 9505 4129
rect 10431 4103 10457 4129
rect 11775 4103 11801 4129
rect 12951 4103 12977 4129
rect 13231 4103 13257 4129
rect 14407 4103 14433 4129
rect 15751 4103 15777 4129
rect 16255 4103 16281 4129
rect 16423 4103 16449 4129
rect 17487 4103 17513 4129
rect 18383 4103 18409 4129
rect 19055 4103 19081 4129
rect 19951 4103 19977 4129
rect 20511 4103 20537 4129
rect 21351 4103 21377 4129
rect 22751 4103 22777 4129
rect 23871 4103 23897 4129
rect 24487 4103 24513 4129
rect 25383 4103 25409 4129
rect 26839 4103 26865 4129
rect 27511 4103 27537 4129
rect 28463 4103 28489 4129
rect 28687 4103 28713 4129
rect 28911 4103 28937 4129
rect 30087 4103 30113 4129
rect 30983 4103 31009 4129
rect 31879 4103 31905 4129
rect 32159 4103 32185 4129
rect 33335 4103 33361 4129
rect 33671 4103 33697 4129
rect 34679 4103 34705 4129
rect 35855 4103 35881 4129
rect 36135 4103 36161 4129
rect 37087 4103 37113 4129
rect 38823 4103 38849 4129
rect 38935 4103 38961 4129
rect 4999 4047 5025 4073
rect 6455 4047 6481 4073
rect 7799 4047 7825 4073
rect 10431 4047 10457 4073
rect 11775 4047 11801 4073
rect 14407 4047 14433 4073
rect 18383 4047 18409 4073
rect 19951 4047 19977 4073
rect 21351 4047 21377 4073
rect 23871 4047 23897 4073
rect 25383 4047 25409 4073
rect 27679 4047 27705 4073
rect 30143 4047 30169 4073
rect 30311 4047 30337 4073
rect 31879 4047 31905 4073
rect 33335 4047 33361 4073
rect 33727 4047 33753 4073
rect 33895 4047 33921 4073
rect 35855 4047 35881 4073
rect 37087 4047 37113 4073
rect 37591 4047 37617 4073
rect 37703 4047 37729 4073
rect 37871 4047 37897 4073
rect 38655 4047 38681 4073
rect 4574 3907 4600 3933
rect 4636 3907 4662 3933
rect 4698 3907 4724 3933
rect 4760 3907 4786 3933
rect 4822 3907 4848 3933
rect 4884 3907 4910 3933
rect 4946 3907 4972 3933
rect 5008 3907 5034 3933
rect 9574 3907 9600 3933
rect 9636 3907 9662 3933
rect 9698 3907 9724 3933
rect 9760 3907 9786 3933
rect 9822 3907 9848 3933
rect 9884 3907 9910 3933
rect 9946 3907 9972 3933
rect 10008 3907 10034 3933
rect 14574 3907 14600 3933
rect 14636 3907 14662 3933
rect 14698 3907 14724 3933
rect 14760 3907 14786 3933
rect 14822 3907 14848 3933
rect 14884 3907 14910 3933
rect 14946 3907 14972 3933
rect 15008 3907 15034 3933
rect 19574 3907 19600 3933
rect 19636 3907 19662 3933
rect 19698 3907 19724 3933
rect 19760 3907 19786 3933
rect 19822 3907 19848 3933
rect 19884 3907 19910 3933
rect 19946 3907 19972 3933
rect 20008 3907 20034 3933
rect 24574 3907 24600 3933
rect 24636 3907 24662 3933
rect 24698 3907 24724 3933
rect 24760 3907 24786 3933
rect 24822 3907 24848 3933
rect 24884 3907 24910 3933
rect 24946 3907 24972 3933
rect 25008 3907 25034 3933
rect 29574 3907 29600 3933
rect 29636 3907 29662 3933
rect 29698 3907 29724 3933
rect 29760 3907 29786 3933
rect 29822 3907 29848 3933
rect 29884 3907 29910 3933
rect 29946 3907 29972 3933
rect 30008 3907 30034 3933
rect 34574 3907 34600 3933
rect 34636 3907 34662 3933
rect 34698 3907 34724 3933
rect 34760 3907 34786 3933
rect 34822 3907 34848 3933
rect 34884 3907 34910 3933
rect 34946 3907 34972 3933
rect 35008 3907 35034 3933
rect 4495 3767 4521 3793
rect 7015 3767 7041 3793
rect 10879 3767 10905 3793
rect 14967 3767 14993 3793
rect 16423 3767 16449 3793
rect 18383 3767 18409 3793
rect 20007 3767 20033 3793
rect 25943 3767 25969 3793
rect 27175 3767 27201 3793
rect 29695 3767 29721 3793
rect 31375 3767 31401 3793
rect 33895 3767 33921 3793
rect 35351 3767 35377 3793
rect 35743 3767 35769 3793
rect 37647 3767 37673 3793
rect 2367 3711 2393 3737
rect 2479 3711 2505 3737
rect 2983 3711 3009 3737
rect 3599 3711 3625 3737
rect 4495 3711 4521 3737
rect 6063 3711 6089 3737
rect 7015 3711 7041 3737
rect 7799 3711 7825 3737
rect 8023 3711 8049 3737
rect 8471 3711 8497 3737
rect 9815 3711 9841 3737
rect 10879 3711 10905 3737
rect 11383 3711 11409 3737
rect 11831 3711 11857 3737
rect 11943 3711 11969 3737
rect 13791 3711 13817 3737
rect 14967 3711 14993 3737
rect 15247 3711 15273 3737
rect 16423 3711 16449 3737
rect 17599 3711 17625 3737
rect 18383 3711 18409 3737
rect 19111 3711 19137 3737
rect 20007 3711 20033 3737
rect 20959 3711 20985 3737
rect 21351 3711 21377 3737
rect 21463 3711 21489 3737
rect 22527 3711 22553 3737
rect 22695 3711 22721 3737
rect 22919 3711 22945 3737
rect 24767 3711 24793 3737
rect 25943 3711 25969 3737
rect 26223 3711 26249 3737
rect 27175 3711 27201 3737
rect 28015 3711 28041 3737
rect 28183 3711 28209 3737
rect 28295 3711 28321 3737
rect 28967 3711 28993 3737
rect 29471 3711 29497 3737
rect 30479 3711 30505 3737
rect 31375 3711 31401 3737
rect 32047 3711 32073 3737
rect 32159 3711 32185 3737
rect 32327 3711 32353 3737
rect 32887 3711 32913 3737
rect 33895 3711 33921 3737
rect 34175 3711 34201 3737
rect 35351 3711 35377 3737
rect 35687 3711 35713 3737
rect 35911 3711 35937 3737
rect 36695 3711 36721 3737
rect 37647 3711 37673 3737
rect 38151 3711 38177 3737
rect 38263 3711 38289 3737
rect 38431 3711 38457 3737
rect 38655 3711 38681 3737
rect 38823 3711 38849 3737
rect 38991 3711 39017 3737
rect 2074 3515 2100 3541
rect 2136 3515 2162 3541
rect 2198 3515 2224 3541
rect 2260 3515 2286 3541
rect 2322 3515 2348 3541
rect 2384 3515 2410 3541
rect 2446 3515 2472 3541
rect 2508 3515 2534 3541
rect 7074 3515 7100 3541
rect 7136 3515 7162 3541
rect 7198 3515 7224 3541
rect 7260 3515 7286 3541
rect 7322 3515 7348 3541
rect 7384 3515 7410 3541
rect 7446 3515 7472 3541
rect 7508 3515 7534 3541
rect 12074 3515 12100 3541
rect 12136 3515 12162 3541
rect 12198 3515 12224 3541
rect 12260 3515 12286 3541
rect 12322 3515 12348 3541
rect 12384 3515 12410 3541
rect 12446 3515 12472 3541
rect 12508 3515 12534 3541
rect 17074 3515 17100 3541
rect 17136 3515 17162 3541
rect 17198 3515 17224 3541
rect 17260 3515 17286 3541
rect 17322 3515 17348 3541
rect 17384 3515 17410 3541
rect 17446 3515 17472 3541
rect 17508 3515 17534 3541
rect 22074 3515 22100 3541
rect 22136 3515 22162 3541
rect 22198 3515 22224 3541
rect 22260 3515 22286 3541
rect 22322 3515 22348 3541
rect 22384 3515 22410 3541
rect 22446 3515 22472 3541
rect 22508 3515 22534 3541
rect 27074 3515 27100 3541
rect 27136 3515 27162 3541
rect 27198 3515 27224 3541
rect 27260 3515 27286 3541
rect 27322 3515 27348 3541
rect 27384 3515 27410 3541
rect 27446 3515 27472 3541
rect 27508 3515 27534 3541
rect 32074 3515 32100 3541
rect 32136 3515 32162 3541
rect 32198 3515 32224 3541
rect 32260 3515 32286 3541
rect 32322 3515 32348 3541
rect 32384 3515 32410 3541
rect 32446 3515 32472 3541
rect 32508 3515 32534 3541
rect 37074 3515 37100 3541
rect 37136 3515 37162 3541
rect 37198 3515 37224 3541
rect 37260 3515 37286 3541
rect 37322 3515 37348 3541
rect 37384 3515 37410 3541
rect 37446 3515 37472 3541
rect 37508 3515 37534 3541
rect 1359 3319 1385 3345
rect 2479 3319 2505 3345
rect 4103 3319 4129 3345
rect 4383 3319 4409 3345
rect 4495 3319 4521 3345
rect 5727 3319 5753 3345
rect 6007 3319 6033 3345
rect 6455 3319 6481 3345
rect 8303 3319 8329 3345
rect 8415 3319 8441 3345
rect 8975 3319 9001 3345
rect 9479 3319 9505 3345
rect 10431 3319 10457 3345
rect 11999 3319 12025 3345
rect 12335 3319 12361 3345
rect 12447 3319 12473 3345
rect 13231 3319 13257 3345
rect 14407 3319 14433 3345
rect 15751 3319 15777 3345
rect 16759 3319 16785 3345
rect 17487 3319 17513 3345
rect 18383 3319 18409 3345
rect 19055 3319 19081 3345
rect 19951 3319 19977 3345
rect 20511 3319 20537 3345
rect 21351 3319 21377 3345
rect 22751 3319 22777 3345
rect 23871 3319 23897 3345
rect 24431 3319 24457 3345
rect 25383 3319 25409 3345
rect 26895 3319 26921 3345
rect 27679 3319 27705 3345
rect 28463 3319 28489 3345
rect 29359 3319 29385 3345
rect 30703 3319 30729 3345
rect 31879 3319 31905 3345
rect 32439 3319 32465 3345
rect 32719 3319 32745 3345
rect 32831 3319 32857 3345
rect 33671 3319 33697 3345
rect 33895 3319 33921 3345
rect 34679 3319 34705 3345
rect 35631 3319 35657 3345
rect 36135 3319 36161 3345
rect 37311 3319 37337 3345
rect 1359 3263 1385 3289
rect 10431 3263 10457 3289
rect 14407 3263 14433 3289
rect 16759 3263 16785 3289
rect 18383 3263 18409 3289
rect 19951 3263 19977 3289
rect 21351 3263 21377 3289
rect 23871 3263 23897 3289
rect 25383 3263 25409 3289
rect 27679 3263 27705 3289
rect 29359 3263 29385 3289
rect 30031 3263 30057 3289
rect 30143 3263 30169 3289
rect 30311 3263 30337 3289
rect 31879 3263 31905 3289
rect 33727 3263 33753 3289
rect 35631 3263 35657 3289
rect 37311 3263 37337 3289
rect 37591 3263 37617 3289
rect 37703 3263 37729 3289
rect 37871 3263 37897 3289
rect 38655 3263 38681 3289
rect 38823 3263 38849 3289
rect 38935 3263 38961 3289
rect 4574 3123 4600 3149
rect 4636 3123 4662 3149
rect 4698 3123 4724 3149
rect 4760 3123 4786 3149
rect 4822 3123 4848 3149
rect 4884 3123 4910 3149
rect 4946 3123 4972 3149
rect 5008 3123 5034 3149
rect 9574 3123 9600 3149
rect 9636 3123 9662 3149
rect 9698 3123 9724 3149
rect 9760 3123 9786 3149
rect 9822 3123 9848 3149
rect 9884 3123 9910 3149
rect 9946 3123 9972 3149
rect 10008 3123 10034 3149
rect 14574 3123 14600 3149
rect 14636 3123 14662 3149
rect 14698 3123 14724 3149
rect 14760 3123 14786 3149
rect 14822 3123 14848 3149
rect 14884 3123 14910 3149
rect 14946 3123 14972 3149
rect 15008 3123 15034 3149
rect 19574 3123 19600 3149
rect 19636 3123 19662 3149
rect 19698 3123 19724 3149
rect 19760 3123 19786 3149
rect 19822 3123 19848 3149
rect 19884 3123 19910 3149
rect 19946 3123 19972 3149
rect 20008 3123 20034 3149
rect 24574 3123 24600 3149
rect 24636 3123 24662 3149
rect 24698 3123 24724 3149
rect 24760 3123 24786 3149
rect 24822 3123 24848 3149
rect 24884 3123 24910 3149
rect 24946 3123 24972 3149
rect 25008 3123 25034 3149
rect 29574 3123 29600 3149
rect 29636 3123 29662 3149
rect 29698 3123 29724 3149
rect 29760 3123 29786 3149
rect 29822 3123 29848 3149
rect 29884 3123 29910 3149
rect 29946 3123 29972 3149
rect 30008 3123 30034 3149
rect 34574 3123 34600 3149
rect 34636 3123 34662 3149
rect 34698 3123 34724 3149
rect 34760 3123 34786 3149
rect 34822 3123 34848 3149
rect 34884 3123 34910 3149
rect 34946 3123 34972 3149
rect 35008 3123 35034 3149
rect 1975 2983 2001 3009
rect 4495 2983 4521 3009
rect 8471 2983 8497 3009
rect 12447 2983 12473 3009
rect 14967 2983 14993 3009
rect 18383 2983 18409 3009
rect 20007 2983 20033 3009
rect 23423 2983 23449 3009
rect 25943 2983 25969 3009
rect 27399 2983 27425 3009
rect 28071 2983 28097 3009
rect 28351 2983 28377 3009
rect 29919 2983 29945 3009
rect 31263 2983 31289 3009
rect 32159 2983 32185 3009
rect 32327 2983 32353 3009
rect 35351 2983 35377 3009
rect 35743 2983 35769 3009
rect 35911 2983 35937 3009
rect 38431 2983 38457 3009
rect 1975 2927 2001 2953
rect 3039 2927 3065 2953
rect 3599 2927 3625 2953
rect 4495 2927 4521 2953
rect 6343 2927 6369 2953
rect 6455 2927 6481 2953
rect 7015 2927 7041 2953
rect 7575 2927 7601 2953
rect 8471 2927 8497 2953
rect 10319 2927 10345 2953
rect 10487 2927 10513 2953
rect 10879 2927 10905 2953
rect 11383 2927 11409 2953
rect 12447 2927 12473 2953
rect 14071 2927 14097 2953
rect 14967 2927 14993 2953
rect 15247 2927 15273 2953
rect 15695 2927 15721 2953
rect 16423 2927 16449 2953
rect 17599 2927 17625 2953
rect 18383 2927 18409 2953
rect 19111 2927 19137 2953
rect 20007 2927 20033 2953
rect 20959 2927 20985 2953
rect 21351 2927 21377 2953
rect 21463 2927 21489 2953
rect 22527 2927 22553 2953
rect 23423 2927 23449 2953
rect 24767 2927 24793 2953
rect 25943 2927 25969 2953
rect 26223 2927 26249 2953
rect 27399 2927 27425 2953
rect 28183 2927 28209 2953
rect 28743 2927 28769 2953
rect 29919 2927 29945 2953
rect 30367 2927 30393 2953
rect 31263 2927 31289 2953
rect 32047 2927 32073 2953
rect 32999 2927 33025 2953
rect 33167 2927 33193 2953
rect 33391 2927 33417 2953
rect 34175 2927 34201 2953
rect 35351 2927 35377 2953
rect 35687 2927 35713 2953
rect 36751 2927 36777 2953
rect 37143 2927 37169 2953
rect 37367 2927 37393 2953
rect 38207 2927 38233 2953
rect 38263 2927 38289 2953
rect 38655 2927 38681 2953
rect 38823 2927 38849 2953
rect 38935 2927 38961 2953
rect 2074 2731 2100 2757
rect 2136 2731 2162 2757
rect 2198 2731 2224 2757
rect 2260 2731 2286 2757
rect 2322 2731 2348 2757
rect 2384 2731 2410 2757
rect 2446 2731 2472 2757
rect 2508 2731 2534 2757
rect 7074 2731 7100 2757
rect 7136 2731 7162 2757
rect 7198 2731 7224 2757
rect 7260 2731 7286 2757
rect 7322 2731 7348 2757
rect 7384 2731 7410 2757
rect 7446 2731 7472 2757
rect 7508 2731 7534 2757
rect 12074 2731 12100 2757
rect 12136 2731 12162 2757
rect 12198 2731 12224 2757
rect 12260 2731 12286 2757
rect 12322 2731 12348 2757
rect 12384 2731 12410 2757
rect 12446 2731 12472 2757
rect 12508 2731 12534 2757
rect 17074 2731 17100 2757
rect 17136 2731 17162 2757
rect 17198 2731 17224 2757
rect 17260 2731 17286 2757
rect 17322 2731 17348 2757
rect 17384 2731 17410 2757
rect 17446 2731 17472 2757
rect 17508 2731 17534 2757
rect 22074 2731 22100 2757
rect 22136 2731 22162 2757
rect 22198 2731 22224 2757
rect 22260 2731 22286 2757
rect 22322 2731 22348 2757
rect 22384 2731 22410 2757
rect 22446 2731 22472 2757
rect 22508 2731 22534 2757
rect 27074 2731 27100 2757
rect 27136 2731 27162 2757
rect 27198 2731 27224 2757
rect 27260 2731 27286 2757
rect 27322 2731 27348 2757
rect 27384 2731 27410 2757
rect 27446 2731 27472 2757
rect 27508 2731 27534 2757
rect 32074 2731 32100 2757
rect 32136 2731 32162 2757
rect 32198 2731 32224 2757
rect 32260 2731 32286 2757
rect 32322 2731 32348 2757
rect 32384 2731 32410 2757
rect 32446 2731 32472 2757
rect 32508 2731 32534 2757
rect 37074 2731 37100 2757
rect 37136 2731 37162 2757
rect 37198 2731 37224 2757
rect 37260 2731 37286 2757
rect 37322 2731 37348 2757
rect 37384 2731 37410 2757
rect 37446 2731 37472 2757
rect 37508 2731 37534 2757
rect 1639 2535 1665 2561
rect 2479 2535 2505 2561
rect 4047 2535 4073 2561
rect 4999 2535 5025 2561
rect 5727 2535 5753 2561
rect 6455 2535 6481 2561
rect 8079 2535 8105 2561
rect 8975 2535 9001 2561
rect 9479 2535 9505 2561
rect 10431 2535 10457 2561
rect 12223 2535 12249 2561
rect 13175 2535 13201 2561
rect 15751 2535 15777 2561
rect 16759 2535 16785 2561
rect 17375 2535 17401 2561
rect 18271 2535 18297 2561
rect 19055 2535 19081 2561
rect 19951 2535 19977 2561
rect 20511 2535 20537 2561
rect 21351 2535 21377 2561
rect 22751 2535 22777 2561
rect 23871 2535 23897 2561
rect 24431 2535 24457 2561
rect 25383 2535 25409 2561
rect 26727 2535 26753 2561
rect 27679 2535 27705 2561
rect 28463 2535 28489 2561
rect 29359 2535 29385 2561
rect 30087 2535 30113 2561
rect 30143 2535 30169 2561
rect 30311 2535 30337 2561
rect 30815 2535 30841 2561
rect 31879 2535 31905 2561
rect 32159 2535 32185 2561
rect 33335 2535 33361 2561
rect 33671 2535 33697 2561
rect 33895 2535 33921 2561
rect 34679 2535 34705 2561
rect 35855 2535 35881 2561
rect 36135 2535 36161 2561
rect 36975 2535 37001 2561
rect 38655 2535 38681 2561
rect 38767 2535 38793 2561
rect 1527 2479 1553 2505
rect 4999 2479 5025 2505
rect 5503 2479 5529 2505
rect 8975 2479 9001 2505
rect 10431 2479 10457 2505
rect 13175 2479 13201 2505
rect 16759 2479 16785 2505
rect 18271 2479 18297 2505
rect 19951 2479 19977 2505
rect 21351 2479 21377 2505
rect 23871 2479 23897 2505
rect 25383 2479 25409 2505
rect 27679 2479 27705 2505
rect 29359 2479 29385 2505
rect 31879 2479 31905 2505
rect 33335 2479 33361 2505
rect 33727 2479 33753 2505
rect 35855 2479 35881 2505
rect 37087 2479 37113 2505
rect 37591 2479 37617 2505
rect 37703 2479 37729 2505
rect 37871 2479 37897 2505
rect 38935 2479 38961 2505
rect 4574 2339 4600 2365
rect 4636 2339 4662 2365
rect 4698 2339 4724 2365
rect 4760 2339 4786 2365
rect 4822 2339 4848 2365
rect 4884 2339 4910 2365
rect 4946 2339 4972 2365
rect 5008 2339 5034 2365
rect 9574 2339 9600 2365
rect 9636 2339 9662 2365
rect 9698 2339 9724 2365
rect 9760 2339 9786 2365
rect 9822 2339 9848 2365
rect 9884 2339 9910 2365
rect 9946 2339 9972 2365
rect 10008 2339 10034 2365
rect 14574 2339 14600 2365
rect 14636 2339 14662 2365
rect 14698 2339 14724 2365
rect 14760 2339 14786 2365
rect 14822 2339 14848 2365
rect 14884 2339 14910 2365
rect 14946 2339 14972 2365
rect 15008 2339 15034 2365
rect 19574 2339 19600 2365
rect 19636 2339 19662 2365
rect 19698 2339 19724 2365
rect 19760 2339 19786 2365
rect 19822 2339 19848 2365
rect 19884 2339 19910 2365
rect 19946 2339 19972 2365
rect 20008 2339 20034 2365
rect 24574 2339 24600 2365
rect 24636 2339 24662 2365
rect 24698 2339 24724 2365
rect 24760 2339 24786 2365
rect 24822 2339 24848 2365
rect 24884 2339 24910 2365
rect 24946 2339 24972 2365
rect 25008 2339 25034 2365
rect 29574 2339 29600 2365
rect 29636 2339 29662 2365
rect 29698 2339 29724 2365
rect 29760 2339 29786 2365
rect 29822 2339 29848 2365
rect 29884 2339 29910 2365
rect 29946 2339 29972 2365
rect 30008 2339 30034 2365
rect 34574 2339 34600 2365
rect 34636 2339 34662 2365
rect 34698 2339 34724 2365
rect 34760 2339 34786 2365
rect 34822 2339 34848 2365
rect 34884 2339 34910 2365
rect 34946 2339 34972 2365
rect 35008 2339 35034 2365
rect 4495 2199 4521 2225
rect 5839 2199 5865 2225
rect 8359 2199 8385 2225
rect 10823 2199 10849 2225
rect 18271 2199 18297 2225
rect 19503 2199 19529 2225
rect 21799 2199 21825 2225
rect 23423 2199 23449 2225
rect 25943 2199 25969 2225
rect 27399 2199 27425 2225
rect 28071 2199 28097 2225
rect 29919 2199 29945 2225
rect 31375 2199 31401 2225
rect 32159 2199 32185 2225
rect 32327 2199 32353 2225
rect 33839 2199 33865 2225
rect 35183 2199 35209 2225
rect 35743 2199 35769 2225
rect 35911 2199 35937 2225
rect 37647 2199 37673 2225
rect 38151 2199 38177 2225
rect 38431 2199 38457 2225
rect 38711 2199 38737 2225
rect 38879 2199 38905 2225
rect 2367 2143 2393 2169
rect 2479 2143 2505 2169
rect 3039 2143 3065 2169
rect 3543 2143 3569 2169
rect 4439 2143 4465 2169
rect 5839 2143 5865 2169
rect 7015 2143 7041 2169
rect 7519 2143 7545 2169
rect 8359 2143 8385 2169
rect 10039 2143 10065 2169
rect 10823 2143 10849 2169
rect 11383 2143 11409 2169
rect 11775 2143 11801 2169
rect 11943 2143 11969 2169
rect 13791 2143 13817 2169
rect 14239 2143 14265 2169
rect 14463 2143 14489 2169
rect 15247 2143 15273 2169
rect 15695 2143 15721 2169
rect 15919 2143 15945 2169
rect 17375 2143 17401 2169
rect 18271 2143 18297 2169
rect 18831 2143 18857 2169
rect 19503 2143 19529 2169
rect 20791 2143 20817 2169
rect 21799 2143 21825 2169
rect 22247 2143 22273 2169
rect 23423 2143 23449 2169
rect 24767 2143 24793 2169
rect 25943 2143 25969 2169
rect 26223 2143 26249 2169
rect 27399 2143 27425 2169
rect 28183 2143 28209 2169
rect 28351 2143 28377 2169
rect 28743 2143 28769 2169
rect 29919 2143 29945 2169
rect 30311 2143 30337 2169
rect 31375 2143 31401 2169
rect 32103 2143 32129 2169
rect 32719 2143 32745 2169
rect 33839 2143 33865 2169
rect 34231 2143 34257 2169
rect 35183 2143 35209 2169
rect 35687 2143 35713 2169
rect 36695 2143 36721 2169
rect 37647 2143 37673 2169
rect 38319 2143 38345 2169
rect 38935 2143 38961 2169
rect 2074 1947 2100 1973
rect 2136 1947 2162 1973
rect 2198 1947 2224 1973
rect 2260 1947 2286 1973
rect 2322 1947 2348 1973
rect 2384 1947 2410 1973
rect 2446 1947 2472 1973
rect 2508 1947 2534 1973
rect 7074 1947 7100 1973
rect 7136 1947 7162 1973
rect 7198 1947 7224 1973
rect 7260 1947 7286 1973
rect 7322 1947 7348 1973
rect 7384 1947 7410 1973
rect 7446 1947 7472 1973
rect 7508 1947 7534 1973
rect 12074 1947 12100 1973
rect 12136 1947 12162 1973
rect 12198 1947 12224 1973
rect 12260 1947 12286 1973
rect 12322 1947 12348 1973
rect 12384 1947 12410 1973
rect 12446 1947 12472 1973
rect 12508 1947 12534 1973
rect 17074 1947 17100 1973
rect 17136 1947 17162 1973
rect 17198 1947 17224 1973
rect 17260 1947 17286 1973
rect 17322 1947 17348 1973
rect 17384 1947 17410 1973
rect 17446 1947 17472 1973
rect 17508 1947 17534 1973
rect 22074 1947 22100 1973
rect 22136 1947 22162 1973
rect 22198 1947 22224 1973
rect 22260 1947 22286 1973
rect 22322 1947 22348 1973
rect 22384 1947 22410 1973
rect 22446 1947 22472 1973
rect 22508 1947 22534 1973
rect 27074 1947 27100 1973
rect 27136 1947 27162 1973
rect 27198 1947 27224 1973
rect 27260 1947 27286 1973
rect 27322 1947 27348 1973
rect 27384 1947 27410 1973
rect 27446 1947 27472 1973
rect 27508 1947 27534 1973
rect 32074 1947 32100 1973
rect 32136 1947 32162 1973
rect 32198 1947 32224 1973
rect 32260 1947 32286 1973
rect 32322 1947 32348 1973
rect 32384 1947 32410 1973
rect 32446 1947 32472 1973
rect 32508 1947 32534 1973
rect 37074 1947 37100 1973
rect 37136 1947 37162 1973
rect 37198 1947 37224 1973
rect 37260 1947 37286 1973
rect 37322 1947 37348 1973
rect 37384 1947 37410 1973
rect 37446 1947 37472 1973
rect 37508 1947 37534 1973
rect 1191 1751 1217 1777
rect 1919 1751 1945 1777
rect 3543 1751 3569 1777
rect 4439 1751 4465 1777
rect 5503 1751 5529 1777
rect 6399 1751 6425 1777
rect 7463 1751 7489 1777
rect 8359 1751 8385 1777
rect 9367 1751 9393 1777
rect 9703 1751 9729 1777
rect 9815 1751 9841 1777
rect 11383 1751 11409 1777
rect 11663 1751 11689 1777
rect 11775 1751 11801 1777
rect 13063 1751 13089 1777
rect 13511 1751 13537 1777
rect 13735 1751 13761 1777
rect 15247 1751 15273 1777
rect 15583 1751 15609 1777
rect 15695 1751 15721 1777
rect 17263 1751 17289 1777
rect 18159 1751 18185 1777
rect 18831 1751 18857 1777
rect 19503 1751 19529 1777
rect 20511 1751 20537 1777
rect 21687 1751 21713 1777
rect 22471 1751 22497 1777
rect 23647 1751 23673 1777
rect 24431 1751 24457 1777
rect 25607 1751 25633 1777
rect 26391 1751 26417 1777
rect 27567 1751 27593 1777
rect 28519 1751 28545 1777
rect 29359 1751 29385 1777
rect 30311 1751 30337 1777
rect 31487 1751 31513 1777
rect 32551 1751 32577 1777
rect 33447 1751 33473 1777
rect 34231 1751 34257 1777
rect 35183 1751 35209 1777
rect 36191 1751 36217 1777
rect 36975 1751 37001 1777
rect 38151 1751 38177 1777
rect 38263 1751 38289 1777
rect 38431 1751 38457 1777
rect 38655 1751 38681 1777
rect 38823 1751 38849 1777
rect 38935 1751 38961 1777
rect 1919 1695 1945 1721
rect 4439 1695 4465 1721
rect 6399 1695 6425 1721
rect 8359 1695 8385 1721
rect 18159 1695 18185 1721
rect 19503 1695 19529 1721
rect 21687 1695 21713 1721
rect 23647 1695 23673 1721
rect 25607 1695 25633 1721
rect 27567 1695 27593 1721
rect 29359 1695 29385 1721
rect 31487 1695 31513 1721
rect 33447 1695 33473 1721
rect 35183 1695 35209 1721
rect 37143 1695 37169 1721
rect 4574 1555 4600 1581
rect 4636 1555 4662 1581
rect 4698 1555 4724 1581
rect 4760 1555 4786 1581
rect 4822 1555 4848 1581
rect 4884 1555 4910 1581
rect 4946 1555 4972 1581
rect 5008 1555 5034 1581
rect 9574 1555 9600 1581
rect 9636 1555 9662 1581
rect 9698 1555 9724 1581
rect 9760 1555 9786 1581
rect 9822 1555 9848 1581
rect 9884 1555 9910 1581
rect 9946 1555 9972 1581
rect 10008 1555 10034 1581
rect 14574 1555 14600 1581
rect 14636 1555 14662 1581
rect 14698 1555 14724 1581
rect 14760 1555 14786 1581
rect 14822 1555 14848 1581
rect 14884 1555 14910 1581
rect 14946 1555 14972 1581
rect 15008 1555 15034 1581
rect 19574 1555 19600 1581
rect 19636 1555 19662 1581
rect 19698 1555 19724 1581
rect 19760 1555 19786 1581
rect 19822 1555 19848 1581
rect 19884 1555 19910 1581
rect 19946 1555 19972 1581
rect 20008 1555 20034 1581
rect 24574 1555 24600 1581
rect 24636 1555 24662 1581
rect 24698 1555 24724 1581
rect 24760 1555 24786 1581
rect 24822 1555 24848 1581
rect 24884 1555 24910 1581
rect 24946 1555 24972 1581
rect 25008 1555 25034 1581
rect 29574 1555 29600 1581
rect 29636 1555 29662 1581
rect 29698 1555 29724 1581
rect 29760 1555 29786 1581
rect 29822 1555 29848 1581
rect 29884 1555 29910 1581
rect 29946 1555 29972 1581
rect 30008 1555 30034 1581
rect 34574 1555 34600 1581
rect 34636 1555 34662 1581
rect 34698 1555 34724 1581
rect 34760 1555 34786 1581
rect 34822 1555 34848 1581
rect 34884 1555 34910 1581
rect 34946 1555 34972 1581
rect 35008 1555 35034 1581
<< metal2 >>
rect 2520 19600 2576 20000
rect 7014 19614 7378 19642
rect 2534 18522 2562 19600
rect 2534 18494 2674 18522
rect 2073 18438 2535 18443
rect 2073 18437 2082 18438
rect 2073 18411 2074 18437
rect 2073 18410 2082 18411
rect 2110 18410 2134 18438
rect 2162 18410 2186 18438
rect 2214 18437 2238 18438
rect 2266 18437 2290 18438
rect 2224 18411 2238 18437
rect 2286 18411 2290 18437
rect 2214 18410 2238 18411
rect 2266 18410 2290 18411
rect 2318 18437 2342 18438
rect 2370 18437 2394 18438
rect 2318 18411 2322 18437
rect 2370 18411 2384 18437
rect 2318 18410 2342 18411
rect 2370 18410 2394 18411
rect 2422 18410 2446 18438
rect 2474 18410 2498 18438
rect 2526 18437 2535 18438
rect 2534 18411 2535 18437
rect 2526 18410 2535 18411
rect 2073 18405 2535 18410
rect 2073 17654 2535 17659
rect 2073 17653 2082 17654
rect 2073 17627 2074 17653
rect 2073 17626 2082 17627
rect 2110 17626 2134 17654
rect 2162 17626 2186 17654
rect 2214 17653 2238 17654
rect 2266 17653 2290 17654
rect 2224 17627 2238 17653
rect 2286 17627 2290 17653
rect 2214 17626 2238 17627
rect 2266 17626 2290 17627
rect 2318 17653 2342 17654
rect 2370 17653 2394 17654
rect 2318 17627 2322 17653
rect 2370 17627 2384 17653
rect 2318 17626 2342 17627
rect 2370 17626 2394 17627
rect 2422 17626 2446 17654
rect 2474 17626 2498 17654
rect 2526 17653 2535 17654
rect 2534 17627 2535 17653
rect 2526 17626 2535 17627
rect 2073 17621 2535 17626
rect 2073 16870 2535 16875
rect 2073 16869 2082 16870
rect 2073 16843 2074 16869
rect 2073 16842 2082 16843
rect 2110 16842 2134 16870
rect 2162 16842 2186 16870
rect 2214 16869 2238 16870
rect 2266 16869 2290 16870
rect 2224 16843 2238 16869
rect 2286 16843 2290 16869
rect 2214 16842 2238 16843
rect 2266 16842 2290 16843
rect 2318 16869 2342 16870
rect 2370 16869 2394 16870
rect 2318 16843 2322 16869
rect 2370 16843 2384 16869
rect 2318 16842 2342 16843
rect 2370 16842 2394 16843
rect 2422 16842 2446 16870
rect 2474 16842 2498 16870
rect 2526 16869 2535 16870
rect 2534 16843 2535 16869
rect 2526 16842 2535 16843
rect 2073 16837 2535 16842
rect 2073 16086 2535 16091
rect 2073 16085 2082 16086
rect 2073 16059 2074 16085
rect 2073 16058 2082 16059
rect 2110 16058 2134 16086
rect 2162 16058 2186 16086
rect 2214 16085 2238 16086
rect 2266 16085 2290 16086
rect 2224 16059 2238 16085
rect 2286 16059 2290 16085
rect 2214 16058 2238 16059
rect 2266 16058 2290 16059
rect 2318 16085 2342 16086
rect 2370 16085 2394 16086
rect 2318 16059 2322 16085
rect 2370 16059 2384 16085
rect 2318 16058 2342 16059
rect 2370 16058 2394 16059
rect 2422 16058 2446 16086
rect 2474 16058 2498 16086
rect 2526 16085 2535 16086
rect 2534 16059 2535 16085
rect 2526 16058 2535 16059
rect 2073 16053 2535 16058
rect 2073 15302 2535 15307
rect 2073 15301 2082 15302
rect 2073 15275 2074 15301
rect 2073 15274 2082 15275
rect 2110 15274 2134 15302
rect 2162 15274 2186 15302
rect 2214 15301 2238 15302
rect 2266 15301 2290 15302
rect 2224 15275 2238 15301
rect 2286 15275 2290 15301
rect 2214 15274 2238 15275
rect 2266 15274 2290 15275
rect 2318 15301 2342 15302
rect 2370 15301 2394 15302
rect 2318 15275 2322 15301
rect 2370 15275 2384 15301
rect 2318 15274 2342 15275
rect 2370 15274 2394 15275
rect 2422 15274 2446 15302
rect 2474 15274 2498 15302
rect 2526 15301 2535 15302
rect 2534 15275 2535 15301
rect 2526 15274 2535 15275
rect 2073 15269 2535 15274
rect 1806 15106 1834 15111
rect 1918 15106 1946 15111
rect 1806 15105 1946 15106
rect 1806 15079 1807 15105
rect 1833 15079 1919 15105
rect 1945 15079 1946 15105
rect 1806 15078 1946 15079
rect 1806 15073 1834 15078
rect 1862 14769 1890 15078
rect 1918 15073 1946 15078
rect 2422 15105 2450 15111
rect 2422 15079 2423 15105
rect 2449 15079 2450 15105
rect 1862 14743 1863 14769
rect 1889 14743 1890 14769
rect 1862 14713 1890 14743
rect 1862 14687 1863 14713
rect 1889 14687 1890 14713
rect 1806 14322 1834 14327
rect 1862 14322 1890 14687
rect 2422 14714 2450 15079
rect 2422 14681 2450 14686
rect 2590 14714 2618 14719
rect 2073 14518 2535 14523
rect 2073 14517 2082 14518
rect 2073 14491 2074 14517
rect 2073 14490 2082 14491
rect 2110 14490 2134 14518
rect 2162 14490 2186 14518
rect 2214 14517 2238 14518
rect 2266 14517 2290 14518
rect 2224 14491 2238 14517
rect 2286 14491 2290 14517
rect 2214 14490 2238 14491
rect 2266 14490 2290 14491
rect 2318 14517 2342 14518
rect 2370 14517 2394 14518
rect 2318 14491 2322 14517
rect 2370 14491 2384 14517
rect 2318 14490 2342 14491
rect 2370 14490 2394 14491
rect 2422 14490 2446 14518
rect 2474 14490 2498 14518
rect 2526 14517 2535 14518
rect 2534 14491 2535 14517
rect 2526 14490 2535 14491
rect 2073 14485 2535 14490
rect 2478 14378 2506 14383
rect 1918 14322 1946 14327
rect 1806 14321 1946 14322
rect 1806 14295 1807 14321
rect 1833 14295 1919 14321
rect 1945 14295 1946 14321
rect 1806 14294 1946 14295
rect 1806 13538 1834 14294
rect 1918 14289 1946 14294
rect 2422 14322 2450 14327
rect 2422 14275 2450 14294
rect 2366 13930 2394 13935
rect 2478 13930 2506 14350
rect 2366 13929 2506 13930
rect 2366 13903 2367 13929
rect 2393 13903 2479 13929
rect 2505 13903 2506 13929
rect 2366 13902 2506 13903
rect 2366 13897 2394 13902
rect 2478 13897 2506 13902
rect 2590 14322 2618 14686
rect 2073 13734 2535 13739
rect 2073 13733 2082 13734
rect 2073 13707 2074 13733
rect 2073 13706 2082 13707
rect 2110 13706 2134 13734
rect 2162 13706 2186 13734
rect 2214 13733 2238 13734
rect 2266 13733 2290 13734
rect 2224 13707 2238 13733
rect 2286 13707 2290 13733
rect 2214 13706 2238 13707
rect 2266 13706 2290 13707
rect 2318 13733 2342 13734
rect 2370 13733 2394 13734
rect 2318 13707 2322 13733
rect 2370 13707 2384 13733
rect 2318 13706 2342 13707
rect 2370 13706 2394 13707
rect 2422 13706 2446 13734
rect 2474 13706 2498 13734
rect 2526 13733 2535 13734
rect 2534 13707 2535 13733
rect 2526 13706 2535 13707
rect 2073 13701 2535 13706
rect 1918 13538 1946 13543
rect 1638 13537 1946 13538
rect 1638 13511 1807 13537
rect 1833 13511 1919 13537
rect 1945 13511 1946 13537
rect 1638 13510 1946 13511
rect 1638 12586 1666 13510
rect 1806 13505 1834 13510
rect 1918 13505 1946 13510
rect 2478 13538 2506 13543
rect 2590 13538 2618 14294
rect 2478 13537 2618 13538
rect 2478 13511 2479 13537
rect 2505 13511 2618 13537
rect 2478 13510 2618 13511
rect 2478 13505 2506 13510
rect 1974 13146 2002 13151
rect 1806 12754 1834 12759
rect 1974 12754 2002 13118
rect 2366 13146 2394 13151
rect 2590 13146 2618 13151
rect 2646 13146 2674 18494
rect 4573 18046 5035 18051
rect 4573 18045 4582 18046
rect 4573 18019 4574 18045
rect 4573 18018 4582 18019
rect 4610 18018 4634 18046
rect 4662 18018 4686 18046
rect 4714 18045 4738 18046
rect 4766 18045 4790 18046
rect 4724 18019 4738 18045
rect 4786 18019 4790 18045
rect 4714 18018 4738 18019
rect 4766 18018 4790 18019
rect 4818 18045 4842 18046
rect 4870 18045 4894 18046
rect 4818 18019 4822 18045
rect 4870 18019 4884 18045
rect 4818 18018 4842 18019
rect 4870 18018 4894 18019
rect 4922 18018 4946 18046
rect 4974 18018 4998 18046
rect 5026 18045 5035 18046
rect 5034 18019 5035 18045
rect 5026 18018 5035 18019
rect 4573 18013 5035 18018
rect 4573 17262 5035 17267
rect 4573 17261 4582 17262
rect 4573 17235 4574 17261
rect 4573 17234 4582 17235
rect 4610 17234 4634 17262
rect 4662 17234 4686 17262
rect 4714 17261 4738 17262
rect 4766 17261 4790 17262
rect 4724 17235 4738 17261
rect 4786 17235 4790 17261
rect 4714 17234 4738 17235
rect 4766 17234 4790 17235
rect 4818 17261 4842 17262
rect 4870 17261 4894 17262
rect 4818 17235 4822 17261
rect 4870 17235 4884 17261
rect 4818 17234 4842 17235
rect 4870 17234 4894 17235
rect 4922 17234 4946 17262
rect 4974 17234 4998 17262
rect 5026 17261 5035 17262
rect 5034 17235 5035 17261
rect 5026 17234 5035 17235
rect 4573 17229 5035 17234
rect 4573 16478 5035 16483
rect 4573 16477 4582 16478
rect 4573 16451 4574 16477
rect 4573 16450 4582 16451
rect 4610 16450 4634 16478
rect 4662 16450 4686 16478
rect 4714 16477 4738 16478
rect 4766 16477 4790 16478
rect 4724 16451 4738 16477
rect 4786 16451 4790 16477
rect 4714 16450 4738 16451
rect 4766 16450 4790 16451
rect 4818 16477 4842 16478
rect 4870 16477 4894 16478
rect 4818 16451 4822 16477
rect 4870 16451 4884 16477
rect 4818 16450 4842 16451
rect 4870 16450 4894 16451
rect 4922 16450 4946 16478
rect 4974 16450 4998 16478
rect 5026 16477 5035 16478
rect 5034 16451 5035 16477
rect 5026 16450 5035 16451
rect 4573 16445 5035 16450
rect 7014 16337 7042 19614
rect 7350 19530 7378 19614
rect 7504 19600 7560 20000
rect 12488 19600 12544 20000
rect 16870 19614 17346 19642
rect 7518 19530 7546 19600
rect 7350 19502 7546 19530
rect 12502 18522 12530 19600
rect 12502 18494 12642 18522
rect 7073 18438 7535 18443
rect 7073 18437 7082 18438
rect 7073 18411 7074 18437
rect 7073 18410 7082 18411
rect 7110 18410 7134 18438
rect 7162 18410 7186 18438
rect 7214 18437 7238 18438
rect 7266 18437 7290 18438
rect 7224 18411 7238 18437
rect 7286 18411 7290 18437
rect 7214 18410 7238 18411
rect 7266 18410 7290 18411
rect 7318 18437 7342 18438
rect 7370 18437 7394 18438
rect 7318 18411 7322 18437
rect 7370 18411 7384 18437
rect 7318 18410 7342 18411
rect 7370 18410 7394 18411
rect 7422 18410 7446 18438
rect 7474 18410 7498 18438
rect 7526 18437 7535 18438
rect 7534 18411 7535 18437
rect 7526 18410 7535 18411
rect 7073 18405 7535 18410
rect 12073 18438 12535 18443
rect 12073 18437 12082 18438
rect 12073 18411 12074 18437
rect 12073 18410 12082 18411
rect 12110 18410 12134 18438
rect 12162 18410 12186 18438
rect 12214 18437 12238 18438
rect 12266 18437 12290 18438
rect 12224 18411 12238 18437
rect 12286 18411 12290 18437
rect 12214 18410 12238 18411
rect 12266 18410 12290 18411
rect 12318 18437 12342 18438
rect 12370 18437 12394 18438
rect 12318 18411 12322 18437
rect 12370 18411 12384 18437
rect 12318 18410 12342 18411
rect 12370 18410 12394 18411
rect 12422 18410 12446 18438
rect 12474 18410 12498 18438
rect 12526 18437 12535 18438
rect 12534 18411 12535 18437
rect 12526 18410 12535 18411
rect 12073 18405 12535 18410
rect 12614 18354 12642 18494
rect 12558 18326 12642 18354
rect 9573 18046 10035 18051
rect 9573 18045 9582 18046
rect 9573 18019 9574 18045
rect 9573 18018 9582 18019
rect 9610 18018 9634 18046
rect 9662 18018 9686 18046
rect 9714 18045 9738 18046
rect 9766 18045 9790 18046
rect 9724 18019 9738 18045
rect 9786 18019 9790 18045
rect 9714 18018 9738 18019
rect 9766 18018 9790 18019
rect 9818 18045 9842 18046
rect 9870 18045 9894 18046
rect 9818 18019 9822 18045
rect 9870 18019 9884 18045
rect 9818 18018 9842 18019
rect 9870 18018 9894 18019
rect 9922 18018 9946 18046
rect 9974 18018 9998 18046
rect 10026 18045 10035 18046
rect 10034 18019 10035 18045
rect 10026 18018 10035 18019
rect 9573 18013 10035 18018
rect 12558 17738 12586 18326
rect 14573 18046 15035 18051
rect 14573 18045 14582 18046
rect 14573 18019 14574 18045
rect 14573 18018 14582 18019
rect 14610 18018 14634 18046
rect 14662 18018 14686 18046
rect 14714 18045 14738 18046
rect 14766 18045 14790 18046
rect 14724 18019 14738 18045
rect 14786 18019 14790 18045
rect 14714 18018 14738 18019
rect 14766 18018 14790 18019
rect 14818 18045 14842 18046
rect 14870 18045 14894 18046
rect 14818 18019 14822 18045
rect 14870 18019 14884 18045
rect 14818 18018 14842 18019
rect 14870 18018 14894 18019
rect 14922 18018 14946 18046
rect 14974 18018 14998 18046
rect 15026 18045 15035 18046
rect 15034 18019 15035 18045
rect 15026 18018 15035 18019
rect 14573 18013 15035 18018
rect 12558 17710 12642 17738
rect 7073 17654 7535 17659
rect 7073 17653 7082 17654
rect 7073 17627 7074 17653
rect 7073 17626 7082 17627
rect 7110 17626 7134 17654
rect 7162 17626 7186 17654
rect 7214 17653 7238 17654
rect 7266 17653 7290 17654
rect 7224 17627 7238 17653
rect 7286 17627 7290 17653
rect 7214 17626 7238 17627
rect 7266 17626 7290 17627
rect 7318 17653 7342 17654
rect 7370 17653 7394 17654
rect 7318 17627 7322 17653
rect 7370 17627 7384 17653
rect 7318 17626 7342 17627
rect 7370 17626 7394 17627
rect 7422 17626 7446 17654
rect 7474 17626 7498 17654
rect 7526 17653 7535 17654
rect 7534 17627 7535 17653
rect 7526 17626 7535 17627
rect 7073 17621 7535 17626
rect 12073 17654 12535 17659
rect 12073 17653 12082 17654
rect 12073 17627 12074 17653
rect 12073 17626 12082 17627
rect 12110 17626 12134 17654
rect 12162 17626 12186 17654
rect 12214 17653 12238 17654
rect 12266 17653 12290 17654
rect 12224 17627 12238 17653
rect 12286 17627 12290 17653
rect 12214 17626 12238 17627
rect 12266 17626 12290 17627
rect 12318 17653 12342 17654
rect 12370 17653 12394 17654
rect 12318 17627 12322 17653
rect 12370 17627 12384 17653
rect 12318 17626 12342 17627
rect 12370 17626 12394 17627
rect 12422 17626 12446 17654
rect 12474 17626 12498 17654
rect 12526 17653 12535 17654
rect 12534 17627 12535 17653
rect 12526 17626 12535 17627
rect 12073 17621 12535 17626
rect 12502 17457 12530 17463
rect 12502 17431 12503 17457
rect 12529 17431 12530 17457
rect 9573 17262 10035 17267
rect 9573 17261 9582 17262
rect 9573 17235 9574 17261
rect 9573 17234 9582 17235
rect 9610 17234 9634 17262
rect 9662 17234 9686 17262
rect 9714 17261 9738 17262
rect 9766 17261 9790 17262
rect 9724 17235 9738 17261
rect 9786 17235 9790 17261
rect 9714 17234 9738 17235
rect 9766 17234 9790 17235
rect 9818 17261 9842 17262
rect 9870 17261 9894 17262
rect 9818 17235 9822 17261
rect 9870 17235 9884 17261
rect 9818 17234 9842 17235
rect 9870 17234 9894 17235
rect 9922 17234 9946 17262
rect 9974 17234 9998 17262
rect 10026 17261 10035 17262
rect 10034 17235 10035 17261
rect 10026 17234 10035 17235
rect 9573 17229 10035 17234
rect 10598 17121 10626 17127
rect 10598 17095 10599 17121
rect 10625 17095 10626 17121
rect 9646 17065 9674 17071
rect 9646 17039 9647 17065
rect 9673 17039 9674 17065
rect 7073 16870 7535 16875
rect 7073 16869 7082 16870
rect 7073 16843 7074 16869
rect 7073 16842 7082 16843
rect 7110 16842 7134 16870
rect 7162 16842 7186 16870
rect 7214 16869 7238 16870
rect 7266 16869 7290 16870
rect 7224 16843 7238 16869
rect 7286 16843 7290 16869
rect 7214 16842 7238 16843
rect 7266 16842 7290 16843
rect 7318 16869 7342 16870
rect 7370 16869 7394 16870
rect 7318 16843 7322 16869
rect 7370 16843 7384 16869
rect 7318 16842 7342 16843
rect 7370 16842 7394 16843
rect 7422 16842 7446 16870
rect 7474 16842 7498 16870
rect 7526 16869 7535 16870
rect 7534 16843 7535 16869
rect 7526 16842 7535 16843
rect 7073 16837 7535 16842
rect 9534 16674 9562 16679
rect 9646 16674 9674 17039
rect 9310 16673 9674 16674
rect 9310 16647 9535 16673
rect 9561 16647 9674 16673
rect 9310 16646 9674 16647
rect 10430 17065 10458 17071
rect 10430 17039 10431 17065
rect 10457 17039 10458 17065
rect 10430 16673 10458 17039
rect 10430 16647 10431 16673
rect 10457 16647 10458 16673
rect 7014 16311 7015 16337
rect 7041 16311 7042 16337
rect 5894 16282 5922 16287
rect 5894 15974 5922 16254
rect 6118 16282 6146 16287
rect 6118 16235 6146 16254
rect 7014 16281 7042 16311
rect 8358 16337 8386 16343
rect 8358 16311 8359 16337
rect 8385 16311 8386 16337
rect 7014 16255 7015 16281
rect 7041 16255 7042 16281
rect 7014 15974 7042 16255
rect 7518 16282 7546 16287
rect 7518 16170 7546 16254
rect 8358 16281 8386 16311
rect 8358 16255 8359 16281
rect 8385 16255 8386 16281
rect 7518 16142 7602 16170
rect 7073 16086 7535 16091
rect 7073 16085 7082 16086
rect 7073 16059 7074 16085
rect 7073 16058 7082 16059
rect 7110 16058 7134 16086
rect 7162 16058 7186 16086
rect 7214 16085 7238 16086
rect 7266 16085 7290 16086
rect 7224 16059 7238 16085
rect 7286 16059 7290 16085
rect 7214 16058 7238 16059
rect 7266 16058 7290 16059
rect 7318 16085 7342 16086
rect 7370 16085 7394 16086
rect 7318 16059 7322 16085
rect 7370 16059 7384 16085
rect 7318 16058 7342 16059
rect 7370 16058 7394 16059
rect 7422 16058 7446 16086
rect 7474 16058 7498 16086
rect 7526 16085 7535 16086
rect 7534 16059 7535 16085
rect 7526 16058 7535 16059
rect 7073 16053 7535 16058
rect 5838 15946 5922 15974
rect 6902 15946 7042 15974
rect 5278 15889 5306 15895
rect 5278 15863 5279 15889
rect 5305 15863 5306 15889
rect 4573 15694 5035 15699
rect 4573 15693 4582 15694
rect 4573 15667 4574 15693
rect 4573 15666 4582 15667
rect 4610 15666 4634 15694
rect 4662 15666 4686 15694
rect 4714 15693 4738 15694
rect 4766 15693 4790 15694
rect 4724 15667 4738 15693
rect 4786 15667 4790 15693
rect 4714 15666 4738 15667
rect 4766 15666 4790 15667
rect 4818 15693 4842 15694
rect 4870 15693 4894 15694
rect 4818 15667 4822 15693
rect 4870 15667 4884 15693
rect 4818 15666 4842 15667
rect 4870 15666 4894 15667
rect 4922 15666 4946 15694
rect 4974 15666 4998 15694
rect 5026 15693 5035 15694
rect 5034 15667 5035 15693
rect 5026 15666 5035 15667
rect 4573 15661 5035 15666
rect 3822 15105 3850 15111
rect 3822 15079 3823 15105
rect 3849 15079 3850 15105
rect 3038 14714 3066 14719
rect 3038 13929 3066 14686
rect 3598 14714 3626 14719
rect 3822 14714 3850 15079
rect 4382 15106 4410 15111
rect 4494 15106 4522 15111
rect 4382 15105 4522 15106
rect 4382 15079 4383 15105
rect 4409 15079 4495 15105
rect 4521 15079 4522 15105
rect 4382 15078 4522 15079
rect 4382 15073 4410 15078
rect 3626 14686 3850 14714
rect 3598 14648 3626 14686
rect 3822 14658 3850 14686
rect 3822 14625 3850 14630
rect 4494 14769 4522 15078
rect 5278 15105 5306 15863
rect 5278 15079 5279 15105
rect 5305 15079 5306 15105
rect 4573 14910 5035 14915
rect 4573 14909 4582 14910
rect 4573 14883 4574 14909
rect 4573 14882 4582 14883
rect 4610 14882 4634 14910
rect 4662 14882 4686 14910
rect 4714 14909 4738 14910
rect 4766 14909 4790 14910
rect 4724 14883 4738 14909
rect 4786 14883 4790 14909
rect 4714 14882 4738 14883
rect 4766 14882 4790 14883
rect 4818 14909 4842 14910
rect 4870 14909 4894 14910
rect 4818 14883 4822 14909
rect 4870 14883 4884 14909
rect 4818 14882 4842 14883
rect 4870 14882 4894 14883
rect 4922 14882 4946 14910
rect 4974 14882 4998 14910
rect 5026 14909 5035 14910
rect 5034 14883 5035 14909
rect 5026 14882 5035 14883
rect 4573 14877 5035 14882
rect 4494 14743 4495 14769
rect 4521 14743 4522 14769
rect 4494 14713 4522 14743
rect 4494 14687 4495 14713
rect 4521 14687 4522 14713
rect 4494 14378 4522 14687
rect 5278 14714 5306 15079
rect 3822 14322 3850 14327
rect 3038 13903 3039 13929
rect 3065 13903 3066 13929
rect 3038 13897 3066 13903
rect 3374 13929 3402 13935
rect 3374 13903 3375 13929
rect 3401 13903 3402 13929
rect 3374 13426 3402 13903
rect 2394 13145 2674 13146
rect 2394 13119 2591 13145
rect 2617 13119 2674 13145
rect 2394 13118 2674 13119
rect 2366 13080 2394 13118
rect 2590 13113 2618 13118
rect 2073 12950 2535 12955
rect 2073 12949 2082 12950
rect 2073 12923 2074 12949
rect 2073 12922 2082 12923
rect 2110 12922 2134 12950
rect 2162 12922 2186 12950
rect 2214 12949 2238 12950
rect 2266 12949 2290 12950
rect 2224 12923 2238 12949
rect 2286 12923 2290 12949
rect 2214 12922 2238 12923
rect 2266 12922 2290 12923
rect 2318 12949 2342 12950
rect 2370 12949 2394 12950
rect 2318 12923 2322 12949
rect 2370 12923 2384 12949
rect 2318 12922 2342 12923
rect 2370 12922 2394 12923
rect 2422 12922 2446 12950
rect 2474 12922 2498 12950
rect 2526 12949 2535 12950
rect 2534 12923 2535 12949
rect 2526 12922 2535 12923
rect 2073 12917 2535 12922
rect 1806 12753 2002 12754
rect 1806 12727 1807 12753
rect 1833 12727 1975 12753
rect 2001 12727 2002 12753
rect 1806 12726 2002 12727
rect 1806 12721 1834 12726
rect 1974 12721 2002 12726
rect 2198 12753 2226 12759
rect 2198 12727 2199 12753
rect 2225 12727 2226 12753
rect 2198 12698 2226 12727
rect 2198 12642 2226 12670
rect 1974 12614 2226 12642
rect 2646 12642 2674 13118
rect 1638 12558 1890 12586
rect 1862 12417 1890 12558
rect 1862 12391 1863 12417
rect 1889 12391 1890 12417
rect 1862 12361 1890 12391
rect 1862 12335 1863 12361
rect 1889 12335 1890 12361
rect 1806 11970 1834 11975
rect 1862 11970 1890 12335
rect 1918 11970 1946 11975
rect 1806 11969 1946 11970
rect 1806 11943 1807 11969
rect 1833 11943 1919 11969
rect 1945 11943 1946 11969
rect 1806 11942 1946 11943
rect 1806 11937 1834 11942
rect 1862 11633 1890 11942
rect 1918 11937 1946 11942
rect 1974 11970 2002 12614
rect 2646 12609 2674 12614
rect 2758 13146 2786 13151
rect 2758 12698 2786 13118
rect 3318 13146 3346 13151
rect 3374 13146 3402 13398
rect 3822 13537 3850 14294
rect 4494 13985 4522 14350
rect 4998 14378 5026 14383
rect 4998 14321 5026 14350
rect 4998 14295 4999 14321
rect 5025 14295 5026 14321
rect 4998 14265 5026 14295
rect 5278 14322 5306 14686
rect 5838 15497 5866 15946
rect 5838 15471 5839 15497
rect 5865 15471 5866 15497
rect 5838 14714 5866 15471
rect 6454 15889 6482 15895
rect 6454 15863 6455 15889
rect 6481 15863 6482 15889
rect 6454 15833 6482 15863
rect 6454 15807 6455 15833
rect 6481 15807 6482 15833
rect 6398 15105 6426 15111
rect 6398 15079 6399 15105
rect 6425 15079 6426 15105
rect 6398 15049 6426 15079
rect 6398 15023 6399 15049
rect 6425 15023 6426 15049
rect 5838 14667 5866 14686
rect 6006 14770 6034 14775
rect 5278 14275 5306 14294
rect 4998 14239 4999 14265
rect 5025 14239 5026 14265
rect 4998 14233 5026 14239
rect 4573 14126 5035 14131
rect 4573 14125 4582 14126
rect 4573 14099 4574 14125
rect 4573 14098 4582 14099
rect 4610 14098 4634 14126
rect 4662 14098 4686 14126
rect 4714 14125 4738 14126
rect 4766 14125 4790 14126
rect 4724 14099 4738 14125
rect 4786 14099 4790 14125
rect 4714 14098 4738 14099
rect 4766 14098 4790 14099
rect 4818 14125 4842 14126
rect 4870 14125 4894 14126
rect 4818 14099 4822 14125
rect 4870 14099 4884 14125
rect 4818 14098 4842 14099
rect 4870 14098 4894 14099
rect 4922 14098 4946 14126
rect 4974 14098 4998 14126
rect 5026 14125 5035 14126
rect 5034 14099 5035 14125
rect 5026 14098 5035 14099
rect 4573 14093 5035 14098
rect 4494 13959 4495 13985
rect 4521 13959 4522 13985
rect 4494 13929 4522 13959
rect 4494 13903 4495 13929
rect 4521 13903 4522 13929
rect 3822 13511 3823 13537
rect 3849 13511 3850 13537
rect 3822 13426 3850 13511
rect 3822 13393 3850 13398
rect 4102 13538 4130 13543
rect 3346 13118 3402 13146
rect 3318 13099 3346 13118
rect 2758 12361 2786 12670
rect 4102 12753 4130 13510
rect 4382 13538 4410 13543
rect 4494 13538 4522 13903
rect 5838 13930 5866 13935
rect 4382 13537 4522 13538
rect 4382 13511 4383 13537
rect 4409 13511 4495 13537
rect 4521 13511 4522 13537
rect 4382 13510 4522 13511
rect 4382 13505 4410 13510
rect 4494 13201 4522 13510
rect 5278 13538 5306 13543
rect 5278 13491 5306 13510
rect 5838 13538 5866 13902
rect 5838 13505 5866 13510
rect 4573 13342 5035 13347
rect 4573 13341 4582 13342
rect 4573 13315 4574 13341
rect 4573 13314 4582 13315
rect 4610 13314 4634 13342
rect 4662 13314 4686 13342
rect 4714 13341 4738 13342
rect 4766 13341 4790 13342
rect 4724 13315 4738 13341
rect 4786 13315 4790 13341
rect 4714 13314 4738 13315
rect 4766 13314 4790 13315
rect 4818 13341 4842 13342
rect 4870 13341 4894 13342
rect 4818 13315 4822 13341
rect 4870 13315 4884 13341
rect 4818 13314 4842 13315
rect 4870 13314 4894 13315
rect 4922 13314 4946 13342
rect 4974 13314 4998 13342
rect 5026 13341 5035 13342
rect 5034 13315 5035 13341
rect 5026 13314 5035 13315
rect 4573 13309 5035 13314
rect 4494 13175 4495 13201
rect 4521 13175 4522 13201
rect 4494 13145 4522 13175
rect 4494 13119 4495 13145
rect 4521 13119 4522 13145
rect 4102 12727 4103 12753
rect 4129 12727 4130 12753
rect 2758 12335 2759 12361
rect 2785 12335 2786 12361
rect 2758 12329 2786 12335
rect 3038 12362 3066 12367
rect 2073 12166 2535 12171
rect 2073 12165 2082 12166
rect 2073 12139 2074 12165
rect 2073 12138 2082 12139
rect 2110 12138 2134 12166
rect 2162 12138 2186 12166
rect 2214 12165 2238 12166
rect 2266 12165 2290 12166
rect 2224 12139 2238 12165
rect 2286 12139 2290 12165
rect 2214 12138 2238 12139
rect 2266 12138 2290 12139
rect 2318 12165 2342 12166
rect 2370 12165 2394 12166
rect 2318 12139 2322 12165
rect 2370 12139 2384 12165
rect 2318 12138 2342 12139
rect 2370 12138 2394 12139
rect 2422 12138 2446 12166
rect 2474 12138 2498 12166
rect 2526 12165 2535 12166
rect 2534 12139 2535 12165
rect 2526 12138 2535 12139
rect 2073 12133 2535 12138
rect 2198 11970 2226 11975
rect 1974 11969 2226 11970
rect 1974 11943 2199 11969
rect 2225 11943 2226 11969
rect 1974 11942 2226 11943
rect 1862 11607 1863 11633
rect 1889 11607 1890 11633
rect 1862 11577 1890 11607
rect 1862 11551 1863 11577
rect 1889 11551 1890 11577
rect 1806 11186 1834 11191
rect 1862 11186 1890 11551
rect 1918 11186 1946 11191
rect 1638 11185 1946 11186
rect 1638 11159 1807 11185
rect 1833 11159 1919 11185
rect 1945 11159 1946 11185
rect 1638 11158 1946 11159
rect 1638 10402 1666 11158
rect 1806 11153 1834 11158
rect 1918 11153 1946 11158
rect 1526 10401 1666 10402
rect 1526 10375 1639 10401
rect 1665 10375 1666 10401
rect 1526 10374 1666 10375
rect 1526 10345 1554 10374
rect 1526 10319 1527 10345
rect 1553 10319 1554 10345
rect 1526 10313 1554 10319
rect 1638 9226 1666 10374
rect 1862 10794 1890 10799
rect 1862 10065 1890 10766
rect 1862 10039 1863 10065
rect 1889 10039 1890 10065
rect 1862 10009 1890 10039
rect 1862 9983 1863 10009
rect 1889 9983 1890 10009
rect 1638 9193 1666 9198
rect 1806 9618 1834 9623
rect 1862 9618 1890 9983
rect 1806 9617 1890 9618
rect 1806 9591 1807 9617
rect 1833 9591 1890 9617
rect 1806 9590 1890 9591
rect 1414 8833 1442 8839
rect 1414 8807 1415 8833
rect 1441 8807 1442 8833
rect 1414 8777 1442 8807
rect 1414 8751 1415 8777
rect 1441 8751 1442 8777
rect 1414 8442 1442 8751
rect 1358 3346 1386 3351
rect 1414 3346 1442 8414
rect 1806 8049 1834 9590
rect 1918 9338 1946 9343
rect 1862 9281 1890 9287
rect 1862 9255 1863 9281
rect 1889 9255 1890 9281
rect 1862 9226 1890 9255
rect 1862 8497 1890 9198
rect 1862 8471 1863 8497
rect 1889 8471 1890 8497
rect 1862 8442 1890 8471
rect 1862 8395 1890 8414
rect 1806 8023 1807 8049
rect 1833 8023 1834 8049
rect 1526 7994 1554 7999
rect 1806 7994 1834 8023
rect 1526 7993 1834 7994
rect 1526 7967 1527 7993
rect 1553 7967 1834 7993
rect 1526 7966 1834 7967
rect 1526 7209 1554 7966
rect 1526 7183 1527 7209
rect 1553 7183 1554 7209
rect 1526 6425 1554 7183
rect 1526 6399 1527 6425
rect 1553 6399 1554 6425
rect 1526 6393 1554 6399
rect 1806 7714 1834 7966
rect 1862 7714 1890 7719
rect 1806 7713 1890 7714
rect 1806 7687 1863 7713
rect 1889 7687 1890 7713
rect 1806 7686 1890 7687
rect 1806 7265 1834 7686
rect 1862 7657 1890 7686
rect 1862 7631 1863 7657
rect 1889 7631 1890 7657
rect 1862 7625 1890 7631
rect 1806 7239 1807 7265
rect 1833 7239 1834 7265
rect 1806 6930 1834 7239
rect 1862 6930 1890 6935
rect 1806 6929 1890 6930
rect 1806 6903 1863 6929
rect 1889 6903 1890 6929
rect 1806 6902 1890 6903
rect 1806 6481 1834 6902
rect 1862 6873 1890 6902
rect 1862 6847 1863 6873
rect 1889 6847 1890 6873
rect 1862 6841 1890 6847
rect 1806 6455 1807 6481
rect 1833 6455 1834 6481
rect 1806 6146 1834 6455
rect 1918 6482 1946 9310
rect 1918 6449 1946 6454
rect 1862 6146 1890 6151
rect 1806 6145 1890 6146
rect 1806 6119 1863 6145
rect 1889 6119 1890 6145
rect 1806 6118 1890 6119
rect 1806 5698 1834 6118
rect 1862 6089 1890 6118
rect 1862 6063 1863 6089
rect 1889 6063 1890 6089
rect 1862 6057 1890 6063
rect 1918 5698 1946 5703
rect 1806 5697 1946 5698
rect 1806 5671 1807 5697
rect 1833 5671 1919 5697
rect 1945 5671 1946 5697
rect 1806 5670 1946 5671
rect 1806 5665 1834 5670
rect 1862 5361 1890 5670
rect 1918 5665 1946 5670
rect 1862 5335 1863 5361
rect 1889 5335 1890 5361
rect 1862 5306 1890 5335
rect 1806 5305 1890 5306
rect 1806 5279 1863 5305
rect 1889 5279 1890 5305
rect 1806 5278 1890 5279
rect 1806 4914 1834 5278
rect 1862 5273 1890 5278
rect 1918 4914 1946 4919
rect 1806 4913 1946 4914
rect 1806 4887 1807 4913
rect 1833 4887 1919 4913
rect 1945 4887 1946 4913
rect 1806 4886 1946 4887
rect 1806 4881 1834 4886
rect 1862 4577 1890 4886
rect 1918 4881 1946 4886
rect 1862 4551 1863 4577
rect 1889 4551 1890 4577
rect 1862 4522 1890 4551
rect 1862 4521 1946 4522
rect 1862 4495 1863 4521
rect 1889 4495 1946 4521
rect 1862 4494 1946 4495
rect 1862 4489 1890 4494
rect 1806 4130 1834 4135
rect 1806 4083 1834 4102
rect 1918 4130 1946 4494
rect 1918 4097 1946 4102
rect 1358 3345 1442 3346
rect 1358 3319 1359 3345
rect 1385 3319 1442 3345
rect 1358 3318 1442 3319
rect 1918 3626 1946 3631
rect 1358 3289 1386 3318
rect 1358 3263 1359 3289
rect 1385 3263 1386 3289
rect 1358 3257 1386 3263
rect 1190 2674 1218 2679
rect 1190 1777 1218 2646
rect 1638 2561 1666 2567
rect 1638 2535 1639 2561
rect 1665 2535 1666 2561
rect 1526 2506 1554 2511
rect 1638 2506 1666 2535
rect 1526 2505 1666 2506
rect 1526 2479 1527 2505
rect 1553 2479 1666 2505
rect 1526 2478 1666 2479
rect 1526 2473 1554 2478
rect 1638 2226 1666 2478
rect 1638 2193 1666 2198
rect 1190 1751 1191 1777
rect 1217 1751 1218 1777
rect 854 462 1050 490
rect 854 400 882 462
rect 840 0 896 400
rect 1022 378 1050 462
rect 1190 378 1218 1751
rect 1918 1777 1946 3598
rect 1974 3346 2002 11942
rect 2198 11937 2226 11942
rect 3038 11577 3066 12334
rect 3598 12362 3626 12367
rect 3598 12315 3626 12334
rect 4102 12362 4130 12727
rect 4382 12754 4410 12759
rect 4494 12754 4522 13119
rect 5838 13145 5866 13151
rect 5838 13119 5839 13145
rect 5865 13119 5866 13145
rect 4382 12753 4522 12754
rect 4382 12727 4383 12753
rect 4409 12727 4495 12753
rect 4521 12727 4522 12753
rect 4382 12726 4522 12727
rect 4382 12721 4410 12726
rect 4102 12329 4130 12334
rect 4326 12586 4354 12591
rect 4102 11970 4130 11975
rect 4102 11923 4130 11942
rect 4326 11970 4354 12558
rect 4494 12417 4522 12726
rect 5278 12753 5306 12759
rect 5278 12727 5279 12753
rect 5305 12727 5306 12753
rect 4573 12558 5035 12563
rect 4573 12557 4582 12558
rect 4573 12531 4574 12557
rect 4573 12530 4582 12531
rect 4610 12530 4634 12558
rect 4662 12530 4686 12558
rect 4714 12557 4738 12558
rect 4766 12557 4790 12558
rect 4724 12531 4738 12557
rect 4786 12531 4790 12557
rect 4714 12530 4738 12531
rect 4766 12530 4790 12531
rect 4818 12557 4842 12558
rect 4870 12557 4894 12558
rect 4818 12531 4822 12557
rect 4870 12531 4884 12557
rect 4818 12530 4842 12531
rect 4870 12530 4894 12531
rect 4922 12530 4946 12558
rect 4974 12530 4998 12558
rect 5026 12557 5035 12558
rect 5034 12531 5035 12557
rect 5026 12530 5035 12531
rect 4573 12525 5035 12530
rect 4494 12391 4495 12417
rect 4521 12391 4522 12417
rect 4494 12361 4522 12391
rect 4494 12335 4495 12361
rect 4521 12335 4522 12361
rect 4494 12329 4522 12335
rect 4494 11970 4522 11975
rect 4326 11969 4522 11970
rect 4326 11943 4327 11969
rect 4353 11943 4495 11969
rect 4521 11943 4522 11969
rect 4326 11942 4522 11943
rect 4326 11937 4354 11942
rect 4438 11633 4466 11942
rect 4494 11937 4522 11942
rect 5278 11970 5306 12727
rect 4573 11774 5035 11779
rect 4573 11773 4582 11774
rect 4573 11747 4574 11773
rect 4573 11746 4582 11747
rect 4610 11746 4634 11774
rect 4662 11746 4686 11774
rect 4714 11773 4738 11774
rect 4766 11773 4790 11774
rect 4724 11747 4738 11773
rect 4786 11747 4790 11773
rect 4714 11746 4738 11747
rect 4766 11746 4790 11747
rect 4818 11773 4842 11774
rect 4870 11773 4894 11774
rect 4818 11747 4822 11773
rect 4870 11747 4884 11773
rect 4818 11746 4842 11747
rect 4870 11746 4894 11747
rect 4922 11746 4946 11774
rect 4974 11746 4998 11774
rect 5026 11773 5035 11774
rect 5034 11747 5035 11773
rect 5026 11746 5035 11747
rect 4573 11741 5035 11746
rect 4438 11607 4439 11633
rect 4465 11607 4466 11633
rect 3038 11551 3039 11577
rect 3065 11551 3066 11577
rect 2073 11382 2535 11387
rect 2073 11381 2082 11382
rect 2073 11355 2074 11381
rect 2073 11354 2082 11355
rect 2110 11354 2134 11382
rect 2162 11354 2186 11382
rect 2214 11381 2238 11382
rect 2266 11381 2290 11382
rect 2224 11355 2238 11381
rect 2286 11355 2290 11381
rect 2214 11354 2238 11355
rect 2266 11354 2290 11355
rect 2318 11381 2342 11382
rect 2370 11381 2394 11382
rect 2318 11355 2322 11381
rect 2370 11355 2384 11381
rect 2318 11354 2342 11355
rect 2370 11354 2394 11355
rect 2422 11354 2446 11382
rect 2474 11354 2498 11382
rect 2526 11381 2535 11382
rect 2534 11355 2535 11381
rect 2526 11354 2535 11355
rect 2073 11349 2535 11354
rect 2478 11185 2506 11191
rect 2478 11159 2479 11185
rect 2505 11159 2506 11185
rect 2478 10906 2506 11159
rect 2478 10873 2506 10878
rect 2590 10906 2618 10911
rect 2086 10849 2114 10855
rect 2086 10823 2087 10849
rect 2113 10823 2114 10849
rect 2086 10794 2114 10823
rect 2086 10728 2114 10766
rect 2073 10598 2535 10603
rect 2073 10597 2082 10598
rect 2073 10571 2074 10597
rect 2073 10570 2082 10571
rect 2110 10570 2134 10598
rect 2162 10570 2186 10598
rect 2214 10597 2238 10598
rect 2266 10597 2290 10598
rect 2224 10571 2238 10597
rect 2286 10571 2290 10597
rect 2214 10570 2238 10571
rect 2266 10570 2290 10571
rect 2318 10597 2342 10598
rect 2370 10597 2394 10598
rect 2318 10571 2322 10597
rect 2370 10571 2384 10597
rect 2318 10570 2342 10571
rect 2370 10570 2394 10571
rect 2422 10570 2446 10598
rect 2474 10570 2498 10598
rect 2526 10597 2535 10598
rect 2534 10571 2535 10597
rect 2526 10570 2535 10571
rect 2073 10565 2535 10570
rect 2478 10402 2506 10407
rect 2590 10402 2618 10878
rect 3038 10906 3066 11551
rect 3038 10793 3066 10878
rect 3038 10767 3039 10793
rect 3065 10767 3066 10793
rect 3038 10761 3066 10767
rect 3598 11577 3626 11583
rect 3598 11551 3599 11577
rect 3625 11551 3626 11577
rect 3598 11186 3626 11551
rect 4438 11577 4466 11607
rect 4438 11551 4439 11577
rect 4465 11551 4466 11577
rect 3822 11186 3850 11191
rect 3598 11185 3850 11186
rect 3598 11159 3823 11185
rect 3849 11159 3850 11185
rect 3598 11158 3850 11159
rect 3598 10793 3626 11158
rect 3598 10767 3599 10793
rect 3625 10767 3626 10793
rect 2478 10401 2618 10402
rect 2478 10375 2479 10401
rect 2505 10375 2618 10401
rect 2478 10374 2618 10375
rect 2478 10369 2506 10374
rect 2590 10094 2618 10374
rect 2590 10066 2786 10094
rect 2073 9814 2535 9819
rect 2073 9813 2082 9814
rect 2073 9787 2074 9813
rect 2073 9786 2082 9787
rect 2110 9786 2134 9814
rect 2162 9786 2186 9814
rect 2214 9813 2238 9814
rect 2266 9813 2290 9814
rect 2224 9787 2238 9813
rect 2286 9787 2290 9813
rect 2214 9786 2238 9787
rect 2266 9786 2290 9787
rect 2318 9813 2342 9814
rect 2370 9813 2394 9814
rect 2318 9787 2322 9813
rect 2370 9787 2384 9813
rect 2318 9786 2342 9787
rect 2370 9786 2394 9787
rect 2422 9786 2446 9814
rect 2474 9786 2498 9814
rect 2526 9813 2535 9814
rect 2534 9787 2535 9813
rect 2526 9786 2535 9787
rect 2073 9781 2535 9786
rect 2030 9617 2058 9623
rect 2030 9591 2031 9617
rect 2057 9591 2058 9617
rect 2030 9282 2058 9591
rect 2478 9618 2506 9623
rect 2590 9618 2618 10066
rect 2758 10009 2786 10066
rect 2758 9983 2759 10009
rect 2785 9983 2786 10009
rect 2758 9977 2786 9983
rect 3598 10009 3626 10767
rect 3822 10402 3850 11158
rect 4382 11186 4410 11191
rect 4438 11186 4466 11551
rect 4494 11186 4522 11191
rect 4382 11185 4522 11186
rect 4382 11159 4383 11185
rect 4409 11159 4495 11185
rect 4521 11159 4522 11185
rect 4382 11158 4522 11159
rect 4382 11153 4410 11158
rect 4438 10849 4466 11158
rect 4494 11153 4522 11158
rect 5278 11185 5306 11942
rect 5278 11159 5279 11185
rect 5305 11159 5306 11185
rect 4573 10990 5035 10995
rect 4573 10989 4582 10990
rect 4573 10963 4574 10989
rect 4573 10962 4582 10963
rect 4610 10962 4634 10990
rect 4662 10962 4686 10990
rect 4714 10989 4738 10990
rect 4766 10989 4790 10990
rect 4724 10963 4738 10989
rect 4786 10963 4790 10989
rect 4714 10962 4738 10963
rect 4766 10962 4790 10963
rect 4818 10989 4842 10990
rect 4870 10989 4894 10990
rect 4818 10963 4822 10989
rect 4870 10963 4884 10989
rect 4818 10962 4842 10963
rect 4870 10962 4894 10963
rect 4922 10962 4946 10990
rect 4974 10962 4998 10990
rect 5026 10989 5035 10990
rect 5034 10963 5035 10989
rect 5026 10962 5035 10963
rect 4573 10957 5035 10962
rect 4438 10823 4439 10849
rect 4465 10823 4466 10849
rect 4438 10793 4466 10823
rect 4438 10767 4439 10793
rect 4465 10767 4466 10793
rect 4382 10402 4410 10407
rect 4438 10402 4466 10767
rect 5278 10794 5306 11159
rect 4494 10402 4522 10407
rect 3822 10336 3850 10374
rect 4214 10401 4522 10402
rect 4214 10375 4383 10401
rect 4409 10375 4495 10401
rect 4521 10375 4522 10401
rect 4214 10374 4522 10375
rect 4214 10066 4242 10374
rect 4382 10369 4410 10374
rect 4494 10369 4522 10374
rect 5278 10402 5306 10766
rect 5838 12361 5866 13119
rect 5838 12335 5839 12361
rect 5865 12335 5866 12361
rect 5838 11577 5866 12335
rect 5838 11551 5839 11577
rect 5865 11551 5866 11577
rect 5838 10962 5866 11551
rect 5838 10794 5866 10934
rect 5838 10747 5866 10766
rect 4573 10206 5035 10211
rect 4573 10205 4582 10206
rect 4573 10179 4574 10205
rect 4573 10178 4582 10179
rect 4610 10178 4634 10206
rect 4662 10178 4686 10206
rect 4714 10205 4738 10206
rect 4766 10205 4790 10206
rect 4724 10179 4738 10205
rect 4786 10179 4790 10205
rect 4714 10178 4738 10179
rect 4766 10178 4790 10179
rect 4818 10205 4842 10206
rect 4870 10205 4894 10206
rect 4818 10179 4822 10205
rect 4870 10179 4884 10205
rect 4818 10178 4842 10179
rect 4870 10178 4894 10179
rect 4922 10178 4946 10206
rect 4974 10178 4998 10206
rect 5026 10205 5035 10206
rect 5034 10179 5035 10205
rect 5026 10178 5035 10179
rect 4573 10173 5035 10178
rect 3990 10038 4242 10066
rect 3598 9983 3599 10009
rect 3625 9983 3626 10009
rect 3598 9977 3626 9983
rect 3822 10010 3850 10015
rect 3990 10010 4018 10038
rect 3822 10009 4018 10010
rect 3822 9983 3823 10009
rect 3849 9983 3991 10009
rect 4017 9983 4018 10009
rect 3822 9982 4018 9983
rect 2478 9617 2618 9618
rect 2478 9591 2479 9617
rect 2505 9591 2618 9617
rect 2478 9590 2618 9591
rect 3822 9618 3850 9982
rect 3990 9977 4018 9982
rect 2478 9338 2506 9590
rect 2478 9305 2506 9310
rect 3822 9561 3850 9590
rect 3822 9535 3823 9561
rect 3849 9535 3850 9561
rect 2030 9249 2058 9254
rect 3374 9282 3402 9287
rect 3038 9225 3066 9231
rect 3038 9199 3039 9225
rect 3065 9199 3066 9225
rect 2073 9030 2535 9035
rect 2073 9029 2082 9030
rect 2073 9003 2074 9029
rect 2073 9002 2082 9003
rect 2110 9002 2134 9030
rect 2162 9002 2186 9030
rect 2214 9029 2238 9030
rect 2266 9029 2290 9030
rect 2224 9003 2238 9029
rect 2286 9003 2290 9029
rect 2214 9002 2238 9003
rect 2266 9002 2290 9003
rect 2318 9029 2342 9030
rect 2370 9029 2394 9030
rect 2318 9003 2322 9029
rect 2370 9003 2384 9029
rect 2318 9002 2342 9003
rect 2370 9002 2394 9003
rect 2422 9002 2446 9030
rect 2474 9002 2498 9030
rect 2526 9029 2535 9030
rect 2534 9003 2535 9029
rect 2526 9002 2535 9003
rect 2073 8997 2535 9002
rect 2478 8834 2506 8839
rect 2478 8833 2618 8834
rect 2478 8807 2479 8833
rect 2505 8807 2618 8833
rect 2478 8806 2618 8807
rect 2478 8801 2506 8806
rect 2073 8246 2535 8251
rect 2073 8245 2082 8246
rect 2073 8219 2074 8245
rect 2073 8218 2082 8219
rect 2110 8218 2134 8246
rect 2162 8218 2186 8246
rect 2214 8245 2238 8246
rect 2266 8245 2290 8246
rect 2224 8219 2238 8245
rect 2286 8219 2290 8245
rect 2214 8218 2238 8219
rect 2266 8218 2290 8219
rect 2318 8245 2342 8246
rect 2370 8245 2394 8246
rect 2318 8219 2322 8245
rect 2370 8219 2384 8245
rect 2318 8218 2342 8219
rect 2370 8218 2394 8219
rect 2422 8218 2446 8246
rect 2474 8218 2498 8246
rect 2526 8245 2535 8246
rect 2534 8219 2535 8245
rect 2526 8218 2535 8219
rect 2073 8213 2535 8218
rect 2478 8050 2506 8055
rect 2590 8050 2618 8806
rect 2478 8049 2618 8050
rect 2478 8023 2479 8049
rect 2505 8023 2618 8049
rect 2478 8022 2618 8023
rect 2478 8017 2506 8022
rect 2073 7462 2535 7467
rect 2073 7461 2082 7462
rect 2073 7435 2074 7461
rect 2073 7434 2082 7435
rect 2110 7434 2134 7462
rect 2162 7434 2186 7462
rect 2214 7461 2238 7462
rect 2266 7461 2290 7462
rect 2224 7435 2238 7461
rect 2286 7435 2290 7461
rect 2214 7434 2238 7435
rect 2266 7434 2290 7435
rect 2318 7461 2342 7462
rect 2370 7461 2394 7462
rect 2318 7435 2322 7461
rect 2370 7435 2384 7461
rect 2318 7434 2342 7435
rect 2370 7434 2394 7435
rect 2422 7434 2446 7462
rect 2474 7434 2498 7462
rect 2526 7461 2535 7462
rect 2534 7435 2535 7461
rect 2526 7434 2535 7435
rect 2073 7429 2535 7434
rect 2478 7266 2506 7271
rect 2478 7219 2506 7238
rect 2590 7266 2618 8022
rect 2590 7233 2618 7238
rect 3038 8441 3066 9199
rect 3374 9225 3402 9254
rect 3374 9199 3375 9225
rect 3401 9199 3402 9225
rect 3374 9193 3402 9199
rect 3822 9282 3850 9535
rect 3822 8833 3850 9254
rect 3822 8807 3823 8833
rect 3849 8807 3850 8833
rect 3822 8777 3850 8807
rect 3822 8751 3823 8777
rect 3849 8751 3850 8777
rect 3038 8415 3039 8441
rect 3065 8415 3066 8441
rect 3038 7657 3066 8415
rect 3038 7631 3039 7657
rect 3065 7631 3066 7657
rect 3038 7266 3066 7631
rect 3038 6874 3066 7238
rect 3038 6827 3066 6846
rect 3598 8441 3626 8447
rect 3598 8415 3599 8441
rect 3625 8415 3626 8441
rect 3598 7657 3626 8415
rect 3598 7631 3599 7657
rect 3625 7631 3626 7657
rect 3598 6874 3626 7631
rect 2073 6678 2535 6683
rect 2073 6677 2082 6678
rect 2073 6651 2074 6677
rect 2073 6650 2082 6651
rect 2110 6650 2134 6678
rect 2162 6650 2186 6678
rect 2214 6677 2238 6678
rect 2266 6677 2290 6678
rect 2224 6651 2238 6677
rect 2286 6651 2290 6677
rect 2214 6650 2238 6651
rect 2266 6650 2290 6651
rect 2318 6677 2342 6678
rect 2370 6677 2394 6678
rect 2318 6651 2322 6677
rect 2370 6651 2384 6677
rect 2318 6650 2342 6651
rect 2370 6650 2394 6651
rect 2422 6650 2446 6678
rect 2474 6650 2498 6678
rect 2526 6677 2535 6678
rect 2534 6651 2535 6677
rect 2526 6650 2535 6651
rect 2073 6645 2535 6650
rect 2198 6482 2226 6487
rect 2198 6435 2226 6454
rect 2758 6482 2786 6487
rect 2758 6090 2786 6454
rect 2590 6089 2786 6090
rect 2590 6063 2759 6089
rect 2785 6063 2786 6089
rect 2590 6062 2786 6063
rect 2073 5894 2535 5899
rect 2073 5893 2082 5894
rect 2073 5867 2074 5893
rect 2073 5866 2082 5867
rect 2110 5866 2134 5894
rect 2162 5866 2186 5894
rect 2214 5893 2238 5894
rect 2266 5893 2290 5894
rect 2224 5867 2238 5893
rect 2286 5867 2290 5893
rect 2214 5866 2238 5867
rect 2266 5866 2290 5867
rect 2318 5893 2342 5894
rect 2370 5893 2394 5894
rect 2318 5867 2322 5893
rect 2370 5867 2384 5893
rect 2318 5866 2342 5867
rect 2370 5866 2394 5867
rect 2422 5866 2446 5894
rect 2474 5866 2498 5894
rect 2526 5893 2535 5894
rect 2534 5867 2535 5893
rect 2526 5866 2535 5867
rect 2073 5861 2535 5866
rect 2478 5698 2506 5703
rect 2590 5698 2618 6062
rect 2478 5697 2618 5698
rect 2478 5671 2479 5697
rect 2505 5671 2618 5697
rect 2478 5670 2618 5671
rect 2478 5665 2506 5670
rect 2073 5110 2535 5115
rect 2073 5109 2082 5110
rect 2073 5083 2074 5109
rect 2073 5082 2082 5083
rect 2110 5082 2134 5110
rect 2162 5082 2186 5110
rect 2214 5109 2238 5110
rect 2266 5109 2290 5110
rect 2224 5083 2238 5109
rect 2286 5083 2290 5109
rect 2214 5082 2238 5083
rect 2266 5082 2290 5083
rect 2318 5109 2342 5110
rect 2370 5109 2394 5110
rect 2318 5083 2322 5109
rect 2370 5083 2384 5109
rect 2318 5082 2342 5083
rect 2370 5082 2394 5083
rect 2422 5082 2446 5110
rect 2474 5082 2498 5110
rect 2526 5109 2535 5110
rect 2534 5083 2535 5109
rect 2526 5082 2535 5083
rect 2073 5077 2535 5082
rect 2478 4914 2506 4919
rect 2590 4914 2618 5670
rect 2478 4913 2618 4914
rect 2478 4887 2479 4913
rect 2505 4887 2618 4913
rect 2478 4886 2618 4887
rect 2478 4881 2506 4886
rect 2073 4326 2535 4331
rect 2073 4325 2082 4326
rect 2073 4299 2074 4325
rect 2073 4298 2082 4299
rect 2110 4298 2134 4326
rect 2162 4298 2186 4326
rect 2214 4325 2238 4326
rect 2266 4325 2290 4326
rect 2224 4299 2238 4325
rect 2286 4299 2290 4325
rect 2214 4298 2238 4299
rect 2266 4298 2290 4299
rect 2318 4325 2342 4326
rect 2370 4325 2394 4326
rect 2318 4299 2322 4325
rect 2370 4299 2384 4325
rect 2318 4298 2342 4299
rect 2370 4298 2394 4299
rect 2422 4298 2446 4326
rect 2474 4298 2498 4326
rect 2526 4325 2535 4326
rect 2534 4299 2535 4325
rect 2526 4298 2535 4299
rect 2073 4293 2535 4298
rect 2590 4214 2618 4886
rect 2758 5305 2786 6062
rect 3598 6089 3626 6846
rect 3822 6874 3850 8751
rect 4046 9954 4074 9959
rect 3990 6874 4018 6879
rect 3822 6873 4018 6874
rect 3822 6847 3823 6873
rect 3849 6847 3991 6873
rect 4017 6847 4018 6873
rect 3822 6846 4018 6847
rect 3822 6841 3850 6846
rect 3990 6538 4018 6846
rect 3598 6063 3599 6089
rect 3625 6063 3626 6089
rect 3598 6057 3626 6063
rect 3878 6090 3906 6095
rect 3990 6090 4018 6510
rect 3878 6089 4018 6090
rect 3878 6063 3879 6089
rect 3905 6063 3991 6089
rect 4017 6063 4018 6089
rect 3878 6062 4018 6063
rect 3878 6057 3906 6062
rect 3990 6057 4018 6062
rect 2758 5279 2759 5305
rect 2785 5279 2786 5305
rect 2758 4522 2786 5279
rect 3598 5306 3626 5311
rect 3598 5259 3626 5278
rect 2758 4456 2786 4494
rect 2982 4522 3010 4527
rect 2478 4186 2618 4214
rect 2030 4130 2058 4135
rect 2030 3626 2058 4102
rect 2478 4129 2506 4186
rect 2478 4103 2479 4129
rect 2505 4103 2506 4129
rect 2478 4097 2506 4103
rect 2366 3738 2394 3743
rect 2478 3738 2506 3743
rect 2366 3737 2506 3738
rect 2366 3711 2367 3737
rect 2393 3711 2479 3737
rect 2505 3711 2506 3737
rect 2366 3710 2506 3711
rect 2366 3705 2394 3710
rect 2030 3593 2058 3598
rect 2478 3626 2506 3710
rect 2982 3737 3010 4494
rect 3318 4522 3346 4527
rect 3318 4475 3346 4494
rect 3598 4522 3626 4527
rect 2982 3711 2983 3737
rect 3009 3711 3010 3737
rect 2982 3705 3010 3711
rect 3262 3794 3290 3799
rect 2478 3593 2506 3598
rect 2073 3542 2535 3547
rect 2073 3541 2082 3542
rect 2073 3515 2074 3541
rect 2073 3514 2082 3515
rect 2110 3514 2134 3542
rect 2162 3514 2186 3542
rect 2214 3541 2238 3542
rect 2266 3541 2290 3542
rect 2224 3515 2238 3541
rect 2286 3515 2290 3541
rect 2214 3514 2238 3515
rect 2266 3514 2290 3515
rect 2318 3541 2342 3542
rect 2370 3541 2394 3542
rect 2318 3515 2322 3541
rect 2370 3515 2384 3541
rect 2318 3514 2342 3515
rect 2370 3514 2394 3515
rect 2422 3514 2446 3542
rect 2474 3514 2498 3542
rect 2526 3541 2535 3542
rect 2534 3515 2535 3541
rect 2526 3514 2535 3515
rect 2073 3509 2535 3514
rect 2478 3346 2506 3351
rect 1974 3345 2506 3346
rect 1974 3319 2479 3345
rect 2505 3319 2506 3345
rect 1974 3318 2506 3319
rect 1974 3009 2002 3015
rect 1974 2983 1975 3009
rect 2001 2983 2002 3009
rect 1974 2953 2002 2983
rect 1974 2927 1975 2953
rect 2001 2927 2002 2953
rect 1974 2562 2002 2927
rect 2478 2842 2506 3318
rect 3038 2953 3066 2959
rect 3038 2927 3039 2953
rect 3065 2927 3066 2953
rect 2478 2814 2618 2842
rect 2073 2758 2535 2763
rect 2073 2757 2082 2758
rect 2073 2731 2074 2757
rect 2073 2730 2082 2731
rect 2110 2730 2134 2758
rect 2162 2730 2186 2758
rect 2214 2757 2238 2758
rect 2266 2757 2290 2758
rect 2224 2731 2238 2757
rect 2286 2731 2290 2757
rect 2214 2730 2238 2731
rect 2266 2730 2290 2731
rect 2318 2757 2342 2758
rect 2370 2757 2394 2758
rect 2318 2731 2322 2757
rect 2370 2731 2384 2757
rect 2318 2730 2342 2731
rect 2370 2730 2394 2731
rect 2422 2730 2446 2758
rect 2474 2730 2498 2758
rect 2526 2757 2535 2758
rect 2534 2731 2535 2757
rect 2526 2730 2535 2731
rect 2073 2725 2535 2730
rect 2478 2618 2506 2623
rect 1974 2529 2002 2534
rect 2366 2562 2394 2567
rect 2366 2170 2394 2534
rect 2478 2561 2506 2590
rect 2478 2535 2479 2561
rect 2505 2535 2506 2561
rect 2478 2529 2506 2535
rect 2590 2282 2618 2814
rect 3038 2618 3066 2927
rect 3038 2585 3066 2590
rect 2590 2249 2618 2254
rect 2478 2170 2506 2175
rect 2366 2169 2506 2170
rect 2366 2143 2367 2169
rect 2393 2143 2479 2169
rect 2505 2143 2506 2169
rect 2366 2142 2506 2143
rect 2366 2137 2394 2142
rect 2478 2137 2506 2142
rect 3038 2170 3066 2175
rect 3038 2123 3066 2142
rect 2073 1974 2535 1979
rect 2073 1973 2082 1974
rect 2073 1947 2074 1973
rect 2073 1946 2082 1947
rect 2110 1946 2134 1974
rect 2162 1946 2186 1974
rect 2214 1973 2238 1974
rect 2266 1973 2290 1974
rect 2224 1947 2238 1973
rect 2286 1947 2290 1973
rect 2214 1946 2238 1947
rect 2266 1946 2290 1947
rect 2318 1973 2342 1974
rect 2370 1973 2394 1974
rect 2318 1947 2322 1973
rect 2370 1947 2384 1973
rect 2318 1946 2342 1947
rect 2370 1946 2394 1947
rect 2422 1946 2446 1974
rect 2474 1946 2498 1974
rect 2526 1973 2535 1974
rect 2534 1947 2535 1973
rect 2526 1946 2535 1947
rect 2073 1941 2535 1946
rect 1918 1751 1919 1777
rect 1945 1751 1946 1777
rect 1918 1721 1946 1751
rect 1918 1695 1919 1721
rect 1945 1695 1946 1721
rect 1918 1689 1946 1695
rect 2086 1890 2114 1895
rect 3262 1890 3290 3766
rect 3598 3737 3626 4494
rect 4046 4214 4074 9926
rect 4998 9617 5026 9623
rect 4998 9591 4999 9617
rect 5025 9591 5026 9617
rect 4998 9506 5026 9591
rect 5278 9617 5306 10374
rect 5278 9591 5279 9617
rect 5305 9591 5306 9617
rect 5278 9585 5306 9591
rect 5446 10738 5474 10743
rect 4998 9478 5138 9506
rect 4573 9422 5035 9427
rect 4573 9421 4582 9422
rect 4573 9395 4574 9421
rect 4573 9394 4582 9395
rect 4610 9394 4634 9422
rect 4662 9394 4686 9422
rect 4714 9421 4738 9422
rect 4766 9421 4790 9422
rect 4724 9395 4738 9421
rect 4786 9395 4790 9421
rect 4714 9394 4738 9395
rect 4766 9394 4790 9395
rect 4818 9421 4842 9422
rect 4870 9421 4894 9422
rect 4818 9395 4822 9421
rect 4870 9395 4884 9421
rect 4818 9394 4842 9395
rect 4870 9394 4894 9395
rect 4922 9394 4946 9422
rect 4974 9394 4998 9422
rect 5026 9421 5035 9422
rect 5034 9395 5035 9421
rect 5026 9394 5035 9395
rect 4573 9389 5035 9394
rect 4494 9226 4522 9231
rect 4494 9179 4522 9198
rect 5110 9226 5138 9478
rect 4998 8834 5026 8839
rect 4998 8787 5026 8806
rect 5110 8834 5138 9198
rect 5110 8801 5138 8806
rect 4573 8638 5035 8643
rect 4573 8637 4582 8638
rect 4573 8611 4574 8637
rect 4573 8610 4582 8611
rect 4610 8610 4634 8638
rect 4662 8610 4686 8638
rect 4714 8637 4738 8638
rect 4766 8637 4790 8638
rect 4724 8611 4738 8637
rect 4786 8611 4790 8637
rect 4714 8610 4738 8611
rect 4766 8610 4790 8611
rect 4818 8637 4842 8638
rect 4870 8637 4894 8638
rect 4818 8611 4822 8637
rect 4870 8611 4884 8637
rect 4818 8610 4842 8611
rect 4870 8610 4894 8611
rect 4922 8610 4946 8638
rect 4974 8610 4998 8638
rect 5026 8637 5035 8638
rect 5034 8611 5035 8637
rect 5026 8610 5035 8611
rect 4573 8605 5035 8610
rect 4494 8497 4522 8503
rect 4494 8471 4495 8497
rect 4521 8471 4522 8497
rect 4494 8442 4522 8471
rect 4102 8049 4130 8055
rect 4102 8023 4103 8049
rect 4129 8023 4130 8049
rect 4102 7265 4130 8023
rect 4382 8050 4410 8055
rect 4494 8050 4522 8414
rect 4382 8049 4522 8050
rect 4382 8023 4383 8049
rect 4409 8023 4495 8049
rect 4521 8023 4522 8049
rect 4382 8022 4522 8023
rect 4382 8017 4410 8022
rect 4102 7239 4103 7265
rect 4129 7239 4130 7265
rect 4102 6874 4130 7239
rect 4494 7713 4522 8022
rect 4573 7854 5035 7859
rect 4573 7853 4582 7854
rect 4573 7827 4574 7853
rect 4573 7826 4582 7827
rect 4610 7826 4634 7854
rect 4662 7826 4686 7854
rect 4714 7853 4738 7854
rect 4766 7853 4790 7854
rect 4724 7827 4738 7853
rect 4786 7827 4790 7853
rect 4714 7826 4738 7827
rect 4766 7826 4790 7827
rect 4818 7853 4842 7854
rect 4870 7853 4894 7854
rect 4818 7827 4822 7853
rect 4870 7827 4884 7853
rect 4818 7826 4842 7827
rect 4870 7826 4894 7827
rect 4922 7826 4946 7854
rect 4974 7826 4998 7854
rect 5026 7853 5035 7854
rect 5034 7827 5035 7853
rect 5026 7826 5035 7827
rect 4573 7821 5035 7826
rect 4494 7687 4495 7713
rect 4521 7687 4522 7713
rect 4494 7657 4522 7687
rect 4494 7631 4495 7657
rect 4521 7631 4522 7657
rect 4494 7210 4522 7631
rect 4494 7177 4522 7182
rect 4998 7265 5026 7271
rect 4998 7239 4999 7265
rect 5025 7239 5026 7265
rect 4998 7210 5026 7239
rect 4998 7163 5026 7182
rect 4573 7070 5035 7075
rect 4573 7069 4582 7070
rect 4573 7043 4574 7069
rect 4573 7042 4582 7043
rect 4610 7042 4634 7070
rect 4662 7042 4686 7070
rect 4714 7069 4738 7070
rect 4766 7069 4790 7070
rect 4724 7043 4738 7069
rect 4786 7043 4790 7069
rect 4714 7042 4738 7043
rect 4766 7042 4790 7043
rect 4818 7069 4842 7070
rect 4870 7069 4894 7070
rect 4818 7043 4822 7069
rect 4870 7043 4884 7069
rect 4818 7042 4842 7043
rect 4870 7042 4894 7043
rect 4922 7042 4946 7070
rect 4974 7042 4998 7070
rect 5026 7069 5035 7070
rect 5034 7043 5035 7069
rect 5026 7042 5035 7043
rect 4573 7037 5035 7042
rect 4102 6482 4130 6846
rect 4102 6435 4130 6454
rect 4270 6538 4298 6543
rect 4270 6482 4298 6510
rect 4494 6482 4522 6487
rect 4270 6481 4522 6482
rect 4270 6455 4271 6481
rect 4297 6455 4495 6481
rect 4521 6455 4522 6481
rect 4270 6454 4522 6455
rect 4270 6449 4298 6454
rect 4102 5697 4130 5703
rect 4102 5671 4103 5697
rect 4129 5671 4130 5697
rect 4102 5306 4130 5671
rect 4382 5698 4410 6454
rect 4494 6449 4522 6454
rect 4573 6286 5035 6291
rect 4573 6285 4582 6286
rect 4573 6259 4574 6285
rect 4573 6258 4582 6259
rect 4610 6258 4634 6286
rect 4662 6258 4686 6286
rect 4714 6285 4738 6286
rect 4766 6285 4790 6286
rect 4724 6259 4738 6285
rect 4786 6259 4790 6285
rect 4714 6258 4738 6259
rect 4766 6258 4790 6259
rect 4818 6285 4842 6286
rect 4870 6285 4894 6286
rect 4818 6259 4822 6285
rect 4870 6259 4884 6285
rect 4818 6258 4842 6259
rect 4870 6258 4894 6259
rect 4922 6258 4946 6286
rect 4974 6258 4998 6286
rect 5026 6285 5035 6286
rect 5034 6259 5035 6285
rect 5026 6258 5035 6259
rect 4573 6253 5035 6258
rect 4494 5698 4522 5703
rect 4382 5697 4522 5698
rect 4382 5671 4383 5697
rect 4409 5671 4495 5697
rect 4521 5671 4522 5697
rect 4382 5670 4522 5671
rect 4382 5665 4410 5670
rect 4102 5082 4130 5278
rect 4102 4913 4130 5054
rect 4438 5361 4466 5670
rect 4494 5665 4522 5670
rect 4573 5502 5035 5507
rect 4573 5501 4582 5502
rect 4573 5475 4574 5501
rect 4573 5474 4582 5475
rect 4610 5474 4634 5502
rect 4662 5474 4686 5502
rect 4714 5501 4738 5502
rect 4766 5501 4790 5502
rect 4724 5475 4738 5501
rect 4786 5475 4790 5501
rect 4714 5474 4738 5475
rect 4766 5474 4790 5475
rect 4818 5501 4842 5502
rect 4870 5501 4894 5502
rect 4818 5475 4822 5501
rect 4870 5475 4884 5501
rect 4818 5474 4842 5475
rect 4870 5474 4894 5475
rect 4922 5474 4946 5502
rect 4974 5474 4998 5502
rect 5026 5501 5035 5502
rect 5034 5475 5035 5501
rect 5026 5474 5035 5475
rect 4573 5469 5035 5474
rect 4438 5335 4439 5361
rect 4465 5335 4466 5361
rect 4438 5305 4466 5335
rect 4438 5279 4439 5305
rect 4465 5279 4466 5305
rect 4102 4887 4103 4913
rect 4129 4887 4130 4913
rect 4102 4881 4130 4887
rect 4382 4914 4410 4919
rect 4438 4914 4466 5279
rect 4494 4914 4522 4919
rect 4382 4913 4522 4914
rect 4382 4887 4383 4913
rect 4409 4887 4495 4913
rect 4521 4887 4522 4913
rect 4382 4886 4522 4887
rect 4382 4881 4410 4886
rect 4438 4577 4466 4886
rect 4494 4881 4522 4886
rect 4573 4718 5035 4723
rect 4573 4717 4582 4718
rect 4573 4691 4574 4717
rect 4573 4690 4582 4691
rect 4610 4690 4634 4718
rect 4662 4690 4686 4718
rect 4714 4717 4738 4718
rect 4766 4717 4790 4718
rect 4724 4691 4738 4717
rect 4786 4691 4790 4717
rect 4714 4690 4738 4691
rect 4766 4690 4790 4691
rect 4818 4717 4842 4718
rect 4870 4717 4894 4718
rect 4818 4691 4822 4717
rect 4870 4691 4884 4717
rect 4818 4690 4842 4691
rect 4870 4690 4894 4691
rect 4922 4690 4946 4718
rect 4974 4690 4998 4718
rect 5026 4717 5035 4718
rect 5034 4691 5035 4717
rect 5026 4690 5035 4691
rect 4573 4685 5035 4690
rect 4438 4551 4439 4577
rect 4465 4551 4466 4577
rect 4438 4522 4466 4551
rect 3598 3711 3599 3737
rect 3625 3711 3626 3737
rect 3598 2953 3626 3711
rect 3598 2927 3599 2953
rect 3625 2927 3626 2953
rect 3542 2618 3570 2623
rect 3542 2169 3570 2590
rect 3598 2450 3626 2927
rect 3598 2417 3626 2422
rect 3934 4186 4074 4214
rect 4270 4521 4466 4522
rect 4270 4495 4439 4521
rect 4465 4495 4466 4521
rect 4270 4494 4466 4495
rect 4270 4186 4298 4494
rect 4438 4489 4466 4494
rect 5278 4242 5306 4247
rect 3542 2143 3543 2169
rect 3569 2143 3570 2169
rect 3262 1862 3346 1890
rect 2086 400 2114 1862
rect 3318 400 3346 1862
rect 3542 1777 3570 2143
rect 3934 1890 3962 4186
rect 4270 4153 4298 4158
rect 4494 4186 4522 4191
rect 4102 4129 4130 4135
rect 4102 4103 4103 4129
rect 4129 4103 4130 4129
rect 4102 3345 4130 4103
rect 4494 3793 4522 4158
rect 4998 4186 5026 4191
rect 4998 4129 5026 4158
rect 4998 4103 4999 4129
rect 5025 4103 5026 4129
rect 4998 4073 5026 4103
rect 5278 4129 5306 4214
rect 5278 4103 5279 4129
rect 5305 4103 5306 4129
rect 5278 4097 5306 4103
rect 4998 4047 4999 4073
rect 5025 4047 5026 4073
rect 4998 4041 5026 4047
rect 4573 3934 5035 3939
rect 4573 3933 4582 3934
rect 4573 3907 4574 3933
rect 4573 3906 4582 3907
rect 4610 3906 4634 3934
rect 4662 3906 4686 3934
rect 4714 3933 4738 3934
rect 4766 3933 4790 3934
rect 4724 3907 4738 3933
rect 4786 3907 4790 3933
rect 4714 3906 4738 3907
rect 4766 3906 4790 3907
rect 4818 3933 4842 3934
rect 4870 3933 4894 3934
rect 4818 3907 4822 3933
rect 4870 3907 4884 3933
rect 4818 3906 4842 3907
rect 4870 3906 4894 3907
rect 4922 3906 4946 3934
rect 4974 3906 4998 3934
rect 5026 3933 5035 3934
rect 5034 3907 5035 3933
rect 5026 3906 5035 3907
rect 4573 3901 5035 3906
rect 4494 3767 4495 3793
rect 4521 3767 4522 3793
rect 4494 3737 4522 3767
rect 4494 3711 4495 3737
rect 4521 3711 4522 3737
rect 4494 3626 4522 3711
rect 4102 3319 4103 3345
rect 4129 3319 4130 3345
rect 4046 2618 4074 2623
rect 4046 2561 4074 2590
rect 4046 2535 4047 2561
rect 4073 2535 4074 2561
rect 4046 2529 4074 2535
rect 4102 2450 4130 3319
rect 4382 3346 4410 3351
rect 4494 3346 4522 3598
rect 4382 3345 4522 3346
rect 4382 3319 4383 3345
rect 4409 3319 4495 3345
rect 4521 3319 4522 3345
rect 4382 3318 4522 3319
rect 4382 3313 4410 3318
rect 4494 3009 4522 3318
rect 4573 3150 5035 3155
rect 4573 3149 4582 3150
rect 4573 3123 4574 3149
rect 4573 3122 4582 3123
rect 4610 3122 4634 3150
rect 4662 3122 4686 3150
rect 4714 3149 4738 3150
rect 4766 3149 4790 3150
rect 4724 3123 4738 3149
rect 4786 3123 4790 3149
rect 4714 3122 4738 3123
rect 4766 3122 4790 3123
rect 4818 3149 4842 3150
rect 4870 3149 4894 3150
rect 4818 3123 4822 3149
rect 4870 3123 4884 3149
rect 4818 3122 4842 3123
rect 4870 3122 4894 3123
rect 4922 3122 4946 3150
rect 4974 3122 4998 3150
rect 5026 3149 5035 3150
rect 5034 3123 5035 3149
rect 5026 3122 5035 3123
rect 4573 3117 5035 3122
rect 4494 2983 4495 3009
rect 4521 2983 4522 3009
rect 4494 2953 4522 2983
rect 4494 2927 4495 2953
rect 4521 2927 4522 2953
rect 4494 2921 4522 2927
rect 5446 2674 5474 10710
rect 5894 10009 5922 10015
rect 5894 9983 5895 10009
rect 5921 9983 5922 10009
rect 5558 8834 5586 8839
rect 5558 8049 5586 8806
rect 5894 8834 5922 9983
rect 5950 9618 5978 9623
rect 5950 9571 5978 9590
rect 5894 8801 5922 8806
rect 5558 8023 5559 8049
rect 5585 8023 5586 8049
rect 5558 7658 5586 8023
rect 5558 7625 5586 7630
rect 5558 7265 5586 7271
rect 5558 7239 5559 7265
rect 5585 7239 5586 7265
rect 5558 7154 5586 7239
rect 6006 7154 6034 14742
rect 6398 14378 6426 15023
rect 6398 14321 6426 14350
rect 6398 14295 6399 14321
rect 6425 14295 6426 14321
rect 6398 14265 6426 14295
rect 6398 14239 6399 14265
rect 6425 14239 6426 14265
rect 6398 13538 6426 14239
rect 6398 13481 6426 13510
rect 6398 13455 6399 13481
rect 6425 13455 6426 13481
rect 6398 13449 6426 13455
rect 6454 13482 6482 15807
rect 6902 15553 6930 15946
rect 6902 15527 6903 15553
rect 6929 15527 6930 15553
rect 6902 15497 6930 15527
rect 6902 15471 6903 15497
rect 6929 15471 6930 15497
rect 6902 14769 6930 15471
rect 6902 14743 6903 14769
rect 6929 14743 6930 14769
rect 6902 14713 6930 14743
rect 6902 14687 6903 14713
rect 6929 14687 6930 14713
rect 6454 12753 6482 13454
rect 6454 12727 6455 12753
rect 6481 12727 6482 12753
rect 6454 12697 6482 12727
rect 6454 12671 6455 12697
rect 6481 12671 6482 12697
rect 6398 11969 6426 11975
rect 6398 11943 6399 11969
rect 6425 11943 6426 11969
rect 6398 11913 6426 11943
rect 6398 11887 6399 11913
rect 6425 11887 6426 11913
rect 6398 11802 6426 11887
rect 6398 11769 6426 11774
rect 6454 11185 6482 12671
rect 6454 11159 6455 11185
rect 6481 11159 6482 11185
rect 6454 11129 6482 11159
rect 6454 11103 6455 11129
rect 6481 11103 6482 11129
rect 6454 10401 6482 11103
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 6454 10345 6482 10375
rect 6454 10319 6455 10345
rect 6481 10319 6482 10345
rect 6230 9618 6258 9623
rect 6230 9562 6258 9590
rect 6230 9561 6314 9562
rect 6230 9535 6231 9561
rect 6257 9535 6314 9561
rect 6230 9534 6314 9535
rect 6230 9529 6258 9534
rect 6118 9225 6146 9231
rect 6118 9199 6119 9225
rect 6145 9199 6146 9225
rect 6118 8442 6146 9199
rect 6286 9226 6314 9534
rect 6454 9226 6482 10319
rect 6846 14658 6874 14663
rect 6846 10094 6874 14630
rect 6902 13985 6930 14687
rect 7014 15498 7042 15503
rect 7014 14714 7042 15470
rect 7294 15498 7322 15503
rect 7294 15451 7322 15470
rect 7073 15302 7535 15307
rect 7073 15301 7082 15302
rect 7073 15275 7074 15301
rect 7073 15274 7082 15275
rect 7110 15274 7134 15302
rect 7162 15274 7186 15302
rect 7214 15301 7238 15302
rect 7266 15301 7290 15302
rect 7224 15275 7238 15301
rect 7286 15275 7290 15301
rect 7214 15274 7238 15275
rect 7266 15274 7290 15275
rect 7318 15301 7342 15302
rect 7370 15301 7394 15302
rect 7318 15275 7322 15301
rect 7370 15275 7384 15301
rect 7318 15274 7342 15275
rect 7370 15274 7394 15275
rect 7422 15274 7446 15302
rect 7474 15274 7498 15302
rect 7526 15301 7535 15302
rect 7534 15275 7535 15301
rect 7526 15274 7535 15275
rect 7073 15269 7535 15274
rect 7574 15050 7602 16142
rect 7798 15890 7826 15895
rect 7798 15498 7826 15862
rect 7798 15465 7826 15470
rect 8358 15890 8386 16255
rect 8470 15890 8498 15895
rect 8358 15889 8498 15890
rect 8358 15863 8359 15889
rect 8385 15863 8471 15889
rect 8497 15863 8498 15889
rect 8358 15862 8498 15863
rect 8358 15553 8386 15862
rect 8470 15857 8498 15862
rect 9254 15889 9282 15895
rect 9254 15863 9255 15889
rect 9281 15863 9282 15889
rect 8358 15527 8359 15553
rect 8385 15527 8386 15553
rect 8358 15497 8386 15527
rect 8358 15471 8359 15497
rect 8385 15471 8386 15497
rect 7574 15017 7602 15022
rect 7798 15105 7826 15111
rect 7798 15079 7799 15105
rect 7825 15079 7826 15105
rect 7294 14714 7322 14719
rect 7014 14713 7322 14714
rect 7014 14687 7295 14713
rect 7321 14687 7322 14713
rect 7014 14686 7322 14687
rect 6902 13959 6903 13985
rect 6929 13959 6930 13985
rect 6902 13929 6930 13959
rect 6902 13903 6903 13929
rect 6929 13903 6930 13929
rect 6902 13538 6930 13903
rect 6902 12418 6930 13510
rect 6958 13986 6986 13991
rect 6958 13482 6986 13958
rect 7014 13930 7042 14686
rect 7294 14681 7322 14686
rect 7073 14518 7535 14523
rect 7073 14517 7082 14518
rect 7073 14491 7074 14517
rect 7073 14490 7082 14491
rect 7110 14490 7134 14518
rect 7162 14490 7186 14518
rect 7214 14517 7238 14518
rect 7266 14517 7290 14518
rect 7224 14491 7238 14517
rect 7286 14491 7290 14517
rect 7214 14490 7238 14491
rect 7266 14490 7290 14491
rect 7318 14517 7342 14518
rect 7370 14517 7394 14518
rect 7318 14491 7322 14517
rect 7370 14491 7384 14517
rect 7318 14490 7342 14491
rect 7370 14490 7394 14491
rect 7422 14490 7446 14518
rect 7474 14490 7498 14518
rect 7526 14517 7535 14518
rect 7534 14491 7535 14517
rect 7526 14490 7535 14491
rect 7073 14485 7535 14490
rect 7798 14321 7826 15079
rect 8358 14769 8386 15471
rect 9254 15498 9282 15863
rect 9310 15890 9338 16646
rect 9534 16641 9562 16646
rect 10430 16618 10458 16647
rect 10598 16618 10626 17095
rect 12054 17121 12082 17127
rect 12054 17095 12055 17121
rect 12081 17095 12082 17121
rect 11102 17065 11130 17071
rect 11102 17039 11103 17065
rect 11129 17039 11130 17065
rect 10934 16673 10962 16679
rect 10934 16647 10935 16673
rect 10961 16647 10962 16673
rect 10430 16617 10906 16618
rect 10430 16591 10431 16617
rect 10457 16591 10906 16617
rect 10430 16590 10906 16591
rect 10430 16585 10458 16590
rect 9573 16478 10035 16483
rect 9573 16477 9582 16478
rect 9573 16451 9574 16477
rect 9573 16450 9582 16451
rect 9610 16450 9634 16478
rect 9662 16450 9686 16478
rect 9714 16477 9738 16478
rect 9766 16477 9790 16478
rect 9724 16451 9738 16477
rect 9786 16451 9790 16477
rect 9714 16450 9738 16451
rect 9766 16450 9790 16451
rect 9818 16477 9842 16478
rect 9870 16477 9894 16478
rect 9818 16451 9822 16477
rect 9870 16451 9884 16477
rect 9818 16450 9842 16451
rect 9870 16450 9894 16451
rect 9922 16450 9946 16478
rect 9974 16450 9998 16478
rect 10026 16477 10035 16478
rect 10034 16451 10035 16477
rect 10026 16450 10035 16451
rect 9573 16445 10035 16450
rect 10150 16338 10178 16343
rect 9310 15857 9338 15862
rect 9478 16282 9506 16287
rect 9478 15498 9506 16254
rect 9982 16282 10010 16287
rect 9982 16235 10010 16254
rect 10150 15889 10178 16310
rect 10822 16338 10850 16343
rect 10822 16281 10850 16310
rect 10822 16255 10823 16281
rect 10849 16255 10850 16281
rect 10822 16249 10850 16255
rect 10150 15863 10151 15889
rect 10177 15863 10178 15889
rect 10150 15834 10178 15863
rect 10206 15834 10234 15839
rect 10150 15833 10234 15834
rect 10150 15807 10207 15833
rect 10233 15807 10234 15833
rect 10150 15806 10234 15807
rect 9573 15694 10035 15699
rect 9573 15693 9582 15694
rect 9573 15667 9574 15693
rect 9573 15666 9582 15667
rect 9610 15666 9634 15694
rect 9662 15666 9686 15694
rect 9714 15693 9738 15694
rect 9766 15693 9790 15694
rect 9724 15667 9738 15693
rect 9786 15667 9790 15693
rect 9714 15666 9738 15667
rect 9766 15666 9790 15667
rect 9818 15693 9842 15694
rect 9870 15693 9894 15694
rect 9818 15667 9822 15693
rect 9870 15667 9884 15693
rect 9818 15666 9842 15667
rect 9870 15666 9894 15667
rect 9922 15666 9946 15694
rect 9974 15666 9998 15694
rect 10026 15693 10035 15694
rect 10034 15667 10035 15693
rect 10026 15666 10035 15667
rect 9573 15661 10035 15666
rect 9814 15498 9842 15503
rect 9254 15497 9842 15498
rect 9254 15471 9815 15497
rect 9841 15471 9842 15497
rect 9254 15470 9842 15471
rect 8358 14743 8359 14769
rect 8385 14743 8386 14769
rect 8358 14714 8386 14743
rect 8974 15106 9002 15111
rect 8974 15049 9002 15078
rect 8974 15023 8975 15049
rect 9001 15023 9002 15049
rect 8358 14713 8442 14714
rect 8358 14687 8359 14713
rect 8385 14687 8442 14713
rect 8358 14686 8442 14687
rect 8358 14681 8386 14686
rect 7798 14295 7799 14321
rect 7825 14295 7826 14321
rect 7014 13897 7042 13902
rect 7574 13929 7602 13935
rect 7574 13903 7575 13929
rect 7601 13903 7602 13929
rect 7073 13734 7535 13739
rect 7073 13733 7082 13734
rect 7073 13707 7074 13733
rect 7073 13706 7082 13707
rect 7110 13706 7134 13734
rect 7162 13706 7186 13734
rect 7214 13733 7238 13734
rect 7266 13733 7290 13734
rect 7224 13707 7238 13733
rect 7286 13707 7290 13733
rect 7214 13706 7238 13707
rect 7266 13706 7290 13707
rect 7318 13733 7342 13734
rect 7370 13733 7394 13734
rect 7318 13707 7322 13733
rect 7370 13707 7384 13733
rect 7318 13706 7342 13707
rect 7370 13706 7394 13707
rect 7422 13706 7446 13734
rect 7474 13706 7498 13734
rect 7526 13733 7535 13734
rect 7534 13707 7535 13733
rect 7526 13706 7535 13707
rect 7073 13701 7535 13706
rect 6958 13201 6986 13454
rect 6958 13175 6959 13201
rect 6985 13175 6986 13201
rect 6958 13145 6986 13175
rect 6958 13119 6959 13145
rect 6985 13119 6986 13145
rect 6958 13113 6986 13119
rect 7574 13145 7602 13903
rect 7574 13119 7575 13145
rect 7601 13119 7602 13145
rect 7073 12950 7535 12955
rect 7073 12949 7082 12950
rect 7073 12923 7074 12949
rect 7073 12922 7082 12923
rect 7110 12922 7134 12950
rect 7162 12922 7186 12950
rect 7214 12949 7238 12950
rect 7266 12949 7290 12950
rect 7224 12923 7238 12949
rect 7286 12923 7290 12949
rect 7214 12922 7238 12923
rect 7266 12922 7290 12923
rect 7318 12949 7342 12950
rect 7370 12949 7394 12950
rect 7318 12923 7322 12949
rect 7370 12923 7384 12949
rect 7318 12922 7342 12923
rect 7370 12922 7394 12923
rect 7422 12922 7446 12950
rect 7474 12922 7498 12950
rect 7526 12949 7535 12950
rect 7534 12923 7535 12949
rect 7526 12922 7535 12923
rect 7073 12917 7535 12922
rect 7574 12754 7602 13119
rect 7798 13537 7826 14295
rect 7798 13511 7799 13537
rect 7825 13511 7826 13537
rect 7798 12754 7826 13511
rect 7574 12753 7826 12754
rect 7574 12727 7799 12753
rect 7825 12727 7826 12753
rect 7574 12726 7826 12727
rect 7014 12418 7042 12423
rect 6902 12417 7042 12418
rect 6902 12391 7015 12417
rect 7041 12391 7042 12417
rect 6902 12390 7042 12391
rect 7014 12361 7042 12390
rect 7014 12335 7015 12361
rect 7041 12335 7042 12361
rect 7014 11802 7042 12335
rect 7574 12361 7602 12726
rect 7798 12721 7826 12726
rect 8358 13538 8386 13543
rect 8414 13538 8442 14686
rect 8974 14321 9002 15023
rect 8974 14295 8975 14321
rect 9001 14295 9002 14321
rect 8974 14265 9002 14295
rect 8974 14239 8975 14265
rect 9001 14239 9002 14265
rect 8470 13986 8498 13991
rect 8470 13929 8498 13958
rect 8974 13986 9002 14239
rect 8974 13953 9002 13958
rect 9254 15105 9282 15470
rect 9814 15465 9842 15470
rect 10150 15162 10178 15806
rect 10206 15801 10234 15806
rect 10150 15129 10178 15134
rect 10878 15553 10906 16590
rect 10934 16282 10962 16647
rect 10934 16249 10962 16254
rect 11102 15890 11130 17039
rect 11998 17066 12026 17071
rect 12054 17066 12082 17095
rect 11998 17065 12082 17066
rect 11998 17039 11999 17065
rect 12025 17039 12082 17065
rect 11998 17038 12082 17039
rect 12502 17066 12530 17431
rect 12614 17346 12642 17710
rect 12614 17313 12642 17318
rect 13286 17457 13314 17463
rect 13286 17431 13287 17457
rect 13313 17431 13314 17457
rect 13286 17401 13314 17431
rect 13286 17375 13287 17401
rect 13313 17375 13314 17401
rect 12838 17066 12866 17071
rect 12502 17065 12866 17066
rect 12502 17039 12839 17065
rect 12865 17039 12866 17065
rect 12502 17038 12866 17039
rect 11382 16674 11410 16679
rect 11494 16674 11522 16679
rect 11382 16673 11522 16674
rect 11382 16647 11383 16673
rect 11409 16647 11495 16673
rect 11521 16647 11522 16673
rect 11382 16646 11522 16647
rect 11382 16338 11410 16646
rect 11494 16641 11522 16646
rect 11998 16618 12026 17038
rect 12073 16870 12535 16875
rect 12073 16869 12082 16870
rect 12073 16843 12074 16869
rect 12073 16842 12082 16843
rect 12110 16842 12134 16870
rect 12162 16842 12186 16870
rect 12214 16869 12238 16870
rect 12266 16869 12290 16870
rect 12224 16843 12238 16869
rect 12286 16843 12290 16869
rect 12214 16842 12238 16843
rect 12266 16842 12290 16843
rect 12318 16869 12342 16870
rect 12370 16869 12394 16870
rect 12318 16843 12322 16869
rect 12370 16843 12384 16869
rect 12318 16842 12342 16843
rect 12370 16842 12394 16843
rect 12422 16842 12446 16870
rect 12474 16842 12498 16870
rect 12526 16869 12535 16870
rect 12534 16843 12535 16869
rect 12526 16842 12535 16843
rect 12073 16837 12535 16842
rect 12558 16674 12586 16679
rect 12614 16674 12642 17038
rect 12558 16673 12642 16674
rect 12558 16647 12559 16673
rect 12585 16647 12642 16673
rect 12558 16646 12642 16647
rect 12558 16641 12586 16646
rect 11998 16585 12026 16590
rect 12334 16618 12362 16623
rect 11382 16305 11410 16310
rect 12334 16337 12362 16590
rect 12334 16311 12335 16337
rect 12361 16311 12362 16337
rect 11158 16282 11186 16287
rect 11158 16235 11186 16254
rect 12334 16281 12362 16311
rect 12334 16255 12335 16281
rect 12361 16255 12362 16281
rect 12334 16249 12362 16255
rect 12614 16562 12642 16567
rect 12073 16086 12535 16091
rect 12073 16085 12082 16086
rect 12073 16059 12074 16085
rect 12073 16058 12082 16059
rect 12110 16058 12134 16086
rect 12162 16058 12186 16086
rect 12214 16085 12238 16086
rect 12266 16085 12290 16086
rect 12224 16059 12238 16085
rect 12286 16059 12290 16085
rect 12214 16058 12238 16059
rect 12266 16058 12290 16059
rect 12318 16085 12342 16086
rect 12370 16085 12394 16086
rect 12318 16059 12322 16085
rect 12370 16059 12384 16085
rect 12318 16058 12342 16059
rect 12370 16058 12394 16059
rect 12422 16058 12446 16086
rect 12474 16058 12498 16086
rect 12526 16085 12535 16086
rect 12534 16059 12535 16085
rect 12526 16058 12535 16059
rect 12073 16053 12535 16058
rect 12614 15974 12642 16534
rect 12838 16282 12866 17038
rect 13286 17066 13314 17375
rect 14573 17262 15035 17267
rect 14573 17261 14582 17262
rect 14573 17235 14574 17261
rect 14573 17234 14582 17235
rect 14610 17234 14634 17262
rect 14662 17234 14686 17262
rect 14714 17261 14738 17262
rect 14766 17261 14790 17262
rect 14724 17235 14738 17261
rect 14786 17235 14790 17261
rect 14714 17234 14738 17235
rect 14766 17234 14790 17235
rect 14818 17261 14842 17262
rect 14870 17261 14894 17262
rect 14818 17235 14822 17261
rect 14870 17235 14884 17261
rect 14818 17234 14842 17235
rect 14870 17234 14894 17235
rect 14922 17234 14946 17262
rect 14974 17234 14998 17262
rect 15026 17261 15035 17262
rect 15034 17235 15035 17261
rect 15026 17234 15035 17235
rect 14573 17229 15035 17234
rect 13510 17066 13538 17071
rect 13286 17065 13538 17066
rect 13286 17039 13287 17065
rect 13313 17039 13511 17065
rect 13537 17039 13538 17065
rect 13286 17038 13538 17039
rect 12838 16281 13090 16282
rect 12838 16255 12839 16281
rect 12865 16255 13090 16281
rect 12838 16254 13090 16255
rect 12838 16249 12866 16254
rect 12446 15946 12642 15974
rect 12950 16170 12978 16175
rect 11662 15890 11690 15895
rect 11102 15857 11130 15862
rect 11550 15889 11690 15890
rect 11550 15863 11663 15889
rect 11689 15863 11690 15889
rect 11550 15862 11690 15863
rect 10878 15527 10879 15553
rect 10905 15527 10906 15553
rect 10878 15497 10906 15527
rect 10878 15471 10879 15497
rect 10905 15471 10906 15497
rect 9254 15079 9255 15105
rect 9281 15079 9282 15105
rect 9254 14714 9282 15079
rect 10430 15105 10458 15111
rect 10430 15079 10431 15105
rect 10457 15079 10458 15105
rect 10430 15049 10458 15079
rect 10430 15023 10431 15049
rect 10457 15023 10458 15049
rect 9573 14910 10035 14915
rect 9573 14909 9582 14910
rect 9573 14883 9574 14909
rect 9573 14882 9582 14883
rect 9610 14882 9634 14910
rect 9662 14882 9686 14910
rect 9714 14909 9738 14910
rect 9766 14909 9790 14910
rect 9724 14883 9738 14909
rect 9786 14883 9790 14909
rect 9714 14882 9738 14883
rect 9766 14882 9790 14883
rect 9818 14909 9842 14910
rect 9870 14909 9894 14910
rect 9818 14883 9822 14909
rect 9870 14883 9884 14909
rect 9818 14882 9842 14883
rect 9870 14882 9894 14883
rect 9922 14882 9946 14910
rect 9974 14882 9998 14910
rect 10026 14909 10035 14910
rect 10034 14883 10035 14909
rect 10026 14882 10035 14883
rect 9573 14877 10035 14882
rect 9814 14714 9842 14719
rect 9254 14713 9842 14714
rect 9254 14687 9815 14713
rect 9841 14687 9842 14713
rect 9254 14686 9842 14687
rect 9254 14321 9282 14686
rect 9814 14681 9842 14686
rect 9254 14295 9255 14321
rect 9281 14295 9282 14321
rect 8470 13903 8471 13929
rect 8497 13903 8498 13929
rect 8470 13897 8498 13903
rect 9254 13930 9282 14295
rect 10430 14321 10458 15023
rect 10430 14295 10431 14321
rect 10457 14295 10458 14321
rect 10430 14265 10458 14295
rect 10430 14239 10431 14265
rect 10457 14239 10458 14265
rect 9573 14126 10035 14131
rect 9573 14125 9582 14126
rect 9573 14099 9574 14125
rect 9573 14098 9582 14099
rect 9610 14098 9634 14126
rect 9662 14098 9686 14126
rect 9714 14125 9738 14126
rect 9766 14125 9790 14126
rect 9724 14099 9738 14125
rect 9786 14099 9790 14125
rect 9714 14098 9738 14099
rect 9766 14098 9790 14099
rect 9818 14125 9842 14126
rect 9870 14125 9894 14126
rect 9818 14099 9822 14125
rect 9870 14099 9884 14125
rect 9818 14098 9842 14099
rect 9870 14098 9894 14099
rect 9922 14098 9946 14126
rect 9974 14098 9998 14126
rect 10026 14125 10035 14126
rect 10034 14099 10035 14125
rect 10026 14098 10035 14099
rect 9573 14093 10035 14098
rect 9814 13930 9842 13935
rect 9254 13929 9842 13930
rect 9254 13903 9815 13929
rect 9841 13903 9842 13929
rect 9254 13902 9842 13903
rect 8470 13538 8498 13543
rect 8358 13537 8498 13538
rect 8358 13511 8359 13537
rect 8385 13511 8471 13537
rect 8497 13511 8498 13537
rect 8358 13510 8498 13511
rect 8358 13201 8386 13510
rect 8470 13505 8498 13510
rect 9254 13537 9282 13902
rect 9814 13897 9842 13902
rect 9254 13511 9255 13537
rect 9281 13511 9282 13537
rect 8358 13175 8359 13201
rect 8385 13175 8386 13201
rect 8358 13145 8386 13175
rect 8358 13119 8359 13145
rect 8385 13119 8386 13145
rect 8358 12754 8386 13119
rect 9254 13146 9282 13511
rect 10430 13537 10458 14239
rect 10430 13511 10431 13537
rect 10457 13511 10458 13537
rect 10430 13481 10458 13511
rect 10430 13455 10431 13481
rect 10457 13455 10458 13481
rect 9573 13342 10035 13347
rect 9573 13341 9582 13342
rect 9573 13315 9574 13341
rect 9573 13314 9582 13315
rect 9610 13314 9634 13342
rect 9662 13314 9686 13342
rect 9714 13341 9738 13342
rect 9766 13341 9790 13342
rect 9724 13315 9738 13341
rect 9786 13315 9790 13341
rect 9714 13314 9738 13315
rect 9766 13314 9790 13315
rect 9818 13341 9842 13342
rect 9870 13341 9894 13342
rect 9818 13315 9822 13341
rect 9870 13315 9884 13341
rect 9818 13314 9842 13315
rect 9870 13314 9894 13315
rect 9922 13314 9946 13342
rect 9974 13314 9998 13342
rect 10026 13341 10035 13342
rect 10034 13315 10035 13341
rect 10026 13314 10035 13315
rect 9573 13309 10035 13314
rect 9814 13146 9842 13151
rect 9254 13145 9842 13146
rect 9254 13119 9815 13145
rect 9841 13119 9842 13145
rect 9254 13118 9842 13119
rect 8470 12754 8498 12759
rect 8358 12753 8498 12754
rect 8358 12727 8359 12753
rect 8385 12727 8471 12753
rect 8497 12727 8498 12753
rect 8358 12726 8498 12727
rect 7574 12335 7575 12361
rect 7601 12335 7602 12361
rect 7073 12166 7535 12171
rect 7073 12165 7082 12166
rect 7073 12139 7074 12165
rect 7073 12138 7082 12139
rect 7110 12138 7134 12166
rect 7162 12138 7186 12166
rect 7214 12165 7238 12166
rect 7266 12165 7290 12166
rect 7224 12139 7238 12165
rect 7286 12139 7290 12165
rect 7214 12138 7238 12139
rect 7266 12138 7290 12139
rect 7318 12165 7342 12166
rect 7370 12165 7394 12166
rect 7318 12139 7322 12165
rect 7370 12139 7384 12165
rect 7318 12138 7342 12139
rect 7370 12138 7394 12139
rect 7422 12138 7446 12166
rect 7474 12138 7498 12166
rect 7526 12165 7535 12166
rect 7534 12139 7535 12165
rect 7526 12138 7535 12139
rect 7073 12133 7535 12138
rect 7014 11633 7042 11774
rect 7014 11607 7015 11633
rect 7041 11607 7042 11633
rect 7014 11577 7042 11607
rect 7014 11551 7015 11577
rect 7041 11551 7042 11577
rect 7014 10849 7042 11551
rect 7574 11970 7602 12335
rect 8358 12417 8386 12726
rect 8470 12721 8498 12726
rect 9254 12753 9282 13118
rect 9814 13113 9842 13118
rect 9254 12727 9255 12753
rect 9281 12727 9282 12753
rect 8358 12391 8359 12417
rect 8385 12391 8386 12417
rect 8358 12361 8386 12391
rect 8358 12335 8359 12361
rect 8385 12335 8386 12361
rect 7798 11970 7826 11975
rect 7574 11969 7826 11970
rect 7574 11943 7799 11969
rect 7825 11943 7826 11969
rect 7574 11942 7826 11943
rect 7574 11577 7602 11942
rect 7798 11937 7826 11942
rect 8358 11970 8386 12335
rect 9254 12362 9282 12727
rect 10430 12753 10458 13455
rect 10430 12727 10431 12753
rect 10457 12727 10458 12753
rect 10430 12697 10458 12727
rect 10430 12671 10431 12697
rect 10457 12671 10458 12697
rect 9573 12558 10035 12563
rect 9573 12557 9582 12558
rect 9573 12531 9574 12557
rect 9573 12530 9582 12531
rect 9610 12530 9634 12558
rect 9662 12530 9686 12558
rect 9714 12557 9738 12558
rect 9766 12557 9790 12558
rect 9724 12531 9738 12557
rect 9786 12531 9790 12557
rect 9714 12530 9738 12531
rect 9766 12530 9790 12531
rect 9818 12557 9842 12558
rect 9870 12557 9894 12558
rect 9818 12531 9822 12557
rect 9870 12531 9884 12557
rect 9818 12530 9842 12531
rect 9870 12530 9894 12531
rect 9922 12530 9946 12558
rect 9974 12530 9998 12558
rect 10026 12557 10035 12558
rect 10034 12531 10035 12557
rect 10026 12530 10035 12531
rect 9573 12525 10035 12530
rect 9814 12362 9842 12367
rect 9254 12361 9842 12362
rect 9254 12335 9815 12361
rect 9841 12335 9842 12361
rect 9254 12334 9842 12335
rect 8470 11970 8498 11975
rect 8358 11969 8470 11970
rect 8358 11943 8359 11969
rect 8385 11943 8470 11969
rect 8358 11942 8470 11943
rect 7574 11551 7575 11577
rect 7601 11551 7602 11577
rect 7073 11382 7535 11387
rect 7073 11381 7082 11382
rect 7073 11355 7074 11381
rect 7073 11354 7082 11355
rect 7110 11354 7134 11382
rect 7162 11354 7186 11382
rect 7214 11381 7238 11382
rect 7266 11381 7290 11382
rect 7224 11355 7238 11381
rect 7286 11355 7290 11381
rect 7214 11354 7238 11355
rect 7266 11354 7290 11355
rect 7318 11381 7342 11382
rect 7370 11381 7394 11382
rect 7318 11355 7322 11381
rect 7370 11355 7384 11381
rect 7318 11354 7342 11355
rect 7370 11354 7394 11355
rect 7422 11354 7446 11382
rect 7474 11354 7498 11382
rect 7526 11381 7535 11382
rect 7534 11355 7535 11381
rect 7526 11354 7535 11355
rect 7073 11349 7535 11354
rect 7574 11186 7602 11551
rect 8358 11802 8386 11942
rect 8470 11904 8498 11942
rect 9254 11969 9282 12334
rect 9814 12329 9842 12334
rect 10430 12362 10458 12671
rect 10878 14769 10906 15471
rect 10878 14743 10879 14769
rect 10905 14743 10906 14769
rect 10878 14713 10906 14743
rect 10878 14687 10879 14713
rect 10905 14687 10906 14713
rect 10878 14322 10906 14687
rect 10878 13985 10906 14294
rect 10878 13959 10879 13985
rect 10905 13959 10906 13985
rect 10878 13929 10906 13959
rect 10878 13903 10879 13929
rect 10905 13903 10906 13929
rect 10878 13201 10906 13903
rect 11550 15497 11578 15862
rect 11662 15857 11690 15862
rect 11550 15471 11551 15497
rect 11577 15471 11578 15497
rect 11550 14713 11578 15471
rect 12446 15553 12474 15946
rect 12446 15527 12447 15553
rect 12473 15527 12474 15553
rect 12446 15498 12474 15527
rect 12838 15889 12866 15895
rect 12838 15863 12839 15889
rect 12865 15863 12866 15889
rect 12838 15833 12866 15863
rect 12838 15807 12839 15833
rect 12865 15807 12866 15833
rect 12838 15498 12866 15807
rect 12446 15497 12866 15498
rect 12446 15471 12447 15497
rect 12473 15471 12866 15497
rect 12446 15470 12866 15471
rect 12446 15465 12474 15470
rect 12073 15302 12535 15307
rect 12073 15301 12082 15302
rect 12073 15275 12074 15301
rect 12073 15274 12082 15275
rect 12110 15274 12134 15302
rect 12162 15274 12186 15302
rect 12214 15301 12238 15302
rect 12266 15301 12290 15302
rect 12224 15275 12238 15301
rect 12286 15275 12290 15301
rect 12214 15274 12238 15275
rect 12266 15274 12290 15275
rect 12318 15301 12342 15302
rect 12370 15301 12394 15302
rect 12318 15275 12322 15301
rect 12370 15275 12384 15301
rect 12318 15274 12342 15275
rect 12370 15274 12394 15275
rect 12422 15274 12446 15302
rect 12474 15274 12498 15302
rect 12526 15301 12535 15302
rect 12534 15275 12535 15301
rect 12526 15274 12535 15275
rect 12073 15269 12535 15274
rect 11942 15106 11970 15111
rect 11942 15105 12026 15106
rect 11942 15079 11943 15105
rect 11969 15079 12026 15105
rect 11942 15078 12026 15079
rect 11942 15073 11970 15078
rect 11550 14687 11551 14713
rect 11577 14687 11578 14713
rect 11550 13929 11578 14687
rect 11550 13903 11551 13929
rect 11577 13903 11578 13929
rect 11214 13537 11242 13543
rect 11214 13511 11215 13537
rect 11241 13511 11242 13537
rect 11214 13426 11242 13511
rect 11214 13393 11242 13398
rect 11550 13426 11578 13903
rect 10878 13175 10879 13201
rect 10905 13175 10906 13201
rect 10878 13145 10906 13175
rect 10878 13119 10879 13145
rect 10905 13119 10906 13145
rect 10878 12417 10906 13119
rect 10878 12391 10879 12417
rect 10905 12391 10906 12417
rect 10878 12362 10906 12391
rect 10430 12361 10906 12362
rect 10430 12335 10879 12361
rect 10905 12335 10906 12361
rect 10430 12334 10906 12335
rect 9254 11943 9255 11969
rect 9281 11943 9282 11969
rect 8358 11633 8386 11774
rect 8358 11607 8359 11633
rect 8385 11607 8386 11633
rect 8358 11577 8386 11607
rect 8358 11551 8359 11577
rect 8385 11551 8386 11577
rect 7798 11186 7826 11191
rect 7574 11185 7826 11186
rect 7574 11159 7799 11185
rect 7825 11159 7826 11185
rect 7574 11158 7826 11159
rect 7014 10823 7015 10849
rect 7041 10823 7042 10849
rect 7014 10793 7042 10823
rect 7014 10767 7015 10793
rect 7041 10767 7042 10793
rect 6846 10066 6930 10094
rect 6510 9226 6538 9231
rect 6286 9225 6538 9226
rect 6286 9199 6287 9225
rect 6313 9199 6511 9225
rect 6537 9199 6538 9225
rect 6286 9198 6538 9199
rect 6286 9193 6314 9198
rect 6454 8833 6482 9198
rect 6510 9193 6538 9198
rect 6454 8807 6455 8833
rect 6481 8807 6482 8833
rect 6454 8778 6482 8807
rect 6454 8777 6538 8778
rect 6454 8751 6455 8777
rect 6481 8751 6538 8777
rect 6454 8750 6538 8751
rect 6454 8745 6482 8750
rect 6118 8376 6146 8414
rect 6398 8442 6426 8447
rect 6510 8442 6538 8750
rect 6398 8441 6538 8442
rect 6398 8415 6399 8441
rect 6425 8415 6511 8441
rect 6537 8415 6538 8441
rect 6398 8414 6538 8415
rect 6398 8409 6426 8414
rect 6454 8049 6482 8414
rect 6510 8409 6538 8414
rect 6454 8023 6455 8049
rect 6481 8023 6482 8049
rect 6454 7993 6482 8023
rect 6454 7967 6455 7993
rect 6481 7967 6482 7993
rect 6118 7658 6146 7663
rect 6118 7611 6146 7630
rect 6398 7658 6426 7663
rect 6454 7658 6482 7967
rect 6510 7714 6538 7719
rect 6510 7658 6538 7686
rect 6398 7657 6538 7658
rect 6398 7631 6399 7657
rect 6425 7631 6511 7657
rect 6537 7631 6538 7657
rect 6398 7630 6538 7631
rect 6398 7625 6426 7630
rect 6510 7625 6538 7630
rect 5558 7126 6034 7154
rect 5558 6482 5586 7126
rect 5558 5697 5586 6454
rect 5558 5671 5559 5697
rect 5585 5671 5586 5697
rect 5558 5082 5586 5671
rect 5558 4913 5586 5054
rect 5558 4887 5559 4913
rect 5585 4887 5586 4913
rect 5558 4881 5586 4887
rect 6006 6873 6034 7126
rect 6006 6847 6007 6873
rect 6033 6847 6034 6873
rect 6006 6089 6034 6847
rect 6454 7265 6482 7271
rect 6454 7239 6455 7265
rect 6481 7239 6482 7265
rect 6454 7210 6482 7239
rect 6454 6481 6482 7182
rect 6454 6455 6455 6481
rect 6481 6455 6482 6481
rect 6454 6425 6482 6455
rect 6454 6399 6455 6425
rect 6481 6399 6482 6425
rect 6006 6063 6007 6089
rect 6033 6063 6034 6089
rect 6006 5305 6034 6063
rect 6398 6090 6426 6095
rect 6454 6090 6482 6399
rect 6510 6090 6538 6095
rect 6398 6089 6538 6090
rect 6398 6063 6399 6089
rect 6425 6063 6511 6089
rect 6537 6063 6538 6089
rect 6398 6062 6538 6063
rect 6398 6057 6426 6062
rect 6454 5697 6482 6062
rect 6510 6057 6538 6062
rect 6454 5671 6455 5697
rect 6481 5671 6482 5697
rect 6454 5641 6482 5671
rect 6454 5615 6455 5641
rect 6481 5615 6482 5641
rect 6006 5279 6007 5305
rect 6033 5279 6034 5305
rect 5782 4634 5810 4639
rect 5446 2641 5474 2646
rect 5726 3346 5754 3351
rect 4998 2562 5026 2567
rect 5726 2562 5754 3318
rect 4998 2505 5026 2534
rect 4998 2479 4999 2505
rect 5025 2479 5026 2505
rect 4998 2473 5026 2479
rect 5502 2534 5726 2562
rect 5502 2505 5530 2534
rect 5502 2479 5503 2505
rect 5529 2479 5530 2505
rect 5726 2496 5754 2534
rect 5502 2473 5530 2479
rect 4102 2417 4130 2422
rect 4573 2366 5035 2371
rect 4573 2365 4582 2366
rect 4573 2339 4574 2365
rect 4573 2338 4582 2339
rect 4610 2338 4634 2366
rect 4662 2338 4686 2366
rect 4714 2365 4738 2366
rect 4766 2365 4790 2366
rect 4724 2339 4738 2365
rect 4786 2339 4790 2365
rect 4714 2338 4738 2339
rect 4766 2338 4790 2339
rect 4818 2365 4842 2366
rect 4870 2365 4894 2366
rect 4818 2339 4822 2365
rect 4870 2339 4884 2365
rect 4818 2338 4842 2339
rect 4870 2338 4894 2339
rect 4922 2338 4946 2366
rect 4974 2338 4998 2366
rect 5026 2365 5035 2366
rect 5034 2339 5035 2365
rect 5026 2338 5035 2339
rect 4573 2333 5035 2338
rect 4494 2226 4522 2245
rect 3934 1857 3962 1862
rect 4438 2198 4494 2226
rect 4438 2169 4466 2198
rect 4494 2193 4522 2198
rect 4438 2143 4439 2169
rect 4465 2143 4466 2169
rect 3542 1751 3543 1777
rect 3569 1751 3570 1777
rect 3542 1745 3570 1751
rect 4438 1777 4466 2143
rect 5502 2170 5530 2175
rect 4438 1751 4439 1777
rect 4465 1751 4466 1777
rect 4438 1721 4466 1751
rect 4438 1695 4439 1721
rect 4465 1695 4466 1721
rect 4438 1689 4466 1695
rect 4494 2114 4522 2119
rect 4494 1050 4522 2086
rect 5502 1777 5530 2142
rect 5502 1751 5503 1777
rect 5529 1751 5530 1777
rect 5502 1666 5530 1751
rect 5502 1633 5530 1638
rect 4573 1582 5035 1587
rect 4573 1581 4582 1582
rect 4573 1555 4574 1581
rect 4573 1554 4582 1555
rect 4610 1554 4634 1582
rect 4662 1554 4686 1582
rect 4714 1581 4738 1582
rect 4766 1581 4790 1582
rect 4724 1555 4738 1581
rect 4786 1555 4790 1581
rect 4714 1554 4738 1555
rect 4766 1554 4790 1555
rect 4818 1581 4842 1582
rect 4870 1581 4894 1582
rect 4818 1555 4822 1581
rect 4870 1555 4884 1581
rect 4818 1554 4842 1555
rect 4870 1554 4894 1555
rect 4922 1554 4946 1582
rect 4974 1554 4998 1582
rect 5026 1581 5035 1582
rect 5034 1555 5035 1581
rect 5026 1554 5035 1555
rect 4573 1549 5035 1554
rect 4494 1022 4578 1050
rect 4550 400 4578 1022
rect 5782 400 5810 4606
rect 6006 4522 6034 5279
rect 6398 5306 6426 5311
rect 6454 5306 6482 5615
rect 6510 5306 6538 5311
rect 6398 5305 6510 5306
rect 6398 5279 6399 5305
rect 6425 5279 6510 5305
rect 6398 5278 6510 5279
rect 6398 5273 6426 5278
rect 6510 5240 6538 5278
rect 6006 4242 6034 4494
rect 6398 4913 6426 4919
rect 6398 4887 6399 4913
rect 6425 4887 6426 4913
rect 6398 4857 6426 4887
rect 6398 4831 6399 4857
rect 6425 4831 6426 4857
rect 6398 4214 6426 4831
rect 6006 4186 6090 4214
rect 6398 4186 6482 4214
rect 6062 3737 6090 4186
rect 6454 4129 6482 4158
rect 6454 4103 6455 4129
rect 6481 4103 6482 4129
rect 6454 4073 6482 4103
rect 6454 4047 6455 4073
rect 6481 4047 6482 4073
rect 6454 4041 6482 4047
rect 6062 3711 6063 3737
rect 6089 3711 6090 3737
rect 6062 3705 6090 3711
rect 6006 3346 6034 3351
rect 6006 3299 6034 3318
rect 6454 3346 6482 3351
rect 6454 3345 6538 3346
rect 6454 3319 6455 3345
rect 6481 3319 6538 3345
rect 6454 3318 6538 3319
rect 6454 3313 6482 3318
rect 6342 2954 6370 2959
rect 6454 2954 6482 2959
rect 6342 2953 6482 2954
rect 6342 2927 6343 2953
rect 6369 2927 6455 2953
rect 6481 2927 6482 2953
rect 6342 2926 6482 2927
rect 5838 2562 5866 2567
rect 5838 2225 5866 2534
rect 5838 2199 5839 2225
rect 5865 2199 5866 2225
rect 5838 2169 5866 2199
rect 5838 2143 5839 2169
rect 5865 2143 5866 2169
rect 5838 2137 5866 2143
rect 6342 2226 6370 2926
rect 6454 2921 6482 2926
rect 6454 2562 6482 2567
rect 6510 2562 6538 3318
rect 6482 2534 6538 2562
rect 6454 2515 6482 2534
rect 6342 1778 6370 2198
rect 6398 1778 6426 1783
rect 6342 1777 6426 1778
rect 6342 1751 6399 1777
rect 6425 1751 6426 1777
rect 6342 1750 6426 1751
rect 6398 1722 6426 1750
rect 6398 1675 6426 1694
rect 6902 490 6930 10066
rect 7014 10065 7042 10767
rect 7294 10962 7322 10967
rect 7294 10793 7322 10934
rect 7294 10767 7295 10793
rect 7321 10767 7322 10793
rect 7294 10761 7322 10767
rect 7574 10962 7602 11158
rect 7798 11153 7826 11158
rect 8358 11186 8386 11551
rect 8470 11186 8498 11191
rect 8358 11185 8498 11186
rect 8358 11159 8359 11185
rect 8385 11159 8471 11185
rect 8497 11159 8498 11185
rect 8358 11158 8498 11159
rect 8358 11153 8386 11158
rect 7073 10598 7535 10603
rect 7073 10597 7082 10598
rect 7073 10571 7074 10597
rect 7073 10570 7082 10571
rect 7110 10570 7134 10598
rect 7162 10570 7186 10598
rect 7214 10597 7238 10598
rect 7266 10597 7290 10598
rect 7224 10571 7238 10597
rect 7286 10571 7290 10597
rect 7214 10570 7238 10571
rect 7266 10570 7290 10571
rect 7318 10597 7342 10598
rect 7370 10597 7394 10598
rect 7318 10571 7322 10597
rect 7370 10571 7384 10597
rect 7318 10570 7342 10571
rect 7370 10570 7394 10571
rect 7422 10570 7446 10598
rect 7474 10570 7498 10598
rect 7526 10597 7535 10598
rect 7534 10571 7535 10597
rect 7526 10570 7535 10571
rect 7073 10565 7535 10570
rect 7014 10039 7015 10065
rect 7041 10039 7042 10065
rect 7014 10010 7042 10039
rect 6958 9982 7014 10010
rect 6958 7210 6986 9982
rect 7014 9963 7042 9982
rect 7574 10402 7602 10934
rect 8470 10849 8498 11158
rect 8470 10823 8471 10849
rect 8497 10823 8498 10849
rect 8470 10793 8498 10823
rect 8470 10767 8471 10793
rect 8497 10767 8498 10793
rect 7798 10402 7826 10407
rect 7574 10401 7826 10402
rect 7574 10375 7799 10401
rect 7825 10375 7826 10401
rect 7574 10374 7826 10375
rect 7574 10009 7602 10374
rect 7574 9983 7575 10009
rect 7601 9983 7602 10009
rect 7574 9977 7602 9983
rect 7073 9814 7535 9819
rect 7073 9813 7082 9814
rect 7073 9787 7074 9813
rect 7073 9786 7082 9787
rect 7110 9786 7134 9814
rect 7162 9786 7186 9814
rect 7214 9813 7238 9814
rect 7266 9813 7290 9814
rect 7224 9787 7238 9813
rect 7286 9787 7290 9813
rect 7214 9786 7238 9787
rect 7266 9786 7290 9787
rect 7318 9813 7342 9814
rect 7370 9813 7394 9814
rect 7318 9787 7322 9813
rect 7370 9787 7384 9813
rect 7318 9786 7342 9787
rect 7370 9786 7394 9787
rect 7422 9786 7446 9814
rect 7474 9786 7498 9814
rect 7526 9813 7535 9814
rect 7534 9787 7535 9813
rect 7526 9786 7535 9787
rect 7073 9781 7535 9786
rect 7798 9617 7826 10374
rect 8470 10094 8498 10767
rect 9254 11185 9282 11943
rect 10430 11970 10458 12334
rect 10878 12329 10906 12334
rect 11550 13145 11578 13398
rect 11550 13119 11551 13145
rect 11577 13119 11578 13145
rect 11550 12361 11578 13119
rect 11550 12335 11551 12361
rect 11577 12335 11578 12361
rect 10430 11913 10458 11942
rect 10430 11887 10431 11913
rect 10457 11887 10458 11913
rect 10430 11881 10458 11887
rect 9573 11774 10035 11779
rect 9573 11773 9582 11774
rect 9573 11747 9574 11773
rect 9573 11746 9582 11747
rect 9610 11746 9634 11774
rect 9662 11746 9686 11774
rect 9714 11773 9738 11774
rect 9766 11773 9790 11774
rect 9724 11747 9738 11773
rect 9786 11747 9790 11773
rect 9714 11746 9738 11747
rect 9766 11746 9790 11747
rect 9818 11773 9842 11774
rect 9870 11773 9894 11774
rect 9818 11747 9822 11773
rect 9870 11747 9884 11773
rect 9818 11746 9842 11747
rect 9870 11746 9894 11747
rect 9922 11746 9946 11774
rect 9974 11746 9998 11774
rect 10026 11773 10035 11774
rect 10034 11747 10035 11773
rect 10026 11746 10035 11747
rect 9573 11741 10035 11746
rect 10766 11633 10794 11639
rect 10766 11607 10767 11633
rect 10793 11607 10794 11633
rect 9254 11159 9255 11185
rect 9281 11159 9282 11185
rect 9254 10962 9282 11159
rect 10038 11577 10066 11583
rect 10038 11551 10039 11577
rect 10065 11551 10066 11577
rect 10038 11074 10066 11551
rect 10766 11577 10794 11607
rect 10766 11551 10767 11577
rect 10793 11551 10794 11577
rect 10430 11186 10458 11191
rect 10766 11186 10794 11551
rect 10430 11185 10794 11186
rect 10430 11159 10431 11185
rect 10457 11159 10794 11185
rect 10430 11158 10794 11159
rect 10430 11129 10458 11158
rect 10430 11103 10431 11129
rect 10457 11103 10458 11129
rect 10038 11046 10122 11074
rect 9573 10990 10035 10995
rect 9573 10989 9582 10990
rect 9573 10963 9574 10989
rect 9573 10962 9582 10963
rect 9610 10962 9634 10990
rect 9662 10962 9686 10990
rect 9714 10989 9738 10990
rect 9766 10989 9790 10990
rect 9724 10963 9738 10989
rect 9786 10963 9790 10989
rect 9714 10962 9738 10963
rect 9766 10962 9790 10963
rect 9818 10989 9842 10990
rect 9870 10989 9894 10990
rect 9818 10963 9822 10989
rect 9870 10963 9884 10989
rect 9818 10962 9842 10963
rect 9870 10962 9894 10963
rect 9922 10962 9946 10990
rect 9974 10962 9998 10990
rect 10026 10989 10035 10990
rect 10034 10963 10035 10989
rect 10026 10962 10035 10963
rect 9573 10957 10035 10962
rect 8750 10401 8778 10407
rect 8750 10375 8751 10401
rect 8777 10375 8778 10401
rect 8750 10345 8778 10375
rect 8750 10319 8751 10345
rect 8777 10319 8778 10345
rect 8750 10094 8778 10319
rect 9254 10401 9282 10934
rect 10094 10906 10122 11046
rect 9254 10375 9255 10401
rect 9281 10375 9282 10401
rect 8470 10066 8778 10094
rect 8806 10122 8834 10127
rect 8470 10065 8498 10066
rect 8470 10039 8471 10065
rect 8497 10039 8498 10065
rect 8470 10010 8498 10039
rect 7798 9591 7799 9617
rect 7825 9591 7826 9617
rect 7798 9585 7826 9591
rect 8414 10009 8498 10010
rect 8414 9983 8471 10009
rect 8497 9983 8498 10009
rect 8414 9982 8498 9983
rect 8414 9281 8442 9982
rect 8470 9977 8498 9982
rect 8750 10010 8778 10015
rect 8414 9255 8415 9281
rect 8441 9255 8442 9281
rect 7574 9225 7602 9231
rect 7574 9199 7575 9225
rect 7601 9199 7602 9225
rect 7073 9030 7535 9035
rect 7073 9029 7082 9030
rect 7073 9003 7074 9029
rect 7073 9002 7082 9003
rect 7110 9002 7134 9030
rect 7162 9002 7186 9030
rect 7214 9029 7238 9030
rect 7266 9029 7290 9030
rect 7224 9003 7238 9029
rect 7286 9003 7290 9029
rect 7214 9002 7238 9003
rect 7266 9002 7290 9003
rect 7318 9029 7342 9030
rect 7370 9029 7394 9030
rect 7318 9003 7322 9029
rect 7370 9003 7384 9029
rect 7318 9002 7342 9003
rect 7370 9002 7394 9003
rect 7422 9002 7446 9030
rect 7474 9002 7498 9030
rect 7526 9029 7535 9030
rect 7534 9003 7535 9029
rect 7526 9002 7535 9003
rect 7073 8997 7535 9002
rect 7014 8442 7042 8447
rect 7014 7658 7042 8414
rect 7574 8441 7602 9199
rect 8414 9225 8442 9255
rect 8414 9199 8415 9225
rect 8441 9199 8442 9225
rect 7574 8415 7575 8441
rect 7601 8415 7602 8441
rect 7073 8246 7535 8251
rect 7073 8245 7082 8246
rect 7073 8219 7074 8245
rect 7073 8218 7082 8219
rect 7110 8218 7134 8246
rect 7162 8218 7186 8246
rect 7214 8245 7238 8246
rect 7266 8245 7290 8246
rect 7224 8219 7238 8245
rect 7286 8219 7290 8245
rect 7214 8218 7238 8219
rect 7266 8218 7290 8219
rect 7318 8245 7342 8246
rect 7370 8245 7394 8246
rect 7318 8219 7322 8245
rect 7370 8219 7384 8245
rect 7318 8218 7342 8219
rect 7370 8218 7394 8219
rect 7422 8218 7446 8246
rect 7474 8218 7498 8246
rect 7526 8245 7535 8246
rect 7534 8219 7535 8245
rect 7526 8218 7535 8219
rect 7073 8213 7535 8218
rect 7574 8050 7602 8415
rect 7798 8833 7826 8839
rect 7798 8807 7799 8833
rect 7825 8807 7826 8833
rect 7798 8050 7826 8807
rect 8414 8497 8442 9199
rect 8414 8471 8415 8497
rect 8441 8471 8442 8497
rect 8414 8441 8442 8471
rect 8414 8415 8415 8441
rect 8441 8415 8442 8441
rect 8414 8409 8442 8415
rect 8750 9617 8778 9982
rect 8750 9591 8751 9617
rect 8777 9591 8778 9617
rect 8750 9561 8778 9591
rect 8750 9535 8751 9561
rect 8777 9535 8778 9561
rect 8750 8833 8778 9535
rect 8750 8807 8751 8833
rect 8777 8807 8778 8833
rect 8750 8777 8778 8807
rect 8750 8751 8751 8777
rect 8777 8751 8778 8777
rect 7574 8049 7826 8050
rect 7574 8023 7799 8049
rect 7825 8023 7826 8049
rect 7574 8022 7826 8023
rect 7294 7658 7322 7663
rect 7014 7657 7322 7658
rect 7014 7631 7295 7657
rect 7321 7631 7322 7657
rect 7014 7630 7322 7631
rect 7294 7546 7322 7630
rect 7294 7513 7322 7518
rect 7574 7658 7602 8022
rect 7798 8017 7826 8022
rect 8750 8050 8778 8751
rect 8750 7993 8778 8022
rect 8750 7967 8751 7993
rect 8777 7967 8778 7993
rect 8750 7961 8778 7967
rect 7073 7462 7535 7467
rect 7073 7461 7082 7462
rect 7073 7435 7074 7461
rect 7073 7434 7082 7435
rect 7110 7434 7134 7462
rect 7162 7434 7186 7462
rect 7214 7461 7238 7462
rect 7266 7461 7290 7462
rect 7224 7435 7238 7461
rect 7286 7435 7290 7461
rect 7214 7434 7238 7435
rect 7266 7434 7290 7435
rect 7318 7461 7342 7462
rect 7370 7461 7394 7462
rect 7318 7435 7322 7461
rect 7370 7435 7384 7461
rect 7318 7434 7342 7435
rect 7370 7434 7394 7435
rect 7422 7434 7446 7462
rect 7474 7434 7498 7462
rect 7526 7461 7535 7462
rect 7534 7435 7535 7461
rect 7526 7434 7535 7435
rect 7073 7429 7535 7434
rect 7574 7378 7602 7630
rect 7742 7714 7770 7719
rect 7742 7658 7770 7686
rect 7966 7658 7994 7663
rect 7742 7657 8274 7658
rect 7742 7631 7743 7657
rect 7769 7631 7967 7657
rect 7993 7631 8274 7657
rect 7742 7630 8274 7631
rect 7742 7625 7770 7630
rect 7966 7625 7994 7630
rect 6958 6929 6986 7182
rect 6958 6903 6959 6929
rect 6985 6903 6986 6929
rect 6958 6873 6986 6903
rect 6958 6847 6959 6873
rect 6985 6847 6986 6873
rect 6958 6841 6986 6847
rect 7518 7350 7602 7378
rect 7798 7546 7826 7551
rect 7518 6873 7546 7350
rect 7798 7265 7826 7518
rect 7798 7239 7799 7265
rect 7825 7239 7826 7265
rect 7798 7233 7826 7239
rect 8246 7266 8274 7630
rect 8470 7490 8498 7495
rect 8470 7266 8498 7462
rect 8246 7265 8498 7266
rect 8246 7239 8247 7265
rect 8273 7239 8471 7265
rect 8497 7239 8498 7265
rect 8246 7238 8498 7239
rect 7518 6847 7519 6873
rect 7545 6847 7546 6873
rect 7518 6762 7546 6847
rect 8246 6929 8274 7238
rect 8470 7233 8498 7238
rect 8246 6903 8247 6929
rect 8273 6903 8274 6929
rect 8246 6873 8274 6903
rect 8246 6847 8247 6873
rect 8273 6847 8274 6873
rect 7518 6734 7602 6762
rect 7073 6678 7535 6683
rect 7073 6677 7082 6678
rect 7073 6651 7074 6677
rect 7073 6650 7082 6651
rect 7110 6650 7134 6678
rect 7162 6650 7186 6678
rect 7214 6677 7238 6678
rect 7266 6677 7290 6678
rect 7224 6651 7238 6677
rect 7286 6651 7290 6677
rect 7214 6650 7238 6651
rect 7266 6650 7290 6651
rect 7318 6677 7342 6678
rect 7370 6677 7394 6678
rect 7318 6651 7322 6677
rect 7370 6651 7384 6677
rect 7318 6650 7342 6651
rect 7370 6650 7394 6651
rect 7422 6650 7446 6678
rect 7474 6650 7498 6678
rect 7526 6677 7535 6678
rect 7534 6651 7535 6677
rect 7526 6650 7535 6651
rect 7073 6645 7535 6650
rect 7574 6090 7602 6734
rect 7574 6043 7602 6062
rect 8078 6481 8106 6487
rect 8078 6455 8079 6481
rect 8105 6455 8106 6481
rect 8078 6090 8106 6455
rect 7073 5894 7535 5899
rect 7073 5893 7082 5894
rect 7073 5867 7074 5893
rect 7073 5866 7082 5867
rect 7110 5866 7134 5894
rect 7162 5866 7186 5894
rect 7214 5893 7238 5894
rect 7266 5893 7290 5894
rect 7224 5867 7238 5893
rect 7286 5867 7290 5893
rect 7214 5866 7238 5867
rect 7266 5866 7290 5867
rect 7318 5893 7342 5894
rect 7370 5893 7394 5894
rect 7318 5867 7322 5893
rect 7370 5867 7384 5893
rect 7318 5866 7342 5867
rect 7370 5866 7394 5867
rect 7422 5866 7446 5894
rect 7474 5866 7498 5894
rect 7526 5893 7535 5894
rect 7534 5867 7535 5893
rect 7526 5866 7535 5867
rect 7073 5861 7535 5866
rect 8078 5866 8106 6062
rect 8246 6482 8274 6847
rect 8470 6482 8498 6487
rect 8246 6481 8498 6482
rect 8246 6455 8247 6481
rect 8273 6455 8471 6481
rect 8497 6455 8498 6481
rect 8246 6454 8498 6455
rect 8246 6145 8274 6454
rect 8470 6449 8498 6454
rect 8246 6119 8247 6145
rect 8273 6119 8274 6145
rect 8246 6089 8274 6119
rect 8246 6063 8247 6089
rect 8273 6063 8274 6089
rect 8246 6057 8274 6063
rect 8078 5697 8106 5838
rect 8078 5671 8079 5697
rect 8105 5671 8106 5697
rect 8078 5665 8106 5671
rect 7518 5305 7546 5311
rect 7518 5279 7519 5305
rect 7545 5279 7546 5305
rect 7518 5194 7546 5279
rect 7742 5306 7770 5311
rect 7742 5259 7770 5278
rect 7966 5306 7994 5311
rect 7966 5259 7994 5278
rect 8246 5306 8274 5311
rect 7518 5166 7602 5194
rect 7073 5110 7535 5115
rect 7073 5109 7082 5110
rect 7073 5083 7074 5109
rect 7073 5082 7082 5083
rect 7110 5082 7134 5110
rect 7162 5082 7186 5110
rect 7214 5109 7238 5110
rect 7266 5109 7290 5110
rect 7224 5083 7238 5109
rect 7286 5083 7290 5109
rect 7214 5082 7238 5083
rect 7266 5082 7290 5083
rect 7318 5109 7342 5110
rect 7370 5109 7394 5110
rect 7318 5083 7322 5109
rect 7370 5083 7384 5109
rect 7318 5082 7342 5083
rect 7370 5082 7394 5083
rect 7422 5082 7446 5110
rect 7474 5082 7498 5110
rect 7526 5109 7535 5110
rect 7534 5083 7535 5109
rect 7526 5082 7535 5083
rect 7073 5077 7535 5082
rect 7574 4914 7602 5166
rect 7798 4914 7826 4919
rect 7574 4913 7826 4914
rect 7574 4887 7799 4913
rect 7825 4887 7826 4913
rect 7574 4886 7826 4887
rect 6958 4577 6986 4583
rect 6958 4551 6959 4577
rect 6985 4551 6986 4577
rect 6958 4521 6986 4551
rect 6958 4495 6959 4521
rect 6985 4495 6986 4521
rect 6958 4214 6986 4495
rect 7294 4522 7322 4527
rect 7294 4475 7322 4494
rect 7574 4522 7602 4886
rect 7798 4881 7826 4886
rect 8246 4914 8274 5278
rect 8470 4914 8498 4919
rect 8246 4913 8498 4914
rect 8246 4887 8247 4913
rect 8273 4887 8471 4913
rect 8497 4887 8498 4913
rect 8246 4886 8498 4887
rect 7073 4326 7535 4331
rect 7073 4325 7082 4326
rect 7073 4299 7074 4325
rect 7073 4298 7082 4299
rect 7110 4298 7134 4326
rect 7162 4298 7186 4326
rect 7214 4325 7238 4326
rect 7266 4325 7290 4326
rect 7224 4299 7238 4325
rect 7286 4299 7290 4325
rect 7214 4298 7238 4299
rect 7266 4298 7290 4299
rect 7318 4325 7342 4326
rect 7370 4325 7394 4326
rect 7318 4299 7322 4325
rect 7370 4299 7384 4325
rect 7318 4298 7342 4299
rect 7370 4298 7394 4299
rect 7422 4298 7446 4326
rect 7474 4298 7498 4326
rect 7526 4325 7535 4326
rect 7534 4299 7535 4325
rect 7526 4298 7535 4299
rect 7073 4293 7535 4298
rect 6958 4186 7042 4214
rect 7014 3793 7042 4158
rect 7014 3767 7015 3793
rect 7041 3767 7042 3793
rect 7014 3737 7042 3767
rect 7014 3711 7015 3737
rect 7041 3711 7042 3737
rect 7014 3705 7042 3711
rect 7073 3542 7535 3547
rect 7073 3541 7082 3542
rect 7073 3515 7074 3541
rect 7073 3514 7082 3515
rect 7110 3514 7134 3542
rect 7162 3514 7186 3542
rect 7214 3541 7238 3542
rect 7266 3541 7290 3542
rect 7224 3515 7238 3541
rect 7286 3515 7290 3541
rect 7214 3514 7238 3515
rect 7266 3514 7290 3515
rect 7318 3541 7342 3542
rect 7370 3541 7394 3542
rect 7318 3515 7322 3541
rect 7370 3515 7384 3541
rect 7318 3514 7342 3515
rect 7370 3514 7394 3515
rect 7422 3514 7446 3542
rect 7474 3514 7498 3542
rect 7526 3541 7535 3542
rect 7534 3515 7535 3541
rect 7526 3514 7535 3515
rect 7073 3509 7535 3514
rect 7014 2953 7042 2959
rect 7014 2927 7015 2953
rect 7041 2927 7042 2953
rect 7014 2562 7042 2927
rect 7574 2953 7602 4494
rect 8246 4577 8274 4886
rect 8470 4881 8498 4886
rect 8246 4551 8247 4577
rect 8273 4551 8274 4577
rect 8246 4521 8274 4551
rect 8246 4495 8247 4521
rect 8273 4495 8274 4521
rect 8246 4489 8274 4495
rect 7798 4129 7826 4135
rect 7798 4103 7799 4129
rect 7825 4103 7826 4129
rect 7798 4073 7826 4103
rect 7798 4047 7799 4073
rect 7825 4047 7826 4073
rect 7798 3738 7826 4047
rect 8806 3794 8834 10094
rect 9254 9617 9282 10375
rect 10038 10878 10122 10906
rect 10038 10793 10066 10878
rect 10038 10767 10039 10793
rect 10065 10767 10066 10793
rect 10038 10290 10066 10767
rect 10430 10401 10458 11103
rect 10766 10849 10794 11158
rect 10766 10823 10767 10849
rect 10793 10823 10794 10849
rect 10766 10793 10794 10823
rect 10766 10767 10767 10793
rect 10793 10767 10794 10793
rect 10766 10761 10794 10767
rect 11550 11577 11578 12335
rect 11550 11551 11551 11577
rect 11577 11551 11578 11577
rect 11550 10794 11578 11551
rect 11998 14321 12026 15078
rect 12838 15105 12866 15470
rect 12838 15079 12839 15105
rect 12865 15079 12866 15105
rect 12838 15049 12866 15079
rect 12838 15023 12839 15049
rect 12865 15023 12866 15049
rect 12446 14769 12474 14775
rect 12446 14743 12447 14769
rect 12473 14743 12474 14769
rect 12446 14714 12474 14743
rect 12446 14667 12474 14686
rect 12838 14714 12866 15023
rect 12073 14518 12535 14523
rect 12073 14517 12082 14518
rect 12073 14491 12074 14517
rect 12073 14490 12082 14491
rect 12110 14490 12134 14518
rect 12162 14490 12186 14518
rect 12214 14517 12238 14518
rect 12266 14517 12290 14518
rect 12224 14491 12238 14517
rect 12286 14491 12290 14517
rect 12214 14490 12238 14491
rect 12266 14490 12290 14491
rect 12318 14517 12342 14518
rect 12370 14517 12394 14518
rect 12318 14491 12322 14517
rect 12370 14491 12384 14517
rect 12318 14490 12342 14491
rect 12370 14490 12394 14491
rect 12422 14490 12446 14518
rect 12474 14490 12498 14518
rect 12526 14517 12535 14518
rect 12534 14491 12535 14517
rect 12526 14490 12535 14491
rect 12073 14485 12535 14490
rect 11998 14295 11999 14321
rect 12025 14295 12026 14321
rect 11998 12753 12026 14295
rect 12446 14322 12474 14327
rect 12838 14322 12866 14686
rect 12894 14322 12922 14327
rect 12838 14294 12894 14322
rect 12446 13985 12474 14294
rect 12894 14265 12922 14294
rect 12894 14239 12895 14265
rect 12921 14239 12922 14265
rect 12894 14233 12922 14239
rect 12446 13959 12447 13985
rect 12473 13959 12474 13985
rect 12446 13930 12474 13959
rect 12446 13929 12642 13930
rect 12446 13903 12447 13929
rect 12473 13903 12642 13929
rect 12446 13902 12642 13903
rect 12446 13897 12474 13902
rect 12073 13734 12535 13739
rect 12073 13733 12082 13734
rect 12073 13707 12074 13733
rect 12073 13706 12082 13707
rect 12110 13706 12134 13734
rect 12162 13706 12186 13734
rect 12214 13733 12238 13734
rect 12266 13733 12290 13734
rect 12224 13707 12238 13733
rect 12286 13707 12290 13733
rect 12214 13706 12238 13707
rect 12266 13706 12290 13707
rect 12318 13733 12342 13734
rect 12370 13733 12394 13734
rect 12318 13707 12322 13733
rect 12370 13707 12384 13733
rect 12318 13706 12342 13707
rect 12370 13706 12394 13707
rect 12422 13706 12446 13734
rect 12474 13706 12498 13734
rect 12526 13733 12535 13734
rect 12534 13707 12535 13733
rect 12526 13706 12535 13707
rect 12073 13701 12535 13706
rect 12614 13650 12642 13902
rect 12446 13622 12642 13650
rect 12110 13538 12138 13543
rect 12446 13538 12474 13622
rect 12110 13537 12474 13538
rect 12110 13511 12111 13537
rect 12137 13511 12474 13537
rect 12110 13510 12474 13511
rect 12110 13481 12138 13510
rect 12110 13455 12111 13481
rect 12137 13455 12138 13481
rect 12110 13449 12138 13455
rect 12446 13201 12474 13510
rect 12670 13537 12698 13543
rect 12670 13511 12671 13537
rect 12697 13511 12698 13537
rect 12670 13426 12698 13511
rect 12670 13393 12698 13398
rect 12446 13175 12447 13201
rect 12473 13175 12474 13201
rect 12446 13145 12474 13175
rect 12446 13119 12447 13145
rect 12473 13119 12474 13145
rect 12446 13113 12474 13119
rect 12950 13146 12978 16142
rect 13062 15974 13090 16254
rect 13286 16170 13314 17038
rect 13510 17033 13538 17038
rect 13454 16673 13482 16679
rect 13454 16647 13455 16673
rect 13481 16647 13482 16673
rect 13454 16618 13482 16647
rect 13454 16571 13482 16590
rect 13790 16618 13818 16623
rect 13790 16337 13818 16590
rect 14573 16478 15035 16483
rect 14573 16477 14582 16478
rect 14573 16451 14574 16477
rect 14573 16450 14582 16451
rect 14610 16450 14634 16478
rect 14662 16450 14686 16478
rect 14714 16477 14738 16478
rect 14766 16477 14790 16478
rect 14724 16451 14738 16477
rect 14786 16451 14790 16477
rect 14714 16450 14738 16451
rect 14766 16450 14790 16451
rect 14818 16477 14842 16478
rect 14870 16477 14894 16478
rect 14818 16451 14822 16477
rect 14870 16451 14884 16477
rect 14818 16450 14842 16451
rect 14870 16450 14894 16451
rect 14922 16450 14946 16478
rect 14974 16450 14998 16478
rect 15026 16477 15035 16478
rect 15034 16451 15035 16477
rect 15026 16450 15035 16451
rect 14573 16445 15035 16450
rect 13790 16311 13791 16337
rect 13817 16311 13818 16337
rect 13790 16281 13818 16311
rect 15470 16337 15498 16343
rect 15470 16311 15471 16337
rect 15497 16311 15498 16337
rect 13790 16255 13791 16281
rect 13817 16255 13818 16281
rect 13790 16249 13818 16255
rect 14294 16281 14322 16287
rect 14294 16255 14295 16281
rect 14321 16255 14322 16281
rect 13286 16137 13314 16142
rect 13062 15946 13146 15974
rect 13062 15106 13090 15946
rect 13118 15889 13146 15946
rect 13118 15863 13119 15889
rect 13145 15863 13146 15889
rect 13118 15857 13146 15863
rect 14014 15889 14042 15895
rect 14014 15863 14015 15889
rect 14041 15863 14042 15889
rect 14014 15834 14042 15863
rect 14070 15834 14098 15839
rect 14014 15833 14098 15834
rect 14014 15807 14071 15833
rect 14097 15807 14098 15833
rect 14014 15806 14098 15807
rect 14014 15553 14042 15806
rect 14070 15801 14098 15806
rect 14014 15527 14015 15553
rect 14041 15527 14042 15553
rect 13062 14770 13090 15078
rect 13062 14737 13090 14742
rect 13118 15497 13146 15503
rect 13118 15471 13119 15497
rect 13145 15471 13146 15497
rect 13118 15105 13146 15471
rect 13118 15079 13119 15105
rect 13145 15079 13146 15105
rect 13118 14713 13146 15079
rect 13118 14687 13119 14713
rect 13145 14687 13146 14713
rect 13118 14322 13146 14687
rect 14014 15497 14042 15527
rect 14014 15471 14015 15497
rect 14041 15471 14042 15497
rect 14014 15105 14042 15471
rect 14014 15079 14015 15105
rect 14041 15079 14042 15105
rect 14014 15050 14042 15079
rect 14294 15497 14322 16255
rect 15470 16281 15498 16311
rect 15470 16255 15471 16281
rect 15497 16255 15498 16281
rect 15470 15974 15498 16255
rect 15414 15946 15498 15974
rect 16814 15946 16842 15951
rect 15302 15918 15414 15946
rect 15078 15890 15106 15895
rect 15078 15843 15106 15862
rect 14573 15694 15035 15699
rect 14573 15693 14582 15694
rect 14573 15667 14574 15693
rect 14573 15666 14582 15667
rect 14610 15666 14634 15694
rect 14662 15666 14686 15694
rect 14714 15693 14738 15694
rect 14766 15693 14790 15694
rect 14724 15667 14738 15693
rect 14786 15667 14790 15693
rect 14714 15666 14738 15667
rect 14766 15666 14790 15667
rect 14818 15693 14842 15694
rect 14870 15693 14894 15694
rect 14818 15667 14822 15693
rect 14870 15667 14884 15693
rect 14818 15666 14842 15667
rect 14870 15666 14894 15667
rect 14922 15666 14946 15694
rect 14974 15666 14998 15694
rect 15026 15693 15035 15694
rect 15034 15667 15035 15693
rect 15026 15666 15035 15667
rect 14573 15661 15035 15666
rect 14294 15471 14295 15497
rect 14321 15471 14322 15497
rect 14294 15106 14322 15471
rect 14294 15073 14322 15078
rect 14798 15106 14826 15111
rect 14798 15059 14826 15078
rect 14070 15050 14098 15055
rect 14014 15049 14098 15050
rect 14014 15023 14071 15049
rect 14097 15023 14098 15049
rect 14014 15022 14098 15023
rect 14014 14769 14042 15022
rect 14070 15017 14098 15022
rect 14573 14910 15035 14915
rect 14573 14909 14582 14910
rect 14573 14883 14574 14909
rect 14573 14882 14582 14883
rect 14610 14882 14634 14910
rect 14662 14882 14686 14910
rect 14714 14909 14738 14910
rect 14766 14909 14790 14910
rect 14724 14883 14738 14909
rect 14786 14883 14790 14909
rect 14714 14882 14738 14883
rect 14766 14882 14790 14883
rect 14818 14909 14842 14910
rect 14870 14909 14894 14910
rect 14818 14883 14822 14909
rect 14870 14883 14884 14909
rect 14818 14882 14842 14883
rect 14870 14882 14894 14883
rect 14922 14882 14946 14910
rect 14974 14882 14998 14910
rect 15026 14909 15035 14910
rect 15034 14883 15035 14909
rect 15026 14882 15035 14883
rect 14573 14877 15035 14882
rect 14014 14743 14015 14769
rect 14041 14743 14042 14769
rect 14014 14713 14042 14743
rect 15302 14769 15330 15918
rect 15414 15913 15442 15918
rect 15526 15889 15554 15895
rect 15526 15863 15527 15889
rect 15553 15863 15554 15889
rect 15526 15834 15554 15863
rect 16478 15889 16506 15895
rect 16478 15863 16479 15889
rect 16505 15863 16506 15889
rect 15750 15834 15778 15839
rect 15526 15833 15778 15834
rect 15526 15807 15751 15833
rect 15777 15807 15778 15833
rect 15526 15806 15778 15807
rect 15358 15553 15386 15559
rect 15358 15527 15359 15553
rect 15385 15527 15386 15553
rect 15358 15497 15386 15527
rect 15358 15471 15359 15497
rect 15385 15471 15386 15497
rect 15358 15106 15386 15471
rect 15526 15106 15554 15806
rect 15750 15801 15778 15806
rect 15358 15105 15554 15106
rect 15358 15079 15359 15105
rect 15385 15079 15527 15105
rect 15553 15079 15554 15105
rect 15358 15078 15554 15079
rect 15358 15073 15386 15078
rect 15302 14743 15303 14769
rect 15329 14743 15330 14769
rect 14014 14687 14015 14713
rect 14041 14687 14042 14713
rect 13230 14322 13258 14327
rect 13118 14321 13258 14322
rect 13118 14295 13231 14321
rect 13257 14295 13258 14321
rect 13118 14294 13258 14295
rect 12073 12950 12535 12955
rect 12073 12949 12082 12950
rect 12073 12923 12074 12949
rect 12073 12922 12082 12923
rect 12110 12922 12134 12950
rect 12162 12922 12186 12950
rect 12214 12949 12238 12950
rect 12266 12949 12290 12950
rect 12224 12923 12238 12949
rect 12286 12923 12290 12949
rect 12214 12922 12238 12923
rect 12266 12922 12290 12923
rect 12318 12949 12342 12950
rect 12370 12949 12394 12950
rect 12318 12923 12322 12949
rect 12370 12923 12384 12949
rect 12318 12922 12342 12923
rect 12370 12922 12394 12923
rect 12422 12922 12446 12950
rect 12474 12922 12498 12950
rect 12526 12949 12535 12950
rect 12534 12923 12535 12949
rect 12526 12922 12535 12923
rect 12073 12917 12535 12922
rect 11998 12727 11999 12753
rect 12025 12727 12026 12753
rect 11998 11969 12026 12727
rect 12894 12753 12922 12759
rect 12894 12727 12895 12753
rect 12921 12727 12922 12753
rect 12894 12698 12922 12727
rect 12950 12698 12978 13118
rect 13118 13930 13146 13935
rect 13230 13930 13258 14294
rect 13118 13929 13258 13930
rect 13118 13903 13119 13929
rect 13145 13903 13258 13929
rect 13118 13902 13258 13903
rect 14014 14322 14042 14687
rect 14014 13985 14042 14294
rect 14350 14713 14378 14719
rect 14350 14687 14351 14713
rect 14377 14687 14378 14713
rect 14350 14322 14378 14687
rect 15302 14713 15330 14743
rect 15302 14687 15303 14713
rect 15329 14687 15330 14713
rect 14798 14322 14826 14327
rect 14350 14321 14826 14322
rect 14350 14295 14799 14321
rect 14825 14295 14826 14321
rect 14350 14294 14826 14295
rect 14014 13959 14015 13985
rect 14041 13959 14042 13985
rect 14014 13930 14042 13959
rect 14182 14265 14210 14271
rect 14182 14239 14183 14265
rect 14209 14239 14210 14265
rect 14182 13930 14210 14239
rect 14014 13929 14266 13930
rect 14014 13903 14015 13929
rect 14041 13903 14266 13929
rect 14014 13902 14266 13903
rect 13118 13426 13146 13902
rect 14014 13897 14042 13902
rect 13118 13145 13146 13398
rect 13118 13119 13119 13145
rect 13145 13119 13146 13145
rect 13118 12754 13146 13119
rect 13398 13537 13426 13543
rect 13398 13511 13399 13537
rect 13425 13511 13426 13537
rect 13398 13481 13426 13511
rect 13398 13455 13399 13481
rect 13425 13455 13426 13481
rect 13398 13146 13426 13455
rect 13398 13113 13426 13118
rect 14014 13201 14042 13207
rect 14014 13175 14015 13201
rect 14041 13175 14042 13201
rect 14014 13146 14042 13175
rect 14014 13099 14042 13118
rect 13342 12754 13370 12759
rect 13118 12753 13370 12754
rect 13118 12727 13343 12753
rect 13369 12727 13370 12753
rect 13118 12726 13370 12727
rect 12894 12697 12978 12698
rect 12894 12671 12895 12697
rect 12921 12671 12978 12697
rect 12894 12670 12978 12671
rect 12894 12665 12922 12670
rect 12446 12417 12474 12423
rect 12446 12391 12447 12417
rect 12473 12391 12474 12417
rect 12446 12362 12474 12391
rect 12446 12361 12642 12362
rect 12446 12335 12447 12361
rect 12473 12335 12642 12361
rect 12446 12334 12642 12335
rect 12446 12329 12474 12334
rect 12073 12166 12535 12171
rect 12073 12165 12082 12166
rect 12073 12139 12074 12165
rect 12073 12138 12082 12139
rect 12110 12138 12134 12166
rect 12162 12138 12186 12166
rect 12214 12165 12238 12166
rect 12266 12165 12290 12166
rect 12224 12139 12238 12165
rect 12286 12139 12290 12165
rect 12214 12138 12238 12139
rect 12266 12138 12290 12139
rect 12318 12165 12342 12166
rect 12370 12165 12394 12166
rect 12318 12139 12322 12165
rect 12370 12139 12384 12165
rect 12318 12138 12342 12139
rect 12370 12138 12394 12139
rect 12422 12138 12446 12166
rect 12474 12138 12498 12166
rect 12526 12165 12535 12166
rect 12534 12139 12535 12165
rect 12526 12138 12535 12139
rect 12073 12133 12535 12138
rect 11998 11943 11999 11969
rect 12025 11943 12026 11969
rect 11998 11802 12026 11943
rect 11998 11186 12026 11774
rect 12446 11633 12474 11639
rect 12446 11607 12447 11633
rect 12473 11607 12474 11633
rect 12446 11578 12474 11607
rect 12614 11578 12642 12334
rect 12950 11969 12978 12670
rect 12950 11943 12951 11969
rect 12977 11943 12978 11969
rect 12950 11913 12978 11943
rect 12950 11887 12951 11913
rect 12977 11887 12978 11913
rect 12950 11578 12978 11887
rect 12446 11577 12978 11578
rect 12446 11551 12447 11577
rect 12473 11551 12978 11577
rect 12446 11550 12978 11551
rect 12446 11545 12474 11550
rect 12073 11382 12535 11387
rect 12073 11381 12082 11382
rect 12073 11355 12074 11381
rect 12073 11354 12082 11355
rect 12110 11354 12134 11382
rect 12162 11354 12186 11382
rect 12214 11381 12238 11382
rect 12266 11381 12290 11382
rect 12224 11355 12238 11381
rect 12286 11355 12290 11381
rect 12214 11354 12238 11355
rect 12266 11354 12290 11355
rect 12318 11381 12342 11382
rect 12370 11381 12394 11382
rect 12318 11355 12322 11381
rect 12370 11355 12384 11381
rect 12318 11354 12342 11355
rect 12370 11354 12394 11355
rect 12422 11354 12446 11382
rect 12474 11354 12498 11382
rect 12526 11381 12535 11382
rect 12534 11355 12535 11381
rect 12526 11354 12535 11355
rect 12073 11349 12535 11354
rect 11942 11185 12026 11186
rect 11942 11159 11999 11185
rect 12025 11159 12026 11185
rect 11942 11158 12026 11159
rect 11550 10793 11634 10794
rect 11550 10767 11551 10793
rect 11577 10767 11634 10793
rect 11550 10766 11634 10767
rect 11550 10761 11578 10766
rect 10430 10375 10431 10401
rect 10457 10375 10458 10401
rect 10430 10345 10458 10375
rect 10430 10319 10431 10345
rect 10457 10319 10458 10345
rect 10038 10262 10122 10290
rect 9573 10206 10035 10211
rect 9573 10205 9582 10206
rect 9573 10179 9574 10205
rect 9573 10178 9582 10179
rect 9610 10178 9634 10206
rect 9662 10178 9686 10206
rect 9714 10205 9738 10206
rect 9766 10205 9790 10206
rect 9724 10179 9738 10205
rect 9786 10179 9790 10205
rect 9714 10178 9738 10179
rect 9766 10178 9790 10179
rect 9818 10205 9842 10206
rect 9870 10205 9894 10206
rect 9818 10179 9822 10205
rect 9870 10179 9884 10205
rect 9818 10178 9842 10179
rect 9870 10178 9894 10179
rect 9922 10178 9946 10206
rect 9974 10178 9998 10206
rect 10026 10205 10035 10206
rect 10034 10179 10035 10205
rect 10026 10178 10035 10179
rect 9573 10173 10035 10178
rect 10094 10122 10122 10262
rect 9254 9591 9255 9617
rect 9281 9591 9282 9617
rect 9254 8833 9282 9591
rect 10038 10094 10122 10122
rect 10038 10009 10066 10094
rect 10038 9983 10039 10009
rect 10065 9983 10066 10009
rect 10038 9506 10066 9983
rect 10374 10010 10402 10015
rect 10430 10010 10458 10319
rect 11606 10402 11634 10766
rect 11942 10402 11970 11158
rect 11998 11153 12026 11158
rect 12950 11185 12978 11550
rect 12950 11159 12951 11185
rect 12977 11159 12978 11185
rect 12950 11129 12978 11159
rect 12950 11103 12951 11129
rect 12977 11103 12978 11129
rect 12222 10849 12250 10855
rect 12222 10823 12223 10849
rect 12249 10823 12250 10849
rect 12222 10794 12250 10823
rect 11606 10401 11970 10402
rect 11606 10375 11943 10401
rect 11969 10375 11970 10401
rect 11606 10374 11970 10375
rect 10542 10010 10570 10015
rect 10374 10009 10570 10010
rect 10374 9983 10375 10009
rect 10401 9983 10543 10009
rect 10569 9983 10570 10009
rect 10374 9982 10570 9983
rect 10374 9977 10402 9982
rect 10430 9617 10458 9623
rect 10430 9591 10431 9617
rect 10457 9591 10458 9617
rect 10430 9562 10458 9591
rect 10318 9561 10458 9562
rect 10318 9535 10431 9561
rect 10457 9535 10458 9561
rect 10318 9534 10458 9535
rect 10038 9478 10122 9506
rect 9573 9422 10035 9427
rect 9573 9421 9582 9422
rect 9573 9395 9574 9421
rect 9573 9394 9582 9395
rect 9610 9394 9634 9422
rect 9662 9394 9686 9422
rect 9714 9421 9738 9422
rect 9766 9421 9790 9422
rect 9724 9395 9738 9421
rect 9786 9395 9790 9421
rect 9714 9394 9738 9395
rect 9766 9394 9790 9395
rect 9818 9421 9842 9422
rect 9870 9421 9894 9422
rect 9818 9395 9822 9421
rect 9870 9395 9884 9421
rect 9818 9394 9842 9395
rect 9870 9394 9894 9395
rect 9922 9394 9946 9422
rect 9974 9394 9998 9422
rect 10026 9421 10035 9422
rect 10034 9395 10035 9421
rect 10026 9394 10035 9395
rect 9573 9389 10035 9394
rect 10094 9338 10122 9478
rect 9254 8807 9255 8833
rect 9281 8807 9282 8833
rect 9254 8442 9282 8807
rect 10038 9310 10122 9338
rect 10038 9225 10066 9310
rect 10038 9199 10039 9225
rect 10065 9199 10066 9225
rect 10038 8722 10066 9199
rect 10318 9226 10346 9534
rect 10430 9529 10458 9534
rect 10542 9282 10570 9982
rect 11550 10010 11578 10015
rect 11606 10010 11634 10374
rect 11942 10369 11970 10374
rect 11998 10793 12250 10794
rect 11998 10767 12223 10793
rect 12249 10767 12250 10793
rect 11998 10766 12250 10767
rect 11998 10094 12026 10766
rect 12222 10761 12250 10766
rect 12073 10598 12535 10603
rect 12073 10597 12082 10598
rect 12073 10571 12074 10597
rect 12073 10570 12082 10571
rect 12110 10570 12134 10598
rect 12162 10570 12186 10598
rect 12214 10597 12238 10598
rect 12266 10597 12290 10598
rect 12224 10571 12238 10597
rect 12286 10571 12290 10597
rect 12214 10570 12238 10571
rect 12266 10570 12290 10571
rect 12318 10597 12342 10598
rect 12370 10597 12394 10598
rect 12318 10571 12322 10597
rect 12370 10571 12384 10597
rect 12318 10570 12342 10571
rect 12370 10570 12394 10571
rect 12422 10570 12446 10598
rect 12474 10570 12498 10598
rect 12526 10597 12535 10598
rect 12534 10571 12535 10597
rect 12526 10570 12535 10571
rect 12073 10565 12535 10570
rect 12670 10401 12698 10407
rect 12670 10375 12671 10401
rect 12697 10375 12698 10401
rect 12670 10346 12698 10375
rect 11942 10066 12026 10094
rect 11550 10009 11634 10010
rect 11550 9983 11551 10009
rect 11577 9983 11634 10009
rect 11550 9982 11634 9983
rect 11550 9977 11578 9982
rect 10318 8833 10346 9198
rect 10486 9226 10514 9231
rect 10486 9179 10514 9198
rect 10318 8807 10319 8833
rect 10345 8807 10346 8833
rect 10318 8777 10346 8807
rect 10318 8751 10319 8777
rect 10345 8751 10346 8777
rect 10038 8694 10122 8722
rect 9573 8638 10035 8643
rect 9573 8637 9582 8638
rect 9573 8611 9574 8637
rect 9573 8610 9582 8611
rect 9610 8610 9634 8638
rect 9662 8610 9686 8638
rect 9714 8637 9738 8638
rect 9766 8637 9790 8638
rect 9724 8611 9738 8637
rect 9786 8611 9790 8637
rect 9714 8610 9738 8611
rect 9766 8610 9790 8611
rect 9818 8637 9842 8638
rect 9870 8637 9894 8638
rect 9818 8611 9822 8637
rect 9870 8611 9884 8637
rect 9818 8610 9842 8611
rect 9870 8610 9894 8611
rect 9922 8610 9946 8638
rect 9974 8610 9998 8638
rect 10026 8637 10035 8638
rect 10034 8611 10035 8637
rect 10026 8610 10035 8611
rect 9573 8605 10035 8610
rect 10094 8554 10122 8694
rect 10038 8526 10122 8554
rect 10318 8554 10346 8751
rect 10318 8526 10514 8554
rect 9814 8442 9842 8447
rect 9254 8414 9814 8442
rect 9254 8049 9282 8414
rect 9254 8023 9255 8049
rect 9281 8023 9282 8049
rect 9254 7546 9282 8023
rect 9814 7938 9842 8414
rect 10038 8442 10066 8526
rect 10038 8409 10066 8414
rect 10318 8441 10346 8526
rect 10318 8415 10319 8441
rect 10345 8415 10346 8441
rect 10150 8050 10178 8055
rect 9814 7910 10122 7938
rect 9573 7854 10035 7859
rect 9573 7853 9582 7854
rect 9573 7827 9574 7853
rect 9573 7826 9582 7827
rect 9610 7826 9634 7854
rect 9662 7826 9686 7854
rect 9714 7853 9738 7854
rect 9766 7853 9790 7854
rect 9724 7827 9738 7853
rect 9786 7827 9790 7853
rect 9714 7826 9738 7827
rect 9766 7826 9790 7827
rect 9818 7853 9842 7854
rect 9870 7853 9894 7854
rect 9818 7827 9822 7853
rect 9870 7827 9884 7853
rect 9818 7826 9842 7827
rect 9870 7826 9894 7827
rect 9922 7826 9946 7854
rect 9974 7826 9998 7854
rect 10026 7853 10035 7854
rect 10034 7827 10035 7853
rect 10026 7826 10035 7827
rect 9573 7821 10035 7826
rect 10094 7770 10122 7910
rect 10038 7742 10122 7770
rect 10038 7657 10066 7742
rect 10038 7631 10039 7657
rect 10065 7631 10066 7657
rect 10038 7625 10066 7631
rect 9254 7513 9282 7518
rect 9478 7265 9506 7271
rect 9478 7239 9479 7265
rect 9505 7239 9506 7265
rect 9478 6874 9506 7239
rect 10150 7265 10178 8022
rect 10318 8050 10346 8415
rect 10486 8441 10514 8526
rect 10486 8415 10487 8441
rect 10513 8415 10514 8441
rect 10486 8409 10514 8415
rect 10542 8330 10570 9254
rect 11606 9617 11634 9982
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 10318 8017 10346 8022
rect 10430 8302 10570 8330
rect 11438 9225 11466 9231
rect 11438 9199 11439 9225
rect 11465 9199 11466 9225
rect 11438 8834 11466 9199
rect 11606 8834 11634 9591
rect 11774 10010 11802 10015
rect 11942 10010 11970 10066
rect 11774 10009 11970 10010
rect 11774 9983 11775 10009
rect 11801 9983 11943 10009
rect 11969 9983 11970 10009
rect 11774 9982 11970 9983
rect 11774 9282 11802 9982
rect 11942 9977 11970 9982
rect 11998 9618 12026 10038
rect 12502 10345 12698 10346
rect 12502 10319 12671 10345
rect 12697 10319 12698 10345
rect 12502 10318 12698 10319
rect 12502 10066 12530 10318
rect 12670 10313 12698 10318
rect 12502 10033 12530 10038
rect 12950 10066 12978 11103
rect 12950 10033 12978 10038
rect 13342 12361 13370 12726
rect 14238 12753 14266 13902
rect 14238 12727 14239 12753
rect 14265 12727 14266 12753
rect 14238 12697 14266 12727
rect 14238 12671 14239 12697
rect 14265 12671 14266 12697
rect 14238 12418 14266 12671
rect 14238 12385 14266 12390
rect 13342 12335 13343 12361
rect 13369 12335 13370 12361
rect 13342 11969 13370 12335
rect 13342 11943 13343 11969
rect 13369 11943 13370 11969
rect 13342 11802 13370 11943
rect 13342 11578 13370 11774
rect 13454 11578 13482 11583
rect 13342 11577 13482 11578
rect 13342 11551 13455 11577
rect 13481 11551 13482 11577
rect 13342 11550 13482 11551
rect 13342 11185 13370 11550
rect 13454 11545 13482 11550
rect 13342 11159 13343 11185
rect 13369 11159 13370 11185
rect 13342 10794 13370 11159
rect 14294 11074 14322 11079
rect 13454 10794 13482 10799
rect 13342 10793 13482 10794
rect 13342 10767 13455 10793
rect 13481 10767 13482 10793
rect 13342 10766 13482 10767
rect 13342 10401 13370 10766
rect 13454 10761 13482 10766
rect 13342 10375 13343 10401
rect 13369 10375 13370 10401
rect 13342 10010 13370 10375
rect 14294 10401 14322 11046
rect 14294 10375 14295 10401
rect 14321 10375 14322 10401
rect 14294 10345 14322 10375
rect 14294 10319 14295 10345
rect 14321 10319 14322 10345
rect 14294 10313 14322 10319
rect 14350 10094 14378 14294
rect 14798 14289 14826 14294
rect 15302 14322 15330 14687
rect 15470 14322 15498 14327
rect 15302 14321 15498 14322
rect 15302 14295 15303 14321
rect 15329 14295 15471 14321
rect 15497 14295 15498 14321
rect 15302 14294 15498 14295
rect 14573 14126 15035 14131
rect 14573 14125 14582 14126
rect 14573 14099 14574 14125
rect 14573 14098 14582 14099
rect 14610 14098 14634 14126
rect 14662 14098 14686 14126
rect 14714 14125 14738 14126
rect 14766 14125 14790 14126
rect 14724 14099 14738 14125
rect 14786 14099 14790 14125
rect 14714 14098 14738 14099
rect 14766 14098 14790 14099
rect 14818 14125 14842 14126
rect 14870 14125 14894 14126
rect 14818 14099 14822 14125
rect 14870 14099 14884 14125
rect 14818 14098 14842 14099
rect 14870 14098 14894 14099
rect 14922 14098 14946 14126
rect 14974 14098 14998 14126
rect 15026 14125 15035 14126
rect 15034 14099 15035 14125
rect 15026 14098 15035 14099
rect 14573 14093 15035 14098
rect 14574 13929 14602 13935
rect 14574 13903 14575 13929
rect 14601 13903 14602 13929
rect 14574 13538 14602 13903
rect 14798 13538 14826 13543
rect 14462 13537 14826 13538
rect 14462 13511 14799 13537
rect 14825 13511 14826 13537
rect 14462 13510 14826 13511
rect 14462 13145 14490 13510
rect 14798 13505 14826 13510
rect 14573 13342 15035 13347
rect 14573 13341 14582 13342
rect 14573 13315 14574 13341
rect 14573 13314 14582 13315
rect 14610 13314 14634 13342
rect 14662 13314 14686 13342
rect 14714 13341 14738 13342
rect 14766 13341 14790 13342
rect 14724 13315 14738 13341
rect 14786 13315 14790 13341
rect 14714 13314 14738 13315
rect 14766 13314 14790 13315
rect 14818 13341 14842 13342
rect 14870 13341 14894 13342
rect 14818 13315 14822 13341
rect 14870 13315 14884 13341
rect 14818 13314 14842 13315
rect 14870 13314 14894 13315
rect 14922 13314 14946 13342
rect 14974 13314 14998 13342
rect 15026 13341 15035 13342
rect 15034 13315 15035 13341
rect 15026 13314 15035 13315
rect 14573 13309 15035 13314
rect 14462 13119 14463 13145
rect 14489 13119 14490 13145
rect 14462 12754 14490 13119
rect 15302 13201 15330 14294
rect 15470 14289 15498 14294
rect 15470 13986 15498 13991
rect 15526 13986 15554 15078
rect 16478 15105 16506 15863
rect 16814 15889 16842 15918
rect 16814 15863 16815 15889
rect 16841 15863 16842 15889
rect 16814 15857 16842 15863
rect 16478 15079 16479 15105
rect 16505 15079 16506 15105
rect 16478 15050 16506 15079
rect 16478 14714 16506 15022
rect 16478 14681 16506 14686
rect 16534 15106 16562 15111
rect 15470 13985 15554 13986
rect 15470 13959 15471 13985
rect 15497 13959 15554 13985
rect 15470 13958 15554 13959
rect 16534 14321 16562 15078
rect 16534 14295 16535 14321
rect 16561 14295 16562 14321
rect 15470 13929 15498 13958
rect 15470 13903 15471 13929
rect 15497 13903 15498 13929
rect 15470 13482 15498 13903
rect 16366 13930 16394 13935
rect 15470 13449 15498 13454
rect 15862 13537 15890 13543
rect 15862 13511 15863 13537
rect 15889 13511 15890 13537
rect 15862 13482 15890 13511
rect 15302 13175 15303 13201
rect 15329 13175 15330 13201
rect 15302 13146 15330 13175
rect 14798 12754 14826 12759
rect 14462 12753 14826 12754
rect 14462 12727 14799 12753
rect 14825 12727 14826 12753
rect 14462 12726 14826 12727
rect 14406 12418 14434 12423
rect 14406 12361 14434 12390
rect 14406 12335 14407 12361
rect 14433 12335 14434 12361
rect 14406 11969 14434 12335
rect 14462 12362 14490 12726
rect 14798 12721 14826 12726
rect 15302 12754 15330 13118
rect 15470 12754 15498 12759
rect 15302 12753 15498 12754
rect 15302 12727 15303 12753
rect 15329 12727 15471 12753
rect 15497 12727 15498 12753
rect 15302 12726 15498 12727
rect 14573 12558 15035 12563
rect 14573 12557 14582 12558
rect 14573 12531 14574 12557
rect 14573 12530 14582 12531
rect 14610 12530 14634 12558
rect 14662 12530 14686 12558
rect 14714 12557 14738 12558
rect 14766 12557 14790 12558
rect 14724 12531 14738 12557
rect 14786 12531 14790 12557
rect 14714 12530 14738 12531
rect 14766 12530 14790 12531
rect 14818 12557 14842 12558
rect 14870 12557 14894 12558
rect 14818 12531 14822 12557
rect 14870 12531 14884 12557
rect 14818 12530 14842 12531
rect 14870 12530 14894 12531
rect 14922 12530 14946 12558
rect 14974 12530 14998 12558
rect 15026 12557 15035 12558
rect 15034 12531 15035 12557
rect 15026 12530 15035 12531
rect 14573 12525 15035 12530
rect 14742 12362 14770 12367
rect 14462 12361 14770 12362
rect 14462 12335 14743 12361
rect 14769 12335 14770 12361
rect 14462 12334 14770 12335
rect 14406 11943 14407 11969
rect 14433 11943 14434 11969
rect 14406 11913 14434 11943
rect 14742 11970 14770 12334
rect 15302 12362 15330 12726
rect 15470 12721 15498 12726
rect 15414 12362 15442 12367
rect 15302 12361 15442 12362
rect 15302 12335 15303 12361
rect 15329 12335 15415 12361
rect 15441 12335 15442 12361
rect 15302 12334 15442 12335
rect 14798 11970 14826 11975
rect 14742 11969 15106 11970
rect 14742 11943 14799 11969
rect 14825 11943 15106 11969
rect 14742 11942 15106 11943
rect 14798 11937 14826 11942
rect 14406 11887 14407 11913
rect 14433 11887 14434 11913
rect 14406 11634 14434 11887
rect 14573 11774 15035 11779
rect 14573 11773 14582 11774
rect 14573 11747 14574 11773
rect 14573 11746 14582 11747
rect 14610 11746 14634 11774
rect 14662 11746 14686 11774
rect 14714 11773 14738 11774
rect 14766 11773 14790 11774
rect 14724 11747 14738 11773
rect 14786 11747 14790 11773
rect 14714 11746 14738 11747
rect 14766 11746 14790 11747
rect 14818 11773 14842 11774
rect 14870 11773 14894 11774
rect 14818 11747 14822 11773
rect 14870 11747 14884 11773
rect 14818 11746 14842 11747
rect 14870 11746 14894 11747
rect 14922 11746 14946 11774
rect 14974 11746 14998 11774
rect 15026 11773 15035 11774
rect 15034 11747 15035 11773
rect 15026 11746 15035 11747
rect 14573 11741 15035 11746
rect 15078 11746 15106 11942
rect 14462 11634 14490 11639
rect 14406 11633 14490 11634
rect 14406 11607 14463 11633
rect 14489 11607 14490 11633
rect 14406 11606 14490 11607
rect 14462 11577 14490 11606
rect 14462 11551 14463 11577
rect 14489 11551 14490 11577
rect 14406 11186 14434 11191
rect 14462 11186 14490 11551
rect 14406 11185 14490 11186
rect 14406 11159 14407 11185
rect 14433 11159 14490 11185
rect 14406 11158 14490 11159
rect 14406 11129 14434 11158
rect 14406 11103 14407 11129
rect 14433 11103 14434 11129
rect 14406 11097 14434 11103
rect 14462 11074 14490 11158
rect 14462 10849 14490 11046
rect 15078 11577 15106 11718
rect 15078 11551 15079 11577
rect 15105 11551 15106 11577
rect 15078 11185 15106 11551
rect 15078 11159 15079 11185
rect 15105 11159 15106 11185
rect 14573 10990 15035 10995
rect 14573 10989 14582 10990
rect 14573 10963 14574 10989
rect 14573 10962 14582 10963
rect 14610 10962 14634 10990
rect 14662 10962 14686 10990
rect 14714 10989 14738 10990
rect 14766 10989 14790 10990
rect 14724 10963 14738 10989
rect 14786 10963 14790 10989
rect 14714 10962 14738 10963
rect 14766 10962 14790 10963
rect 14818 10989 14842 10990
rect 14870 10989 14894 10990
rect 14818 10963 14822 10989
rect 14870 10963 14884 10989
rect 14818 10962 14842 10963
rect 14870 10962 14894 10963
rect 14922 10962 14946 10990
rect 14974 10962 14998 10990
rect 15026 10989 15035 10990
rect 15034 10963 15035 10989
rect 15026 10962 15035 10963
rect 14573 10957 15035 10962
rect 14462 10823 14463 10849
rect 14489 10823 14490 10849
rect 14462 10793 14490 10823
rect 14462 10767 14463 10793
rect 14489 10767 14490 10793
rect 14462 10761 14490 10767
rect 15078 10793 15106 11159
rect 15302 11186 15330 12334
rect 15414 12329 15442 12334
rect 15862 11969 15890 13454
rect 15862 11943 15863 11969
rect 15889 11943 15890 11969
rect 15862 11913 15890 11943
rect 15862 11887 15863 11913
rect 15889 11887 15890 11913
rect 15862 11633 15890 11887
rect 15862 11607 15863 11633
rect 15889 11607 15890 11633
rect 15862 11577 15890 11607
rect 15862 11551 15863 11577
rect 15889 11551 15890 11577
rect 15470 11186 15498 11191
rect 15302 11185 15498 11186
rect 15302 11159 15303 11185
rect 15329 11159 15471 11185
rect 15497 11159 15498 11185
rect 15302 11158 15498 11159
rect 15302 11153 15330 11158
rect 15078 10767 15079 10793
rect 15105 10767 15106 10793
rect 15078 10401 15106 10767
rect 15078 10375 15079 10401
rect 15105 10375 15106 10401
rect 14573 10206 15035 10211
rect 14573 10205 14582 10206
rect 14573 10179 14574 10205
rect 14573 10178 14582 10179
rect 14610 10178 14634 10206
rect 14662 10178 14686 10206
rect 14714 10205 14738 10206
rect 14766 10205 14790 10206
rect 14724 10179 14738 10205
rect 14786 10179 14790 10205
rect 14714 10178 14738 10179
rect 14766 10178 14790 10179
rect 14818 10205 14842 10206
rect 14870 10205 14894 10206
rect 14818 10179 14822 10205
rect 14870 10179 14884 10205
rect 14818 10178 14842 10179
rect 14870 10178 14894 10179
rect 14922 10178 14946 10206
rect 14974 10178 14998 10206
rect 15026 10205 15035 10206
rect 15034 10179 15035 10205
rect 15026 10178 15035 10179
rect 14573 10173 15035 10178
rect 14350 10066 14434 10094
rect 12073 9814 12535 9819
rect 12073 9813 12082 9814
rect 12073 9787 12074 9813
rect 12073 9786 12082 9787
rect 12110 9786 12134 9814
rect 12162 9786 12186 9814
rect 12214 9813 12238 9814
rect 12266 9813 12290 9814
rect 12224 9787 12238 9813
rect 12286 9787 12290 9813
rect 12214 9786 12238 9787
rect 12266 9786 12290 9787
rect 12318 9813 12342 9814
rect 12370 9813 12394 9814
rect 12318 9787 12322 9813
rect 12370 9787 12384 9813
rect 12318 9786 12342 9787
rect 12370 9786 12394 9787
rect 12422 9786 12446 9814
rect 12474 9786 12498 9814
rect 12526 9813 12535 9814
rect 12534 9787 12535 9813
rect 12526 9786 12535 9787
rect 12073 9781 12535 9786
rect 12054 9618 12082 9623
rect 12278 9618 12306 9623
rect 11998 9617 12306 9618
rect 11998 9591 12055 9617
rect 12081 9591 12279 9617
rect 12305 9591 12306 9617
rect 11998 9590 12306 9591
rect 12054 9585 12082 9590
rect 12278 9585 12306 9590
rect 13342 9617 13370 9982
rect 13622 10010 13650 10015
rect 14070 10010 14098 10015
rect 14294 10010 14322 10015
rect 13622 9963 13650 9982
rect 14014 10009 14322 10010
rect 14014 9983 14071 10009
rect 14097 9983 14295 10009
rect 14321 9983 14322 10009
rect 14014 9982 14322 9983
rect 13342 9591 13343 9617
rect 13369 9591 13370 9617
rect 11774 9225 11802 9254
rect 11774 9199 11775 9225
rect 11801 9199 11802 9225
rect 11774 9193 11802 9199
rect 11942 9282 11970 9287
rect 11942 9225 11970 9254
rect 13342 9282 13370 9591
rect 13342 9226 13370 9254
rect 14014 9617 14042 9982
rect 14070 9977 14098 9982
rect 14294 9977 14322 9982
rect 14014 9591 14015 9617
rect 14041 9591 14042 9617
rect 14014 9561 14042 9591
rect 14014 9535 14015 9561
rect 14041 9535 14042 9561
rect 14014 9338 14042 9535
rect 11942 9199 11943 9225
rect 11969 9199 11970 9225
rect 11942 9193 11970 9199
rect 13062 9225 13370 9226
rect 13062 9199 13343 9225
rect 13369 9199 13370 9225
rect 13062 9198 13370 9199
rect 12073 9030 12535 9035
rect 12073 9029 12082 9030
rect 12073 9003 12074 9029
rect 12073 9002 12082 9003
rect 12110 9002 12134 9030
rect 12162 9002 12186 9030
rect 12214 9029 12238 9030
rect 12266 9029 12290 9030
rect 12224 9003 12238 9029
rect 12286 9003 12290 9029
rect 12214 9002 12238 9003
rect 12266 9002 12290 9003
rect 12318 9029 12342 9030
rect 12370 9029 12394 9030
rect 12318 9003 12322 9029
rect 12370 9003 12384 9029
rect 12318 9002 12342 9003
rect 12370 9002 12394 9003
rect 12422 9002 12446 9030
rect 12474 9002 12498 9030
rect 12526 9029 12535 9030
rect 12534 9003 12535 9029
rect 12526 9002 12535 9003
rect 12073 8997 12535 9002
rect 12054 8834 12082 8839
rect 12278 8834 12306 8839
rect 13062 8834 13090 9198
rect 13342 9193 13370 9198
rect 13790 9226 13818 9231
rect 14014 9226 14042 9310
rect 13790 9225 14042 9226
rect 13790 9199 13791 9225
rect 13817 9199 14015 9225
rect 14041 9199 14042 9225
rect 13790 9198 14042 9199
rect 11438 8833 11634 8834
rect 11438 8807 11607 8833
rect 11633 8807 11634 8833
rect 11438 8806 11634 8807
rect 11438 8442 11466 8806
rect 11606 8801 11634 8806
rect 11998 8833 12306 8834
rect 11998 8807 12055 8833
rect 12081 8807 12279 8833
rect 12305 8807 12306 8833
rect 11998 8806 12306 8807
rect 10430 8049 10458 8302
rect 10430 8023 10431 8049
rect 10457 8023 10458 8049
rect 10430 7993 10458 8023
rect 11438 8049 11466 8414
rect 11438 8023 11439 8049
rect 11465 8023 11466 8049
rect 10430 7967 10431 7993
rect 10457 7967 10458 7993
rect 10206 7658 10234 7663
rect 10430 7658 10458 7967
rect 10206 7657 10458 7658
rect 10206 7631 10207 7657
rect 10233 7631 10431 7657
rect 10457 7631 10458 7657
rect 10206 7630 10458 7631
rect 10206 7602 10234 7630
rect 10430 7625 10458 7630
rect 10542 7994 10570 7999
rect 10206 7569 10234 7574
rect 10150 7239 10151 7265
rect 10177 7239 10178 7265
rect 10150 7210 10178 7239
rect 10206 7210 10234 7215
rect 10150 7209 10234 7210
rect 10150 7183 10207 7209
rect 10233 7183 10234 7209
rect 10150 7182 10234 7183
rect 9573 7070 10035 7075
rect 9573 7069 9582 7070
rect 9573 7043 9574 7069
rect 9573 7042 9582 7043
rect 9610 7042 9634 7070
rect 9662 7042 9686 7070
rect 9714 7069 9738 7070
rect 9766 7069 9790 7070
rect 9724 7043 9738 7069
rect 9786 7043 9790 7069
rect 9714 7042 9738 7043
rect 9766 7042 9790 7043
rect 9818 7069 9842 7070
rect 9870 7069 9894 7070
rect 9818 7043 9822 7069
rect 9870 7043 9884 7069
rect 9818 7042 9842 7043
rect 9870 7042 9894 7043
rect 9922 7042 9946 7070
rect 9974 7042 9998 7070
rect 10026 7069 10035 7070
rect 10034 7043 10035 7069
rect 10026 7042 10035 7043
rect 9573 7037 10035 7042
rect 9702 6874 9730 6879
rect 9478 6873 9730 6874
rect 9478 6847 9703 6873
rect 9729 6847 9730 6873
rect 9478 6846 9730 6847
rect 9478 6481 9506 6846
rect 9702 6841 9730 6846
rect 10206 6874 10234 7182
rect 10374 6874 10402 6879
rect 10206 6873 10402 6874
rect 10206 6847 10207 6873
rect 10233 6847 10375 6873
rect 10401 6847 10402 6873
rect 10206 6846 10402 6847
rect 10206 6841 10234 6846
rect 9478 6455 9479 6481
rect 9505 6455 9506 6481
rect 9478 5866 9506 6455
rect 10374 6706 10402 6846
rect 10374 6481 10402 6678
rect 10374 6455 10375 6481
rect 10401 6455 10402 6481
rect 10374 6425 10402 6455
rect 10374 6399 10375 6425
rect 10401 6399 10402 6425
rect 9573 6286 10035 6291
rect 9573 6285 9582 6286
rect 9573 6259 9574 6285
rect 9573 6258 9582 6259
rect 9610 6258 9634 6286
rect 9662 6258 9686 6286
rect 9714 6285 9738 6286
rect 9766 6285 9790 6286
rect 9724 6259 9738 6285
rect 9786 6259 9790 6285
rect 9714 6258 9738 6259
rect 9766 6258 9790 6259
rect 9818 6285 9842 6286
rect 9870 6285 9894 6286
rect 9818 6259 9822 6285
rect 9870 6259 9884 6285
rect 9818 6258 9842 6259
rect 9870 6258 9894 6259
rect 9922 6258 9946 6286
rect 9974 6258 9998 6286
rect 10026 6285 10035 6286
rect 10034 6259 10035 6285
rect 10026 6258 10035 6259
rect 9573 6253 10035 6258
rect 10038 6089 10066 6095
rect 10038 6063 10039 6089
rect 10065 6063 10066 6089
rect 9534 5866 9562 5871
rect 9478 5838 9534 5866
rect 8974 5697 9002 5703
rect 8974 5671 8975 5697
rect 9001 5671 9002 5697
rect 8974 5642 9002 5671
rect 9534 5697 9562 5838
rect 10038 5866 10066 6063
rect 10374 6090 10402 6399
rect 10486 6090 10514 6095
rect 10374 6089 10514 6090
rect 10374 6063 10375 6089
rect 10401 6063 10487 6089
rect 10513 6063 10514 6089
rect 10374 6062 10514 6063
rect 10374 6057 10402 6062
rect 10486 6057 10514 6062
rect 10038 5833 10066 5838
rect 9534 5671 9535 5697
rect 9561 5671 9562 5697
rect 9534 5665 9562 5671
rect 10430 5697 10458 5703
rect 10430 5671 10431 5697
rect 10457 5671 10458 5697
rect 8974 5641 9058 5642
rect 8974 5615 8975 5641
rect 9001 5615 9058 5641
rect 8974 5614 9058 5615
rect 8974 5609 9002 5614
rect 9030 4522 9058 5614
rect 10430 5641 10458 5671
rect 10430 5615 10431 5641
rect 10457 5615 10458 5641
rect 9573 5502 10035 5507
rect 9573 5501 9582 5502
rect 9573 5475 9574 5501
rect 9573 5474 9582 5475
rect 9610 5474 9634 5502
rect 9662 5474 9686 5502
rect 9714 5501 9738 5502
rect 9766 5501 9790 5502
rect 9724 5475 9738 5501
rect 9786 5475 9790 5501
rect 9714 5474 9738 5475
rect 9766 5474 9790 5475
rect 9818 5501 9842 5502
rect 9870 5501 9894 5502
rect 9818 5475 9822 5501
rect 9870 5475 9884 5501
rect 9818 5474 9842 5475
rect 9870 5474 9894 5475
rect 9922 5474 9946 5502
rect 9974 5474 9998 5502
rect 10026 5501 10035 5502
rect 10034 5475 10035 5501
rect 10026 5474 10035 5475
rect 9573 5469 10035 5474
rect 9534 5306 9562 5311
rect 9534 4913 9562 5278
rect 9814 5306 9842 5311
rect 9814 5259 9842 5278
rect 10262 5306 10290 5311
rect 10430 5306 10458 5615
rect 10486 5306 10514 5311
rect 10262 5305 10514 5306
rect 10262 5279 10263 5305
rect 10289 5279 10487 5305
rect 10513 5279 10514 5305
rect 10262 5278 10514 5279
rect 9534 4887 9535 4913
rect 9561 4887 9562 4913
rect 9534 4881 9562 4887
rect 10038 5250 10066 5255
rect 10038 4802 10066 5222
rect 10262 4913 10290 5278
rect 10486 5273 10514 5278
rect 10262 4887 10263 4913
rect 10289 4887 10290 4913
rect 10262 4857 10290 4887
rect 10262 4831 10263 4857
rect 10289 4831 10290 4857
rect 10038 4774 10122 4802
rect 9573 4718 10035 4723
rect 9573 4717 9582 4718
rect 9573 4691 9574 4717
rect 9573 4690 9582 4691
rect 9610 4690 9634 4718
rect 9662 4690 9686 4718
rect 9714 4717 9738 4718
rect 9766 4717 9790 4718
rect 9724 4691 9738 4717
rect 9786 4691 9790 4717
rect 9714 4690 9738 4691
rect 9766 4690 9790 4691
rect 9818 4717 9842 4718
rect 9870 4717 9894 4718
rect 9818 4691 9822 4717
rect 9870 4691 9884 4717
rect 9818 4690 9842 4691
rect 9870 4690 9894 4691
rect 9922 4690 9946 4718
rect 9974 4690 9998 4718
rect 10026 4717 10035 4718
rect 10034 4691 10035 4717
rect 10026 4690 10035 4691
rect 9573 4685 10035 4690
rect 10094 4634 10122 4774
rect 8806 3761 8834 3766
rect 8974 4129 9002 4135
rect 8974 4103 8975 4129
rect 9001 4103 9002 4129
rect 8022 3738 8050 3743
rect 7798 3737 8050 3738
rect 7798 3711 7799 3737
rect 7825 3711 8023 3737
rect 8049 3711 8050 3737
rect 7798 3710 8050 3711
rect 7798 3705 7826 3710
rect 8022 3458 8050 3710
rect 8470 3738 8498 3743
rect 8470 3691 8498 3710
rect 8974 3738 9002 4103
rect 8022 3425 8050 3430
rect 8302 3458 8330 3463
rect 8302 3346 8330 3430
rect 8974 3402 9002 3710
rect 8414 3346 8442 3351
rect 8302 3345 8442 3346
rect 8302 3319 8303 3345
rect 8329 3319 8415 3345
rect 8441 3319 8442 3345
rect 8302 3318 8442 3319
rect 8302 3313 8330 3318
rect 8414 3313 8442 3318
rect 8974 3345 9002 3374
rect 8974 3319 8975 3345
rect 9001 3319 9002 3345
rect 8974 3313 9002 3319
rect 7574 2927 7575 2953
rect 7601 2927 7602 2953
rect 7073 2758 7535 2763
rect 7073 2757 7082 2758
rect 7073 2731 7074 2757
rect 7073 2730 7082 2731
rect 7110 2730 7134 2758
rect 7162 2730 7186 2758
rect 7214 2757 7238 2758
rect 7266 2757 7290 2758
rect 7224 2731 7238 2757
rect 7286 2731 7290 2757
rect 7214 2730 7238 2731
rect 7266 2730 7290 2731
rect 7318 2757 7342 2758
rect 7370 2757 7394 2758
rect 7318 2731 7322 2757
rect 7370 2731 7384 2757
rect 7318 2730 7342 2731
rect 7370 2730 7394 2731
rect 7422 2730 7446 2758
rect 7474 2730 7498 2758
rect 7526 2757 7535 2758
rect 7534 2731 7535 2757
rect 7526 2730 7535 2731
rect 7073 2725 7535 2730
rect 7014 2169 7042 2534
rect 7574 2562 7602 2927
rect 8470 3009 8498 3015
rect 8470 2983 8471 3009
rect 8497 2983 8498 3009
rect 8470 2953 8498 2983
rect 8470 2927 8471 2953
rect 8497 2927 8498 2953
rect 7574 2529 7602 2534
rect 8078 2562 8106 2567
rect 8078 2515 8106 2534
rect 8470 2506 8498 2927
rect 8470 2473 8498 2478
rect 8974 2562 9002 2567
rect 9030 2562 9058 4494
rect 10038 4606 10122 4634
rect 10038 4521 10066 4606
rect 10038 4495 10039 4521
rect 10065 4495 10066 4521
rect 10038 4489 10066 4495
rect 10262 4522 10290 4831
rect 10262 4475 10290 4494
rect 10486 4522 10514 4527
rect 10486 4475 10514 4494
rect 9478 4129 9506 4135
rect 9478 4103 9479 4129
rect 9505 4103 9506 4129
rect 9478 3738 9506 4103
rect 10430 4129 10458 4135
rect 10430 4103 10431 4129
rect 10457 4103 10458 4129
rect 10430 4074 10458 4103
rect 10430 4073 10514 4074
rect 10430 4047 10431 4073
rect 10457 4047 10514 4073
rect 10430 4046 10514 4047
rect 10430 4041 10458 4046
rect 9573 3934 10035 3939
rect 9573 3933 9582 3934
rect 9573 3907 9574 3933
rect 9573 3906 9582 3907
rect 9610 3906 9634 3934
rect 9662 3906 9686 3934
rect 9714 3933 9738 3934
rect 9766 3933 9790 3934
rect 9724 3907 9738 3933
rect 9786 3907 9790 3933
rect 9714 3906 9738 3907
rect 9766 3906 9790 3907
rect 9818 3933 9842 3934
rect 9870 3933 9894 3934
rect 9818 3907 9822 3933
rect 9870 3907 9884 3933
rect 9818 3906 9842 3907
rect 9870 3906 9894 3907
rect 9922 3906 9946 3934
rect 9974 3906 9998 3934
rect 10026 3933 10035 3934
rect 10034 3907 10035 3933
rect 10026 3906 10035 3907
rect 9573 3901 10035 3906
rect 9478 3402 9506 3710
rect 9814 3738 9842 3743
rect 9814 3691 9842 3710
rect 10486 3738 10514 4046
rect 9478 3345 9506 3374
rect 10486 3458 10514 3710
rect 9478 3319 9479 3345
rect 9505 3319 9506 3345
rect 8974 2561 9058 2562
rect 8974 2535 8975 2561
rect 9001 2535 9058 2561
rect 8974 2534 9058 2535
rect 9366 2562 9394 2567
rect 8974 2506 9002 2534
rect 8246 2282 8274 2287
rect 7014 2143 7015 2169
rect 7041 2143 7042 2169
rect 7014 2058 7042 2143
rect 7014 2025 7042 2030
rect 7518 2169 7546 2175
rect 7518 2143 7519 2169
rect 7545 2143 7546 2169
rect 7518 2058 7546 2143
rect 7518 2025 7546 2030
rect 7073 1974 7535 1979
rect 7073 1973 7082 1974
rect 7073 1947 7074 1973
rect 7073 1946 7082 1947
rect 7110 1946 7134 1974
rect 7162 1946 7186 1974
rect 7214 1973 7238 1974
rect 7266 1973 7290 1974
rect 7224 1947 7238 1973
rect 7286 1947 7290 1973
rect 7214 1946 7238 1947
rect 7266 1946 7290 1947
rect 7318 1973 7342 1974
rect 7370 1973 7394 1974
rect 7318 1947 7322 1973
rect 7370 1947 7384 1973
rect 7318 1946 7342 1947
rect 7370 1946 7394 1947
rect 7422 1946 7446 1974
rect 7474 1946 7498 1974
rect 7526 1973 7535 1974
rect 7534 1947 7535 1973
rect 7526 1946 7535 1947
rect 7073 1941 7535 1946
rect 7462 1890 7490 1895
rect 7462 1777 7490 1862
rect 7462 1751 7463 1777
rect 7489 1751 7490 1777
rect 7462 1745 7490 1751
rect 6902 462 7042 490
rect 7014 400 7042 462
rect 8246 400 8274 2254
rect 8358 2225 8386 2231
rect 8358 2199 8359 2225
rect 8385 2199 8386 2225
rect 8358 2169 8386 2199
rect 8358 2143 8359 2169
rect 8385 2143 8386 2169
rect 8358 1777 8386 2143
rect 8358 1751 8359 1777
rect 8385 1751 8386 1777
rect 8358 1722 8386 1751
rect 8974 1778 9002 2478
rect 8974 1745 9002 1750
rect 9366 1834 9394 2534
rect 9478 2561 9506 3319
rect 10430 3345 10458 3351
rect 10430 3319 10431 3345
rect 10457 3319 10458 3345
rect 10430 3290 10458 3319
rect 10486 3290 10514 3430
rect 10430 3289 10514 3290
rect 10430 3263 10431 3289
rect 10457 3263 10514 3289
rect 10430 3262 10514 3263
rect 10430 3257 10458 3262
rect 9573 3150 10035 3155
rect 9573 3149 9582 3150
rect 9573 3123 9574 3149
rect 9573 3122 9582 3123
rect 9610 3122 9634 3150
rect 9662 3122 9686 3150
rect 9714 3149 9738 3150
rect 9766 3149 9790 3150
rect 9724 3123 9738 3149
rect 9786 3123 9790 3149
rect 9714 3122 9738 3123
rect 9766 3122 9790 3123
rect 9818 3149 9842 3150
rect 9870 3149 9894 3150
rect 9818 3123 9822 3149
rect 9870 3123 9884 3149
rect 9818 3122 9842 3123
rect 9870 3122 9894 3123
rect 9922 3122 9946 3150
rect 9974 3122 9998 3150
rect 10026 3149 10035 3150
rect 10034 3123 10035 3149
rect 10026 3122 10035 3123
rect 9573 3117 10035 3122
rect 10318 2954 10346 2959
rect 10486 2954 10514 3262
rect 10318 2953 10514 2954
rect 10318 2927 10319 2953
rect 10345 2927 10487 2953
rect 10513 2927 10514 2953
rect 10318 2926 10514 2927
rect 10318 2921 10346 2926
rect 9478 2535 9479 2561
rect 9505 2535 9506 2561
rect 9366 1777 9394 1806
rect 9366 1751 9367 1777
rect 9393 1751 9394 1777
rect 9366 1745 9394 1751
rect 9422 2450 9450 2455
rect 8358 1675 8386 1694
rect 9422 1218 9450 2422
rect 9478 2226 9506 2535
rect 10430 2561 10458 2567
rect 10430 2535 10431 2561
rect 10457 2535 10458 2561
rect 10430 2506 10458 2535
rect 10486 2506 10514 2926
rect 10430 2505 10514 2506
rect 10430 2479 10431 2505
rect 10457 2479 10514 2505
rect 10430 2478 10514 2479
rect 10430 2473 10458 2478
rect 9573 2366 10035 2371
rect 9573 2365 9582 2366
rect 9573 2339 9574 2365
rect 9573 2338 9582 2339
rect 9610 2338 9634 2366
rect 9662 2338 9686 2366
rect 9714 2365 9738 2366
rect 9766 2365 9790 2366
rect 9724 2339 9738 2365
rect 9786 2339 9790 2365
rect 9714 2338 9738 2339
rect 9766 2338 9790 2339
rect 9818 2365 9842 2366
rect 9870 2365 9894 2366
rect 9818 2339 9822 2365
rect 9870 2339 9884 2365
rect 9818 2338 9842 2339
rect 9870 2338 9894 2339
rect 9922 2338 9946 2366
rect 9974 2338 9998 2366
rect 10026 2365 10035 2366
rect 10034 2339 10035 2365
rect 10026 2338 10035 2339
rect 9573 2333 10035 2338
rect 9478 2193 9506 2198
rect 10038 2226 10066 2231
rect 10038 2169 10066 2198
rect 10038 2143 10039 2169
rect 10065 2143 10066 2169
rect 10038 2137 10066 2143
rect 10542 2114 10570 7966
rect 11438 7657 11466 8023
rect 11438 7631 11439 7657
rect 11465 7631 11466 7657
rect 11438 7265 11466 7631
rect 11438 7239 11439 7265
rect 11465 7239 11466 7265
rect 11438 6874 11466 7239
rect 11774 8442 11802 8447
rect 11942 8442 11970 8447
rect 11774 8441 11970 8442
rect 11774 8415 11775 8441
rect 11801 8415 11943 8441
rect 11969 8415 11970 8441
rect 11774 8414 11970 8415
rect 11774 8050 11802 8414
rect 11942 8409 11970 8414
rect 11886 8050 11914 8055
rect 11774 8049 11914 8050
rect 11774 8023 11775 8049
rect 11801 8023 11887 8049
rect 11913 8023 11914 8049
rect 11774 8022 11914 8023
rect 11774 7658 11802 8022
rect 11886 8017 11914 8022
rect 11886 7658 11914 7663
rect 11774 7657 11914 7658
rect 11774 7631 11775 7657
rect 11801 7631 11887 7657
rect 11913 7631 11914 7657
rect 11774 7630 11914 7631
rect 11774 7266 11802 7630
rect 11886 7625 11914 7630
rect 11886 7266 11914 7271
rect 11774 7265 11914 7266
rect 11774 7239 11775 7265
rect 11801 7239 11887 7265
rect 11913 7239 11914 7265
rect 11774 7238 11914 7239
rect 11718 6874 11746 6879
rect 11774 6874 11802 7238
rect 11886 7233 11914 7238
rect 11998 7266 12026 8806
rect 12054 8801 12082 8806
rect 12278 8801 12306 8806
rect 13006 8833 13090 8834
rect 13006 8807 13063 8833
rect 13089 8807 13090 8833
rect 13006 8806 13090 8807
rect 13006 8442 13034 8806
rect 13062 8801 13090 8806
rect 13510 8833 13538 8839
rect 13734 8834 13762 8839
rect 13790 8834 13818 9198
rect 14014 9193 14042 9198
rect 13510 8807 13511 8833
rect 13537 8807 13538 8833
rect 12894 8441 13034 8442
rect 12894 8415 13007 8441
rect 13033 8415 13034 8441
rect 12894 8414 13034 8415
rect 12073 8246 12535 8251
rect 12073 8245 12082 8246
rect 12073 8219 12074 8245
rect 12073 8218 12082 8219
rect 12110 8218 12134 8246
rect 12162 8218 12186 8246
rect 12214 8245 12238 8246
rect 12266 8245 12290 8246
rect 12224 8219 12238 8245
rect 12286 8219 12290 8245
rect 12214 8218 12238 8219
rect 12266 8218 12290 8219
rect 12318 8245 12342 8246
rect 12370 8245 12394 8246
rect 12318 8219 12322 8245
rect 12370 8219 12384 8245
rect 12318 8218 12342 8219
rect 12370 8218 12394 8219
rect 12422 8218 12446 8246
rect 12474 8218 12498 8246
rect 12526 8245 12535 8246
rect 12534 8219 12535 8245
rect 12526 8218 12535 8219
rect 12073 8213 12535 8218
rect 12894 8050 12922 8414
rect 13006 8409 13034 8414
rect 13454 8442 13482 8447
rect 13510 8442 13538 8807
rect 13678 8833 13818 8834
rect 13678 8807 13735 8833
rect 13761 8807 13818 8833
rect 13678 8806 13818 8807
rect 13678 8442 13706 8806
rect 13734 8801 13762 8806
rect 13454 8441 13706 8442
rect 13454 8415 13455 8441
rect 13481 8415 13679 8441
rect 13705 8415 13706 8441
rect 13454 8414 13706 8415
rect 12838 8049 12922 8050
rect 12838 8023 12895 8049
rect 12921 8023 12922 8049
rect 12838 8022 12922 8023
rect 12838 7658 12866 8022
rect 12894 8017 12922 8022
rect 13454 8050 13482 8414
rect 13678 8409 13706 8414
rect 14406 8442 14434 10066
rect 15078 10009 15106 10375
rect 15358 10794 15386 11158
rect 15470 11153 15498 11158
rect 15862 11074 15890 11551
rect 15582 10794 15610 10799
rect 15358 10793 15610 10794
rect 15358 10767 15359 10793
rect 15385 10767 15583 10793
rect 15609 10767 15610 10793
rect 15358 10766 15610 10767
rect 15358 10402 15386 10766
rect 15582 10761 15610 10766
rect 15470 10402 15498 10407
rect 15358 10401 15498 10402
rect 15358 10375 15359 10401
rect 15385 10375 15471 10401
rect 15497 10375 15498 10401
rect 15358 10374 15498 10375
rect 15358 10094 15386 10374
rect 15470 10369 15498 10374
rect 15078 9983 15079 10009
rect 15105 9983 15106 10009
rect 13566 8050 13594 8055
rect 13454 8049 13594 8050
rect 13454 8023 13455 8049
rect 13481 8023 13567 8049
rect 13593 8023 13594 8049
rect 13454 8022 13594 8023
rect 12782 7657 12866 7658
rect 12782 7631 12839 7657
rect 12865 7631 12866 7657
rect 12782 7630 12866 7631
rect 12073 7462 12535 7467
rect 12073 7461 12082 7462
rect 12073 7435 12074 7461
rect 12073 7434 12082 7435
rect 12110 7434 12134 7462
rect 12162 7434 12186 7462
rect 12214 7461 12238 7462
rect 12266 7461 12290 7462
rect 12224 7435 12238 7461
rect 12286 7435 12290 7461
rect 12214 7434 12238 7435
rect 12266 7434 12290 7435
rect 12318 7461 12342 7462
rect 12370 7461 12394 7462
rect 12318 7435 12322 7461
rect 12370 7435 12384 7461
rect 12318 7434 12342 7435
rect 12370 7434 12394 7435
rect 12422 7434 12446 7462
rect 12474 7434 12498 7462
rect 12526 7461 12535 7462
rect 12534 7435 12535 7461
rect 12526 7434 12535 7435
rect 12073 7429 12535 7434
rect 11830 6874 11858 6879
rect 11438 6873 11522 6874
rect 11438 6847 11439 6873
rect 11465 6847 11522 6873
rect 11438 6846 11522 6847
rect 11438 6841 11466 6846
rect 11494 6481 11522 6846
rect 11718 6873 11858 6874
rect 11718 6847 11719 6873
rect 11745 6847 11831 6873
rect 11857 6847 11858 6873
rect 11718 6846 11858 6847
rect 11718 6841 11746 6846
rect 11494 6455 11495 6481
rect 11521 6455 11522 6481
rect 11494 4521 11522 6455
rect 11830 6706 11858 6846
rect 11550 6089 11578 6095
rect 11550 6063 11551 6089
rect 11577 6063 11578 6089
rect 11550 5866 11578 6063
rect 11830 6090 11858 6678
rect 11998 6482 12026 7238
rect 12782 7265 12810 7630
rect 12838 7625 12866 7630
rect 13398 7658 13426 7663
rect 13454 7658 13482 8022
rect 13566 8017 13594 8022
rect 13510 7658 13538 7663
rect 13398 7657 13538 7658
rect 13398 7631 13399 7657
rect 13425 7631 13511 7657
rect 13537 7631 13538 7657
rect 13398 7630 13538 7631
rect 13398 7625 13426 7630
rect 12782 7239 12783 7265
rect 12809 7239 12810 7265
rect 12073 6678 12535 6683
rect 12073 6677 12082 6678
rect 12073 6651 12074 6677
rect 12073 6650 12082 6651
rect 12110 6650 12134 6678
rect 12162 6650 12186 6678
rect 12214 6677 12238 6678
rect 12266 6677 12290 6678
rect 12224 6651 12238 6677
rect 12286 6651 12290 6677
rect 12214 6650 12238 6651
rect 12266 6650 12290 6651
rect 12318 6677 12342 6678
rect 12370 6677 12394 6678
rect 12318 6651 12322 6677
rect 12370 6651 12384 6677
rect 12318 6650 12342 6651
rect 12370 6650 12394 6651
rect 12422 6650 12446 6678
rect 12474 6650 12498 6678
rect 12526 6677 12535 6678
rect 12534 6651 12535 6677
rect 12526 6650 12535 6651
rect 12073 6645 12535 6650
rect 12166 6482 12194 6487
rect 11998 6481 12194 6482
rect 11998 6455 11999 6481
rect 12025 6455 12167 6481
rect 12193 6455 12194 6481
rect 11998 6454 12194 6455
rect 11942 6090 11970 6095
rect 11830 6089 11970 6090
rect 11830 6063 11831 6089
rect 11857 6063 11943 6089
rect 11969 6063 11970 6089
rect 11830 6062 11970 6063
rect 11830 6057 11858 6062
rect 11550 5642 11578 5838
rect 11550 5305 11578 5614
rect 11942 5698 11970 6062
rect 11550 5279 11551 5305
rect 11577 5279 11578 5305
rect 11550 5250 11578 5279
rect 11830 5306 11858 5311
rect 11942 5306 11970 5670
rect 11830 5305 11970 5306
rect 11830 5279 11831 5305
rect 11857 5279 11943 5305
rect 11969 5279 11970 5305
rect 11830 5278 11970 5279
rect 11830 5273 11858 5278
rect 11942 5273 11970 5278
rect 11550 5217 11578 5222
rect 11494 4495 11495 4521
rect 11521 4495 11522 4521
rect 11494 4489 11522 4495
rect 11774 4522 11802 4527
rect 11774 4475 11802 4494
rect 11942 4522 11970 4527
rect 11998 4522 12026 6454
rect 12166 6449 12194 6454
rect 12073 5894 12535 5899
rect 12073 5893 12082 5894
rect 12073 5867 12074 5893
rect 12073 5866 12082 5867
rect 12110 5866 12134 5894
rect 12162 5866 12186 5894
rect 12214 5893 12238 5894
rect 12266 5893 12290 5894
rect 12224 5867 12238 5893
rect 12286 5867 12290 5893
rect 12214 5866 12238 5867
rect 12266 5866 12290 5867
rect 12318 5893 12342 5894
rect 12370 5893 12394 5894
rect 12318 5867 12322 5893
rect 12370 5867 12384 5893
rect 12318 5866 12342 5867
rect 12370 5866 12394 5867
rect 12422 5866 12446 5894
rect 12474 5866 12498 5894
rect 12526 5893 12535 5894
rect 12534 5867 12535 5893
rect 12526 5866 12535 5867
rect 12073 5861 12535 5866
rect 12334 5697 12362 5703
rect 12334 5671 12335 5697
rect 12361 5671 12362 5697
rect 12334 5642 12362 5671
rect 12502 5698 12530 5703
rect 12502 5651 12530 5670
rect 12726 5698 12754 5703
rect 12334 5609 12362 5614
rect 12614 5642 12642 5647
rect 12073 5110 12535 5115
rect 12073 5109 12082 5110
rect 12073 5083 12074 5109
rect 12073 5082 12082 5083
rect 12110 5082 12134 5110
rect 12162 5082 12186 5110
rect 12214 5109 12238 5110
rect 12266 5109 12290 5110
rect 12224 5083 12238 5109
rect 12286 5083 12290 5109
rect 12214 5082 12238 5083
rect 12266 5082 12290 5083
rect 12318 5109 12342 5110
rect 12370 5109 12394 5110
rect 12318 5083 12322 5109
rect 12370 5083 12384 5109
rect 12318 5082 12342 5083
rect 12370 5082 12394 5083
rect 12422 5082 12446 5110
rect 12474 5082 12498 5110
rect 12526 5109 12535 5110
rect 12534 5083 12535 5109
rect 12526 5082 12535 5083
rect 12073 5077 12535 5082
rect 12614 5026 12642 5614
rect 11970 4494 12026 4522
rect 12334 4998 12642 5026
rect 12726 5306 12754 5670
rect 12334 4913 12362 4998
rect 12334 4887 12335 4913
rect 12361 4887 12362 4913
rect 11382 4242 11410 4247
rect 10878 3793 10906 3799
rect 10878 3767 10879 3793
rect 10905 3767 10906 3793
rect 10878 3738 10906 3767
rect 10878 3691 10906 3710
rect 11382 3737 11410 4214
rect 11382 3711 11383 3737
rect 11409 3711 11410 3737
rect 10878 2953 10906 2959
rect 10878 2927 10879 2953
rect 10905 2927 10906 2953
rect 10542 2081 10570 2086
rect 10822 2225 10850 2231
rect 10822 2199 10823 2225
rect 10849 2199 10850 2225
rect 10822 2169 10850 2199
rect 10822 2143 10823 2169
rect 10849 2143 10850 2169
rect 10822 2114 10850 2143
rect 10878 2170 10906 2927
rect 11382 2953 11410 3711
rect 11382 2927 11383 2953
rect 11409 2927 11410 2953
rect 11382 2921 11410 2927
rect 11774 4129 11802 4135
rect 11774 4103 11775 4129
rect 11801 4103 11802 4129
rect 11774 4073 11802 4103
rect 11774 4047 11775 4073
rect 11801 4047 11802 4073
rect 11774 3738 11802 4047
rect 11774 3290 11802 3710
rect 11830 3738 11858 3743
rect 11942 3738 11970 4494
rect 12334 4410 12362 4887
rect 12614 4914 12642 4919
rect 12726 4914 12754 5278
rect 12614 4913 12754 4914
rect 12614 4887 12615 4913
rect 12641 4887 12727 4913
rect 12753 4887 12754 4913
rect 12614 4886 12754 4887
rect 12614 4881 12642 4886
rect 12726 4881 12754 4886
rect 11998 4382 12362 4410
rect 11998 4242 12026 4382
rect 12073 4326 12535 4331
rect 12073 4325 12082 4326
rect 12073 4299 12074 4325
rect 12073 4298 12082 4299
rect 12110 4298 12134 4326
rect 12162 4298 12186 4326
rect 12214 4325 12238 4326
rect 12266 4325 12290 4326
rect 12224 4299 12238 4325
rect 12286 4299 12290 4325
rect 12214 4298 12238 4299
rect 12266 4298 12290 4299
rect 12318 4325 12342 4326
rect 12370 4325 12394 4326
rect 12318 4299 12322 4325
rect 12370 4299 12384 4325
rect 12318 4298 12342 4299
rect 12370 4298 12394 4299
rect 12422 4298 12446 4326
rect 12474 4298 12498 4326
rect 12526 4325 12535 4326
rect 12534 4299 12535 4325
rect 12526 4298 12535 4299
rect 12073 4293 12535 4298
rect 11998 4186 12082 4214
rect 11830 3737 11970 3738
rect 11830 3711 11831 3737
rect 11857 3711 11943 3737
rect 11969 3711 11970 3737
rect 11830 3710 11970 3711
rect 11830 3705 11858 3710
rect 11942 3346 11970 3710
rect 12054 3626 12082 4186
rect 11942 3313 11970 3318
rect 11998 3598 12082 3626
rect 11998 3345 12026 3598
rect 12073 3542 12535 3547
rect 12073 3541 12082 3542
rect 12073 3515 12074 3541
rect 12073 3514 12082 3515
rect 12110 3514 12134 3542
rect 12162 3514 12186 3542
rect 12214 3541 12238 3542
rect 12266 3541 12290 3542
rect 12224 3515 12238 3541
rect 12286 3515 12290 3541
rect 12214 3514 12238 3515
rect 12266 3514 12290 3515
rect 12318 3541 12342 3542
rect 12370 3541 12394 3542
rect 12318 3515 12322 3541
rect 12370 3515 12384 3541
rect 12318 3514 12342 3515
rect 12370 3514 12394 3515
rect 12422 3514 12446 3542
rect 12474 3514 12498 3542
rect 12526 3541 12535 3542
rect 12534 3515 12535 3541
rect 12526 3514 12535 3515
rect 12073 3509 12535 3514
rect 11998 3319 11999 3345
rect 12025 3319 12026 3345
rect 10878 2137 10906 2142
rect 11382 2170 11410 2175
rect 10822 2081 10850 2086
rect 11382 1834 11410 2142
rect 9702 1778 9730 1783
rect 9814 1778 9842 1783
rect 9730 1777 9842 1778
rect 9730 1751 9815 1777
rect 9841 1751 9842 1777
rect 9730 1750 9842 1751
rect 9702 1712 9730 1750
rect 9814 1745 9842 1750
rect 10710 1778 10738 1783
rect 9573 1582 10035 1587
rect 9573 1581 9582 1582
rect 9573 1555 9574 1581
rect 9573 1554 9582 1555
rect 9610 1554 9634 1582
rect 9662 1554 9686 1582
rect 9714 1581 9738 1582
rect 9766 1581 9790 1582
rect 9724 1555 9738 1581
rect 9786 1555 9790 1581
rect 9714 1554 9738 1555
rect 9766 1554 9790 1555
rect 9818 1581 9842 1582
rect 9870 1581 9894 1582
rect 9818 1555 9822 1581
rect 9870 1555 9884 1581
rect 9818 1554 9842 1555
rect 9870 1554 9894 1555
rect 9922 1554 9946 1582
rect 9974 1554 9998 1582
rect 10026 1581 10035 1582
rect 10034 1555 10035 1581
rect 10026 1554 10035 1555
rect 9573 1549 10035 1554
rect 9422 1190 9506 1218
rect 9478 400 9506 1190
rect 10710 400 10738 1750
rect 11382 1777 11410 1806
rect 11774 2170 11802 3262
rect 11382 1751 11383 1777
rect 11409 1751 11410 1777
rect 11382 1745 11410 1751
rect 11662 1778 11690 1783
rect 11774 1778 11802 2142
rect 11942 2170 11970 2175
rect 11942 2123 11970 2142
rect 11998 2058 12026 3319
rect 12334 3346 12362 3351
rect 12446 3346 12474 3351
rect 12362 3345 12474 3346
rect 12362 3319 12447 3345
rect 12473 3319 12474 3345
rect 12362 3318 12474 3319
rect 12334 3280 12362 3318
rect 12446 3009 12474 3318
rect 12446 2983 12447 3009
rect 12473 2983 12474 3009
rect 12446 2954 12474 2983
rect 12446 2907 12474 2926
rect 12073 2758 12535 2763
rect 12073 2757 12082 2758
rect 12073 2731 12074 2757
rect 12073 2730 12082 2731
rect 12110 2730 12134 2758
rect 12162 2730 12186 2758
rect 12214 2757 12238 2758
rect 12266 2757 12290 2758
rect 12224 2731 12238 2757
rect 12286 2731 12290 2757
rect 12214 2730 12238 2731
rect 12266 2730 12290 2731
rect 12318 2757 12342 2758
rect 12370 2757 12394 2758
rect 12318 2731 12322 2757
rect 12370 2731 12384 2757
rect 12318 2730 12342 2731
rect 12370 2730 12394 2731
rect 12422 2730 12446 2758
rect 12474 2730 12498 2758
rect 12526 2757 12535 2758
rect 12534 2731 12535 2757
rect 12526 2730 12535 2731
rect 12073 2725 12535 2730
rect 12222 2561 12250 2567
rect 12222 2535 12223 2561
rect 12249 2535 12250 2561
rect 12222 2058 12250 2535
rect 11662 1777 11802 1778
rect 11662 1751 11663 1777
rect 11689 1751 11775 1777
rect 11801 1751 11802 1777
rect 11662 1750 11802 1751
rect 11662 1745 11690 1750
rect 11774 1745 11802 1750
rect 11942 2030 12250 2058
rect 11942 400 11970 2030
rect 12073 1974 12535 1979
rect 12073 1973 12082 1974
rect 12073 1947 12074 1973
rect 12073 1946 12082 1947
rect 12110 1946 12134 1974
rect 12162 1946 12186 1974
rect 12214 1973 12238 1974
rect 12266 1973 12290 1974
rect 12224 1947 12238 1973
rect 12286 1947 12290 1973
rect 12214 1946 12238 1947
rect 12266 1946 12290 1947
rect 12318 1973 12342 1974
rect 12370 1973 12394 1974
rect 12318 1947 12322 1973
rect 12370 1947 12384 1973
rect 12318 1946 12342 1947
rect 12370 1946 12394 1947
rect 12422 1946 12446 1974
rect 12474 1946 12498 1974
rect 12526 1973 12535 1974
rect 12534 1947 12535 1973
rect 12526 1946 12535 1947
rect 12073 1941 12535 1946
rect 1022 350 1218 378
rect 2072 0 2128 400
rect 3304 0 3360 400
rect 4536 0 4592 400
rect 5768 0 5824 400
rect 7000 0 7056 400
rect 8232 0 8288 400
rect 9464 0 9520 400
rect 10696 0 10752 400
rect 11928 0 11984 400
rect 12782 378 12810 7239
rect 13118 7266 13146 7271
rect 13118 7219 13146 7238
rect 13454 7266 13482 7630
rect 13510 7625 13538 7630
rect 14406 7657 14434 8414
rect 14462 9618 14490 9623
rect 14462 9282 14490 9590
rect 14798 9618 14826 9623
rect 14798 9571 14826 9590
rect 15078 9618 15106 9983
rect 15078 9585 15106 9590
rect 15246 10066 15386 10094
rect 15750 10066 15778 10071
rect 15246 9618 15274 10066
rect 15526 10010 15554 10015
rect 15750 10010 15778 10038
rect 15470 10009 15778 10010
rect 15470 9983 15527 10009
rect 15553 9983 15751 10009
rect 15777 9983 15778 10009
rect 15470 9982 15778 9983
rect 15470 9618 15498 9982
rect 15526 9977 15554 9982
rect 15750 9977 15778 9982
rect 15246 9617 15498 9618
rect 15246 9591 15247 9617
rect 15273 9591 15471 9617
rect 15497 9591 15498 9617
rect 15246 9590 15498 9591
rect 14573 9422 15035 9427
rect 14573 9421 14582 9422
rect 14573 9395 14574 9421
rect 14573 9394 14582 9395
rect 14610 9394 14634 9422
rect 14662 9394 14686 9422
rect 14714 9421 14738 9422
rect 14766 9421 14790 9422
rect 14724 9395 14738 9421
rect 14786 9395 14790 9421
rect 14714 9394 14738 9395
rect 14766 9394 14790 9395
rect 14818 9421 14842 9422
rect 14870 9421 14894 9422
rect 14818 9395 14822 9421
rect 14870 9395 14884 9421
rect 14818 9394 14842 9395
rect 14870 9394 14894 9395
rect 14922 9394 14946 9422
rect 14974 9394 14998 9422
rect 15026 9421 15035 9422
rect 15034 9395 15035 9421
rect 15026 9394 15035 9395
rect 14573 9389 15035 9394
rect 14462 8834 14490 9254
rect 15134 9338 15162 9343
rect 15246 9338 15274 9590
rect 15470 9585 15498 9590
rect 15750 9618 15778 9623
rect 15162 9310 15274 9338
rect 14798 9225 14826 9231
rect 14798 9199 14799 9225
rect 14825 9199 14826 9225
rect 14798 8834 14826 9199
rect 14462 8833 14826 8834
rect 14462 8807 14799 8833
rect 14825 8807 14826 8833
rect 14462 8806 14826 8807
rect 14462 8441 14490 8806
rect 14798 8801 14826 8806
rect 15134 8834 15162 9310
rect 15750 9281 15778 9590
rect 15862 9618 15890 11046
rect 15862 9585 15890 9590
rect 16254 9617 16282 9623
rect 16254 9591 16255 9617
rect 16281 9591 16282 9617
rect 15750 9255 15751 9281
rect 15777 9255 15778 9281
rect 15750 9225 15778 9255
rect 15750 9199 15751 9225
rect 15777 9199 15778 9225
rect 15246 8834 15274 8839
rect 15470 8834 15498 8839
rect 15134 8833 15498 8834
rect 15134 8807 15247 8833
rect 15273 8807 15471 8833
rect 15497 8807 15498 8833
rect 15134 8806 15498 8807
rect 14573 8638 15035 8643
rect 14573 8637 14582 8638
rect 14573 8611 14574 8637
rect 14573 8610 14582 8611
rect 14610 8610 14634 8638
rect 14662 8610 14686 8638
rect 14714 8637 14738 8638
rect 14766 8637 14790 8638
rect 14724 8611 14738 8637
rect 14786 8611 14790 8637
rect 14714 8610 14738 8611
rect 14766 8610 14790 8611
rect 14818 8637 14842 8638
rect 14870 8637 14894 8638
rect 14818 8611 14822 8637
rect 14870 8611 14884 8637
rect 14818 8610 14842 8611
rect 14870 8610 14894 8611
rect 14922 8610 14946 8638
rect 14974 8610 14998 8638
rect 15026 8637 15035 8638
rect 15034 8611 15035 8637
rect 15026 8610 15035 8611
rect 14573 8605 15035 8610
rect 14462 8415 14463 8441
rect 14489 8415 14490 8441
rect 14462 8409 14490 8415
rect 14966 8442 14994 8447
rect 14966 8050 14994 8414
rect 15022 8442 15050 8447
rect 15134 8442 15162 8806
rect 15246 8801 15274 8806
rect 15470 8801 15498 8806
rect 15022 8441 15162 8442
rect 15022 8415 15023 8441
rect 15049 8415 15135 8441
rect 15161 8415 15162 8441
rect 15022 8414 15162 8415
rect 15022 8409 15050 8414
rect 15134 8409 15162 8414
rect 14966 8049 15106 8050
rect 14966 8023 14967 8049
rect 14993 8023 15106 8049
rect 14966 8022 15106 8023
rect 14966 8017 14994 8022
rect 14573 7854 15035 7859
rect 14573 7853 14582 7854
rect 14573 7827 14574 7853
rect 14573 7826 14582 7827
rect 14610 7826 14634 7854
rect 14662 7826 14686 7854
rect 14714 7853 14738 7854
rect 14766 7853 14790 7854
rect 14724 7827 14738 7853
rect 14786 7827 14790 7853
rect 14714 7826 14738 7827
rect 14766 7826 14790 7827
rect 14818 7853 14842 7854
rect 14870 7853 14894 7854
rect 14818 7827 14822 7853
rect 14870 7827 14884 7853
rect 14818 7826 14842 7827
rect 14870 7826 14894 7827
rect 14922 7826 14946 7854
rect 14974 7826 14998 7854
rect 15026 7853 15035 7854
rect 15034 7827 15035 7853
rect 15026 7826 15035 7827
rect 14573 7821 15035 7826
rect 14406 7631 14407 7657
rect 14433 7631 14434 7657
rect 13454 7219 13482 7238
rect 13118 6930 13146 6935
rect 13118 6873 13146 6902
rect 14406 6930 14434 7631
rect 15078 7265 15106 8022
rect 15750 8049 15778 9199
rect 15750 8023 15751 8049
rect 15777 8023 15778 8049
rect 15750 7993 15778 8023
rect 16254 8833 16282 9591
rect 16254 8807 16255 8833
rect 16281 8807 16282 8833
rect 16254 8442 16282 8807
rect 16254 8049 16282 8414
rect 16254 8023 16255 8049
rect 16281 8023 16282 8049
rect 16254 8017 16282 8023
rect 15750 7967 15751 7993
rect 15777 7967 15778 7993
rect 15750 7961 15778 7967
rect 15078 7239 15079 7265
rect 15105 7239 15106 7265
rect 15078 7233 15106 7239
rect 15246 7713 15274 7719
rect 15246 7687 15247 7713
rect 15273 7687 15274 7713
rect 15246 7657 15274 7687
rect 15246 7631 15247 7657
rect 15273 7631 15274 7657
rect 15246 7266 15274 7631
rect 15470 7266 15498 7271
rect 15246 7265 15498 7266
rect 15246 7239 15247 7265
rect 15273 7239 15471 7265
rect 15497 7239 15498 7265
rect 15246 7238 15498 7239
rect 14573 7070 15035 7075
rect 14573 7069 14582 7070
rect 14573 7043 14574 7069
rect 14573 7042 14582 7043
rect 14610 7042 14634 7070
rect 14662 7042 14686 7070
rect 14714 7069 14738 7070
rect 14766 7069 14790 7070
rect 14724 7043 14738 7069
rect 14786 7043 14790 7069
rect 14714 7042 14738 7043
rect 14766 7042 14790 7043
rect 14818 7069 14842 7070
rect 14870 7069 14894 7070
rect 14818 7043 14822 7069
rect 14870 7043 14884 7069
rect 14818 7042 14842 7043
rect 14870 7042 14894 7043
rect 14922 7042 14946 7070
rect 14974 7042 14998 7070
rect 15026 7069 15035 7070
rect 15034 7043 15035 7069
rect 15026 7042 15035 7043
rect 14573 7037 15035 7042
rect 13118 6847 13119 6873
rect 13145 6847 13146 6873
rect 13118 6481 13146 6847
rect 13398 6874 13426 6879
rect 13510 6874 13538 6879
rect 13398 6873 13510 6874
rect 13398 6847 13399 6873
rect 13425 6847 13510 6873
rect 13398 6846 13510 6847
rect 13398 6841 13426 6846
rect 13118 6455 13119 6481
rect 13145 6455 13146 6481
rect 13118 6089 13146 6455
rect 13454 6482 13482 6846
rect 13510 6808 13538 6846
rect 14406 6873 14434 6902
rect 15246 6929 15274 7238
rect 15470 7233 15498 7238
rect 15246 6903 15247 6929
rect 15273 6903 15274 6929
rect 14406 6847 14407 6873
rect 14433 6847 14434 6873
rect 14406 6841 14434 6847
rect 15134 6874 15162 6879
rect 15134 6827 15162 6846
rect 15246 6874 15274 6903
rect 15246 6841 15274 6846
rect 13622 6482 13650 6487
rect 13454 6481 13650 6482
rect 13454 6455 13455 6481
rect 13481 6455 13623 6481
rect 13649 6455 13650 6481
rect 13454 6454 13650 6455
rect 13118 6063 13119 6089
rect 13145 6063 13146 6089
rect 13118 5642 13146 6063
rect 13118 5305 13146 5614
rect 13118 5279 13119 5305
rect 13145 5279 13146 5305
rect 13118 5273 13146 5279
rect 13286 6090 13314 6095
rect 13454 6090 13482 6454
rect 13622 6449 13650 6454
rect 15750 6482 15778 6487
rect 14573 6286 15035 6291
rect 14573 6285 14582 6286
rect 14573 6259 14574 6285
rect 14573 6258 14582 6259
rect 14610 6258 14634 6286
rect 14662 6258 14686 6286
rect 14714 6285 14738 6286
rect 14766 6285 14790 6286
rect 14724 6259 14738 6285
rect 14786 6259 14790 6285
rect 14714 6258 14738 6259
rect 14766 6258 14790 6259
rect 14818 6285 14842 6286
rect 14870 6285 14894 6286
rect 14818 6259 14822 6285
rect 14870 6259 14884 6285
rect 14818 6258 14842 6259
rect 14870 6258 14894 6259
rect 14922 6258 14946 6286
rect 14974 6258 14998 6286
rect 15026 6285 15035 6286
rect 15034 6259 15035 6285
rect 15026 6258 15035 6259
rect 14573 6253 15035 6258
rect 13510 6090 13538 6095
rect 13286 6089 13538 6090
rect 13286 6063 13287 6089
rect 13313 6063 13511 6089
rect 13537 6063 13538 6089
rect 13286 6062 13538 6063
rect 13286 5306 13314 6062
rect 13510 6057 13538 6062
rect 15526 6090 15554 6095
rect 15750 6090 15778 6454
rect 15526 6089 15778 6090
rect 15526 6063 15527 6089
rect 15553 6063 15778 6089
rect 15526 6062 15778 6063
rect 15526 6057 15554 6062
rect 15750 5697 15778 6062
rect 15750 5671 15751 5697
rect 15777 5671 15778 5697
rect 14573 5502 15035 5507
rect 14573 5501 14582 5502
rect 14573 5475 14574 5501
rect 14573 5474 14582 5475
rect 14610 5474 14634 5502
rect 14662 5474 14686 5502
rect 14714 5501 14738 5502
rect 14766 5501 14790 5502
rect 14724 5475 14738 5501
rect 14786 5475 14790 5501
rect 14714 5474 14738 5475
rect 14766 5474 14790 5475
rect 14818 5501 14842 5502
rect 14870 5501 14894 5502
rect 14818 5475 14822 5501
rect 14870 5475 14884 5501
rect 14818 5474 14842 5475
rect 14870 5474 14894 5475
rect 14922 5474 14946 5502
rect 14974 5474 14998 5502
rect 15026 5501 15035 5502
rect 15034 5475 15035 5501
rect 15026 5474 15035 5475
rect 14573 5469 15035 5474
rect 13286 5259 13314 5278
rect 13510 5306 13538 5311
rect 13510 5259 13538 5278
rect 15358 5305 15386 5311
rect 15358 5279 15359 5305
rect 15385 5279 15386 5305
rect 14573 4718 15035 4723
rect 14573 4717 14582 4718
rect 14573 4691 14574 4717
rect 14573 4690 14582 4691
rect 14610 4690 14634 4718
rect 14662 4690 14686 4718
rect 14714 4717 14738 4718
rect 14766 4717 14790 4718
rect 14724 4691 14738 4717
rect 14786 4691 14790 4717
rect 14714 4690 14738 4691
rect 14766 4690 14790 4691
rect 14818 4717 14842 4718
rect 14870 4717 14894 4718
rect 14818 4691 14822 4717
rect 14870 4691 14884 4717
rect 14818 4690 14842 4691
rect 14870 4690 14894 4691
rect 14922 4690 14946 4718
rect 14974 4690 14998 4718
rect 15026 4717 15035 4718
rect 15034 4691 15035 4717
rect 15026 4690 15035 4691
rect 14573 4685 15035 4690
rect 14742 4577 14770 4583
rect 14742 4551 14743 4577
rect 14769 4551 14770 4577
rect 14070 4521 14098 4527
rect 14070 4495 14071 4521
rect 14097 4495 14098 4521
rect 12950 4130 12978 4135
rect 12950 4083 12978 4102
rect 13230 4130 13258 4135
rect 13230 3738 13258 4102
rect 13230 3345 13258 3710
rect 13790 3738 13818 3743
rect 13790 3691 13818 3710
rect 14070 3738 14098 4495
rect 14742 4521 14770 4551
rect 14742 4495 14743 4521
rect 14769 4495 14770 4521
rect 14742 4214 14770 4495
rect 13230 3319 13231 3345
rect 13257 3319 13258 3345
rect 13230 3313 13258 3319
rect 14070 3402 14098 3710
rect 13174 2954 13202 2959
rect 13174 2561 13202 2926
rect 14070 2953 14098 3374
rect 14406 4186 14770 4214
rect 15358 4521 15386 5279
rect 15358 4495 15359 4521
rect 15385 4495 15386 4521
rect 15358 4214 15386 4495
rect 15750 4913 15778 5671
rect 15750 4887 15751 4913
rect 15777 4887 15778 4913
rect 15358 4186 15554 4214
rect 14406 4129 14434 4186
rect 14406 4103 14407 4129
rect 14433 4103 14434 4129
rect 14406 4073 14434 4103
rect 14406 4047 14407 4073
rect 14433 4047 14434 4073
rect 14406 3345 14434 4047
rect 15526 4130 15554 4186
rect 15750 4130 15778 4887
rect 16366 4634 16394 13902
rect 16534 13538 16562 14295
rect 16534 13491 16562 13510
rect 16534 12753 16562 12759
rect 16534 12727 16535 12753
rect 16561 12727 16562 12753
rect 16534 11969 16562 12727
rect 16534 11943 16535 11969
rect 16561 11943 16562 11969
rect 16534 11746 16562 11943
rect 16534 11185 16562 11718
rect 16534 11159 16535 11185
rect 16561 11159 16562 11185
rect 16534 10794 16562 11159
rect 16814 12361 16842 12367
rect 16814 12335 16815 12361
rect 16841 12335 16842 12361
rect 16814 11577 16842 12335
rect 16814 11551 16815 11577
rect 16841 11551 16842 11577
rect 16814 10794 16842 11551
rect 16534 10793 16842 10794
rect 16534 10767 16815 10793
rect 16841 10767 16842 10793
rect 16534 10766 16842 10767
rect 16534 10401 16562 10766
rect 16814 10761 16842 10766
rect 16534 10375 16535 10401
rect 16561 10375 16562 10401
rect 16534 10369 16562 10375
rect 16814 10402 16842 10407
rect 16814 10094 16842 10374
rect 16758 10066 16842 10094
rect 16870 10094 16898 19614
rect 17318 19530 17346 19614
rect 17472 19600 17528 20000
rect 21854 19614 22330 19642
rect 17486 19530 17514 19600
rect 17318 19502 17514 19530
rect 17073 18438 17535 18443
rect 17073 18437 17082 18438
rect 17073 18411 17074 18437
rect 17073 18410 17082 18411
rect 17110 18410 17134 18438
rect 17162 18410 17186 18438
rect 17214 18437 17238 18438
rect 17266 18437 17290 18438
rect 17224 18411 17238 18437
rect 17286 18411 17290 18437
rect 17214 18410 17238 18411
rect 17266 18410 17290 18411
rect 17318 18437 17342 18438
rect 17370 18437 17394 18438
rect 17318 18411 17322 18437
rect 17370 18411 17384 18437
rect 17318 18410 17342 18411
rect 17370 18410 17394 18411
rect 17422 18410 17446 18438
rect 17474 18410 17498 18438
rect 17526 18437 17535 18438
rect 17534 18411 17535 18437
rect 17526 18410 17535 18411
rect 17073 18405 17535 18410
rect 19573 18046 20035 18051
rect 19573 18045 19582 18046
rect 19573 18019 19574 18045
rect 19573 18018 19582 18019
rect 19610 18018 19634 18046
rect 19662 18018 19686 18046
rect 19714 18045 19738 18046
rect 19766 18045 19790 18046
rect 19724 18019 19738 18045
rect 19786 18019 19790 18045
rect 19714 18018 19738 18019
rect 19766 18018 19790 18019
rect 19818 18045 19842 18046
rect 19870 18045 19894 18046
rect 19818 18019 19822 18045
rect 19870 18019 19884 18045
rect 19818 18018 19842 18019
rect 19870 18018 19894 18019
rect 19922 18018 19946 18046
rect 19974 18018 19998 18046
rect 20026 18045 20035 18046
rect 20034 18019 20035 18045
rect 20026 18018 20035 18019
rect 19573 18013 20035 18018
rect 17073 17654 17535 17659
rect 17073 17653 17082 17654
rect 17073 17627 17074 17653
rect 17073 17626 17082 17627
rect 17110 17626 17134 17654
rect 17162 17626 17186 17654
rect 17214 17653 17238 17654
rect 17266 17653 17290 17654
rect 17224 17627 17238 17653
rect 17286 17627 17290 17653
rect 17214 17626 17238 17627
rect 17266 17626 17290 17627
rect 17318 17653 17342 17654
rect 17370 17653 17394 17654
rect 17318 17627 17322 17653
rect 17370 17627 17384 17653
rect 17318 17626 17342 17627
rect 17370 17626 17394 17627
rect 17422 17626 17446 17654
rect 17474 17626 17498 17654
rect 17526 17653 17535 17654
rect 17534 17627 17535 17653
rect 17526 17626 17535 17627
rect 17073 17621 17535 17626
rect 19573 17262 20035 17267
rect 19573 17261 19582 17262
rect 19573 17235 19574 17261
rect 19573 17234 19582 17235
rect 19610 17234 19634 17262
rect 19662 17234 19686 17262
rect 19714 17261 19738 17262
rect 19766 17261 19790 17262
rect 19724 17235 19738 17261
rect 19786 17235 19790 17261
rect 19714 17234 19738 17235
rect 19766 17234 19790 17235
rect 19818 17261 19842 17262
rect 19870 17261 19894 17262
rect 19818 17235 19822 17261
rect 19870 17235 19884 17261
rect 19818 17234 19842 17235
rect 19870 17234 19894 17235
rect 19922 17234 19946 17262
rect 19974 17234 19998 17262
rect 20026 17261 20035 17262
rect 20034 17235 20035 17261
rect 20026 17234 20035 17235
rect 19573 17229 20035 17234
rect 17073 16870 17535 16875
rect 17073 16869 17082 16870
rect 17073 16843 17074 16869
rect 17073 16842 17082 16843
rect 17110 16842 17134 16870
rect 17162 16842 17186 16870
rect 17214 16869 17238 16870
rect 17266 16869 17290 16870
rect 17224 16843 17238 16869
rect 17286 16843 17290 16869
rect 17214 16842 17238 16843
rect 17266 16842 17290 16843
rect 17318 16869 17342 16870
rect 17370 16869 17394 16870
rect 17318 16843 17322 16869
rect 17370 16843 17384 16869
rect 17318 16842 17342 16843
rect 17370 16842 17394 16843
rect 17422 16842 17446 16870
rect 17474 16842 17498 16870
rect 17526 16869 17535 16870
rect 17534 16843 17535 16869
rect 17526 16842 17535 16843
rect 17073 16837 17535 16842
rect 19573 16478 20035 16483
rect 19573 16477 19582 16478
rect 19573 16451 19574 16477
rect 19573 16450 19582 16451
rect 19610 16450 19634 16478
rect 19662 16450 19686 16478
rect 19714 16477 19738 16478
rect 19766 16477 19790 16478
rect 19724 16451 19738 16477
rect 19786 16451 19790 16477
rect 19714 16450 19738 16451
rect 19766 16450 19790 16451
rect 19818 16477 19842 16478
rect 19870 16477 19894 16478
rect 19818 16451 19822 16477
rect 19870 16451 19884 16477
rect 19818 16450 19842 16451
rect 19870 16450 19894 16451
rect 19922 16450 19946 16478
rect 19974 16450 19998 16478
rect 20026 16477 20035 16478
rect 20034 16451 20035 16477
rect 20026 16450 20035 16451
rect 19573 16445 20035 16450
rect 17073 16086 17535 16091
rect 17073 16085 17082 16086
rect 17073 16059 17074 16085
rect 17073 16058 17082 16059
rect 17110 16058 17134 16086
rect 17162 16058 17186 16086
rect 17214 16085 17238 16086
rect 17266 16085 17290 16086
rect 17224 16059 17238 16085
rect 17286 16059 17290 16085
rect 17214 16058 17238 16059
rect 17266 16058 17290 16059
rect 17318 16085 17342 16086
rect 17370 16085 17394 16086
rect 17318 16059 17322 16085
rect 17370 16059 17384 16085
rect 17318 16058 17342 16059
rect 17370 16058 17394 16059
rect 17422 16058 17446 16086
rect 17474 16058 17498 16086
rect 17526 16085 17535 16086
rect 17534 16059 17535 16085
rect 17526 16058 17535 16059
rect 17073 16053 17535 16058
rect 16926 15946 16954 15951
rect 16926 15889 16954 15918
rect 16926 15863 16927 15889
rect 16953 15863 16954 15889
rect 16926 15857 16954 15863
rect 20286 15890 20314 15895
rect 19573 15694 20035 15699
rect 19573 15693 19582 15694
rect 19573 15667 19574 15693
rect 19573 15666 19582 15667
rect 19610 15666 19634 15694
rect 19662 15666 19686 15694
rect 19714 15693 19738 15694
rect 19766 15693 19790 15694
rect 19724 15667 19738 15693
rect 19786 15667 19790 15693
rect 19714 15666 19738 15667
rect 19766 15666 19790 15667
rect 19818 15693 19842 15694
rect 19870 15693 19894 15694
rect 19818 15667 19822 15693
rect 19870 15667 19884 15693
rect 19818 15666 19842 15667
rect 19870 15666 19894 15667
rect 19922 15666 19946 15694
rect 19974 15666 19998 15694
rect 20026 15693 20035 15694
rect 20034 15667 20035 15693
rect 20026 15666 20035 15667
rect 19573 15661 20035 15666
rect 17073 15302 17535 15307
rect 17073 15301 17082 15302
rect 17073 15275 17074 15301
rect 17073 15274 17082 15275
rect 17110 15274 17134 15302
rect 17162 15274 17186 15302
rect 17214 15301 17238 15302
rect 17266 15301 17290 15302
rect 17224 15275 17238 15301
rect 17286 15275 17290 15301
rect 17214 15274 17238 15275
rect 17266 15274 17290 15275
rect 17318 15301 17342 15302
rect 17370 15301 17394 15302
rect 17318 15275 17322 15301
rect 17370 15275 17384 15301
rect 17318 15274 17342 15275
rect 17370 15274 17394 15275
rect 17422 15274 17446 15302
rect 17474 15274 17498 15302
rect 17526 15301 17535 15302
rect 17534 15275 17535 15301
rect 17526 15274 17535 15275
rect 17073 15269 17535 15274
rect 17430 15105 17458 15111
rect 17430 15079 17431 15105
rect 17457 15079 17458 15105
rect 17430 15049 17458 15079
rect 17430 15023 17431 15049
rect 17457 15023 17458 15049
rect 17430 14770 17458 15023
rect 18774 15105 18802 15111
rect 18774 15079 18775 15105
rect 18801 15079 18802 15105
rect 17766 14770 17794 14775
rect 17430 14769 17794 14770
rect 17430 14743 17767 14769
rect 17793 14743 17794 14769
rect 17430 14742 17794 14743
rect 17094 14714 17122 14719
rect 17094 14667 17122 14686
rect 17766 14713 17794 14742
rect 17766 14687 17767 14713
rect 17793 14687 17794 14713
rect 17073 14518 17535 14523
rect 17073 14517 17082 14518
rect 17073 14491 17074 14517
rect 17073 14490 17082 14491
rect 17110 14490 17134 14518
rect 17162 14490 17186 14518
rect 17214 14517 17238 14518
rect 17266 14517 17290 14518
rect 17224 14491 17238 14517
rect 17286 14491 17290 14517
rect 17214 14490 17238 14491
rect 17266 14490 17290 14491
rect 17318 14517 17342 14518
rect 17370 14517 17394 14518
rect 17318 14491 17322 14517
rect 17370 14491 17384 14517
rect 17318 14490 17342 14491
rect 17370 14490 17394 14491
rect 17422 14490 17446 14518
rect 17474 14490 17498 14518
rect 17526 14517 17535 14518
rect 17534 14491 17535 14517
rect 17526 14490 17535 14491
rect 17073 14485 17535 14490
rect 17430 14321 17458 14327
rect 17430 14295 17431 14321
rect 17457 14295 17458 14321
rect 17430 14266 17458 14295
rect 17430 14219 17458 14238
rect 17766 14266 17794 14687
rect 18270 14713 18298 14719
rect 18270 14687 18271 14713
rect 18297 14687 18298 14713
rect 18270 14658 18298 14687
rect 18270 14625 18298 14630
rect 18438 14714 18466 14719
rect 17766 13985 17794 14238
rect 17766 13959 17767 13985
rect 17793 13959 17794 13985
rect 16982 13929 17010 13935
rect 16982 13903 16983 13929
rect 17009 13903 17010 13929
rect 16982 13538 17010 13903
rect 17766 13929 17794 13959
rect 17766 13903 17767 13929
rect 17793 13903 17794 13929
rect 17073 13734 17535 13739
rect 17073 13733 17082 13734
rect 17073 13707 17074 13733
rect 17073 13706 17082 13707
rect 17110 13706 17134 13734
rect 17162 13706 17186 13734
rect 17214 13733 17238 13734
rect 17266 13733 17290 13734
rect 17224 13707 17238 13733
rect 17286 13707 17290 13733
rect 17214 13706 17238 13707
rect 17266 13706 17290 13707
rect 17318 13733 17342 13734
rect 17370 13733 17394 13734
rect 17318 13707 17322 13733
rect 17370 13707 17384 13733
rect 17318 13706 17342 13707
rect 17370 13706 17394 13707
rect 17422 13706 17446 13734
rect 17474 13706 17498 13734
rect 17526 13733 17535 13734
rect 17534 13707 17535 13733
rect 17526 13706 17535 13707
rect 17073 13701 17535 13706
rect 16982 13146 17010 13510
rect 17430 13537 17458 13543
rect 17430 13511 17431 13537
rect 17457 13511 17458 13537
rect 17430 13482 17458 13511
rect 16982 13113 17010 13118
rect 17094 13146 17122 13151
rect 17430 13146 17458 13454
rect 17766 13201 17794 13903
rect 18438 13930 18466 14686
rect 18718 14713 18746 14719
rect 18718 14687 18719 14713
rect 18745 14687 18746 14713
rect 18718 14266 18746 14687
rect 18774 14658 18802 15079
rect 19334 15106 19362 15111
rect 19446 15106 19474 15111
rect 19334 15105 19474 15106
rect 19334 15079 19335 15105
rect 19361 15079 19447 15105
rect 19473 15079 19474 15105
rect 19334 15078 19474 15079
rect 19334 15073 19362 15078
rect 18774 14322 18802 14630
rect 18774 14256 18802 14294
rect 18942 14713 18970 14719
rect 18942 14687 18943 14713
rect 18969 14687 18970 14713
rect 18942 14266 18970 14687
rect 19334 14322 19362 14327
rect 19446 14322 19474 15078
rect 19573 14910 20035 14915
rect 19573 14909 19582 14910
rect 19573 14883 19574 14909
rect 19573 14882 19582 14883
rect 19610 14882 19634 14910
rect 19662 14882 19686 14910
rect 19714 14909 19738 14910
rect 19766 14909 19790 14910
rect 19724 14883 19738 14909
rect 19786 14883 19790 14909
rect 19714 14882 19738 14883
rect 19766 14882 19790 14883
rect 19818 14909 19842 14910
rect 19870 14909 19894 14910
rect 19818 14883 19822 14909
rect 19870 14883 19884 14909
rect 19818 14882 19842 14883
rect 19870 14882 19894 14883
rect 19922 14882 19946 14910
rect 19974 14882 19998 14910
rect 20026 14909 20035 14910
rect 20034 14883 20035 14909
rect 20026 14882 20035 14883
rect 19573 14877 20035 14882
rect 19334 14321 19474 14322
rect 19334 14295 19335 14321
rect 19361 14295 19447 14321
rect 19473 14295 19474 14321
rect 19334 14294 19474 14295
rect 19334 14289 19362 14294
rect 18718 14233 18746 14238
rect 18942 14233 18970 14238
rect 19446 13985 19474 14294
rect 20230 14322 20258 14327
rect 19573 14126 20035 14131
rect 19573 14125 19582 14126
rect 19573 14099 19574 14125
rect 19573 14098 19582 14099
rect 19610 14098 19634 14126
rect 19662 14098 19686 14126
rect 19714 14125 19738 14126
rect 19766 14125 19790 14126
rect 19724 14099 19738 14125
rect 19786 14099 19790 14125
rect 19714 14098 19738 14099
rect 19766 14098 19790 14099
rect 19818 14125 19842 14126
rect 19870 14125 19894 14126
rect 19818 14099 19822 14125
rect 19870 14099 19884 14125
rect 19818 14098 19842 14099
rect 19870 14098 19894 14099
rect 19922 14098 19946 14126
rect 19974 14098 19998 14126
rect 20026 14125 20035 14126
rect 20034 14099 20035 14125
rect 20026 14098 20035 14099
rect 19573 14093 20035 14098
rect 19446 13959 19447 13985
rect 19473 13959 19474 13985
rect 18550 13930 18578 13935
rect 18438 13929 18578 13930
rect 18438 13903 18551 13929
rect 18577 13903 18578 13929
rect 18438 13902 18578 13903
rect 18550 13538 18578 13902
rect 19446 13929 19474 13959
rect 19446 13903 19447 13929
rect 19473 13903 19474 13929
rect 18550 13505 18578 13510
rect 19054 13538 19082 13543
rect 19054 13491 19082 13510
rect 19334 13538 19362 13543
rect 19446 13538 19474 13903
rect 19334 13537 19474 13538
rect 19334 13511 19335 13537
rect 19361 13511 19447 13537
rect 19473 13511 19474 13537
rect 19334 13510 19474 13511
rect 19334 13505 19362 13510
rect 17766 13175 17767 13201
rect 17793 13175 17794 13201
rect 17598 13146 17626 13151
rect 17766 13146 17794 13175
rect 19446 13201 19474 13510
rect 20230 13537 20258 14294
rect 20230 13511 20231 13537
rect 20257 13511 20258 13537
rect 20230 13505 20258 13511
rect 19573 13342 20035 13347
rect 19573 13341 19582 13342
rect 19573 13315 19574 13341
rect 19573 13314 19582 13315
rect 19610 13314 19634 13342
rect 19662 13314 19686 13342
rect 19714 13341 19738 13342
rect 19766 13341 19790 13342
rect 19724 13315 19738 13341
rect 19786 13315 19790 13341
rect 19714 13314 19738 13315
rect 19766 13314 19790 13315
rect 19818 13341 19842 13342
rect 19870 13341 19894 13342
rect 19818 13315 19822 13341
rect 19870 13315 19884 13341
rect 19818 13314 19842 13315
rect 19870 13314 19894 13315
rect 19922 13314 19946 13342
rect 19974 13314 19998 13342
rect 20026 13341 20035 13342
rect 20034 13315 20035 13341
rect 20026 13314 20035 13315
rect 19573 13309 20035 13314
rect 19446 13175 19447 13201
rect 19473 13175 19474 13201
rect 17430 13145 17794 13146
rect 17430 13119 17599 13145
rect 17625 13119 17794 13145
rect 17430 13118 17794 13119
rect 18550 13146 18578 13151
rect 17094 13099 17122 13118
rect 17073 12950 17535 12955
rect 17073 12949 17082 12950
rect 17073 12923 17074 12949
rect 17073 12922 17082 12923
rect 17110 12922 17134 12950
rect 17162 12922 17186 12950
rect 17214 12949 17238 12950
rect 17266 12949 17290 12950
rect 17224 12923 17238 12949
rect 17286 12923 17290 12949
rect 17214 12922 17238 12923
rect 17266 12922 17290 12923
rect 17318 12949 17342 12950
rect 17370 12949 17394 12950
rect 17318 12923 17322 12949
rect 17370 12923 17384 12949
rect 17318 12922 17342 12923
rect 17370 12922 17394 12923
rect 17422 12922 17446 12950
rect 17474 12922 17498 12950
rect 17526 12949 17535 12950
rect 17534 12923 17535 12949
rect 17526 12922 17535 12923
rect 17073 12917 17535 12922
rect 17430 12753 17458 12759
rect 17430 12727 17431 12753
rect 17457 12727 17458 12753
rect 17430 12697 17458 12727
rect 17430 12671 17431 12697
rect 17457 12671 17458 12697
rect 17430 12642 17458 12671
rect 17598 12642 17626 13118
rect 17430 12614 17626 12642
rect 17073 12166 17535 12171
rect 17073 12165 17082 12166
rect 17073 12139 17074 12165
rect 17073 12138 17082 12139
rect 17110 12138 17134 12166
rect 17162 12138 17186 12166
rect 17214 12165 17238 12166
rect 17266 12165 17290 12166
rect 17224 12139 17238 12165
rect 17286 12139 17290 12165
rect 17214 12138 17238 12139
rect 17266 12138 17290 12139
rect 17318 12165 17342 12166
rect 17370 12165 17394 12166
rect 17318 12139 17322 12165
rect 17370 12139 17384 12165
rect 17318 12138 17342 12139
rect 17370 12138 17394 12139
rect 17422 12138 17446 12166
rect 17474 12138 17498 12166
rect 17526 12165 17535 12166
rect 17534 12139 17535 12165
rect 17526 12138 17535 12139
rect 17073 12133 17535 12138
rect 17430 11970 17458 11975
rect 17430 11913 17458 11942
rect 17598 11970 17626 12614
rect 18550 12642 18578 13118
rect 19446 13145 19474 13175
rect 19446 13119 19447 13145
rect 19473 13119 19474 13145
rect 17598 11937 17626 11942
rect 17990 12417 18018 12423
rect 17990 12391 17991 12417
rect 18017 12391 18018 12417
rect 17990 12361 18018 12391
rect 17990 12335 17991 12361
rect 18017 12335 18018 12361
rect 17990 11970 18018 12335
rect 18550 12361 18578 12614
rect 18550 12335 18551 12361
rect 18577 12335 18578 12361
rect 18550 12329 18578 12335
rect 19054 12753 19082 12759
rect 19054 12727 19055 12753
rect 19081 12727 19082 12753
rect 19054 12642 19082 12727
rect 17430 11887 17431 11913
rect 17457 11887 17458 11913
rect 17430 11881 17458 11887
rect 17990 11633 18018 11942
rect 17990 11607 17991 11633
rect 18017 11607 18018 11633
rect 17990 11577 18018 11607
rect 19054 11969 19082 12614
rect 19054 11943 19055 11969
rect 19081 11943 19082 11969
rect 17990 11551 17991 11577
rect 18017 11551 18018 11577
rect 17073 11382 17535 11387
rect 17073 11381 17082 11382
rect 17073 11355 17074 11381
rect 17073 11354 17082 11355
rect 17110 11354 17134 11382
rect 17162 11354 17186 11382
rect 17214 11381 17238 11382
rect 17266 11381 17290 11382
rect 17224 11355 17238 11381
rect 17286 11355 17290 11381
rect 17214 11354 17238 11355
rect 17266 11354 17290 11355
rect 17318 11381 17342 11382
rect 17370 11381 17394 11382
rect 17318 11355 17322 11381
rect 17370 11355 17384 11381
rect 17318 11354 17342 11355
rect 17370 11354 17394 11355
rect 17422 11354 17446 11382
rect 17474 11354 17498 11382
rect 17526 11381 17535 11382
rect 17534 11355 17535 11381
rect 17526 11354 17535 11355
rect 17073 11349 17535 11354
rect 17262 11185 17290 11191
rect 17262 11159 17263 11185
rect 17289 11159 17290 11185
rect 17262 11129 17290 11159
rect 17262 11103 17263 11129
rect 17289 11103 17290 11129
rect 16926 10794 16954 10799
rect 16926 10402 16954 10766
rect 17262 10794 17290 11103
rect 17262 10747 17290 10766
rect 17486 10794 17514 10799
rect 17486 10747 17514 10766
rect 17073 10598 17535 10603
rect 17073 10597 17082 10598
rect 17073 10571 17074 10597
rect 17073 10570 17082 10571
rect 17110 10570 17134 10598
rect 17162 10570 17186 10598
rect 17214 10597 17238 10598
rect 17266 10597 17290 10598
rect 17224 10571 17238 10597
rect 17286 10571 17290 10597
rect 17214 10570 17238 10571
rect 17266 10570 17290 10571
rect 17318 10597 17342 10598
rect 17370 10597 17394 10598
rect 17318 10571 17322 10597
rect 17370 10571 17384 10597
rect 17318 10570 17342 10571
rect 17370 10570 17394 10571
rect 17422 10570 17446 10598
rect 17474 10570 17498 10598
rect 17526 10597 17535 10598
rect 17534 10571 17535 10597
rect 17526 10570 17535 10571
rect 17073 10565 17535 10570
rect 16926 10355 16954 10374
rect 16870 10066 17010 10094
rect 16758 10033 16786 10038
rect 16814 10009 16842 10015
rect 16814 9983 16815 10009
rect 16841 9983 16842 10009
rect 16814 9730 16842 9983
rect 16758 9702 16842 9730
rect 16758 9226 16786 9702
rect 16814 9618 16842 9623
rect 16926 9618 16954 9623
rect 16842 9617 16954 9618
rect 16842 9591 16927 9617
rect 16953 9591 16954 9617
rect 16842 9590 16954 9591
rect 16814 9571 16842 9590
rect 16814 9226 16842 9231
rect 16758 9225 16842 9226
rect 16758 9199 16815 9225
rect 16841 9199 16842 9225
rect 16758 9198 16842 9199
rect 16758 8442 16786 9198
rect 16814 9193 16842 9198
rect 16814 8834 16842 8839
rect 16926 8834 16954 9590
rect 16814 8833 16954 8834
rect 16814 8807 16815 8833
rect 16841 8807 16927 8833
rect 16953 8807 16954 8833
rect 16814 8806 16954 8807
rect 16814 8801 16842 8806
rect 16814 8442 16842 8447
rect 16758 8414 16814 8442
rect 16814 8395 16842 8414
rect 16814 8050 16842 8055
rect 16926 8050 16954 8806
rect 16814 8049 16954 8050
rect 16814 8023 16815 8049
rect 16841 8023 16927 8049
rect 16953 8023 16954 8049
rect 16814 8022 16954 8023
rect 16814 8017 16842 8022
rect 16926 8017 16954 8022
rect 16758 6481 16786 6487
rect 16758 6455 16759 6481
rect 16785 6455 16786 6481
rect 16758 6425 16786 6455
rect 16758 6399 16759 6425
rect 16785 6399 16786 6425
rect 16366 4601 16394 4606
rect 16422 6145 16450 6151
rect 16422 6119 16423 6145
rect 16449 6119 16450 6145
rect 16422 6089 16450 6119
rect 16422 6063 16423 6089
rect 16449 6063 16450 6089
rect 16422 5361 16450 6063
rect 16422 5335 16423 5361
rect 16449 5335 16450 5361
rect 16422 5305 16450 5335
rect 16422 5279 16423 5305
rect 16449 5279 16450 5305
rect 16422 5194 16450 5279
rect 16422 4577 16450 5166
rect 16758 5697 16786 6399
rect 16758 5671 16759 5697
rect 16785 5671 16786 5697
rect 16758 5641 16786 5671
rect 16758 5615 16759 5641
rect 16785 5615 16786 5641
rect 16758 5194 16786 5615
rect 16758 4913 16786 5166
rect 16758 4887 16759 4913
rect 16785 4887 16786 4913
rect 16758 4857 16786 4887
rect 16758 4831 16759 4857
rect 16785 4831 16786 4857
rect 16758 4825 16786 4831
rect 16870 5586 16898 5591
rect 16422 4551 16423 4577
rect 16449 4551 16450 4577
rect 16422 4521 16450 4551
rect 16422 4495 16423 4521
rect 16449 4495 16450 4521
rect 16422 4214 16450 4495
rect 15526 4129 15778 4130
rect 15526 4103 15751 4129
rect 15777 4103 15778 4129
rect 15526 4102 15778 4103
rect 14573 3934 15035 3939
rect 14573 3933 14582 3934
rect 14573 3907 14574 3933
rect 14573 3906 14582 3907
rect 14610 3906 14634 3934
rect 14662 3906 14686 3934
rect 14714 3933 14738 3934
rect 14766 3933 14790 3934
rect 14724 3907 14738 3933
rect 14786 3907 14790 3933
rect 14714 3906 14738 3907
rect 14766 3906 14790 3907
rect 14818 3933 14842 3934
rect 14870 3933 14894 3934
rect 14818 3907 14822 3933
rect 14870 3907 14884 3933
rect 14818 3906 14842 3907
rect 14870 3906 14894 3907
rect 14922 3906 14946 3934
rect 14974 3906 14998 3934
rect 15026 3933 15035 3934
rect 15034 3907 15035 3933
rect 15026 3906 15035 3907
rect 14573 3901 15035 3906
rect 14966 3793 14994 3799
rect 14966 3767 14967 3793
rect 14993 3767 14994 3793
rect 14966 3738 14994 3767
rect 15246 3738 15274 3743
rect 14966 3737 15106 3738
rect 14966 3711 14967 3737
rect 14993 3711 15106 3737
rect 14966 3710 15106 3711
rect 14966 3705 14994 3710
rect 14406 3319 14407 3345
rect 14433 3319 14434 3345
rect 14406 3290 14434 3319
rect 14406 3243 14434 3262
rect 15078 3290 15106 3710
rect 14573 3150 15035 3155
rect 14573 3149 14582 3150
rect 14573 3123 14574 3149
rect 14573 3122 14582 3123
rect 14610 3122 14634 3150
rect 14662 3122 14686 3150
rect 14714 3149 14738 3150
rect 14766 3149 14790 3150
rect 14724 3123 14738 3149
rect 14786 3123 14790 3149
rect 14714 3122 14738 3123
rect 14766 3122 14790 3123
rect 14818 3149 14842 3150
rect 14870 3149 14894 3150
rect 14818 3123 14822 3149
rect 14870 3123 14884 3149
rect 14818 3122 14842 3123
rect 14870 3122 14894 3123
rect 14922 3122 14946 3150
rect 14974 3122 14998 3150
rect 15026 3149 15035 3150
rect 15034 3123 15035 3149
rect 15026 3122 15035 3123
rect 14573 3117 15035 3122
rect 14070 2927 14071 2953
rect 14097 2927 14098 2953
rect 14070 2921 14098 2927
rect 14406 3010 14434 3015
rect 13174 2535 13175 2561
rect 13201 2535 13202 2561
rect 13174 2505 13202 2535
rect 13174 2479 13175 2505
rect 13201 2479 13202 2505
rect 13174 2473 13202 2479
rect 13062 2226 13090 2231
rect 13062 1777 13090 2198
rect 13790 2226 13818 2231
rect 13790 2169 13818 2198
rect 13790 2143 13791 2169
rect 13817 2143 13818 2169
rect 13790 2114 13818 2143
rect 13790 2081 13818 2086
rect 14238 2170 14266 2175
rect 13062 1751 13063 1777
rect 13089 1751 13090 1777
rect 13062 1745 13090 1751
rect 13510 1777 13538 1783
rect 13510 1751 13511 1777
rect 13537 1751 13538 1777
rect 13510 1722 13538 1751
rect 13510 1689 13538 1694
rect 13734 1777 13762 1783
rect 13734 1751 13735 1777
rect 13761 1751 13762 1777
rect 13734 1722 13762 1751
rect 13734 1689 13762 1694
rect 14238 1722 14266 2142
rect 14238 1689 14266 1694
rect 13006 462 13202 490
rect 13006 378 13034 462
rect 13174 400 13202 462
rect 14406 400 14434 2982
rect 14966 3009 14994 3015
rect 14966 2983 14967 3009
rect 14993 2983 14994 3009
rect 14966 2954 14994 2983
rect 14966 2907 14994 2926
rect 15078 2954 15106 3262
rect 15078 2921 15106 2926
rect 15246 3402 15274 3710
rect 15526 3738 15554 4102
rect 15750 4097 15778 4102
rect 16254 4186 16450 4214
rect 16254 4129 16282 4186
rect 16254 4103 16255 4129
rect 16281 4103 16282 4129
rect 15526 3705 15554 3710
rect 15246 2953 15274 3374
rect 15750 3402 15778 3407
rect 15750 3345 15778 3374
rect 15750 3319 15751 3345
rect 15777 3319 15778 3345
rect 15246 2927 15247 2953
rect 15273 2927 15274 2953
rect 14573 2366 15035 2371
rect 14573 2365 14582 2366
rect 14573 2339 14574 2365
rect 14573 2338 14582 2339
rect 14610 2338 14634 2366
rect 14662 2338 14686 2366
rect 14714 2365 14738 2366
rect 14766 2365 14790 2366
rect 14724 2339 14738 2365
rect 14786 2339 14790 2365
rect 14714 2338 14738 2339
rect 14766 2338 14790 2339
rect 14818 2365 14842 2366
rect 14870 2365 14894 2366
rect 14818 2339 14822 2365
rect 14870 2339 14884 2365
rect 14818 2338 14842 2339
rect 14870 2338 14894 2339
rect 14922 2338 14946 2366
rect 14974 2338 14998 2366
rect 15026 2365 15035 2366
rect 15034 2339 15035 2365
rect 15026 2338 15035 2339
rect 14573 2333 15035 2338
rect 14462 2170 14490 2175
rect 14462 2123 14490 2142
rect 15246 2169 15274 2927
rect 15694 2954 15722 2959
rect 15246 2143 15247 2169
rect 15273 2143 15274 2169
rect 15246 1777 15274 2143
rect 15246 1751 15247 1777
rect 15273 1751 15274 1777
rect 15246 1745 15274 1751
rect 15526 2898 15554 2903
rect 14573 1582 15035 1587
rect 14573 1581 14582 1582
rect 14573 1555 14574 1581
rect 14573 1554 14582 1555
rect 14610 1554 14634 1582
rect 14662 1554 14686 1582
rect 14714 1581 14738 1582
rect 14766 1581 14790 1582
rect 14724 1555 14738 1581
rect 14786 1555 14790 1581
rect 14714 1554 14738 1555
rect 14766 1554 14790 1555
rect 14818 1581 14842 1582
rect 14870 1581 14894 1582
rect 14818 1555 14822 1581
rect 14870 1555 14884 1581
rect 14818 1554 14842 1555
rect 14870 1554 14894 1555
rect 14922 1554 14946 1582
rect 14974 1554 14998 1582
rect 15026 1581 15035 1582
rect 15034 1555 15035 1581
rect 15026 1554 15035 1555
rect 14573 1549 15035 1554
rect 15526 1498 15554 2870
rect 15694 2170 15722 2926
rect 15750 2561 15778 3319
rect 15750 2535 15751 2561
rect 15777 2535 15778 2561
rect 15750 2529 15778 2535
rect 15918 2170 15946 2175
rect 15694 2169 15946 2170
rect 15694 2143 15695 2169
rect 15721 2143 15919 2169
rect 15945 2143 15946 2169
rect 15694 2142 15946 2143
rect 15582 1778 15610 1783
rect 15582 1731 15610 1750
rect 15694 1778 15722 2142
rect 15918 2137 15946 2142
rect 16254 2170 16282 4103
rect 16310 4130 16338 4186
rect 16422 4130 16450 4135
rect 16310 4129 16450 4130
rect 16310 4103 16423 4129
rect 16449 4103 16450 4129
rect 16310 4102 16450 4103
rect 16422 4097 16450 4102
rect 16422 3793 16450 3799
rect 16422 3767 16423 3793
rect 16449 3767 16450 3793
rect 16422 3737 16450 3767
rect 16422 3711 16423 3737
rect 16449 3711 16450 3737
rect 16422 2954 16450 3711
rect 16422 2907 16450 2926
rect 16758 3345 16786 3351
rect 16758 3319 16759 3345
rect 16785 3319 16786 3345
rect 16758 3289 16786 3319
rect 16758 3263 16759 3289
rect 16785 3263 16786 3289
rect 16758 2954 16786 3263
rect 16758 2562 16786 2926
rect 16758 2505 16786 2534
rect 16758 2479 16759 2505
rect 16785 2479 16786 2505
rect 16758 2473 16786 2479
rect 16870 2618 16898 5558
rect 16982 4466 17010 10066
rect 17990 10065 18018 11551
rect 18550 11577 18578 11583
rect 18550 11551 18551 11577
rect 18577 11551 18578 11577
rect 18550 11186 18578 11551
rect 18830 11578 18858 11583
rect 18942 11578 18970 11583
rect 18830 11577 18970 11578
rect 18830 11551 18831 11577
rect 18857 11551 18943 11577
rect 18969 11551 18970 11577
rect 18830 11550 18970 11551
rect 18830 11242 18858 11550
rect 18942 11545 18970 11550
rect 18774 11186 18802 11191
rect 18550 11185 18802 11186
rect 18550 11159 18775 11185
rect 18801 11159 18802 11185
rect 18550 11158 18802 11159
rect 18550 10793 18578 11158
rect 18550 10767 18551 10793
rect 18577 10767 18578 10793
rect 18550 10761 18578 10767
rect 18774 10401 18802 11158
rect 18830 10794 18858 11214
rect 19054 11186 19082 11943
rect 19334 12754 19362 12759
rect 19446 12754 19474 13119
rect 19334 12753 19474 12754
rect 19334 12727 19335 12753
rect 19361 12727 19447 12753
rect 19473 12727 19474 12753
rect 19334 12726 19474 12727
rect 19054 11153 19082 11158
rect 19222 11242 19250 11247
rect 19222 11185 19250 11214
rect 19334 11242 19362 12726
rect 19446 12721 19474 12726
rect 19573 12558 20035 12563
rect 19573 12557 19582 12558
rect 19573 12531 19574 12557
rect 19573 12530 19582 12531
rect 19610 12530 19634 12558
rect 19662 12530 19686 12558
rect 19714 12557 19738 12558
rect 19766 12557 19790 12558
rect 19724 12531 19738 12557
rect 19786 12531 19790 12557
rect 19714 12530 19738 12531
rect 19766 12530 19790 12531
rect 19818 12557 19842 12558
rect 19870 12557 19894 12558
rect 19818 12531 19822 12557
rect 19870 12531 19884 12557
rect 19818 12530 19842 12531
rect 19870 12530 19894 12531
rect 19922 12530 19946 12558
rect 19974 12530 19998 12558
rect 20026 12557 20035 12558
rect 20034 12531 20035 12557
rect 20026 12530 20035 12531
rect 19573 12525 20035 12530
rect 19446 12417 19474 12423
rect 19446 12391 19447 12417
rect 19473 12391 19474 12417
rect 19446 12362 19474 12391
rect 19446 12361 19530 12362
rect 19446 12335 19447 12361
rect 19473 12335 19530 12361
rect 19446 12334 19530 12335
rect 19446 12329 19474 12334
rect 19334 11209 19362 11214
rect 19502 11914 19530 12334
rect 19222 11159 19223 11185
rect 19249 11159 19250 11185
rect 19222 11153 19250 11159
rect 18830 10761 18858 10766
rect 19278 10849 19306 10855
rect 19278 10823 19279 10849
rect 19305 10823 19306 10849
rect 19278 10793 19306 10823
rect 19278 10767 19279 10793
rect 19305 10767 19306 10793
rect 18774 10375 18775 10401
rect 18801 10375 18802 10401
rect 17990 10039 17991 10065
rect 18017 10039 18018 10065
rect 17990 10009 18018 10039
rect 17990 9983 17991 10009
rect 18017 9983 18018 10009
rect 17073 9814 17535 9819
rect 17073 9813 17082 9814
rect 17073 9787 17074 9813
rect 17073 9786 17082 9787
rect 17110 9786 17134 9814
rect 17162 9786 17186 9814
rect 17214 9813 17238 9814
rect 17266 9813 17290 9814
rect 17224 9787 17238 9813
rect 17286 9787 17290 9813
rect 17214 9786 17238 9787
rect 17266 9786 17290 9787
rect 17318 9813 17342 9814
rect 17370 9813 17394 9814
rect 17318 9787 17322 9813
rect 17370 9787 17384 9813
rect 17318 9786 17342 9787
rect 17370 9786 17394 9787
rect 17422 9786 17446 9814
rect 17474 9786 17498 9814
rect 17526 9813 17535 9814
rect 17534 9787 17535 9813
rect 17526 9786 17535 9787
rect 17073 9781 17535 9786
rect 17990 9282 18018 9983
rect 17990 9225 18018 9254
rect 17990 9199 17991 9225
rect 18017 9199 18018 9225
rect 17073 9030 17535 9035
rect 17073 9029 17082 9030
rect 17073 9003 17074 9029
rect 17073 9002 17082 9003
rect 17110 9002 17134 9030
rect 17162 9002 17186 9030
rect 17214 9029 17238 9030
rect 17266 9029 17290 9030
rect 17224 9003 17238 9029
rect 17286 9003 17290 9029
rect 17214 9002 17238 9003
rect 17266 9002 17290 9003
rect 17318 9029 17342 9030
rect 17370 9029 17394 9030
rect 17318 9003 17322 9029
rect 17370 9003 17384 9029
rect 17318 9002 17342 9003
rect 17370 9002 17394 9003
rect 17422 9002 17446 9030
rect 17474 9002 17498 9030
rect 17526 9029 17535 9030
rect 17534 9003 17535 9029
rect 17526 9002 17535 9003
rect 17073 8997 17535 9002
rect 17990 8497 18018 9199
rect 17990 8471 17991 8497
rect 18017 8471 18018 8497
rect 17990 8441 18018 8471
rect 17990 8415 17991 8441
rect 18017 8415 18018 8441
rect 17990 8409 18018 8415
rect 18214 10346 18242 10351
rect 17073 8246 17535 8251
rect 17073 8245 17082 8246
rect 17073 8219 17074 8245
rect 17073 8218 17082 8219
rect 17110 8218 17134 8246
rect 17162 8218 17186 8246
rect 17214 8245 17238 8246
rect 17266 8245 17290 8246
rect 17224 8219 17238 8245
rect 17286 8219 17290 8245
rect 17214 8218 17238 8219
rect 17266 8218 17290 8219
rect 17318 8245 17342 8246
rect 17370 8245 17394 8246
rect 17318 8219 17322 8245
rect 17370 8219 17384 8245
rect 17318 8218 17342 8219
rect 17370 8218 17394 8219
rect 17422 8218 17446 8246
rect 17474 8218 17498 8246
rect 17526 8245 17535 8246
rect 17534 8219 17535 8245
rect 17526 8218 17535 8219
rect 17073 8213 17535 8218
rect 17598 7657 17626 7663
rect 17598 7631 17599 7657
rect 17625 7631 17626 7657
rect 17073 7462 17535 7467
rect 17073 7461 17082 7462
rect 17073 7435 17074 7461
rect 17073 7434 17082 7435
rect 17110 7434 17134 7462
rect 17162 7434 17186 7462
rect 17214 7461 17238 7462
rect 17266 7461 17290 7462
rect 17224 7435 17238 7461
rect 17286 7435 17290 7461
rect 17214 7434 17238 7435
rect 17266 7434 17290 7435
rect 17318 7461 17342 7462
rect 17370 7461 17394 7462
rect 17318 7435 17322 7461
rect 17370 7435 17384 7461
rect 17318 7434 17342 7435
rect 17370 7434 17394 7435
rect 17422 7434 17446 7462
rect 17474 7434 17498 7462
rect 17526 7461 17535 7462
rect 17534 7435 17535 7461
rect 17526 7434 17535 7435
rect 17073 7429 17535 7434
rect 17486 7266 17514 7271
rect 17598 7266 17626 7631
rect 17486 7265 17626 7266
rect 17486 7239 17487 7265
rect 17513 7239 17626 7265
rect 17486 7238 17626 7239
rect 17486 7233 17514 7238
rect 17598 6873 17626 7238
rect 17598 6847 17599 6873
rect 17625 6847 17626 6873
rect 17073 6678 17535 6683
rect 17073 6677 17082 6678
rect 17073 6651 17074 6677
rect 17073 6650 17082 6651
rect 17110 6650 17134 6678
rect 17162 6650 17186 6678
rect 17214 6677 17238 6678
rect 17266 6677 17290 6678
rect 17224 6651 17238 6677
rect 17286 6651 17290 6677
rect 17214 6650 17238 6651
rect 17266 6650 17290 6651
rect 17318 6677 17342 6678
rect 17370 6677 17394 6678
rect 17318 6651 17322 6677
rect 17370 6651 17384 6677
rect 17318 6650 17342 6651
rect 17370 6650 17394 6651
rect 17422 6650 17446 6678
rect 17474 6650 17498 6678
rect 17526 6677 17535 6678
rect 17534 6651 17535 6677
rect 17526 6650 17535 6651
rect 17073 6645 17535 6650
rect 17486 6482 17514 6487
rect 17598 6482 17626 6847
rect 17514 6454 17626 6482
rect 17486 6416 17514 6454
rect 17598 6089 17626 6454
rect 17598 6063 17599 6089
rect 17625 6063 17626 6089
rect 17073 5894 17535 5899
rect 17073 5893 17082 5894
rect 17073 5867 17074 5893
rect 17073 5866 17082 5867
rect 17110 5866 17134 5894
rect 17162 5866 17186 5894
rect 17214 5893 17238 5894
rect 17266 5893 17290 5894
rect 17224 5867 17238 5893
rect 17286 5867 17290 5893
rect 17214 5866 17238 5867
rect 17266 5866 17290 5867
rect 17318 5893 17342 5894
rect 17370 5893 17394 5894
rect 17318 5867 17322 5893
rect 17370 5867 17384 5893
rect 17318 5866 17342 5867
rect 17370 5866 17394 5867
rect 17422 5866 17446 5894
rect 17474 5866 17498 5894
rect 17526 5893 17535 5894
rect 17534 5867 17535 5893
rect 17526 5866 17535 5867
rect 17073 5861 17535 5866
rect 17486 5698 17514 5703
rect 17598 5698 17626 6063
rect 17486 5697 17626 5698
rect 17486 5671 17487 5697
rect 17513 5671 17626 5697
rect 17486 5670 17626 5671
rect 17486 5665 17514 5670
rect 17598 5305 17626 5670
rect 17598 5279 17599 5305
rect 17625 5279 17626 5305
rect 17073 5110 17535 5115
rect 17073 5109 17082 5110
rect 17073 5083 17074 5109
rect 17073 5082 17082 5083
rect 17110 5082 17134 5110
rect 17162 5082 17186 5110
rect 17214 5109 17238 5110
rect 17266 5109 17290 5110
rect 17224 5083 17238 5109
rect 17286 5083 17290 5109
rect 17214 5082 17238 5083
rect 17266 5082 17290 5083
rect 17318 5109 17342 5110
rect 17370 5109 17394 5110
rect 17318 5083 17322 5109
rect 17370 5083 17384 5109
rect 17318 5082 17342 5083
rect 17370 5082 17394 5083
rect 17422 5082 17446 5110
rect 17474 5082 17498 5110
rect 17526 5109 17535 5110
rect 17534 5083 17535 5109
rect 17526 5082 17535 5083
rect 17073 5077 17535 5082
rect 17486 4914 17514 4919
rect 17598 4914 17626 5279
rect 17486 4913 17626 4914
rect 17486 4887 17487 4913
rect 17513 4887 17626 4913
rect 17486 4886 17626 4887
rect 17486 4881 17514 4886
rect 16982 4433 17010 4438
rect 17598 4521 17626 4886
rect 17598 4495 17599 4521
rect 17625 4495 17626 4521
rect 17073 4326 17535 4331
rect 17073 4325 17082 4326
rect 17073 4299 17074 4325
rect 17073 4298 17082 4299
rect 17110 4298 17134 4326
rect 17162 4298 17186 4326
rect 17214 4325 17238 4326
rect 17266 4325 17290 4326
rect 17224 4299 17238 4325
rect 17286 4299 17290 4325
rect 17214 4298 17238 4299
rect 17266 4298 17290 4299
rect 17318 4325 17342 4326
rect 17370 4325 17394 4326
rect 17318 4299 17322 4325
rect 17370 4299 17384 4325
rect 17318 4298 17342 4299
rect 17370 4298 17394 4299
rect 17422 4298 17446 4326
rect 17474 4298 17498 4326
rect 17526 4325 17535 4326
rect 17534 4299 17535 4325
rect 17526 4298 17535 4299
rect 17073 4293 17535 4298
rect 17486 4130 17514 4135
rect 17598 4130 17626 4495
rect 17486 4129 17626 4130
rect 17486 4103 17487 4129
rect 17513 4103 17626 4129
rect 17486 4102 17626 4103
rect 17486 4097 17514 4102
rect 17598 3737 17626 4102
rect 17598 3711 17599 3737
rect 17625 3711 17626 3737
rect 17073 3542 17535 3547
rect 17073 3541 17082 3542
rect 17073 3515 17074 3541
rect 17073 3514 17082 3515
rect 17110 3514 17134 3542
rect 17162 3514 17186 3542
rect 17214 3541 17238 3542
rect 17266 3541 17290 3542
rect 17224 3515 17238 3541
rect 17286 3515 17290 3541
rect 17214 3514 17238 3515
rect 17266 3514 17290 3515
rect 17318 3541 17342 3542
rect 17370 3541 17394 3542
rect 17318 3515 17322 3541
rect 17370 3515 17384 3541
rect 17318 3514 17342 3515
rect 17370 3514 17394 3515
rect 17422 3514 17446 3542
rect 17474 3514 17498 3542
rect 17526 3541 17535 3542
rect 17534 3515 17535 3541
rect 17526 3514 17535 3515
rect 17073 3509 17535 3514
rect 17598 3402 17626 3711
rect 17486 3346 17514 3351
rect 17598 3346 17626 3374
rect 17486 3345 17626 3346
rect 17486 3319 17487 3345
rect 17513 3319 17626 3345
rect 17486 3318 17626 3319
rect 17486 3313 17514 3318
rect 17598 2953 17626 3318
rect 18214 3010 18242 10318
rect 18270 10009 18298 10015
rect 18270 9983 18271 10009
rect 18297 9983 18298 10009
rect 18270 9225 18298 9983
rect 18270 9199 18271 9225
rect 18297 9199 18298 9225
rect 18270 8442 18298 9199
rect 18270 8395 18298 8414
rect 18774 9617 18802 10375
rect 19278 10402 19306 10767
rect 19502 10402 19530 11886
rect 19950 11969 19978 11975
rect 19950 11943 19951 11969
rect 19977 11943 19978 11969
rect 19950 11914 19978 11943
rect 20286 11970 20314 15862
rect 20846 14322 20874 14327
rect 20790 13930 20818 13935
rect 20790 13883 20818 13902
rect 20510 13538 20538 13543
rect 20510 12753 20538 13510
rect 20846 13454 20874 14294
rect 21014 14321 21042 14327
rect 21014 14295 21015 14321
rect 21041 14295 21042 14321
rect 21014 14266 21042 14295
rect 21182 14266 21210 14271
rect 21014 14265 21210 14266
rect 21014 14239 21183 14265
rect 21209 14239 21210 14265
rect 21014 14238 21210 14239
rect 21014 13537 21042 14238
rect 21182 14233 21210 14238
rect 21742 13985 21770 13991
rect 21742 13959 21743 13985
rect 21769 13959 21770 13985
rect 21742 13929 21770 13959
rect 21742 13903 21743 13929
rect 21769 13903 21770 13929
rect 21014 13511 21015 13537
rect 21041 13511 21042 13537
rect 21014 13482 21042 13511
rect 21406 13538 21434 13543
rect 21182 13482 21210 13487
rect 21238 13482 21266 13487
rect 21014 13481 21238 13482
rect 21014 13455 21183 13481
rect 21209 13455 21238 13481
rect 21014 13454 21238 13455
rect 20846 13426 20986 13454
rect 20510 12727 20511 12753
rect 20537 12727 20538 12753
rect 20510 12362 20538 12727
rect 20958 13145 20986 13426
rect 20958 13119 20959 13145
rect 20985 13119 20986 13145
rect 20902 12362 20930 12367
rect 20510 12361 20930 12362
rect 20510 12335 20903 12361
rect 20929 12335 20930 12361
rect 20510 12334 20930 12335
rect 20510 11970 20538 11975
rect 20286 11969 20818 11970
rect 20286 11943 20511 11969
rect 20537 11943 20818 11969
rect 20286 11942 20818 11943
rect 20510 11937 20538 11942
rect 19950 11867 19978 11886
rect 19573 11774 20035 11779
rect 19573 11773 19582 11774
rect 19573 11747 19574 11773
rect 19573 11746 19582 11747
rect 19610 11746 19634 11774
rect 19662 11746 19686 11774
rect 19714 11773 19738 11774
rect 19766 11773 19790 11774
rect 19724 11747 19738 11773
rect 19786 11747 19790 11773
rect 19714 11746 19738 11747
rect 19766 11746 19790 11747
rect 19818 11773 19842 11774
rect 19870 11773 19894 11774
rect 19818 11747 19822 11773
rect 19870 11747 19884 11773
rect 19818 11746 19842 11747
rect 19870 11746 19894 11747
rect 19922 11746 19946 11774
rect 19974 11746 19998 11774
rect 20026 11773 20035 11774
rect 20034 11747 20035 11773
rect 20026 11746 20035 11747
rect 19573 11741 20035 11746
rect 20790 11577 20818 11942
rect 20790 11551 20791 11577
rect 20817 11551 20818 11577
rect 20790 11545 20818 11551
rect 19950 11242 19978 11247
rect 19950 11185 19978 11214
rect 19950 11159 19951 11185
rect 19977 11159 19978 11185
rect 19950 11074 19978 11159
rect 20230 11186 20258 11191
rect 20230 11139 20258 11158
rect 20790 11186 20818 11191
rect 19950 11041 19978 11046
rect 19573 10990 20035 10995
rect 19573 10989 19582 10990
rect 19573 10963 19574 10989
rect 19573 10962 19582 10963
rect 19610 10962 19634 10990
rect 19662 10962 19686 10990
rect 19714 10989 19738 10990
rect 19766 10989 19790 10990
rect 19724 10963 19738 10989
rect 19786 10963 19790 10989
rect 19714 10962 19738 10963
rect 19766 10962 19790 10963
rect 19818 10989 19842 10990
rect 19870 10989 19894 10990
rect 19818 10963 19822 10989
rect 19870 10963 19884 10989
rect 19818 10962 19842 10963
rect 19870 10962 19894 10963
rect 19922 10962 19946 10990
rect 19974 10962 19998 10990
rect 20026 10989 20035 10990
rect 20034 10963 20035 10989
rect 20026 10962 20035 10963
rect 19573 10957 20035 10962
rect 20790 10794 20818 11158
rect 20902 10794 20930 12334
rect 20958 12362 20986 13119
rect 21014 12754 21042 13454
rect 21182 13449 21210 13454
rect 21238 13426 21322 13454
rect 21238 13416 21266 13426
rect 21294 13145 21322 13426
rect 21294 13119 21295 13145
rect 21321 13119 21322 13145
rect 21294 13113 21322 13119
rect 21294 12754 21322 12759
rect 21014 12753 21322 12754
rect 21014 12727 21295 12753
rect 21321 12727 21322 12753
rect 21014 12726 21322 12727
rect 20958 12329 20986 12334
rect 21294 12697 21322 12726
rect 21294 12671 21295 12697
rect 21321 12671 21322 12697
rect 20790 10793 20874 10794
rect 20790 10767 20791 10793
rect 20817 10767 20874 10793
rect 20790 10766 20874 10767
rect 20790 10761 20818 10766
rect 19278 10401 19530 10402
rect 19278 10375 19279 10401
rect 19305 10375 19503 10401
rect 19529 10375 19530 10401
rect 19278 10374 19530 10375
rect 19278 10369 19306 10374
rect 19446 10065 19474 10374
rect 19502 10369 19530 10374
rect 20230 10401 20258 10407
rect 20230 10375 20231 10401
rect 20257 10375 20258 10401
rect 19573 10206 20035 10211
rect 19573 10205 19582 10206
rect 19573 10179 19574 10205
rect 19573 10178 19582 10179
rect 19610 10178 19634 10206
rect 19662 10178 19686 10206
rect 19714 10205 19738 10206
rect 19766 10205 19790 10206
rect 19724 10179 19738 10205
rect 19786 10179 19790 10205
rect 19714 10178 19738 10179
rect 19766 10178 19790 10179
rect 19818 10205 19842 10206
rect 19870 10205 19894 10206
rect 19818 10179 19822 10205
rect 19870 10179 19884 10205
rect 19818 10178 19842 10179
rect 19870 10178 19894 10179
rect 19922 10178 19946 10206
rect 19974 10178 19998 10206
rect 20026 10205 20035 10206
rect 20034 10179 20035 10205
rect 20026 10178 20035 10179
rect 19573 10173 20035 10178
rect 19446 10039 19447 10065
rect 19473 10039 19474 10065
rect 19446 10009 19474 10039
rect 19446 9983 19447 10009
rect 19473 9983 19474 10009
rect 18774 9591 18775 9617
rect 18801 9591 18802 9617
rect 18774 8833 18802 9591
rect 19334 9618 19362 9623
rect 19446 9618 19474 9983
rect 19334 9617 19474 9618
rect 19334 9591 19335 9617
rect 19361 9591 19447 9617
rect 19473 9591 19474 9617
rect 19334 9590 19474 9591
rect 19278 9282 19306 9287
rect 19334 9282 19362 9590
rect 19446 9585 19474 9590
rect 20230 9617 20258 10375
rect 20230 9591 20231 9617
rect 20257 9591 20258 9617
rect 19573 9422 20035 9427
rect 19573 9421 19582 9422
rect 19573 9395 19574 9421
rect 19573 9394 19582 9395
rect 19610 9394 19634 9422
rect 19662 9394 19686 9422
rect 19714 9421 19738 9422
rect 19766 9421 19790 9422
rect 19724 9395 19738 9421
rect 19786 9395 19790 9421
rect 19714 9394 19738 9395
rect 19766 9394 19790 9395
rect 19818 9421 19842 9422
rect 19870 9421 19894 9422
rect 19818 9395 19822 9421
rect 19870 9395 19884 9421
rect 19818 9394 19842 9395
rect 19870 9394 19894 9395
rect 19922 9394 19946 9422
rect 19974 9394 19998 9422
rect 20026 9421 20035 9422
rect 20034 9395 20035 9421
rect 20026 9394 20035 9395
rect 19573 9389 20035 9394
rect 19306 9281 19362 9282
rect 19306 9255 19335 9281
rect 19361 9255 19362 9281
rect 19306 9254 19362 9255
rect 19278 9225 19306 9254
rect 19278 9199 19279 9225
rect 19305 9199 19306 9225
rect 19334 9216 19362 9254
rect 19278 9193 19306 9199
rect 18774 8807 18775 8833
rect 18801 8807 18802 8833
rect 18774 8442 18802 8807
rect 19334 8834 19362 8839
rect 19446 8834 19474 8839
rect 19334 8833 19474 8834
rect 19334 8807 19335 8833
rect 19361 8807 19447 8833
rect 19473 8807 19474 8833
rect 19334 8806 19474 8807
rect 19334 8801 19362 8806
rect 18774 8049 18802 8414
rect 19446 8497 19474 8806
rect 20230 8833 20258 9591
rect 20230 8807 20231 8833
rect 20257 8807 20258 8833
rect 19573 8638 20035 8643
rect 19573 8637 19582 8638
rect 19573 8611 19574 8637
rect 19573 8610 19582 8611
rect 19610 8610 19634 8638
rect 19662 8610 19686 8638
rect 19714 8637 19738 8638
rect 19766 8637 19790 8638
rect 19724 8611 19738 8637
rect 19786 8611 19790 8637
rect 19714 8610 19738 8611
rect 19766 8610 19790 8611
rect 19818 8637 19842 8638
rect 19870 8637 19894 8638
rect 19818 8611 19822 8637
rect 19870 8611 19884 8637
rect 19818 8610 19842 8611
rect 19870 8610 19894 8611
rect 19922 8610 19946 8638
rect 19974 8610 19998 8638
rect 20026 8637 20035 8638
rect 20034 8611 20035 8637
rect 20026 8610 20035 8611
rect 19573 8605 20035 8610
rect 19446 8471 19447 8497
rect 19473 8471 19474 8497
rect 19446 8442 19474 8471
rect 20230 8498 20258 8807
rect 19446 8395 19474 8414
rect 19950 8442 19978 8447
rect 18774 8023 18775 8049
rect 18801 8023 18802 8049
rect 18774 8017 18802 8023
rect 19950 8049 19978 8414
rect 19950 8023 19951 8049
rect 19977 8023 19978 8049
rect 19950 7993 19978 8023
rect 20230 8049 20258 8470
rect 20790 10009 20818 10015
rect 20790 9983 20791 10009
rect 20817 9983 20818 10009
rect 20790 9225 20818 9983
rect 20846 10010 20874 10766
rect 20902 10761 20930 10766
rect 21294 11074 21322 12671
rect 21406 11969 21434 13510
rect 21742 13538 21770 13903
rect 21742 13505 21770 13510
rect 21462 13482 21490 13487
rect 21462 13145 21490 13454
rect 21462 13119 21463 13145
rect 21489 13119 21490 13145
rect 21462 13113 21490 13119
rect 21798 12417 21826 12423
rect 21798 12391 21799 12417
rect 21825 12391 21826 12417
rect 21798 12361 21826 12391
rect 21798 12335 21799 12361
rect 21825 12335 21826 12361
rect 21798 12250 21826 12335
rect 21798 12217 21826 12222
rect 21406 11943 21407 11969
rect 21433 11943 21434 11969
rect 21294 10402 21322 11046
rect 21350 11914 21378 11919
rect 21406 11914 21434 11943
rect 21378 11913 21434 11914
rect 21378 11887 21407 11913
rect 21433 11887 21434 11913
rect 21378 11886 21434 11887
rect 21350 11578 21378 11886
rect 21406 11881 21434 11886
rect 21462 11578 21490 11583
rect 21350 11577 21490 11578
rect 21350 11551 21351 11577
rect 21377 11551 21463 11577
rect 21489 11551 21490 11577
rect 21350 11550 21490 11551
rect 21350 11185 21378 11550
rect 21462 11545 21490 11550
rect 21350 11159 21351 11185
rect 21377 11159 21378 11185
rect 21350 11129 21378 11159
rect 21350 11103 21351 11129
rect 21377 11103 21378 11129
rect 21350 10794 21378 11103
rect 21854 11186 21882 19614
rect 22302 19530 22330 19614
rect 22456 19600 22512 20000
rect 26894 19614 27314 19642
rect 22470 19530 22498 19600
rect 22302 19502 22498 19530
rect 22073 18438 22535 18443
rect 22073 18437 22082 18438
rect 22073 18411 22074 18437
rect 22073 18410 22082 18411
rect 22110 18410 22134 18438
rect 22162 18410 22186 18438
rect 22214 18437 22238 18438
rect 22266 18437 22290 18438
rect 22224 18411 22238 18437
rect 22286 18411 22290 18437
rect 22214 18410 22238 18411
rect 22266 18410 22290 18411
rect 22318 18437 22342 18438
rect 22370 18437 22394 18438
rect 22318 18411 22322 18437
rect 22370 18411 22384 18437
rect 22318 18410 22342 18411
rect 22370 18410 22394 18411
rect 22422 18410 22446 18438
rect 22474 18410 22498 18438
rect 22526 18437 22535 18438
rect 22534 18411 22535 18437
rect 22526 18410 22535 18411
rect 22073 18405 22535 18410
rect 24573 18046 25035 18051
rect 24573 18045 24582 18046
rect 24573 18019 24574 18045
rect 24573 18018 24582 18019
rect 24610 18018 24634 18046
rect 24662 18018 24686 18046
rect 24714 18045 24738 18046
rect 24766 18045 24790 18046
rect 24724 18019 24738 18045
rect 24786 18019 24790 18045
rect 24714 18018 24738 18019
rect 24766 18018 24790 18019
rect 24818 18045 24842 18046
rect 24870 18045 24894 18046
rect 24818 18019 24822 18045
rect 24870 18019 24884 18045
rect 24818 18018 24842 18019
rect 24870 18018 24894 18019
rect 24922 18018 24946 18046
rect 24974 18018 24998 18046
rect 25026 18045 25035 18046
rect 25034 18019 25035 18045
rect 25026 18018 25035 18019
rect 24573 18013 25035 18018
rect 22073 17654 22535 17659
rect 22073 17653 22082 17654
rect 22073 17627 22074 17653
rect 22073 17626 22082 17627
rect 22110 17626 22134 17654
rect 22162 17626 22186 17654
rect 22214 17653 22238 17654
rect 22266 17653 22290 17654
rect 22224 17627 22238 17653
rect 22286 17627 22290 17653
rect 22214 17626 22238 17627
rect 22266 17626 22290 17627
rect 22318 17653 22342 17654
rect 22370 17653 22394 17654
rect 22318 17627 22322 17653
rect 22370 17627 22384 17653
rect 22318 17626 22342 17627
rect 22370 17626 22394 17627
rect 22422 17626 22446 17654
rect 22474 17626 22498 17654
rect 22526 17653 22535 17654
rect 22534 17627 22535 17653
rect 22526 17626 22535 17627
rect 22073 17621 22535 17626
rect 23926 17346 23954 17351
rect 22073 16870 22535 16875
rect 22073 16869 22082 16870
rect 22073 16843 22074 16869
rect 22073 16842 22082 16843
rect 22110 16842 22134 16870
rect 22162 16842 22186 16870
rect 22214 16869 22238 16870
rect 22266 16869 22290 16870
rect 22224 16843 22238 16869
rect 22286 16843 22290 16869
rect 22214 16842 22238 16843
rect 22266 16842 22290 16843
rect 22318 16869 22342 16870
rect 22370 16869 22394 16870
rect 22318 16843 22322 16869
rect 22370 16843 22384 16869
rect 22318 16842 22342 16843
rect 22370 16842 22394 16843
rect 22422 16842 22446 16870
rect 22474 16842 22498 16870
rect 22526 16869 22535 16870
rect 22534 16843 22535 16869
rect 22526 16842 22535 16843
rect 22073 16837 22535 16842
rect 22073 16086 22535 16091
rect 22073 16085 22082 16086
rect 22073 16059 22074 16085
rect 22073 16058 22082 16059
rect 22110 16058 22134 16086
rect 22162 16058 22186 16086
rect 22214 16085 22238 16086
rect 22266 16085 22290 16086
rect 22224 16059 22238 16085
rect 22286 16059 22290 16085
rect 22214 16058 22238 16059
rect 22266 16058 22290 16059
rect 22318 16085 22342 16086
rect 22370 16085 22394 16086
rect 22318 16059 22322 16085
rect 22370 16059 22384 16085
rect 22318 16058 22342 16059
rect 22370 16058 22394 16059
rect 22422 16058 22446 16086
rect 22474 16058 22498 16086
rect 22526 16085 22535 16086
rect 22534 16059 22535 16085
rect 22526 16058 22535 16059
rect 22073 16053 22535 16058
rect 22073 15302 22535 15307
rect 22073 15301 22082 15302
rect 22073 15275 22074 15301
rect 22073 15274 22082 15275
rect 22110 15274 22134 15302
rect 22162 15274 22186 15302
rect 22214 15301 22238 15302
rect 22266 15301 22290 15302
rect 22224 15275 22238 15301
rect 22286 15275 22290 15301
rect 22214 15274 22238 15275
rect 22266 15274 22290 15275
rect 22318 15301 22342 15302
rect 22370 15301 22394 15302
rect 22318 15275 22322 15301
rect 22370 15275 22384 15301
rect 22318 15274 22342 15275
rect 22370 15274 22394 15275
rect 22422 15274 22446 15302
rect 22474 15274 22498 15302
rect 22526 15301 22535 15302
rect 22534 15275 22535 15301
rect 22526 15274 22535 15275
rect 22073 15269 22535 15274
rect 22073 14518 22535 14523
rect 22073 14517 22082 14518
rect 22073 14491 22074 14517
rect 22073 14490 22082 14491
rect 22110 14490 22134 14518
rect 22162 14490 22186 14518
rect 22214 14517 22238 14518
rect 22266 14517 22290 14518
rect 22224 14491 22238 14517
rect 22286 14491 22290 14517
rect 22214 14490 22238 14491
rect 22266 14490 22290 14491
rect 22318 14517 22342 14518
rect 22370 14517 22394 14518
rect 22318 14491 22322 14517
rect 22370 14491 22384 14517
rect 22318 14490 22342 14491
rect 22370 14490 22394 14491
rect 22422 14490 22446 14518
rect 22474 14490 22498 14518
rect 22526 14517 22535 14518
rect 22534 14491 22535 14517
rect 22526 14490 22535 14491
rect 22073 14485 22535 14490
rect 23030 14321 23058 14327
rect 23030 14295 23031 14321
rect 23057 14295 23058 14321
rect 22526 13930 22554 13935
rect 22526 13929 22610 13930
rect 22526 13903 22527 13929
rect 22553 13903 22610 13929
rect 22526 13902 22610 13903
rect 22526 13897 22554 13902
rect 22582 13874 22610 13902
rect 22073 13734 22535 13739
rect 22073 13733 22082 13734
rect 22073 13707 22074 13733
rect 22073 13706 22082 13707
rect 22110 13706 22134 13734
rect 22162 13706 22186 13734
rect 22214 13733 22238 13734
rect 22266 13733 22290 13734
rect 22224 13707 22238 13733
rect 22286 13707 22290 13733
rect 22214 13706 22238 13707
rect 22266 13706 22290 13707
rect 22318 13733 22342 13734
rect 22370 13733 22394 13734
rect 22318 13707 22322 13733
rect 22370 13707 22384 13733
rect 22318 13706 22342 13707
rect 22370 13706 22394 13707
rect 22422 13706 22446 13734
rect 22474 13706 22498 13734
rect 22526 13733 22535 13734
rect 22534 13707 22535 13733
rect 22526 13706 22535 13707
rect 22073 13701 22535 13706
rect 22526 13482 22554 13487
rect 22582 13482 22610 13846
rect 22554 13454 22610 13482
rect 23030 13537 23058 14295
rect 23870 14321 23898 14327
rect 23870 14295 23871 14321
rect 23897 14295 23898 14321
rect 23870 14266 23898 14295
rect 23870 14219 23898 14238
rect 23030 13511 23031 13537
rect 23057 13511 23058 13537
rect 23030 13482 23058 13511
rect 22526 13145 22554 13454
rect 22526 13119 22527 13145
rect 22553 13119 22554 13145
rect 22526 13113 22554 13119
rect 22974 13426 23058 13454
rect 23422 13985 23450 13991
rect 23422 13959 23423 13985
rect 23449 13959 23450 13985
rect 23422 13929 23450 13959
rect 23422 13903 23423 13929
rect 23449 13903 23450 13929
rect 23422 13538 23450 13903
rect 22073 12950 22535 12955
rect 22073 12949 22082 12950
rect 22073 12923 22074 12949
rect 22073 12922 22082 12923
rect 22110 12922 22134 12950
rect 22162 12922 22186 12950
rect 22214 12949 22238 12950
rect 22266 12949 22290 12950
rect 22224 12923 22238 12949
rect 22286 12923 22290 12949
rect 22214 12922 22238 12923
rect 22266 12922 22290 12923
rect 22318 12949 22342 12950
rect 22370 12949 22394 12950
rect 22318 12923 22322 12949
rect 22370 12923 22384 12949
rect 22318 12922 22342 12923
rect 22370 12922 22394 12923
rect 22422 12922 22446 12950
rect 22474 12922 22498 12950
rect 22526 12949 22535 12950
rect 22534 12923 22535 12949
rect 22526 12922 22535 12923
rect 22073 12917 22535 12922
rect 22974 12753 23002 13426
rect 23422 13201 23450 13510
rect 23422 13175 23423 13201
rect 23449 13175 23450 13201
rect 23422 13145 23450 13175
rect 23422 13119 23423 13145
rect 23449 13119 23450 13145
rect 23422 13113 23450 13119
rect 23870 13538 23898 13543
rect 23870 13481 23898 13510
rect 23870 13455 23871 13481
rect 23897 13455 23898 13481
rect 22974 12727 22975 12753
rect 23001 12727 23002 12753
rect 22974 12721 23002 12727
rect 23870 12753 23898 13455
rect 23870 12727 23871 12753
rect 23897 12727 23898 12753
rect 23870 12698 23898 12727
rect 23870 12651 23898 12670
rect 23422 12417 23450 12423
rect 23422 12391 23423 12417
rect 23449 12391 23450 12417
rect 22526 12362 22554 12367
rect 22554 12334 22610 12362
rect 22526 12296 22554 12334
rect 22073 12166 22535 12171
rect 22073 12165 22082 12166
rect 22073 12139 22074 12165
rect 22073 12138 22082 12139
rect 22110 12138 22134 12166
rect 22162 12138 22186 12166
rect 22214 12165 22238 12166
rect 22266 12165 22290 12166
rect 22224 12139 22238 12165
rect 22286 12139 22290 12165
rect 22214 12138 22238 12139
rect 22266 12138 22290 12139
rect 22318 12165 22342 12166
rect 22370 12165 22394 12166
rect 22318 12139 22322 12165
rect 22370 12139 22384 12165
rect 22318 12138 22342 12139
rect 22370 12138 22394 12139
rect 22422 12138 22446 12166
rect 22474 12138 22498 12166
rect 22526 12165 22535 12166
rect 22534 12139 22535 12165
rect 22526 12138 22535 12139
rect 22073 12133 22535 12138
rect 22582 11970 22610 12334
rect 23422 12361 23450 12391
rect 23422 12335 23423 12361
rect 23449 12335 23450 12361
rect 23422 12250 23450 12335
rect 22582 11937 22610 11942
rect 23030 11970 23058 11975
rect 23030 11923 23058 11942
rect 23310 11970 23338 11975
rect 23422 11970 23450 12222
rect 23310 11969 23450 11970
rect 23310 11943 23311 11969
rect 23337 11943 23423 11969
rect 23449 11943 23450 11969
rect 23310 11942 23450 11943
rect 23310 11633 23338 11942
rect 23422 11937 23450 11942
rect 23310 11607 23311 11633
rect 23337 11607 23338 11633
rect 22526 11578 22554 11583
rect 22526 11577 22610 11578
rect 22526 11551 22527 11577
rect 22553 11551 22610 11577
rect 22526 11550 22610 11551
rect 22526 11545 22554 11550
rect 22073 11382 22535 11387
rect 22073 11381 22082 11382
rect 22073 11355 22074 11381
rect 22073 11354 22082 11355
rect 22110 11354 22134 11382
rect 22162 11354 22186 11382
rect 22214 11381 22238 11382
rect 22266 11381 22290 11382
rect 22224 11355 22238 11381
rect 22286 11355 22290 11381
rect 22214 11354 22238 11355
rect 22266 11354 22290 11355
rect 22318 11381 22342 11382
rect 22370 11381 22394 11382
rect 22318 11355 22322 11381
rect 22370 11355 22384 11381
rect 22318 11354 22342 11355
rect 22370 11354 22394 11355
rect 22422 11354 22446 11382
rect 22474 11354 22498 11382
rect 22526 11381 22535 11382
rect 22534 11355 22535 11381
rect 22526 11354 22535 11355
rect 22073 11349 22535 11354
rect 21462 10794 21490 10799
rect 21350 10793 21490 10794
rect 21350 10767 21351 10793
rect 21377 10767 21463 10793
rect 21489 10767 21490 10793
rect 21350 10766 21490 10767
rect 21350 10761 21378 10766
rect 21462 10761 21490 10766
rect 21350 10402 21378 10407
rect 21294 10401 21378 10402
rect 21294 10375 21351 10401
rect 21377 10375 21378 10401
rect 21294 10374 21378 10375
rect 20846 9977 20874 9982
rect 21350 10345 21378 10374
rect 21350 10319 21351 10345
rect 21377 10319 21378 10345
rect 21350 10010 21378 10319
rect 21462 10010 21490 10015
rect 21350 10009 21490 10010
rect 21350 9983 21351 10009
rect 21377 9983 21463 10009
rect 21489 9983 21490 10009
rect 21350 9982 21490 9983
rect 20790 9199 20791 9225
rect 20817 9199 20818 9225
rect 20790 8498 20818 9199
rect 21350 9617 21378 9982
rect 21462 9977 21490 9982
rect 21350 9591 21351 9617
rect 21377 9591 21378 9617
rect 21350 9561 21378 9591
rect 21350 9535 21351 9561
rect 21377 9535 21378 9561
rect 21350 9226 21378 9535
rect 21462 9226 21490 9231
rect 21350 9225 21490 9226
rect 21350 9199 21351 9225
rect 21377 9199 21463 9225
rect 21489 9199 21490 9225
rect 21350 9198 21490 9199
rect 21350 9193 21378 9198
rect 20790 8441 20818 8470
rect 20790 8415 20791 8441
rect 20817 8415 20818 8441
rect 20790 8409 20818 8415
rect 21406 8833 21434 9198
rect 21462 9193 21490 9198
rect 21406 8807 21407 8833
rect 21433 8807 21434 8833
rect 21406 8777 21434 8807
rect 21406 8751 21407 8777
rect 21433 8751 21434 8777
rect 21406 8442 21434 8751
rect 20230 8023 20231 8049
rect 20257 8023 20258 8049
rect 20230 8017 20258 8023
rect 21406 8330 21434 8414
rect 21406 8049 21434 8302
rect 21798 8497 21826 8503
rect 21798 8471 21799 8497
rect 21825 8471 21826 8497
rect 21798 8441 21826 8471
rect 21798 8415 21799 8441
rect 21825 8415 21826 8441
rect 21798 8330 21826 8415
rect 21798 8297 21826 8302
rect 21406 8023 21407 8049
rect 21433 8023 21434 8049
rect 19950 7967 19951 7993
rect 19977 7967 19978 7993
rect 19950 7961 19978 7967
rect 21406 7993 21434 8023
rect 21406 7967 21407 7993
rect 21433 7967 21434 7993
rect 21406 7961 21434 7967
rect 19573 7854 20035 7859
rect 19573 7853 19582 7854
rect 19573 7827 19574 7853
rect 19573 7826 19582 7827
rect 19610 7826 19634 7854
rect 19662 7826 19686 7854
rect 19714 7853 19738 7854
rect 19766 7853 19790 7854
rect 19724 7827 19738 7853
rect 19786 7827 19790 7853
rect 19714 7826 19738 7827
rect 19766 7826 19790 7827
rect 19818 7853 19842 7854
rect 19870 7853 19894 7854
rect 19818 7827 19822 7853
rect 19870 7827 19884 7853
rect 19818 7826 19842 7827
rect 19870 7826 19894 7827
rect 19922 7826 19946 7854
rect 19974 7826 19998 7854
rect 20026 7853 20035 7854
rect 20034 7827 20035 7853
rect 20026 7826 20035 7827
rect 19573 7821 20035 7826
rect 18382 7713 18410 7719
rect 18382 7687 18383 7713
rect 18409 7687 18410 7713
rect 18382 7657 18410 7687
rect 20006 7713 20034 7719
rect 20006 7687 20007 7713
rect 20033 7687 20034 7713
rect 18382 7631 18383 7657
rect 18409 7631 18410 7657
rect 18382 7265 18410 7631
rect 19110 7657 19138 7663
rect 19110 7631 19111 7657
rect 19137 7631 19138 7657
rect 18382 7239 18383 7265
rect 18409 7239 18410 7265
rect 18382 7210 18410 7239
rect 19054 7266 19082 7271
rect 19110 7266 19138 7631
rect 20006 7658 20034 7687
rect 21798 7714 21826 7719
rect 21854 7714 21882 11158
rect 22526 10794 22554 10799
rect 22582 10794 22610 11550
rect 23310 11577 23338 11607
rect 23310 11551 23311 11577
rect 23337 11551 23338 11577
rect 22554 10766 22610 10794
rect 23030 11185 23058 11191
rect 23030 11159 23031 11185
rect 23057 11159 23058 11185
rect 23030 10794 23058 11159
rect 23310 11186 23338 11551
rect 23422 11186 23450 11191
rect 23310 11185 23450 11186
rect 23310 11159 23311 11185
rect 23337 11159 23423 11185
rect 23449 11159 23450 11185
rect 23310 11158 23450 11159
rect 23310 11153 23338 11158
rect 22526 10747 22554 10766
rect 22073 10598 22535 10603
rect 22073 10597 22082 10598
rect 22073 10571 22074 10597
rect 22073 10570 22082 10571
rect 22110 10570 22134 10598
rect 22162 10570 22186 10598
rect 22214 10597 22238 10598
rect 22266 10597 22290 10598
rect 22224 10571 22238 10597
rect 22286 10571 22290 10597
rect 22214 10570 22238 10571
rect 22266 10570 22290 10571
rect 22318 10597 22342 10598
rect 22370 10597 22394 10598
rect 22318 10571 22322 10597
rect 22370 10571 22384 10597
rect 22318 10570 22342 10571
rect 22370 10570 22394 10571
rect 22422 10570 22446 10598
rect 22474 10570 22498 10598
rect 22526 10597 22535 10598
rect 22534 10571 22535 10597
rect 22526 10570 22535 10571
rect 22073 10565 22535 10570
rect 23030 10401 23058 10766
rect 23030 10375 23031 10401
rect 23057 10375 23058 10401
rect 23030 10290 23058 10375
rect 23030 10257 23058 10262
rect 23422 10849 23450 11158
rect 23422 10823 23423 10849
rect 23449 10823 23450 10849
rect 23422 10793 23450 10823
rect 23422 10767 23423 10793
rect 23449 10767 23450 10793
rect 23422 10065 23450 10767
rect 23422 10039 23423 10065
rect 23449 10039 23450 10065
rect 22246 10010 22274 10015
rect 22246 9963 22274 9982
rect 22582 10010 22610 10015
rect 22073 9814 22535 9819
rect 22073 9813 22082 9814
rect 22073 9787 22074 9813
rect 22073 9786 22082 9787
rect 22110 9786 22134 9814
rect 22162 9786 22186 9814
rect 22214 9813 22238 9814
rect 22266 9813 22290 9814
rect 22224 9787 22238 9813
rect 22286 9787 22290 9813
rect 22214 9786 22238 9787
rect 22266 9786 22290 9787
rect 22318 9813 22342 9814
rect 22370 9813 22394 9814
rect 22318 9787 22322 9813
rect 22370 9787 22384 9813
rect 22318 9786 22342 9787
rect 22370 9786 22394 9787
rect 22422 9786 22446 9814
rect 22474 9786 22498 9814
rect 22526 9813 22535 9814
rect 22534 9787 22535 9813
rect 22526 9786 22535 9787
rect 22073 9781 22535 9786
rect 22582 9618 22610 9982
rect 23422 10010 23450 10039
rect 23422 9963 23450 9982
rect 23870 10401 23898 10407
rect 23870 10375 23871 10401
rect 23897 10375 23898 10401
rect 23870 10345 23898 10375
rect 23870 10319 23871 10345
rect 23897 10319 23898 10345
rect 23870 10010 23898 10319
rect 22750 9618 22778 9623
rect 22582 9617 22778 9618
rect 22582 9591 22751 9617
rect 22777 9591 22778 9617
rect 22582 9590 22778 9591
rect 22526 9226 22554 9231
rect 22582 9226 22610 9590
rect 22526 9225 22610 9226
rect 22526 9199 22527 9225
rect 22553 9199 22610 9225
rect 22526 9198 22610 9199
rect 22526 9193 22554 9198
rect 22073 9030 22535 9035
rect 22073 9029 22082 9030
rect 22073 9003 22074 9029
rect 22073 9002 22082 9003
rect 22110 9002 22134 9030
rect 22162 9002 22186 9030
rect 22214 9029 22238 9030
rect 22266 9029 22290 9030
rect 22224 9003 22238 9029
rect 22286 9003 22290 9029
rect 22214 9002 22238 9003
rect 22266 9002 22290 9003
rect 22318 9029 22342 9030
rect 22370 9029 22394 9030
rect 22318 9003 22322 9029
rect 22370 9003 22384 9029
rect 22318 9002 22342 9003
rect 22370 9002 22394 9003
rect 22422 9002 22446 9030
rect 22474 9002 22498 9030
rect 22526 9029 22535 9030
rect 22534 9003 22535 9029
rect 22526 9002 22535 9003
rect 22073 8997 22535 9002
rect 22526 8442 22554 8447
rect 22582 8442 22610 9198
rect 22526 8441 22610 8442
rect 22526 8415 22527 8441
rect 22553 8415 22610 8441
rect 22526 8414 22610 8415
rect 22750 8833 22778 9590
rect 23870 9617 23898 9982
rect 23870 9591 23871 9617
rect 23897 9591 23898 9617
rect 23870 9562 23898 9591
rect 23870 9515 23898 9534
rect 22750 8807 22751 8833
rect 22777 8807 22778 8833
rect 22526 8409 22554 8414
rect 22073 8246 22535 8251
rect 22073 8245 22082 8246
rect 22073 8219 22074 8245
rect 22073 8218 22082 8219
rect 22110 8218 22134 8246
rect 22162 8218 22186 8246
rect 22214 8245 22238 8246
rect 22266 8245 22290 8246
rect 22224 8219 22238 8245
rect 22286 8219 22290 8245
rect 22214 8218 22238 8219
rect 22266 8218 22290 8219
rect 22318 8245 22342 8246
rect 22370 8245 22394 8246
rect 22318 8219 22322 8245
rect 22370 8219 22384 8245
rect 22318 8218 22342 8219
rect 22370 8218 22394 8219
rect 22422 8218 22446 8246
rect 22474 8218 22498 8246
rect 22526 8245 22535 8246
rect 22534 8219 22535 8245
rect 22526 8218 22535 8219
rect 22073 8213 22535 8218
rect 21798 7713 21882 7714
rect 21798 7687 21799 7713
rect 21825 7687 21882 7713
rect 21798 7686 21882 7687
rect 22750 8049 22778 8807
rect 23422 9281 23450 9287
rect 23422 9255 23423 9281
rect 23449 9255 23450 9281
rect 23422 9225 23450 9255
rect 23422 9199 23423 9225
rect 23449 9199 23450 9225
rect 23422 8890 23450 9199
rect 23422 8497 23450 8862
rect 23870 8890 23898 8895
rect 23870 8833 23898 8862
rect 23870 8807 23871 8833
rect 23897 8807 23898 8833
rect 23870 8777 23898 8807
rect 23870 8751 23871 8777
rect 23897 8751 23898 8777
rect 23870 8745 23898 8751
rect 23422 8471 23423 8497
rect 23449 8471 23450 8497
rect 23422 8441 23450 8471
rect 23422 8415 23423 8441
rect 23449 8415 23450 8441
rect 23422 8409 23450 8415
rect 22750 8023 22751 8049
rect 22777 8023 22778 8049
rect 19054 7265 19138 7266
rect 19054 7239 19055 7265
rect 19081 7239 19138 7265
rect 19054 7238 19138 7239
rect 19054 7233 19082 7238
rect 18382 7209 18466 7210
rect 18382 7183 18383 7209
rect 18409 7183 18466 7209
rect 18382 7182 18466 7183
rect 18382 7177 18410 7182
rect 18438 6929 18466 7182
rect 18438 6903 18439 6929
rect 18465 6903 18466 6929
rect 18438 6873 18466 6903
rect 18438 6847 18439 6873
rect 18465 6847 18466 6873
rect 18382 6481 18410 6487
rect 18382 6455 18383 6481
rect 18409 6455 18410 6481
rect 18382 6426 18410 6455
rect 18438 6426 18466 6847
rect 19110 6873 19138 7238
rect 19950 7266 19978 7271
rect 20006 7266 20034 7630
rect 20958 7657 20986 7663
rect 20958 7631 20959 7657
rect 20985 7631 20986 7657
rect 19950 7265 20034 7266
rect 19950 7239 19951 7265
rect 19977 7239 20034 7265
rect 19950 7238 20034 7239
rect 20510 7266 20538 7271
rect 19950 7209 19978 7238
rect 20510 7219 20538 7238
rect 20958 7266 20986 7631
rect 21406 7658 21434 7663
rect 19950 7183 19951 7209
rect 19977 7183 19978 7209
rect 19950 7177 19978 7183
rect 19573 7070 20035 7075
rect 19573 7069 19582 7070
rect 19573 7043 19574 7069
rect 19573 7042 19582 7043
rect 19610 7042 19634 7070
rect 19662 7042 19686 7070
rect 19714 7069 19738 7070
rect 19766 7069 19790 7070
rect 19724 7043 19738 7069
rect 19786 7043 19790 7069
rect 19714 7042 19738 7043
rect 19766 7042 19790 7043
rect 19818 7069 19842 7070
rect 19870 7069 19894 7070
rect 19818 7043 19822 7069
rect 19870 7043 19884 7069
rect 19818 7042 19842 7043
rect 19870 7042 19894 7043
rect 19922 7042 19946 7070
rect 19974 7042 19998 7070
rect 20026 7069 20035 7070
rect 20034 7043 20035 7069
rect 20026 7042 20035 7043
rect 19573 7037 20035 7042
rect 19110 6847 19111 6873
rect 19137 6847 19138 6873
rect 19054 6482 19082 6487
rect 19110 6482 19138 6847
rect 20006 6929 20034 6935
rect 20006 6903 20007 6929
rect 20033 6903 20034 6929
rect 20006 6874 20034 6903
rect 20958 6874 20986 7238
rect 20006 6873 20146 6874
rect 20006 6847 20007 6873
rect 20033 6847 20146 6873
rect 20006 6846 20146 6847
rect 20006 6841 20034 6846
rect 19054 6481 19138 6482
rect 19054 6455 19055 6481
rect 19081 6455 19138 6481
rect 19054 6454 19138 6455
rect 19054 6449 19082 6454
rect 18382 6425 18466 6426
rect 18382 6399 18383 6425
rect 18409 6399 18466 6425
rect 18382 6398 18466 6399
rect 18382 6393 18410 6398
rect 18438 6145 18466 6398
rect 18438 6119 18439 6145
rect 18465 6119 18466 6145
rect 18438 6089 18466 6119
rect 18438 6063 18439 6089
rect 18465 6063 18466 6089
rect 18382 5698 18410 5703
rect 18438 5698 18466 6063
rect 19110 6090 19138 6454
rect 19950 6481 19978 6487
rect 19950 6455 19951 6481
rect 19977 6455 19978 6481
rect 19950 6426 19978 6455
rect 20118 6426 20146 6846
rect 20958 6827 20986 6846
rect 21350 7265 21378 7271
rect 21350 7239 21351 7265
rect 21377 7239 21378 7265
rect 21350 7210 21378 7239
rect 19950 6425 20146 6426
rect 19950 6399 19951 6425
rect 19977 6399 20146 6425
rect 19950 6398 20146 6399
rect 19950 6393 19978 6398
rect 19573 6286 20035 6291
rect 19573 6285 19582 6286
rect 19573 6259 19574 6285
rect 19573 6258 19582 6259
rect 19610 6258 19634 6286
rect 19662 6258 19686 6286
rect 19714 6285 19738 6286
rect 19766 6285 19790 6286
rect 19724 6259 19738 6285
rect 19786 6259 19790 6285
rect 19714 6258 19738 6259
rect 19766 6258 19790 6259
rect 19818 6285 19842 6286
rect 19870 6285 19894 6286
rect 19818 6259 19822 6285
rect 19870 6259 19884 6285
rect 19818 6258 19842 6259
rect 19870 6258 19894 6259
rect 19922 6258 19946 6286
rect 19974 6258 19998 6286
rect 20026 6285 20035 6286
rect 20034 6259 20035 6285
rect 20026 6258 20035 6259
rect 19573 6253 20035 6258
rect 19110 6043 19138 6062
rect 20006 6145 20034 6151
rect 20006 6119 20007 6145
rect 20033 6119 20034 6145
rect 20006 6090 20034 6119
rect 20118 6090 20146 6398
rect 20006 6089 20146 6090
rect 20006 6063 20007 6089
rect 20033 6063 20146 6089
rect 20006 6062 20146 6063
rect 20006 6057 20034 6062
rect 18382 5697 18466 5698
rect 18382 5671 18383 5697
rect 18409 5671 18466 5697
rect 18382 5670 18466 5671
rect 18382 5641 18410 5670
rect 18382 5615 18383 5641
rect 18409 5615 18410 5641
rect 18382 5609 18410 5615
rect 18438 5361 18466 5670
rect 18438 5335 18439 5361
rect 18465 5335 18466 5361
rect 18438 5305 18466 5335
rect 18438 5279 18439 5305
rect 18465 5279 18466 5305
rect 18438 5194 18466 5279
rect 18438 5082 18466 5166
rect 18382 4914 18410 4919
rect 18438 4914 18466 5054
rect 18382 4913 18466 4914
rect 18382 4887 18383 4913
rect 18409 4887 18466 4913
rect 18382 4886 18466 4887
rect 18382 4857 18410 4886
rect 18382 4831 18383 4857
rect 18409 4831 18410 4857
rect 18382 4825 18410 4831
rect 18438 4577 18466 4886
rect 19054 5697 19082 5703
rect 19054 5671 19055 5697
rect 19081 5671 19082 5697
rect 19054 5305 19082 5671
rect 19950 5698 19978 5703
rect 20118 5698 20146 6062
rect 19950 5697 20146 5698
rect 19950 5671 19951 5697
rect 19977 5671 20146 5697
rect 19950 5670 20146 5671
rect 19950 5641 19978 5670
rect 19950 5615 19951 5641
rect 19977 5615 19978 5641
rect 19950 5609 19978 5615
rect 19573 5502 20035 5507
rect 19573 5501 19582 5502
rect 19573 5475 19574 5501
rect 19573 5474 19582 5475
rect 19610 5474 19634 5502
rect 19662 5474 19686 5502
rect 19714 5501 19738 5502
rect 19766 5501 19790 5502
rect 19724 5475 19738 5501
rect 19786 5475 19790 5501
rect 19714 5474 19738 5475
rect 19766 5474 19790 5475
rect 19818 5501 19842 5502
rect 19870 5501 19894 5502
rect 19818 5475 19822 5501
rect 19870 5475 19884 5501
rect 19818 5474 19842 5475
rect 19870 5474 19894 5475
rect 19922 5474 19946 5502
rect 19974 5474 19998 5502
rect 20026 5501 20035 5502
rect 20034 5475 20035 5501
rect 20026 5474 20035 5475
rect 19573 5469 20035 5474
rect 20006 5361 20034 5367
rect 20006 5335 20007 5361
rect 20033 5335 20034 5361
rect 20006 5306 20034 5335
rect 19054 5279 19055 5305
rect 19081 5279 19082 5305
rect 19054 4914 19082 5279
rect 19950 5278 20006 5306
rect 19950 5082 19978 5278
rect 20006 5259 20034 5278
rect 20118 5306 20146 5670
rect 19054 4913 19138 4914
rect 19054 4887 19055 4913
rect 19081 4887 19138 4913
rect 19054 4886 19138 4887
rect 19054 4881 19082 4886
rect 18438 4551 18439 4577
rect 18465 4551 18466 4577
rect 18438 4521 18466 4551
rect 18438 4495 18439 4521
rect 18465 4495 18466 4521
rect 18214 2977 18242 2982
rect 18382 4130 18410 4135
rect 18438 4130 18466 4495
rect 19110 4521 19138 4886
rect 19950 4913 19978 5054
rect 19950 4887 19951 4913
rect 19977 4887 19978 4913
rect 19950 4857 19978 4887
rect 19950 4831 19951 4857
rect 19977 4831 19978 4857
rect 19950 4825 19978 4831
rect 19573 4718 20035 4723
rect 19573 4717 19582 4718
rect 19573 4691 19574 4717
rect 19573 4690 19582 4691
rect 19610 4690 19634 4718
rect 19662 4690 19686 4718
rect 19714 4717 19738 4718
rect 19766 4717 19790 4718
rect 19724 4691 19738 4717
rect 19786 4691 19790 4717
rect 19714 4690 19738 4691
rect 19766 4690 19790 4691
rect 19818 4717 19842 4718
rect 19870 4717 19894 4718
rect 19818 4691 19822 4717
rect 19870 4691 19884 4717
rect 19818 4690 19842 4691
rect 19870 4690 19894 4691
rect 19922 4690 19946 4718
rect 19974 4690 19998 4718
rect 20026 4717 20035 4718
rect 20034 4691 20035 4717
rect 20026 4690 20035 4691
rect 19573 4685 20035 4690
rect 20118 4634 20146 5278
rect 19110 4495 19111 4521
rect 19137 4495 19138 4521
rect 18382 4129 18466 4130
rect 18382 4103 18383 4129
rect 18409 4103 18466 4129
rect 18382 4102 18466 4103
rect 19054 4130 19082 4135
rect 19110 4130 19138 4495
rect 20006 4606 20146 4634
rect 20006 4577 20034 4606
rect 20006 4551 20007 4577
rect 20033 4551 20034 4577
rect 20006 4521 20034 4551
rect 20006 4495 20007 4521
rect 20033 4495 20034 4521
rect 20006 4489 20034 4495
rect 19054 4129 19138 4130
rect 19054 4103 19055 4129
rect 19081 4103 19138 4129
rect 19054 4102 19138 4103
rect 18382 4073 18410 4102
rect 19054 4097 19082 4102
rect 18382 4047 18383 4073
rect 18409 4047 18410 4073
rect 18382 3793 18410 4047
rect 18382 3767 18383 3793
rect 18409 3767 18410 3793
rect 18382 3737 18410 3767
rect 18382 3711 18383 3737
rect 18409 3711 18410 3737
rect 18382 3345 18410 3711
rect 19110 3737 19138 4102
rect 19950 4130 19978 4135
rect 20118 4130 20146 4606
rect 19950 4129 20146 4130
rect 19950 4103 19951 4129
rect 19977 4103 20146 4129
rect 19950 4102 20146 4103
rect 19950 4073 19978 4102
rect 19950 4047 19951 4073
rect 19977 4047 19978 4073
rect 19950 4041 19978 4047
rect 19573 3934 20035 3939
rect 19573 3933 19582 3934
rect 19573 3907 19574 3933
rect 19573 3906 19582 3907
rect 19610 3906 19634 3934
rect 19662 3906 19686 3934
rect 19714 3933 19738 3934
rect 19766 3933 19790 3934
rect 19724 3907 19738 3933
rect 19786 3907 19790 3933
rect 19714 3906 19738 3907
rect 19766 3906 19790 3907
rect 19818 3933 19842 3934
rect 19870 3933 19894 3934
rect 19818 3907 19822 3933
rect 19870 3907 19884 3933
rect 19818 3906 19842 3907
rect 19870 3906 19894 3907
rect 19922 3906 19946 3934
rect 19974 3906 19998 3934
rect 20026 3933 20035 3934
rect 20034 3907 20035 3933
rect 20026 3906 20035 3907
rect 19573 3901 20035 3906
rect 19110 3711 19111 3737
rect 19137 3711 19138 3737
rect 19110 3402 19138 3711
rect 20006 3794 20034 3799
rect 20118 3794 20146 4102
rect 20006 3793 20146 3794
rect 20006 3767 20007 3793
rect 20033 3767 20146 3793
rect 20006 3766 20146 3767
rect 20510 6481 20538 6487
rect 20510 6455 20511 6481
rect 20537 6455 20538 6481
rect 20510 6090 20538 6455
rect 20790 6090 20818 6095
rect 20538 6089 20818 6090
rect 20538 6063 20791 6089
rect 20817 6063 20818 6089
rect 20538 6062 20818 6063
rect 20510 5697 20538 6062
rect 20790 6057 20818 6062
rect 20510 5671 20511 5697
rect 20537 5671 20538 5697
rect 20510 4913 20538 5671
rect 21350 5697 21378 7182
rect 21406 6481 21434 7630
rect 21798 7658 21826 7686
rect 21798 7592 21826 7630
rect 22526 7658 22554 7663
rect 22750 7658 22778 8023
rect 22526 7657 22778 7658
rect 22526 7631 22527 7657
rect 22553 7631 22778 7657
rect 22526 7630 22778 7631
rect 22526 7625 22554 7630
rect 22073 7462 22535 7467
rect 22073 7461 22082 7462
rect 22073 7435 22074 7461
rect 22073 7434 22082 7435
rect 22110 7434 22134 7462
rect 22162 7434 22186 7462
rect 22214 7461 22238 7462
rect 22266 7461 22290 7462
rect 22224 7435 22238 7461
rect 22286 7435 22290 7461
rect 22214 7434 22238 7435
rect 22266 7434 22290 7435
rect 22318 7461 22342 7462
rect 22370 7461 22394 7462
rect 22318 7435 22322 7461
rect 22370 7435 22384 7461
rect 22318 7434 22342 7435
rect 22370 7434 22394 7435
rect 22422 7434 22446 7462
rect 22474 7434 22498 7462
rect 22526 7461 22535 7462
rect 22534 7435 22535 7461
rect 22526 7434 22535 7435
rect 22073 7429 22535 7434
rect 22750 7266 22778 7630
rect 23422 8330 23450 8335
rect 23422 7713 23450 8302
rect 23422 7687 23423 7713
rect 23449 7687 23450 7713
rect 23422 7658 23450 7687
rect 23870 8049 23898 8055
rect 23870 8023 23871 8049
rect 23897 8023 23898 8049
rect 23870 7993 23898 8023
rect 23870 7967 23871 7993
rect 23897 7967 23898 7993
rect 23422 7657 23562 7658
rect 23422 7631 23423 7657
rect 23449 7631 23562 7657
rect 23422 7630 23562 7631
rect 23422 7625 23450 7630
rect 21742 7210 21770 7215
rect 22750 7200 22778 7238
rect 23534 7602 23562 7630
rect 23534 7266 23562 7574
rect 23870 7602 23898 7967
rect 23870 7569 23898 7574
rect 23534 7265 23730 7266
rect 23534 7239 23535 7265
rect 23561 7239 23730 7265
rect 23534 7238 23730 7239
rect 23534 7233 23562 7238
rect 23702 7209 23730 7238
rect 21742 6929 21770 7182
rect 23702 7183 23703 7209
rect 23729 7183 23730 7209
rect 23702 7177 23730 7183
rect 21742 6903 21743 6929
rect 21769 6903 21770 6929
rect 21742 6873 21770 6903
rect 23198 6929 23226 6935
rect 23198 6903 23199 6929
rect 23225 6903 23226 6929
rect 21742 6847 21743 6873
rect 21769 6847 21770 6873
rect 21742 6841 21770 6847
rect 22526 6874 22554 6879
rect 22554 6846 22610 6874
rect 22526 6808 22554 6846
rect 22073 6678 22535 6683
rect 22073 6677 22082 6678
rect 22073 6651 22074 6677
rect 22073 6650 22082 6651
rect 22110 6650 22134 6678
rect 22162 6650 22186 6678
rect 22214 6677 22238 6678
rect 22266 6677 22290 6678
rect 22224 6651 22238 6677
rect 22286 6651 22290 6677
rect 22214 6650 22238 6651
rect 22266 6650 22290 6651
rect 22318 6677 22342 6678
rect 22370 6677 22394 6678
rect 22318 6651 22322 6677
rect 22370 6651 22384 6677
rect 22318 6650 22342 6651
rect 22370 6650 22394 6651
rect 22422 6650 22446 6678
rect 22474 6650 22498 6678
rect 22526 6677 22535 6678
rect 22534 6651 22535 6677
rect 22526 6650 22535 6651
rect 22073 6645 22535 6650
rect 21406 6455 21407 6481
rect 21433 6455 21434 6481
rect 21406 6425 21434 6455
rect 21406 6399 21407 6425
rect 21433 6399 21434 6425
rect 21406 6146 21434 6399
rect 21798 6146 21826 6151
rect 21406 6145 21826 6146
rect 21406 6119 21799 6145
rect 21825 6119 21826 6145
rect 21406 6118 21826 6119
rect 21798 6089 21826 6118
rect 21798 6063 21799 6089
rect 21825 6063 21826 6089
rect 21798 5810 21826 6063
rect 22526 6090 22554 6095
rect 22582 6090 22610 6846
rect 23198 6873 23226 6903
rect 23198 6847 23199 6873
rect 23225 6847 23226 6873
rect 22526 6089 22610 6090
rect 22526 6063 22527 6089
rect 22553 6063 22610 6089
rect 22526 6062 22610 6063
rect 22526 6057 22554 6062
rect 22073 5894 22535 5899
rect 22073 5893 22082 5894
rect 22073 5867 22074 5893
rect 22073 5866 22082 5867
rect 22110 5866 22134 5894
rect 22162 5866 22186 5894
rect 22214 5893 22238 5894
rect 22266 5893 22290 5894
rect 22224 5867 22238 5893
rect 22286 5867 22290 5893
rect 22214 5866 22238 5867
rect 22266 5866 22290 5867
rect 22318 5893 22342 5894
rect 22370 5893 22394 5894
rect 22318 5867 22322 5893
rect 22370 5867 22384 5893
rect 22318 5866 22342 5867
rect 22370 5866 22394 5867
rect 22422 5866 22446 5894
rect 22474 5866 22498 5894
rect 22526 5893 22535 5894
rect 22534 5867 22535 5893
rect 22526 5866 22535 5867
rect 22073 5861 22535 5866
rect 21798 5777 21826 5782
rect 21854 5810 21882 5815
rect 21350 5671 21351 5697
rect 21377 5671 21378 5697
rect 21350 5641 21378 5671
rect 21350 5615 21351 5641
rect 21377 5615 21378 5641
rect 20510 4887 20511 4913
rect 20537 4887 20538 4913
rect 20510 4130 20538 4887
rect 20846 5305 20874 5311
rect 20846 5279 20847 5305
rect 20873 5279 20874 5305
rect 20846 4521 20874 5279
rect 21350 5306 21378 5615
rect 21462 5306 21490 5311
rect 21350 5305 21462 5306
rect 21350 5279 21351 5305
rect 21377 5279 21462 5305
rect 21350 5278 21462 5279
rect 21350 4913 21378 5278
rect 21462 5240 21490 5278
rect 21350 4887 21351 4913
rect 21377 4887 21378 4913
rect 21350 4857 21378 4887
rect 21350 4831 21351 4857
rect 21377 4831 21378 4857
rect 21350 4825 21378 4831
rect 20846 4495 20847 4521
rect 20873 4495 20874 4521
rect 20846 4214 20874 4495
rect 21350 4578 21378 4583
rect 20846 4186 20986 4214
rect 20006 3737 20034 3766
rect 20006 3711 20007 3737
rect 20033 3711 20034 3737
rect 20006 3705 20034 3711
rect 18382 3319 18383 3345
rect 18409 3319 18410 3345
rect 18382 3289 18410 3319
rect 19054 3346 19082 3351
rect 19110 3346 19138 3374
rect 20510 3402 20538 4102
rect 19054 3345 19138 3346
rect 19054 3319 19055 3345
rect 19081 3319 19138 3345
rect 19054 3318 19138 3319
rect 19054 3313 19082 3318
rect 18382 3263 18383 3289
rect 18409 3263 18410 3289
rect 18382 3009 18410 3263
rect 18382 2983 18383 3009
rect 18409 2983 18410 3009
rect 17598 2927 17599 2953
rect 17625 2927 17626 2953
rect 17073 2758 17535 2763
rect 17073 2757 17082 2758
rect 17073 2731 17074 2757
rect 17073 2730 17082 2731
rect 17110 2730 17134 2758
rect 17162 2730 17186 2758
rect 17214 2757 17238 2758
rect 17266 2757 17290 2758
rect 17224 2731 17238 2757
rect 17286 2731 17290 2757
rect 17214 2730 17238 2731
rect 17266 2730 17290 2731
rect 17318 2757 17342 2758
rect 17370 2757 17394 2758
rect 17318 2731 17322 2757
rect 17370 2731 17384 2757
rect 17318 2730 17342 2731
rect 17370 2730 17394 2731
rect 17422 2730 17446 2758
rect 17474 2730 17498 2758
rect 17526 2757 17535 2758
rect 17534 2731 17535 2757
rect 17526 2730 17535 2731
rect 17073 2725 17535 2730
rect 16254 2137 16282 2142
rect 15694 1731 15722 1750
rect 15526 1470 15666 1498
rect 15638 400 15666 1470
rect 16870 400 16898 2590
rect 17374 2561 17402 2567
rect 17374 2535 17375 2561
rect 17401 2535 17402 2561
rect 17374 2170 17402 2535
rect 17598 2170 17626 2927
rect 18382 2953 18410 2983
rect 18382 2927 18383 2953
rect 18409 2927 18410 2953
rect 18382 2921 18410 2927
rect 19110 2953 19138 3318
rect 19950 3345 19978 3351
rect 19950 3319 19951 3345
rect 19977 3319 19978 3345
rect 19950 3290 19978 3319
rect 20510 3345 20538 3374
rect 20510 3319 20511 3345
rect 20537 3319 20538 3345
rect 19950 3289 20146 3290
rect 19950 3263 19951 3289
rect 19977 3263 20146 3289
rect 19950 3262 20146 3263
rect 19950 3257 19978 3262
rect 19573 3150 20035 3155
rect 19573 3149 19582 3150
rect 19573 3123 19574 3149
rect 19573 3122 19582 3123
rect 19610 3122 19634 3150
rect 19662 3122 19686 3150
rect 19714 3149 19738 3150
rect 19766 3149 19790 3150
rect 19724 3123 19738 3149
rect 19786 3123 19790 3149
rect 19714 3122 19738 3123
rect 19766 3122 19790 3123
rect 19818 3149 19842 3150
rect 19870 3149 19894 3150
rect 19818 3123 19822 3149
rect 19870 3123 19884 3149
rect 19818 3122 19842 3123
rect 19870 3122 19894 3123
rect 19922 3122 19946 3150
rect 19974 3122 19998 3150
rect 20026 3149 20035 3150
rect 20034 3123 20035 3149
rect 20026 3122 20035 3123
rect 19573 3117 20035 3122
rect 19110 2927 19111 2953
rect 19137 2927 19138 2953
rect 18270 2562 18298 2567
rect 19054 2562 19082 2567
rect 19110 2562 19138 2927
rect 20006 3009 20034 3015
rect 20006 2983 20007 3009
rect 20033 2983 20034 3009
rect 20006 2954 20034 2983
rect 18270 2505 18298 2534
rect 18270 2479 18271 2505
rect 18297 2479 18298 2505
rect 17374 2169 17626 2170
rect 17374 2143 17375 2169
rect 17401 2143 17626 2169
rect 17374 2142 17626 2143
rect 17374 2137 17402 2142
rect 17073 1974 17535 1979
rect 17073 1973 17082 1974
rect 17073 1947 17074 1973
rect 17073 1946 17082 1947
rect 17110 1946 17134 1974
rect 17162 1946 17186 1974
rect 17214 1973 17238 1974
rect 17266 1973 17290 1974
rect 17224 1947 17238 1973
rect 17286 1947 17290 1973
rect 17214 1946 17238 1947
rect 17266 1946 17290 1947
rect 17318 1973 17342 1974
rect 17370 1973 17394 1974
rect 17318 1947 17322 1973
rect 17370 1947 17384 1973
rect 17318 1946 17342 1947
rect 17370 1946 17394 1947
rect 17422 1946 17446 1974
rect 17474 1946 17498 1974
rect 17526 1973 17535 1974
rect 17534 1947 17535 1973
rect 17526 1946 17535 1947
rect 17073 1941 17535 1946
rect 17262 1778 17290 1783
rect 17598 1778 17626 2142
rect 17262 1777 17626 1778
rect 17262 1751 17263 1777
rect 17289 1751 17626 1777
rect 17262 1750 17626 1751
rect 18102 2282 18130 2287
rect 17262 1745 17290 1750
rect 18102 1666 18130 2254
rect 18270 2225 18298 2479
rect 18270 2199 18271 2225
rect 18297 2199 18298 2225
rect 18270 2170 18298 2199
rect 18158 2169 18298 2170
rect 18158 2143 18271 2169
rect 18297 2143 18298 2169
rect 18158 2142 18298 2143
rect 18158 1777 18186 2142
rect 18270 2137 18298 2142
rect 18830 2561 19138 2562
rect 18830 2535 19055 2561
rect 19081 2535 19138 2561
rect 18830 2534 19138 2535
rect 19502 2562 19530 2567
rect 18830 2169 18858 2534
rect 19054 2529 19082 2534
rect 18830 2143 18831 2169
rect 18857 2143 18858 2169
rect 18158 1751 18159 1777
rect 18185 1751 18186 1777
rect 18158 1721 18186 1751
rect 18830 1777 18858 2143
rect 19502 2225 19530 2534
rect 19950 2562 19978 2567
rect 20006 2562 20034 2926
rect 20118 2954 20146 3262
rect 20118 2921 20146 2926
rect 19978 2534 20034 2562
rect 20510 2561 20538 3319
rect 20958 4130 20986 4186
rect 20958 3738 20986 4102
rect 20958 2953 20986 3710
rect 20958 2927 20959 2953
rect 20985 2927 20986 2953
rect 20958 2921 20986 2927
rect 21350 4129 21378 4550
rect 21798 4578 21826 4583
rect 21798 4521 21826 4550
rect 21798 4495 21799 4521
rect 21825 4495 21826 4521
rect 21798 4489 21826 4495
rect 21854 4522 21882 5782
rect 22526 5418 22554 5423
rect 22582 5418 22610 6062
rect 22554 5390 22610 5418
rect 23030 6481 23058 6487
rect 23030 6455 23031 6481
rect 23057 6455 23058 6481
rect 23030 5697 23058 6455
rect 23030 5671 23031 5697
rect 23057 5671 23058 5697
rect 23030 5418 23058 5671
rect 22526 5305 22554 5390
rect 22526 5279 22527 5305
rect 22553 5279 22554 5305
rect 22526 5273 22554 5279
rect 22073 5110 22535 5115
rect 22073 5109 22082 5110
rect 22073 5083 22074 5109
rect 22073 5082 22082 5083
rect 22110 5082 22134 5110
rect 22162 5082 22186 5110
rect 22214 5109 22238 5110
rect 22266 5109 22290 5110
rect 22224 5083 22238 5109
rect 22286 5083 22290 5109
rect 22214 5082 22238 5083
rect 22266 5082 22290 5083
rect 22318 5109 22342 5110
rect 22370 5109 22394 5110
rect 22318 5083 22322 5109
rect 22370 5083 22384 5109
rect 22318 5082 22342 5083
rect 22370 5082 22394 5083
rect 22422 5082 22446 5110
rect 22474 5082 22498 5110
rect 22526 5109 22535 5110
rect 22534 5083 22535 5109
rect 22526 5082 22535 5083
rect 22073 5077 22535 5082
rect 23030 4914 23058 5390
rect 22750 4913 23058 4914
rect 22750 4887 23031 4913
rect 23057 4887 23058 4913
rect 22750 4886 23058 4887
rect 21854 4489 21882 4494
rect 22526 4522 22554 4527
rect 22694 4522 22722 4527
rect 22526 4521 22610 4522
rect 22526 4495 22527 4521
rect 22553 4495 22610 4521
rect 22526 4494 22610 4495
rect 22526 4489 22554 4494
rect 22073 4326 22535 4331
rect 22073 4325 22082 4326
rect 22073 4299 22074 4325
rect 22073 4298 22082 4299
rect 22110 4298 22134 4326
rect 22162 4298 22186 4326
rect 22214 4325 22238 4326
rect 22266 4325 22290 4326
rect 22224 4299 22238 4325
rect 22286 4299 22290 4325
rect 22214 4298 22238 4299
rect 22266 4298 22290 4299
rect 22318 4325 22342 4326
rect 22370 4325 22394 4326
rect 22318 4299 22322 4325
rect 22370 4299 22384 4325
rect 22318 4298 22342 4299
rect 22370 4298 22394 4299
rect 22422 4298 22446 4326
rect 22474 4298 22498 4326
rect 22526 4325 22535 4326
rect 22534 4299 22535 4325
rect 22526 4298 22535 4299
rect 22073 4293 22535 4298
rect 22582 4214 22610 4494
rect 21350 4103 21351 4129
rect 21377 4103 21378 4129
rect 21350 4073 21378 4103
rect 21350 4047 21351 4073
rect 21377 4047 21378 4073
rect 21350 3738 21378 4047
rect 22526 4186 22610 4214
rect 21462 3738 21490 3743
rect 21350 3737 21490 3738
rect 21350 3711 21351 3737
rect 21377 3711 21463 3737
rect 21489 3711 21490 3737
rect 21350 3710 21490 3711
rect 21350 3345 21378 3710
rect 21462 3705 21490 3710
rect 22526 3738 22554 4186
rect 22526 3691 22554 3710
rect 22694 3737 22722 4494
rect 22694 3711 22695 3737
rect 22721 3711 22722 3737
rect 22694 3705 22722 3711
rect 22750 4129 22778 4886
rect 23030 4881 23058 4886
rect 23198 6482 23226 6847
rect 23198 4914 23226 6454
rect 23534 6482 23562 6487
rect 23534 6435 23562 6454
rect 23422 6145 23450 6151
rect 23422 6119 23423 6145
rect 23449 6119 23450 6145
rect 23422 6089 23450 6119
rect 23422 6063 23423 6089
rect 23449 6063 23450 6089
rect 23422 5810 23450 6063
rect 23422 5361 23450 5782
rect 23422 5335 23423 5361
rect 23449 5335 23450 5361
rect 23422 5306 23450 5335
rect 23422 5240 23450 5278
rect 23870 5810 23898 5815
rect 23870 5697 23898 5782
rect 23870 5671 23871 5697
rect 23897 5671 23898 5697
rect 23870 5641 23898 5671
rect 23870 5615 23871 5641
rect 23897 5615 23898 5641
rect 22750 4103 22751 4129
rect 22777 4103 22778 4129
rect 22073 3542 22535 3547
rect 22073 3541 22082 3542
rect 22073 3515 22074 3541
rect 22073 3514 22082 3515
rect 22110 3514 22134 3542
rect 22162 3514 22186 3542
rect 22214 3541 22238 3542
rect 22266 3541 22290 3542
rect 22224 3515 22238 3541
rect 22286 3515 22290 3541
rect 22214 3514 22238 3515
rect 22266 3514 22290 3515
rect 22318 3541 22342 3542
rect 22370 3541 22394 3542
rect 22318 3515 22322 3541
rect 22370 3515 22384 3541
rect 22318 3514 22342 3515
rect 22370 3514 22394 3515
rect 22422 3514 22446 3542
rect 22474 3514 22498 3542
rect 22526 3541 22535 3542
rect 22534 3515 22535 3541
rect 22526 3514 22535 3515
rect 22073 3509 22535 3514
rect 21350 3319 21351 3345
rect 21377 3319 21378 3345
rect 21350 3289 21378 3319
rect 21350 3263 21351 3289
rect 21377 3263 21378 3289
rect 21350 2954 21378 3263
rect 22750 3345 22778 4103
rect 22918 4522 22946 4527
rect 22918 3737 22946 4494
rect 23198 4522 23226 4886
rect 23198 4489 23226 4494
rect 23870 4913 23898 5615
rect 23870 4887 23871 4913
rect 23897 4887 23898 4913
rect 23870 4857 23898 4887
rect 23870 4831 23871 4857
rect 23897 4831 23898 4857
rect 23870 4129 23898 4831
rect 23870 4103 23871 4129
rect 23897 4103 23898 4129
rect 23870 4073 23898 4103
rect 23870 4047 23871 4073
rect 23897 4047 23898 4073
rect 22918 3711 22919 3737
rect 22945 3711 22946 3737
rect 22918 3705 22946 3711
rect 23030 3738 23058 3743
rect 22750 3319 22751 3345
rect 22777 3319 22778 3345
rect 21462 2954 21490 2959
rect 21378 2953 21490 2954
rect 21378 2927 21463 2953
rect 21489 2927 21490 2953
rect 21378 2926 21490 2927
rect 20510 2535 20511 2561
rect 20537 2535 20538 2561
rect 19950 2505 19978 2534
rect 20510 2529 20538 2535
rect 21350 2561 21378 2926
rect 21462 2921 21490 2926
rect 22526 2954 22554 2959
rect 22526 2953 22610 2954
rect 22526 2927 22527 2953
rect 22553 2927 22610 2953
rect 22526 2926 22610 2927
rect 22526 2921 22554 2926
rect 22073 2758 22535 2763
rect 22073 2757 22082 2758
rect 22073 2731 22074 2757
rect 22073 2730 22082 2731
rect 22110 2730 22134 2758
rect 22162 2730 22186 2758
rect 22214 2757 22238 2758
rect 22266 2757 22290 2758
rect 22224 2731 22238 2757
rect 22286 2731 22290 2757
rect 22214 2730 22238 2731
rect 22266 2730 22290 2731
rect 22318 2757 22342 2758
rect 22370 2757 22394 2758
rect 22318 2731 22322 2757
rect 22370 2731 22384 2757
rect 22318 2730 22342 2731
rect 22370 2730 22394 2731
rect 22422 2730 22446 2758
rect 22474 2730 22498 2758
rect 22526 2757 22535 2758
rect 22534 2731 22535 2757
rect 22526 2730 22535 2731
rect 22073 2725 22535 2730
rect 21350 2535 21351 2561
rect 21377 2535 21378 2561
rect 19950 2479 19951 2505
rect 19977 2479 19978 2505
rect 19950 2473 19978 2479
rect 21350 2505 21378 2535
rect 21350 2479 21351 2505
rect 21377 2479 21378 2505
rect 21350 2473 21378 2479
rect 21798 2562 21826 2567
rect 19573 2366 20035 2371
rect 19573 2365 19582 2366
rect 19573 2339 19574 2365
rect 19573 2338 19582 2339
rect 19610 2338 19634 2366
rect 19662 2338 19686 2366
rect 19714 2365 19738 2366
rect 19766 2365 19790 2366
rect 19724 2339 19738 2365
rect 19786 2339 19790 2365
rect 19714 2338 19738 2339
rect 19766 2338 19790 2339
rect 19818 2365 19842 2366
rect 19870 2365 19894 2366
rect 19818 2339 19822 2365
rect 19870 2339 19884 2365
rect 19818 2338 19842 2339
rect 19870 2338 19894 2339
rect 19922 2338 19946 2366
rect 19974 2338 19998 2366
rect 20026 2365 20035 2366
rect 20034 2339 20035 2365
rect 20026 2338 20035 2339
rect 19573 2333 20035 2338
rect 19502 2199 19503 2225
rect 19529 2199 19530 2225
rect 19502 2169 19530 2199
rect 21798 2225 21826 2534
rect 21798 2199 21799 2225
rect 21825 2199 21826 2225
rect 19502 2143 19503 2169
rect 19529 2143 19530 2169
rect 18830 1751 18831 1777
rect 18857 1751 18858 1777
rect 18830 1745 18858 1751
rect 19334 2058 19362 2063
rect 18158 1695 18159 1721
rect 18185 1695 18186 1721
rect 18158 1689 18186 1695
rect 19334 1722 19362 2030
rect 18102 400 18130 1638
rect 19334 400 19362 1694
rect 19502 1777 19530 2143
rect 20790 2169 20818 2175
rect 20790 2143 20791 2169
rect 20817 2143 20818 2169
rect 19502 1751 19503 1777
rect 19529 1751 19530 1777
rect 19502 1721 19530 1751
rect 20510 2114 20538 2119
rect 20510 1777 20538 2086
rect 20790 2114 20818 2143
rect 21798 2169 21826 2199
rect 22582 2562 22610 2926
rect 22750 2562 22778 3319
rect 22582 2561 22778 2562
rect 22582 2535 22751 2561
rect 22777 2535 22778 2561
rect 22582 2534 22778 2535
rect 21798 2143 21799 2169
rect 21825 2143 21826 2169
rect 20790 2081 20818 2086
rect 21630 2114 21658 2119
rect 20510 1751 20511 1777
rect 20537 1751 20538 1777
rect 20510 1745 20538 1751
rect 20566 1834 20594 1839
rect 19502 1695 19503 1721
rect 19529 1695 19530 1721
rect 19502 1689 19530 1695
rect 19573 1582 20035 1587
rect 19573 1581 19582 1582
rect 19573 1555 19574 1581
rect 19573 1554 19582 1555
rect 19610 1554 19634 1582
rect 19662 1554 19686 1582
rect 19714 1581 19738 1582
rect 19766 1581 19790 1582
rect 19724 1555 19738 1581
rect 19786 1555 19790 1581
rect 19714 1554 19738 1555
rect 19766 1554 19790 1555
rect 19818 1581 19842 1582
rect 19870 1581 19894 1582
rect 19818 1555 19822 1581
rect 19870 1555 19884 1581
rect 19818 1554 19842 1555
rect 19870 1554 19894 1555
rect 19922 1554 19946 1582
rect 19974 1554 19998 1582
rect 20026 1581 20035 1582
rect 20034 1555 20035 1581
rect 20026 1554 20035 1555
rect 19573 1549 20035 1554
rect 20566 400 20594 1806
rect 21630 1610 21658 2086
rect 21686 1778 21714 1783
rect 21798 1778 21826 2143
rect 22246 2169 22274 2175
rect 22246 2143 22247 2169
rect 22273 2143 22274 2169
rect 22246 2114 22274 2143
rect 22246 2081 22274 2086
rect 22582 2114 22610 2534
rect 22750 2529 22778 2534
rect 22582 2081 22610 2086
rect 22073 1974 22535 1979
rect 22073 1973 22082 1974
rect 22073 1947 22074 1973
rect 22073 1946 22082 1947
rect 22110 1946 22134 1974
rect 22162 1946 22186 1974
rect 22214 1973 22238 1974
rect 22266 1973 22290 1974
rect 22224 1947 22238 1973
rect 22286 1947 22290 1973
rect 22214 1946 22238 1947
rect 22266 1946 22290 1947
rect 22318 1973 22342 1974
rect 22370 1973 22394 1974
rect 22318 1947 22322 1973
rect 22370 1947 22384 1973
rect 22318 1946 22342 1947
rect 22370 1946 22394 1947
rect 22422 1946 22446 1974
rect 22474 1946 22498 1974
rect 22526 1973 22535 1974
rect 22534 1947 22535 1973
rect 22526 1946 22535 1947
rect 22073 1941 22535 1946
rect 21686 1777 21826 1778
rect 21686 1751 21687 1777
rect 21713 1751 21826 1777
rect 21686 1750 21826 1751
rect 22470 1834 22498 1839
rect 22470 1777 22498 1806
rect 22470 1751 22471 1777
rect 22497 1751 22498 1777
rect 21686 1721 21714 1750
rect 22470 1745 22498 1751
rect 21686 1695 21687 1721
rect 21713 1695 21714 1721
rect 21686 1689 21714 1695
rect 21630 1582 21826 1610
rect 21798 400 21826 1582
rect 23030 400 23058 3710
rect 23870 3458 23898 4047
rect 23870 3345 23898 3430
rect 23870 3319 23871 3345
rect 23897 3319 23898 3345
rect 23870 3289 23898 3319
rect 23870 3263 23871 3289
rect 23897 3263 23898 3289
rect 23422 3009 23450 3015
rect 23422 2983 23423 3009
rect 23449 2983 23450 3009
rect 23422 2953 23450 2983
rect 23422 2927 23423 2953
rect 23449 2927 23450 2953
rect 23422 2562 23450 2927
rect 23422 2225 23450 2534
rect 23870 2561 23898 3263
rect 23926 2618 23954 17318
rect 24573 17262 25035 17267
rect 24573 17261 24582 17262
rect 24573 17235 24574 17261
rect 24573 17234 24582 17235
rect 24610 17234 24634 17262
rect 24662 17234 24686 17262
rect 24714 17261 24738 17262
rect 24766 17261 24790 17262
rect 24724 17235 24738 17261
rect 24786 17235 24790 17261
rect 24714 17234 24738 17235
rect 24766 17234 24790 17235
rect 24818 17261 24842 17262
rect 24870 17261 24894 17262
rect 24818 17235 24822 17261
rect 24870 17235 24884 17261
rect 24818 17234 24842 17235
rect 24870 17234 24894 17235
rect 24922 17234 24946 17262
rect 24974 17234 24998 17262
rect 25026 17261 25035 17262
rect 25034 17235 25035 17261
rect 25026 17234 25035 17235
rect 24573 17229 25035 17234
rect 24573 16478 25035 16483
rect 24573 16477 24582 16478
rect 24573 16451 24574 16477
rect 24573 16450 24582 16451
rect 24610 16450 24634 16478
rect 24662 16450 24686 16478
rect 24714 16477 24738 16478
rect 24766 16477 24790 16478
rect 24724 16451 24738 16477
rect 24786 16451 24790 16477
rect 24714 16450 24738 16451
rect 24766 16450 24790 16451
rect 24818 16477 24842 16478
rect 24870 16477 24894 16478
rect 24818 16451 24822 16477
rect 24870 16451 24884 16477
rect 24818 16450 24842 16451
rect 24870 16450 24894 16451
rect 24922 16450 24946 16478
rect 24974 16450 24998 16478
rect 25026 16477 25035 16478
rect 25034 16451 25035 16477
rect 25026 16450 25035 16451
rect 24573 16445 25035 16450
rect 24573 15694 25035 15699
rect 24573 15693 24582 15694
rect 24573 15667 24574 15693
rect 24573 15666 24582 15667
rect 24610 15666 24634 15694
rect 24662 15666 24686 15694
rect 24714 15693 24738 15694
rect 24766 15693 24790 15694
rect 24724 15667 24738 15693
rect 24786 15667 24790 15693
rect 24714 15666 24738 15667
rect 24766 15666 24790 15667
rect 24818 15693 24842 15694
rect 24870 15693 24894 15694
rect 24818 15667 24822 15693
rect 24870 15667 24884 15693
rect 24818 15666 24842 15667
rect 24870 15666 24894 15667
rect 24922 15666 24946 15694
rect 24974 15666 24998 15694
rect 25026 15693 25035 15694
rect 25034 15667 25035 15693
rect 25026 15666 25035 15667
rect 24573 15661 25035 15666
rect 24486 15162 24514 15167
rect 24430 14321 24458 14327
rect 24430 14295 24431 14321
rect 24457 14295 24458 14321
rect 24430 13537 24458 14295
rect 24430 13511 24431 13537
rect 24457 13511 24458 13537
rect 24430 13482 24458 13511
rect 24374 13426 24458 13454
rect 24374 12362 24402 13426
rect 24430 13416 24458 13426
rect 24486 13426 24514 15134
rect 26894 15162 26922 19614
rect 27286 19530 27314 19614
rect 27440 19600 27496 20000
rect 31934 19614 32298 19642
rect 27454 19530 27482 19600
rect 27286 19502 27482 19530
rect 27073 18438 27535 18443
rect 27073 18437 27082 18438
rect 27073 18411 27074 18437
rect 27073 18410 27082 18411
rect 27110 18410 27134 18438
rect 27162 18410 27186 18438
rect 27214 18437 27238 18438
rect 27266 18437 27290 18438
rect 27224 18411 27238 18437
rect 27286 18411 27290 18437
rect 27214 18410 27238 18411
rect 27266 18410 27290 18411
rect 27318 18437 27342 18438
rect 27370 18437 27394 18438
rect 27318 18411 27322 18437
rect 27370 18411 27384 18437
rect 27318 18410 27342 18411
rect 27370 18410 27394 18411
rect 27422 18410 27446 18438
rect 27474 18410 27498 18438
rect 27526 18437 27535 18438
rect 27534 18411 27535 18437
rect 27526 18410 27535 18411
rect 27073 18405 27535 18410
rect 29573 18046 30035 18051
rect 29573 18045 29582 18046
rect 29573 18019 29574 18045
rect 29573 18018 29582 18019
rect 29610 18018 29634 18046
rect 29662 18018 29686 18046
rect 29714 18045 29738 18046
rect 29766 18045 29790 18046
rect 29724 18019 29738 18045
rect 29786 18019 29790 18045
rect 29714 18018 29738 18019
rect 29766 18018 29790 18019
rect 29818 18045 29842 18046
rect 29870 18045 29894 18046
rect 29818 18019 29822 18045
rect 29870 18019 29884 18045
rect 29818 18018 29842 18019
rect 29870 18018 29894 18019
rect 29922 18018 29946 18046
rect 29974 18018 29998 18046
rect 30026 18045 30035 18046
rect 30034 18019 30035 18045
rect 30026 18018 30035 18019
rect 29573 18013 30035 18018
rect 27073 17654 27535 17659
rect 27073 17653 27082 17654
rect 27073 17627 27074 17653
rect 27073 17626 27082 17627
rect 27110 17626 27134 17654
rect 27162 17626 27186 17654
rect 27214 17653 27238 17654
rect 27266 17653 27290 17654
rect 27224 17627 27238 17653
rect 27286 17627 27290 17653
rect 27214 17626 27238 17627
rect 27266 17626 27290 17627
rect 27318 17653 27342 17654
rect 27370 17653 27394 17654
rect 27318 17627 27322 17653
rect 27370 17627 27384 17653
rect 27318 17626 27342 17627
rect 27370 17626 27394 17627
rect 27422 17626 27446 17654
rect 27474 17626 27498 17654
rect 27526 17653 27535 17654
rect 27534 17627 27535 17653
rect 27526 17626 27535 17627
rect 27073 17621 27535 17626
rect 29573 17262 30035 17267
rect 29573 17261 29582 17262
rect 29573 17235 29574 17261
rect 29573 17234 29582 17235
rect 29610 17234 29634 17262
rect 29662 17234 29686 17262
rect 29714 17261 29738 17262
rect 29766 17261 29790 17262
rect 29724 17235 29738 17261
rect 29786 17235 29790 17261
rect 29714 17234 29738 17235
rect 29766 17234 29790 17235
rect 29818 17261 29842 17262
rect 29870 17261 29894 17262
rect 29818 17235 29822 17261
rect 29870 17235 29884 17261
rect 29818 17234 29842 17235
rect 29870 17234 29894 17235
rect 29922 17234 29946 17262
rect 29974 17234 29998 17262
rect 30026 17261 30035 17262
rect 30034 17235 30035 17261
rect 30026 17234 30035 17235
rect 29573 17229 30035 17234
rect 27073 16870 27535 16875
rect 27073 16869 27082 16870
rect 27073 16843 27074 16869
rect 27073 16842 27082 16843
rect 27110 16842 27134 16870
rect 27162 16842 27186 16870
rect 27214 16869 27238 16870
rect 27266 16869 27290 16870
rect 27224 16843 27238 16869
rect 27286 16843 27290 16869
rect 27214 16842 27238 16843
rect 27266 16842 27290 16843
rect 27318 16869 27342 16870
rect 27370 16869 27394 16870
rect 27318 16843 27322 16869
rect 27370 16843 27384 16869
rect 27318 16842 27342 16843
rect 27370 16842 27394 16843
rect 27422 16842 27446 16870
rect 27474 16842 27498 16870
rect 27526 16869 27535 16870
rect 27534 16843 27535 16869
rect 27526 16842 27535 16843
rect 27073 16837 27535 16842
rect 29573 16478 30035 16483
rect 29573 16477 29582 16478
rect 29573 16451 29574 16477
rect 29573 16450 29582 16451
rect 29610 16450 29634 16478
rect 29662 16450 29686 16478
rect 29714 16477 29738 16478
rect 29766 16477 29790 16478
rect 29724 16451 29738 16477
rect 29786 16451 29790 16477
rect 29714 16450 29738 16451
rect 29766 16450 29790 16451
rect 29818 16477 29842 16478
rect 29870 16477 29894 16478
rect 29818 16451 29822 16477
rect 29870 16451 29884 16477
rect 29818 16450 29842 16451
rect 29870 16450 29894 16451
rect 29922 16450 29946 16478
rect 29974 16450 29998 16478
rect 30026 16477 30035 16478
rect 30034 16451 30035 16477
rect 30026 16450 30035 16451
rect 29573 16445 30035 16450
rect 27073 16086 27535 16091
rect 27073 16085 27082 16086
rect 27073 16059 27074 16085
rect 27073 16058 27082 16059
rect 27110 16058 27134 16086
rect 27162 16058 27186 16086
rect 27214 16085 27238 16086
rect 27266 16085 27290 16086
rect 27224 16059 27238 16085
rect 27286 16059 27290 16085
rect 27214 16058 27238 16059
rect 27266 16058 27290 16059
rect 27318 16085 27342 16086
rect 27370 16085 27394 16086
rect 27318 16059 27322 16085
rect 27370 16059 27384 16085
rect 27318 16058 27342 16059
rect 27370 16058 27394 16059
rect 27422 16058 27446 16086
rect 27474 16058 27498 16086
rect 27526 16085 27535 16086
rect 27534 16059 27535 16085
rect 27526 16058 27535 16059
rect 27073 16053 27535 16058
rect 29573 15694 30035 15699
rect 29573 15693 29582 15694
rect 29573 15667 29574 15693
rect 29573 15666 29582 15667
rect 29610 15666 29634 15694
rect 29662 15666 29686 15694
rect 29714 15693 29738 15694
rect 29766 15693 29790 15694
rect 29724 15667 29738 15693
rect 29786 15667 29790 15693
rect 29714 15666 29738 15667
rect 29766 15666 29790 15667
rect 29818 15693 29842 15694
rect 29870 15693 29894 15694
rect 29818 15667 29822 15693
rect 29870 15667 29884 15693
rect 29818 15666 29842 15667
rect 29870 15666 29894 15667
rect 29922 15666 29946 15694
rect 29974 15666 29998 15694
rect 30026 15693 30035 15694
rect 30034 15667 30035 15693
rect 30026 15666 30035 15667
rect 29573 15661 30035 15666
rect 27073 15302 27535 15307
rect 27073 15301 27082 15302
rect 27073 15275 27074 15301
rect 27073 15274 27082 15275
rect 27110 15274 27134 15302
rect 27162 15274 27186 15302
rect 27214 15301 27238 15302
rect 27266 15301 27290 15302
rect 27224 15275 27238 15301
rect 27286 15275 27290 15301
rect 27214 15274 27238 15275
rect 27266 15274 27290 15275
rect 27318 15301 27342 15302
rect 27370 15301 27394 15302
rect 27318 15275 27322 15301
rect 27370 15275 27384 15301
rect 27318 15274 27342 15275
rect 27370 15274 27394 15275
rect 27422 15274 27446 15302
rect 27474 15274 27498 15302
rect 27526 15301 27535 15302
rect 27534 15275 27535 15301
rect 27526 15274 27535 15275
rect 27073 15269 27535 15274
rect 26894 15129 26922 15134
rect 24573 14910 25035 14915
rect 24573 14909 24582 14910
rect 24573 14883 24574 14909
rect 24573 14882 24582 14883
rect 24610 14882 24634 14910
rect 24662 14882 24686 14910
rect 24714 14909 24738 14910
rect 24766 14909 24790 14910
rect 24724 14883 24738 14909
rect 24786 14883 24790 14909
rect 24714 14882 24738 14883
rect 24766 14882 24790 14883
rect 24818 14909 24842 14910
rect 24870 14909 24894 14910
rect 24818 14883 24822 14909
rect 24870 14883 24884 14909
rect 24818 14882 24842 14883
rect 24870 14882 24894 14883
rect 24922 14882 24946 14910
rect 24974 14882 24998 14910
rect 25026 14909 25035 14910
rect 25034 14883 25035 14909
rect 25026 14882 25035 14883
rect 24573 14877 25035 14882
rect 29573 14910 30035 14915
rect 29573 14909 29582 14910
rect 29573 14883 29574 14909
rect 29573 14882 29582 14883
rect 29610 14882 29634 14910
rect 29662 14882 29686 14910
rect 29714 14909 29738 14910
rect 29766 14909 29790 14910
rect 29724 14883 29738 14909
rect 29786 14883 29790 14909
rect 29714 14882 29738 14883
rect 29766 14882 29790 14883
rect 29818 14909 29842 14910
rect 29870 14909 29894 14910
rect 29818 14883 29822 14909
rect 29870 14883 29884 14909
rect 29818 14882 29842 14883
rect 29870 14882 29894 14883
rect 29922 14882 29946 14910
rect 29974 14882 29998 14910
rect 30026 14909 30035 14910
rect 30034 14883 30035 14909
rect 30026 14882 30035 14883
rect 29573 14877 30035 14882
rect 27073 14518 27535 14523
rect 27073 14517 27082 14518
rect 27073 14491 27074 14517
rect 27073 14490 27082 14491
rect 27110 14490 27134 14518
rect 27162 14490 27186 14518
rect 27214 14517 27238 14518
rect 27266 14517 27290 14518
rect 27224 14491 27238 14517
rect 27286 14491 27290 14517
rect 27214 14490 27238 14491
rect 27266 14490 27290 14491
rect 27318 14517 27342 14518
rect 27370 14517 27394 14518
rect 27318 14491 27322 14517
rect 27370 14491 27384 14517
rect 27318 14490 27342 14491
rect 27370 14490 27394 14491
rect 27422 14490 27446 14518
rect 27474 14490 27498 14518
rect 27526 14517 27535 14518
rect 27534 14491 27535 14517
rect 27526 14490 27535 14491
rect 27073 14485 27535 14490
rect 25158 14321 25186 14327
rect 25158 14295 25159 14321
rect 25185 14295 25186 14321
rect 25158 14266 25186 14295
rect 25214 14266 25242 14271
rect 25186 14265 25242 14266
rect 25186 14239 25215 14265
rect 25241 14239 25242 14265
rect 25186 14238 25242 14239
rect 25158 14200 25186 14238
rect 24573 14126 25035 14131
rect 24573 14125 24582 14126
rect 24573 14099 24574 14125
rect 24573 14098 24582 14099
rect 24610 14098 24634 14126
rect 24662 14098 24686 14126
rect 24714 14125 24738 14126
rect 24766 14125 24790 14126
rect 24724 14099 24738 14125
rect 24786 14099 24790 14125
rect 24714 14098 24738 14099
rect 24766 14098 24790 14099
rect 24818 14125 24842 14126
rect 24870 14125 24894 14126
rect 24818 14099 24822 14125
rect 24870 14099 24884 14125
rect 24818 14098 24842 14099
rect 24870 14098 24894 14099
rect 24922 14098 24946 14126
rect 24974 14098 24998 14126
rect 25026 14125 25035 14126
rect 25034 14099 25035 14125
rect 25026 14098 25035 14099
rect 24573 14093 25035 14098
rect 25046 13930 25074 13935
rect 25214 13930 25242 14238
rect 29573 14126 30035 14131
rect 29573 14125 29582 14126
rect 29573 14099 29574 14125
rect 29573 14098 29582 14099
rect 29610 14098 29634 14126
rect 29662 14098 29686 14126
rect 29714 14125 29738 14126
rect 29766 14125 29790 14126
rect 29724 14099 29738 14125
rect 29786 14099 29790 14125
rect 29714 14098 29738 14099
rect 29766 14098 29790 14099
rect 29818 14125 29842 14126
rect 29870 14125 29894 14126
rect 29818 14099 29822 14125
rect 29870 14099 29884 14125
rect 29818 14098 29842 14099
rect 29870 14098 29894 14099
rect 29922 14098 29946 14126
rect 29974 14098 29998 14126
rect 30026 14125 30035 14126
rect 30034 14099 30035 14125
rect 30026 14098 30035 14099
rect 29573 14093 30035 14098
rect 25438 13930 25466 13935
rect 25046 13929 25130 13930
rect 25046 13903 25047 13929
rect 25073 13903 25130 13929
rect 25046 13902 25130 13903
rect 25046 13897 25074 13902
rect 24486 13393 24514 13398
rect 24573 13342 25035 13347
rect 24573 13341 24582 13342
rect 24374 12329 24402 12334
rect 24430 13314 24458 13319
rect 24573 13315 24574 13341
rect 24573 13314 24582 13315
rect 24610 13314 24634 13342
rect 24662 13314 24686 13342
rect 24714 13341 24738 13342
rect 24766 13341 24790 13342
rect 24724 13315 24738 13341
rect 24786 13315 24790 13341
rect 24714 13314 24738 13315
rect 24766 13314 24790 13315
rect 24818 13341 24842 13342
rect 24870 13341 24894 13342
rect 24818 13315 24822 13341
rect 24870 13315 24884 13341
rect 24818 13314 24842 13315
rect 24870 13314 24894 13315
rect 24922 13314 24946 13342
rect 24974 13314 24998 13342
rect 25026 13341 25035 13342
rect 25034 13315 25035 13341
rect 25026 13314 25035 13315
rect 24573 13309 25035 13314
rect 24374 11185 24402 11191
rect 24374 11159 24375 11185
rect 24401 11159 24402 11185
rect 24374 10401 24402 11159
rect 24430 10626 24458 13286
rect 25046 13146 25074 13151
rect 25102 13146 25130 13902
rect 25046 13145 25130 13146
rect 25046 13119 25047 13145
rect 25073 13119 25130 13145
rect 25046 13118 25130 13119
rect 25046 13113 25074 13118
rect 24486 12753 24514 12759
rect 24486 12727 24487 12753
rect 24513 12727 24514 12753
rect 24486 12362 24514 12727
rect 24573 12558 25035 12563
rect 24573 12557 24582 12558
rect 24573 12531 24574 12557
rect 24573 12530 24582 12531
rect 24610 12530 24634 12558
rect 24662 12530 24686 12558
rect 24714 12557 24738 12558
rect 24766 12557 24790 12558
rect 24724 12531 24738 12557
rect 24786 12531 24790 12557
rect 24714 12530 24738 12531
rect 24766 12530 24790 12531
rect 24818 12557 24842 12558
rect 24870 12557 24894 12558
rect 24818 12531 24822 12557
rect 24870 12531 24884 12557
rect 24818 12530 24842 12531
rect 24870 12530 24894 12531
rect 24922 12530 24946 12558
rect 24974 12530 24998 12558
rect 25026 12557 25035 12558
rect 25034 12531 25035 12557
rect 25026 12530 25035 12531
rect 24573 12525 25035 12530
rect 24486 11969 24514 12334
rect 24766 12362 24794 12367
rect 24766 12315 24794 12334
rect 25102 12362 25130 13118
rect 25214 13929 25466 13930
rect 25214 13903 25215 13929
rect 25241 13903 25439 13929
rect 25465 13903 25466 13929
rect 25214 13902 25466 13903
rect 25214 13537 25242 13902
rect 25438 13897 25466 13902
rect 27073 13734 27535 13739
rect 27073 13733 27082 13734
rect 27073 13707 27074 13733
rect 27073 13706 27082 13707
rect 27110 13706 27134 13734
rect 27162 13706 27186 13734
rect 27214 13733 27238 13734
rect 27266 13733 27290 13734
rect 27224 13707 27238 13733
rect 27286 13707 27290 13733
rect 27214 13706 27238 13707
rect 27266 13706 27290 13707
rect 27318 13733 27342 13734
rect 27370 13733 27394 13734
rect 27318 13707 27322 13733
rect 27370 13707 27384 13733
rect 27318 13706 27342 13707
rect 27370 13706 27394 13707
rect 27422 13706 27446 13734
rect 27474 13706 27498 13734
rect 27526 13733 27535 13734
rect 27534 13707 27535 13733
rect 27526 13706 27535 13707
rect 27073 13701 27535 13706
rect 25214 13511 25215 13537
rect 25241 13511 25242 13537
rect 25214 13481 25242 13511
rect 25214 13455 25215 13481
rect 25241 13455 25242 13481
rect 25102 12329 25130 12334
rect 25158 12753 25186 12759
rect 25158 12727 25159 12753
rect 25185 12727 25186 12753
rect 25158 12698 25186 12727
rect 24486 11943 24487 11969
rect 24513 11943 24514 11969
rect 24486 11578 24514 11943
rect 25102 11970 25130 11975
rect 24573 11774 25035 11779
rect 24573 11773 24582 11774
rect 24573 11747 24574 11773
rect 24573 11746 24582 11747
rect 24610 11746 24634 11774
rect 24662 11746 24686 11774
rect 24714 11773 24738 11774
rect 24766 11773 24790 11774
rect 24724 11747 24738 11773
rect 24786 11747 24790 11773
rect 24714 11746 24738 11747
rect 24766 11746 24790 11747
rect 24818 11773 24842 11774
rect 24870 11773 24894 11774
rect 24818 11747 24822 11773
rect 24870 11747 24884 11773
rect 24818 11746 24842 11747
rect 24870 11746 24894 11747
rect 24922 11746 24946 11774
rect 24974 11746 24998 11774
rect 25026 11773 25035 11774
rect 25034 11747 25035 11773
rect 25026 11746 25035 11747
rect 24573 11741 25035 11746
rect 24766 11578 24794 11583
rect 24486 11577 24794 11578
rect 24486 11551 24767 11577
rect 24793 11551 24794 11577
rect 24486 11550 24794 11551
rect 24766 11545 24794 11550
rect 24573 10990 25035 10995
rect 24573 10989 24582 10990
rect 24573 10963 24574 10989
rect 24573 10962 24582 10963
rect 24610 10962 24634 10990
rect 24662 10962 24686 10990
rect 24714 10989 24738 10990
rect 24766 10989 24790 10990
rect 24724 10963 24738 10989
rect 24786 10963 24790 10989
rect 24714 10962 24738 10963
rect 24766 10962 24790 10963
rect 24818 10989 24842 10990
rect 24870 10989 24894 10990
rect 24818 10963 24822 10989
rect 24870 10963 24884 10989
rect 24818 10962 24842 10963
rect 24870 10962 24894 10963
rect 24922 10962 24946 10990
rect 24974 10962 24998 10990
rect 25026 10989 25035 10990
rect 25034 10963 25035 10989
rect 25026 10962 25035 10963
rect 24573 10957 25035 10962
rect 25046 10794 25074 10799
rect 25102 10794 25130 11942
rect 25158 11969 25186 12670
rect 25214 12250 25242 13455
rect 29573 13342 30035 13347
rect 29573 13341 29582 13342
rect 29573 13315 29574 13341
rect 29573 13314 29582 13315
rect 29610 13314 29634 13342
rect 29662 13314 29686 13342
rect 29714 13341 29738 13342
rect 29766 13341 29790 13342
rect 29724 13315 29738 13341
rect 29786 13315 29790 13341
rect 29714 13314 29738 13315
rect 29766 13314 29790 13315
rect 29818 13341 29842 13342
rect 29870 13341 29894 13342
rect 29818 13315 29822 13341
rect 29870 13315 29884 13341
rect 29818 13314 29842 13315
rect 29870 13314 29894 13315
rect 29922 13314 29946 13342
rect 29974 13314 29998 13342
rect 30026 13341 30035 13342
rect 30034 13315 30035 13341
rect 30026 13314 30035 13315
rect 29573 13309 30035 13314
rect 25214 12217 25242 12222
rect 25942 13201 25970 13207
rect 25942 13175 25943 13201
rect 25969 13175 25970 13201
rect 25942 13145 25970 13175
rect 25942 13119 25943 13145
rect 25969 13119 25970 13145
rect 25942 12418 25970 13119
rect 27073 12950 27535 12955
rect 27073 12949 27082 12950
rect 27073 12923 27074 12949
rect 27073 12922 27082 12923
rect 27110 12922 27134 12950
rect 27162 12922 27186 12950
rect 27214 12949 27238 12950
rect 27266 12949 27290 12950
rect 27224 12923 27238 12949
rect 27286 12923 27290 12949
rect 27214 12922 27238 12923
rect 27266 12922 27290 12923
rect 27318 12949 27342 12950
rect 27370 12949 27394 12950
rect 27318 12923 27322 12949
rect 27370 12923 27384 12949
rect 27318 12922 27342 12923
rect 27370 12922 27394 12923
rect 27422 12922 27446 12950
rect 27474 12922 27498 12950
rect 27526 12949 27535 12950
rect 27534 12923 27535 12949
rect 27526 12922 27535 12923
rect 27073 12917 27535 12922
rect 29638 12754 29666 12759
rect 29750 12754 29778 12759
rect 29414 12753 29778 12754
rect 29414 12727 29639 12753
rect 29665 12727 29751 12753
rect 29777 12727 29778 12753
rect 29414 12726 29778 12727
rect 25942 12361 25970 12390
rect 27398 12417 27426 12423
rect 27398 12391 27399 12417
rect 27425 12391 27426 12417
rect 25942 12335 25943 12361
rect 25969 12335 25970 12361
rect 25942 12250 25970 12335
rect 26502 12362 26530 12367
rect 27398 12362 27426 12391
rect 26530 12334 26754 12362
rect 26502 12296 26530 12334
rect 25942 12217 25970 12222
rect 25158 11943 25159 11969
rect 25185 11943 25186 11969
rect 25158 11913 25186 11943
rect 26726 11969 26754 12334
rect 27398 12315 27426 12334
rect 27678 12362 27706 12367
rect 27073 12166 27535 12171
rect 27073 12165 27082 12166
rect 27073 12139 27074 12165
rect 27073 12138 27082 12139
rect 27110 12138 27134 12166
rect 27162 12138 27186 12166
rect 27214 12165 27238 12166
rect 27266 12165 27290 12166
rect 27224 12139 27238 12165
rect 27286 12139 27290 12165
rect 27214 12138 27238 12139
rect 27266 12138 27290 12139
rect 27318 12165 27342 12166
rect 27370 12165 27394 12166
rect 27318 12139 27322 12165
rect 27370 12139 27384 12165
rect 27318 12138 27342 12139
rect 27370 12138 27394 12139
rect 27422 12138 27446 12166
rect 27474 12138 27498 12166
rect 27526 12165 27535 12166
rect 27534 12139 27535 12165
rect 27526 12138 27535 12139
rect 27073 12133 27535 12138
rect 26726 11943 26727 11969
rect 26753 11943 26754 11969
rect 26726 11937 26754 11943
rect 27678 11970 27706 12334
rect 25158 11887 25159 11913
rect 25185 11887 25186 11913
rect 25158 11578 25186 11887
rect 27678 11913 27706 11942
rect 27678 11887 27679 11913
rect 27705 11887 27706 11913
rect 27678 11881 27706 11887
rect 28238 11969 28266 11975
rect 28238 11943 28239 11969
rect 28265 11943 28266 11969
rect 25158 11545 25186 11550
rect 25214 11578 25242 11583
rect 25158 11186 25186 11191
rect 25158 11129 25186 11158
rect 25158 11103 25159 11129
rect 25185 11103 25186 11129
rect 25158 11097 25186 11103
rect 25046 10793 25130 10794
rect 25046 10767 25047 10793
rect 25073 10767 25130 10793
rect 25046 10766 25130 10767
rect 25046 10761 25074 10766
rect 24430 10598 24682 10626
rect 24374 10375 24375 10401
rect 24401 10375 24402 10401
rect 24374 10346 24402 10375
rect 24654 10402 24682 10598
rect 24878 10402 24906 10407
rect 24654 10401 25130 10402
rect 24654 10375 24655 10401
rect 24681 10375 24879 10401
rect 24905 10375 25130 10401
rect 24654 10374 25130 10375
rect 24654 10369 24682 10374
rect 24878 10369 24906 10374
rect 24374 10313 24402 10318
rect 24430 10290 24458 10295
rect 24430 9617 24458 10262
rect 24573 10206 25035 10211
rect 24573 10205 24582 10206
rect 24573 10179 24574 10205
rect 24573 10178 24582 10179
rect 24610 10178 24634 10206
rect 24662 10178 24686 10206
rect 24714 10205 24738 10206
rect 24766 10205 24790 10206
rect 24724 10179 24738 10205
rect 24786 10179 24790 10205
rect 24714 10178 24738 10179
rect 24766 10178 24790 10179
rect 24818 10205 24842 10206
rect 24870 10205 24894 10206
rect 24818 10179 24822 10205
rect 24870 10179 24884 10205
rect 24818 10178 24842 10179
rect 24870 10178 24894 10179
rect 24922 10178 24946 10206
rect 24974 10178 24998 10206
rect 25026 10205 25035 10206
rect 25034 10179 25035 10205
rect 25026 10178 25035 10179
rect 24573 10173 25035 10178
rect 24430 9591 24431 9617
rect 24457 9591 24458 9617
rect 24430 8386 24458 9591
rect 24573 9422 25035 9427
rect 24573 9421 24582 9422
rect 24573 9395 24574 9421
rect 24573 9394 24582 9395
rect 24610 9394 24634 9422
rect 24662 9394 24686 9422
rect 24714 9421 24738 9422
rect 24766 9421 24790 9422
rect 24724 9395 24738 9421
rect 24786 9395 24790 9421
rect 24714 9394 24738 9395
rect 24766 9394 24790 9395
rect 24818 9421 24842 9422
rect 24870 9421 24894 9422
rect 24818 9395 24822 9421
rect 24870 9395 24884 9421
rect 24818 9394 24842 9395
rect 24870 9394 24894 9395
rect 24922 9394 24946 9422
rect 24974 9394 24998 9422
rect 25026 9421 25035 9422
rect 25034 9395 25035 9421
rect 25026 9394 25035 9395
rect 24573 9389 25035 9394
rect 25102 9338 25130 10374
rect 24878 9310 25130 9338
rect 24878 8946 24906 9310
rect 25046 9225 25074 9231
rect 25046 9199 25047 9225
rect 25073 9199 25074 9225
rect 25046 9114 25074 9199
rect 25046 9086 25186 9114
rect 24878 8918 25130 8946
rect 24430 8353 24458 8358
rect 24486 8833 24514 8839
rect 24486 8807 24487 8833
rect 24513 8807 24514 8833
rect 24486 8050 24514 8807
rect 24573 8638 25035 8643
rect 24573 8637 24582 8638
rect 24573 8611 24574 8637
rect 24573 8610 24582 8611
rect 24610 8610 24634 8638
rect 24662 8610 24686 8638
rect 24714 8637 24738 8638
rect 24766 8637 24790 8638
rect 24724 8611 24738 8637
rect 24786 8611 24790 8637
rect 24714 8610 24738 8611
rect 24766 8610 24790 8611
rect 24818 8637 24842 8638
rect 24870 8637 24894 8638
rect 24818 8611 24822 8637
rect 24870 8611 24884 8637
rect 24818 8610 24842 8611
rect 24870 8610 24894 8611
rect 24922 8610 24946 8638
rect 24974 8610 24998 8638
rect 25026 8637 25035 8638
rect 25034 8611 25035 8637
rect 25026 8610 25035 8611
rect 24573 8605 25035 8610
rect 24766 8441 24794 8447
rect 24766 8415 24767 8441
rect 24793 8415 24794 8441
rect 24766 8050 24794 8415
rect 24486 8049 24794 8050
rect 24486 8023 24487 8049
rect 24513 8023 24794 8049
rect 24486 8022 24794 8023
rect 24486 7574 24514 8022
rect 24573 7854 25035 7859
rect 24573 7853 24582 7854
rect 24573 7827 24574 7853
rect 24573 7826 24582 7827
rect 24610 7826 24634 7854
rect 24662 7826 24686 7854
rect 24714 7853 24738 7854
rect 24766 7853 24790 7854
rect 24724 7827 24738 7853
rect 24786 7827 24790 7853
rect 24714 7826 24738 7827
rect 24766 7826 24790 7827
rect 24818 7853 24842 7854
rect 24870 7853 24894 7854
rect 24818 7827 24822 7853
rect 24870 7827 24884 7853
rect 24818 7826 24842 7827
rect 24870 7826 24894 7827
rect 24922 7826 24946 7854
rect 24974 7826 24998 7854
rect 25026 7853 25035 7854
rect 25034 7827 25035 7853
rect 25026 7826 25035 7827
rect 24573 7821 25035 7826
rect 24822 7657 24850 7663
rect 24822 7631 24823 7657
rect 24849 7631 24850 7657
rect 24374 7546 24514 7574
rect 24654 7602 24682 7607
rect 24822 7574 24850 7631
rect 24374 7266 24402 7518
rect 24374 7219 24402 7238
rect 24654 7266 24682 7574
rect 24766 7546 24850 7574
rect 25102 7574 25130 8918
rect 25158 8386 25186 9086
rect 25214 8890 25242 11550
rect 25438 11578 25466 11583
rect 25438 11531 25466 11550
rect 27454 11578 27482 11583
rect 28238 11578 28266 11943
rect 29358 11969 29386 11975
rect 29358 11943 29359 11969
rect 29385 11943 29386 11969
rect 28574 11914 28602 11919
rect 28574 11746 28602 11886
rect 29358 11914 29386 11943
rect 29358 11867 29386 11886
rect 28518 11718 28602 11746
rect 27454 11577 28266 11578
rect 27454 11551 27455 11577
rect 27481 11551 28266 11577
rect 27454 11550 28266 11551
rect 28350 11633 28378 11639
rect 28350 11607 28351 11633
rect 28377 11607 28378 11633
rect 28350 11578 28378 11607
rect 27454 11545 27482 11550
rect 27073 11382 27535 11387
rect 27073 11381 27082 11382
rect 27073 11355 27074 11381
rect 27073 11354 27082 11355
rect 27110 11354 27134 11382
rect 27162 11354 27186 11382
rect 27214 11381 27238 11382
rect 27266 11381 27290 11382
rect 27224 11355 27238 11381
rect 27286 11355 27290 11381
rect 27214 11354 27238 11355
rect 27266 11354 27290 11355
rect 27318 11381 27342 11382
rect 27370 11381 27394 11382
rect 27318 11355 27322 11381
rect 27370 11355 27384 11381
rect 27318 11354 27342 11355
rect 27370 11354 27394 11355
rect 27422 11354 27446 11382
rect 27474 11354 27498 11382
rect 27526 11381 27535 11382
rect 27534 11355 27535 11381
rect 27526 11354 27535 11355
rect 27073 11349 27535 11354
rect 27566 11185 27594 11550
rect 27566 11159 27567 11185
rect 27593 11159 27594 11185
rect 25326 10794 25354 10799
rect 25438 10794 25466 10799
rect 25326 10793 25466 10794
rect 25326 10767 25327 10793
rect 25353 10767 25439 10793
rect 25465 10767 25466 10793
rect 25326 10766 25466 10767
rect 25326 10761 25354 10766
rect 25214 8857 25242 8862
rect 25382 9617 25410 10766
rect 25438 10761 25466 10766
rect 27454 10794 27482 10799
rect 27566 10794 27594 11159
rect 27454 10793 27594 10794
rect 27454 10767 27455 10793
rect 27481 10767 27594 10793
rect 27454 10766 27594 10767
rect 27454 10761 27482 10766
rect 27073 10598 27535 10603
rect 27073 10597 27082 10598
rect 27073 10571 27074 10597
rect 27073 10570 27082 10571
rect 27110 10570 27134 10598
rect 27162 10570 27186 10598
rect 27214 10597 27238 10598
rect 27266 10597 27290 10598
rect 27224 10571 27238 10597
rect 27286 10571 27290 10597
rect 27214 10570 27238 10571
rect 27266 10570 27290 10571
rect 27318 10597 27342 10598
rect 27370 10597 27394 10598
rect 27318 10571 27322 10597
rect 27370 10571 27384 10597
rect 27318 10570 27342 10571
rect 27370 10570 27394 10571
rect 27422 10570 27446 10598
rect 27474 10570 27498 10598
rect 27526 10597 27535 10598
rect 27534 10571 27535 10597
rect 27526 10570 27535 10571
rect 27073 10565 27535 10570
rect 25942 10066 25970 10071
rect 25942 10009 25970 10038
rect 25942 9983 25943 10009
rect 25969 9983 25970 10009
rect 25942 9977 25970 9983
rect 26838 10010 26866 10015
rect 26838 9963 26866 9982
rect 27566 10010 27594 10766
rect 28070 10906 28098 10911
rect 27678 10402 27706 10407
rect 27566 9977 27594 9982
rect 27622 10374 27678 10402
rect 27073 9814 27535 9819
rect 27073 9813 27082 9814
rect 27073 9787 27074 9813
rect 27073 9786 27082 9787
rect 27110 9786 27134 9814
rect 27162 9786 27186 9814
rect 27214 9813 27238 9814
rect 27266 9813 27290 9814
rect 27224 9787 27238 9813
rect 27286 9787 27290 9813
rect 27214 9786 27238 9787
rect 27266 9786 27290 9787
rect 27318 9813 27342 9814
rect 27370 9813 27394 9814
rect 27318 9787 27322 9813
rect 27370 9787 27384 9813
rect 27318 9786 27342 9787
rect 27370 9786 27394 9787
rect 27422 9786 27446 9814
rect 27474 9786 27498 9814
rect 27526 9813 27535 9814
rect 27534 9787 27535 9813
rect 27526 9786 27535 9787
rect 27073 9781 27535 9786
rect 25382 9591 25383 9617
rect 25409 9591 25410 9617
rect 25382 9562 25410 9591
rect 25158 8353 25186 8358
rect 25382 8833 25410 9534
rect 25382 8807 25383 8833
rect 25409 8807 25410 8833
rect 25382 8777 25410 8807
rect 25382 8751 25383 8777
rect 25409 8751 25410 8777
rect 25382 8330 25410 8751
rect 25382 8297 25410 8302
rect 25942 9281 25970 9287
rect 25942 9255 25943 9281
rect 25969 9255 25970 9281
rect 25942 9225 25970 9255
rect 27622 9282 27650 10374
rect 27678 10355 27706 10374
rect 28070 10402 28098 10878
rect 28350 10906 28378 11550
rect 28518 11185 28546 11718
rect 28854 11578 28882 11583
rect 28518 11159 28519 11185
rect 28545 11159 28546 11185
rect 28518 11130 28546 11159
rect 28350 10873 28378 10878
rect 28406 11129 28546 11130
rect 28406 11103 28519 11129
rect 28545 11103 28546 11129
rect 28406 11102 28546 11103
rect 28294 10849 28322 10855
rect 28294 10823 28295 10849
rect 28321 10823 28322 10849
rect 28294 10794 28322 10823
rect 28406 10794 28434 11102
rect 28518 11097 28546 11102
rect 28798 11577 28882 11578
rect 28798 11551 28855 11577
rect 28881 11551 28882 11577
rect 28798 11550 28882 11551
rect 28798 11185 28826 11550
rect 28854 11545 28882 11550
rect 29414 11578 29442 12726
rect 29638 12721 29666 12726
rect 29750 12721 29778 12726
rect 30198 12753 30226 12759
rect 30198 12727 30199 12753
rect 30225 12727 30226 12753
rect 29573 12558 30035 12563
rect 29573 12557 29582 12558
rect 29573 12531 29574 12557
rect 29573 12530 29582 12531
rect 29610 12530 29634 12558
rect 29662 12530 29686 12558
rect 29714 12557 29738 12558
rect 29766 12557 29790 12558
rect 29724 12531 29738 12557
rect 29786 12531 29790 12557
rect 29714 12530 29738 12531
rect 29766 12530 29790 12531
rect 29818 12557 29842 12558
rect 29870 12557 29894 12558
rect 29818 12531 29822 12557
rect 29870 12531 29884 12557
rect 29818 12530 29842 12531
rect 29870 12530 29894 12531
rect 29922 12530 29946 12558
rect 29974 12530 29998 12558
rect 30026 12557 30035 12558
rect 30034 12531 30035 12557
rect 30026 12530 30035 12531
rect 29573 12525 30035 12530
rect 29694 12362 29722 12367
rect 29918 12362 29946 12367
rect 29694 12361 29946 12362
rect 29694 12335 29695 12361
rect 29721 12335 29919 12361
rect 29945 12335 29946 12361
rect 29694 12334 29946 12335
rect 29694 12329 29722 12334
rect 29918 11914 29946 12334
rect 30198 12362 30226 12727
rect 31598 12417 31626 12423
rect 31598 12391 31599 12417
rect 31625 12391 31626 12417
rect 30198 12329 30226 12334
rect 30366 12362 30394 12367
rect 30366 12315 30394 12334
rect 30702 12362 30730 12367
rect 29918 11858 29946 11886
rect 30702 11969 30730 12334
rect 31598 12361 31626 12391
rect 31598 12335 31599 12361
rect 31625 12335 31626 12361
rect 31598 11970 31626 12335
rect 30702 11943 30703 11969
rect 30729 11943 30730 11969
rect 29918 11830 30114 11858
rect 29573 11774 30035 11779
rect 29573 11773 29582 11774
rect 29573 11747 29574 11773
rect 29573 11746 29582 11747
rect 29610 11746 29634 11774
rect 29662 11746 29686 11774
rect 29714 11773 29738 11774
rect 29766 11773 29790 11774
rect 29724 11747 29738 11773
rect 29786 11747 29790 11773
rect 29714 11746 29738 11747
rect 29766 11746 29790 11747
rect 29818 11773 29842 11774
rect 29870 11773 29894 11774
rect 29818 11747 29822 11773
rect 29870 11747 29884 11773
rect 29818 11746 29842 11747
rect 29870 11746 29894 11747
rect 29922 11746 29946 11774
rect 29974 11746 29998 11774
rect 30026 11773 30035 11774
rect 30034 11747 30035 11773
rect 30026 11746 30035 11747
rect 29573 11741 30035 11746
rect 29526 11578 29554 11583
rect 29442 11577 29554 11578
rect 29442 11551 29527 11577
rect 29553 11551 29554 11577
rect 29442 11550 29554 11551
rect 29414 11512 29442 11550
rect 28798 11159 28799 11185
rect 28825 11159 28826 11185
rect 28294 10793 28434 10794
rect 28294 10767 28295 10793
rect 28321 10767 28434 10793
rect 28294 10766 28434 10767
rect 28294 10761 28322 10766
rect 28070 10336 28098 10374
rect 27678 10066 27706 10071
rect 27678 10009 27706 10038
rect 27678 9983 27679 10009
rect 27705 9983 27706 10009
rect 27678 9977 27706 9983
rect 27902 10066 27930 10071
rect 27902 10009 27930 10038
rect 28406 10066 28434 10766
rect 28798 10793 28826 11159
rect 28798 10767 28799 10793
rect 28825 10767 28826 10793
rect 28518 10402 28546 10407
rect 28798 10402 28826 10767
rect 28518 10401 28826 10402
rect 28518 10375 28519 10401
rect 28545 10375 28799 10401
rect 28825 10375 28826 10401
rect 28518 10374 28826 10375
rect 28518 10369 28546 10374
rect 27902 9983 27903 10009
rect 27929 9983 27930 10009
rect 27734 9282 27762 9287
rect 27622 9281 27762 9282
rect 27622 9255 27735 9281
rect 27761 9255 27762 9281
rect 27622 9254 27762 9255
rect 25942 9199 25943 9225
rect 25969 9199 25970 9225
rect 25942 8497 25970 9199
rect 25942 8471 25943 8497
rect 25969 8471 25970 8497
rect 25942 8441 25970 8471
rect 26950 9225 26978 9231
rect 26950 9199 26951 9225
rect 26977 9199 26978 9225
rect 25942 8415 25943 8441
rect 25969 8415 25970 8441
rect 25942 8330 25970 8415
rect 25158 8049 25186 8055
rect 25158 8023 25159 8049
rect 25185 8023 25186 8049
rect 25158 7993 25186 8023
rect 25158 7967 25159 7993
rect 25185 7967 25186 7993
rect 25158 7658 25186 7967
rect 25158 7625 25186 7630
rect 25942 7713 25970 8302
rect 25942 7687 25943 7713
rect 25969 7687 25970 7713
rect 25942 7657 25970 7687
rect 25942 7631 25943 7657
rect 25969 7631 25970 7657
rect 25942 7602 25970 7631
rect 26222 8441 26250 8447
rect 26222 8415 26223 8441
rect 26249 8415 26250 8441
rect 26222 8386 26250 8415
rect 26222 8050 26250 8358
rect 26222 7657 26250 8022
rect 26726 8050 26754 8055
rect 26726 8003 26754 8022
rect 26222 7631 26223 7657
rect 26249 7631 26250 7657
rect 26222 7625 26250 7631
rect 25102 7546 25186 7574
rect 25942 7569 25970 7574
rect 24766 7513 24794 7518
rect 24878 7266 24906 7271
rect 24654 7265 24906 7266
rect 24654 7239 24655 7265
rect 24681 7239 24879 7265
rect 24905 7239 24906 7265
rect 24654 7238 24906 7239
rect 24654 7233 24682 7238
rect 24878 7233 24906 7238
rect 24573 7070 25035 7075
rect 24573 7069 24582 7070
rect 24573 7043 24574 7069
rect 24573 7042 24582 7043
rect 24610 7042 24634 7070
rect 24662 7042 24686 7070
rect 24714 7069 24738 7070
rect 24766 7069 24790 7070
rect 24724 7043 24738 7069
rect 24786 7043 24790 7069
rect 24714 7042 24738 7043
rect 24766 7042 24790 7043
rect 24818 7069 24842 7070
rect 24870 7069 24894 7070
rect 24818 7043 24822 7069
rect 24870 7043 24884 7069
rect 24818 7042 24842 7043
rect 24870 7042 24894 7043
rect 24922 7042 24946 7070
rect 24974 7042 24998 7070
rect 25026 7069 25035 7070
rect 25034 7043 25035 7069
rect 25026 7042 25035 7043
rect 24573 7037 25035 7042
rect 24766 6874 24794 6879
rect 24374 6873 24794 6874
rect 24374 6847 24767 6873
rect 24793 6847 24794 6873
rect 24374 6846 24794 6847
rect 23926 2585 23954 2590
rect 24262 3402 24290 3407
rect 23870 2535 23871 2561
rect 23897 2535 23898 2561
rect 23870 2506 23898 2535
rect 23422 2199 23423 2225
rect 23449 2199 23450 2225
rect 23422 2170 23450 2199
rect 23646 2505 23898 2506
rect 23646 2479 23871 2505
rect 23897 2479 23898 2505
rect 23646 2478 23898 2479
rect 23646 2170 23674 2478
rect 23870 2473 23898 2478
rect 23422 2169 23674 2170
rect 23422 2143 23423 2169
rect 23449 2143 23674 2169
rect 23422 2142 23674 2143
rect 23422 2137 23450 2142
rect 23646 1777 23674 2142
rect 23646 1751 23647 1777
rect 23673 1751 23674 1777
rect 23646 1721 23674 1751
rect 23646 1695 23647 1721
rect 23673 1695 23674 1721
rect 23646 1689 23674 1695
rect 24262 400 24290 3374
rect 24374 2450 24402 6846
rect 24766 6841 24794 6846
rect 24486 6481 24514 6487
rect 24486 6455 24487 6481
rect 24513 6455 24514 6481
rect 24430 5697 24458 5703
rect 24430 5671 24431 5697
rect 24457 5671 24458 5697
rect 24430 5418 24458 5671
rect 24486 5642 24514 6455
rect 25158 6481 25186 7546
rect 25158 6455 25159 6481
rect 25185 6455 25186 6481
rect 25158 6425 25186 6455
rect 25158 6399 25159 6425
rect 25185 6399 25186 6425
rect 24573 6286 25035 6291
rect 24573 6285 24582 6286
rect 24573 6259 24574 6285
rect 24573 6258 24582 6259
rect 24610 6258 24634 6286
rect 24662 6258 24686 6286
rect 24714 6285 24738 6286
rect 24766 6285 24790 6286
rect 24724 6259 24738 6285
rect 24786 6259 24790 6285
rect 24714 6258 24738 6259
rect 24766 6258 24790 6259
rect 24818 6285 24842 6286
rect 24870 6285 24894 6286
rect 24818 6259 24822 6285
rect 24870 6259 24884 6285
rect 24818 6258 24842 6259
rect 24870 6258 24894 6259
rect 24922 6258 24946 6286
rect 24974 6258 24998 6286
rect 25026 6285 25035 6286
rect 25034 6259 25035 6285
rect 25026 6258 25035 6259
rect 24573 6253 25035 6258
rect 24486 5609 24514 5614
rect 25046 6089 25074 6095
rect 25046 6063 25047 6089
rect 25073 6063 25074 6089
rect 25046 5642 25074 6063
rect 25158 5810 25186 6399
rect 25158 5777 25186 5782
rect 25214 6874 25242 6879
rect 25438 6874 25466 6879
rect 25214 6873 25466 6874
rect 25214 6847 25215 6873
rect 25241 6847 25439 6873
rect 25465 6847 25466 6873
rect 25214 6846 25466 6847
rect 25214 6090 25242 6846
rect 25438 6841 25466 6846
rect 25438 6090 25466 6095
rect 26222 6090 26250 6095
rect 25214 6089 25466 6090
rect 25214 6063 25215 6089
rect 25241 6063 25439 6089
rect 25465 6063 25466 6089
rect 25214 6062 25466 6063
rect 25046 5609 25074 5614
rect 25158 5698 25186 5703
rect 25214 5698 25242 6062
rect 25438 6057 25466 6062
rect 26166 6089 26250 6090
rect 26166 6063 26223 6089
rect 26249 6063 26250 6089
rect 26166 6062 26250 6063
rect 25158 5697 25242 5698
rect 25158 5671 25159 5697
rect 25185 5671 25242 5697
rect 25158 5670 25242 5671
rect 25158 5641 25186 5670
rect 25158 5615 25159 5641
rect 25185 5615 25186 5641
rect 24573 5502 25035 5507
rect 24573 5501 24582 5502
rect 24573 5475 24574 5501
rect 24573 5474 24582 5475
rect 24610 5474 24634 5502
rect 24662 5474 24686 5502
rect 24714 5501 24738 5502
rect 24766 5501 24790 5502
rect 24724 5475 24738 5501
rect 24786 5475 24790 5501
rect 24714 5474 24738 5475
rect 24766 5474 24790 5475
rect 24818 5501 24842 5502
rect 24870 5501 24894 5502
rect 24818 5475 24822 5501
rect 24870 5475 24884 5501
rect 24818 5474 24842 5475
rect 24870 5474 24894 5475
rect 24922 5474 24946 5502
rect 24974 5474 24998 5502
rect 25026 5501 25035 5502
rect 25034 5475 25035 5501
rect 25026 5474 25035 5475
rect 24573 5469 25035 5474
rect 24430 5385 24458 5390
rect 25046 5418 25074 5423
rect 25046 5306 25074 5390
rect 25158 5306 25186 5615
rect 25214 5306 25242 5311
rect 25438 5306 25466 5311
rect 25046 5305 25130 5306
rect 25046 5279 25047 5305
rect 25073 5279 25130 5305
rect 25046 5278 25130 5279
rect 25046 5273 25074 5278
rect 24486 4913 24514 4919
rect 24486 4887 24487 4913
rect 24513 4887 24514 4913
rect 24486 4522 24514 4887
rect 24654 4914 24682 4919
rect 24654 4867 24682 4886
rect 24878 4914 24906 4919
rect 24878 4867 24906 4886
rect 24573 4718 25035 4723
rect 24573 4717 24582 4718
rect 24573 4691 24574 4717
rect 24573 4690 24582 4691
rect 24610 4690 24634 4718
rect 24662 4690 24686 4718
rect 24714 4717 24738 4718
rect 24766 4717 24790 4718
rect 24724 4691 24738 4717
rect 24786 4691 24790 4717
rect 24714 4690 24738 4691
rect 24766 4690 24790 4691
rect 24818 4717 24842 4718
rect 24870 4717 24894 4718
rect 24818 4691 24822 4717
rect 24870 4691 24884 4717
rect 24818 4690 24842 4691
rect 24870 4690 24894 4691
rect 24922 4690 24946 4718
rect 24974 4690 24998 4718
rect 25026 4717 25035 4718
rect 25034 4691 25035 4717
rect 25026 4690 25035 4691
rect 24573 4685 25035 4690
rect 24766 4522 24794 4527
rect 24486 4521 24794 4522
rect 24486 4495 24767 4521
rect 24793 4495 24794 4521
rect 24486 4494 24794 4495
rect 24486 4214 24514 4494
rect 24766 4489 24794 4494
rect 24374 2282 24402 2422
rect 24374 2249 24402 2254
rect 24430 4186 24514 4214
rect 24430 3346 24458 4186
rect 24486 4130 24514 4135
rect 24486 4083 24514 4102
rect 25102 4130 25130 5278
rect 25158 5305 25466 5306
rect 25158 5279 25215 5305
rect 25241 5279 25439 5305
rect 25465 5279 25466 5305
rect 25158 5278 25466 5279
rect 25158 4914 25186 5278
rect 25214 5273 25242 5278
rect 25438 5273 25466 5278
rect 25186 4886 25242 4914
rect 25158 4881 25186 4886
rect 25214 4522 25242 4886
rect 25438 4522 25466 4527
rect 25214 4521 25438 4522
rect 25214 4495 25215 4521
rect 25241 4495 25438 4521
rect 25214 4494 25438 4495
rect 25214 4489 25242 4494
rect 25438 4456 25466 4494
rect 25102 4097 25130 4102
rect 25382 4129 25410 4135
rect 25382 4103 25383 4129
rect 25409 4103 25410 4129
rect 25382 4073 25410 4103
rect 25382 4047 25383 4073
rect 25409 4047 25410 4073
rect 24573 3934 25035 3939
rect 24573 3933 24582 3934
rect 24573 3907 24574 3933
rect 24573 3906 24582 3907
rect 24610 3906 24634 3934
rect 24662 3906 24686 3934
rect 24714 3933 24738 3934
rect 24766 3933 24790 3934
rect 24724 3907 24738 3933
rect 24786 3907 24790 3933
rect 24714 3906 24738 3907
rect 24766 3906 24790 3907
rect 24818 3933 24842 3934
rect 24870 3933 24894 3934
rect 24818 3907 24822 3933
rect 24870 3907 24884 3933
rect 24818 3906 24842 3907
rect 24870 3906 24894 3907
rect 24922 3906 24946 3934
rect 24974 3906 24998 3934
rect 25026 3933 25035 3934
rect 25034 3907 25035 3933
rect 25026 3906 25035 3907
rect 24573 3901 25035 3906
rect 24766 3737 24794 3743
rect 24766 3711 24767 3737
rect 24793 3711 24794 3737
rect 24766 3346 24794 3711
rect 24430 3345 24794 3346
rect 24430 3319 24431 3345
rect 24457 3319 24794 3345
rect 24430 3318 24794 3319
rect 25382 3458 25410 4047
rect 26166 3850 26194 6062
rect 26222 6057 26250 6062
rect 26894 5697 26922 5703
rect 26894 5671 26895 5697
rect 26921 5671 26922 5697
rect 26502 5642 26530 5647
rect 26502 5305 26530 5614
rect 26894 5586 26922 5671
rect 26894 5553 26922 5558
rect 26502 5279 26503 5305
rect 26529 5279 26530 5305
rect 26502 4746 26530 5279
rect 26782 5306 26810 5311
rect 26894 5306 26922 5311
rect 26782 5305 26922 5306
rect 26782 5279 26783 5305
rect 26809 5279 26895 5305
rect 26921 5279 26922 5305
rect 26782 5278 26922 5279
rect 26782 5273 26810 5278
rect 26894 5026 26922 5278
rect 26894 4993 26922 4998
rect 26502 4713 26530 4718
rect 26894 4913 26922 4919
rect 26894 4887 26895 4913
rect 26921 4887 26922 4913
rect 26894 4746 26922 4887
rect 26894 4713 26922 4718
rect 26502 4521 26530 4527
rect 26502 4495 26503 4521
rect 26529 4495 26530 4521
rect 26502 4130 26530 4495
rect 26894 4522 26922 4527
rect 26894 4242 26922 4494
rect 26502 4097 26530 4102
rect 26838 4130 26866 4135
rect 25382 3345 25410 3430
rect 25382 3319 25383 3345
rect 25409 3319 25410 3345
rect 24430 2561 24458 3318
rect 25382 3289 25410 3319
rect 25382 3263 25383 3289
rect 25409 3263 25410 3289
rect 24573 3150 25035 3155
rect 24573 3149 24582 3150
rect 24573 3123 24574 3149
rect 24573 3122 24582 3123
rect 24610 3122 24634 3150
rect 24662 3122 24686 3150
rect 24714 3149 24738 3150
rect 24766 3149 24790 3150
rect 24724 3123 24738 3149
rect 24786 3123 24790 3149
rect 24714 3122 24738 3123
rect 24766 3122 24790 3123
rect 24818 3149 24842 3150
rect 24870 3149 24894 3150
rect 24818 3123 24822 3149
rect 24870 3123 24884 3149
rect 24818 3122 24842 3123
rect 24870 3122 24894 3123
rect 24922 3122 24946 3150
rect 24974 3122 24998 3150
rect 25026 3149 25035 3150
rect 25034 3123 25035 3149
rect 25026 3122 25035 3123
rect 24573 3117 25035 3122
rect 24430 2535 24431 2561
rect 24457 2535 24458 2561
rect 24430 2506 24458 2535
rect 24430 1834 24458 2478
rect 24766 2953 24794 2959
rect 24766 2927 24767 2953
rect 24793 2927 24794 2953
rect 24766 2506 24794 2927
rect 24766 2473 24794 2478
rect 25382 2561 25410 3263
rect 25382 2535 25383 2561
rect 25409 2535 25410 2561
rect 25382 2505 25410 2535
rect 25382 2479 25383 2505
rect 25409 2479 25410 2505
rect 24573 2366 25035 2371
rect 24573 2365 24582 2366
rect 24573 2339 24574 2365
rect 24573 2338 24582 2339
rect 24610 2338 24634 2366
rect 24662 2338 24686 2366
rect 24714 2365 24738 2366
rect 24766 2365 24790 2366
rect 24724 2339 24738 2365
rect 24786 2339 24790 2365
rect 24714 2338 24738 2339
rect 24766 2338 24790 2339
rect 24818 2365 24842 2366
rect 24870 2365 24894 2366
rect 24818 2339 24822 2365
rect 24870 2339 24884 2365
rect 24818 2338 24842 2339
rect 24870 2338 24894 2339
rect 24922 2338 24946 2366
rect 24974 2338 24998 2366
rect 25026 2365 25035 2366
rect 25034 2339 25035 2365
rect 25026 2338 25035 2339
rect 24573 2333 25035 2338
rect 24430 1777 24458 1806
rect 24766 2170 24794 2175
rect 25382 2170 25410 2479
rect 25942 3793 25970 3799
rect 25942 3767 25943 3793
rect 25969 3767 25970 3793
rect 25942 3737 25970 3767
rect 25942 3711 25943 3737
rect 25969 3711 25970 3737
rect 25942 3009 25970 3711
rect 26166 3402 26194 3822
rect 26166 3369 26194 3374
rect 26222 3737 26250 3743
rect 26222 3711 26223 3737
rect 26249 3711 26250 3737
rect 25942 2983 25943 3009
rect 25969 2983 25970 3009
rect 25942 2953 25970 2983
rect 25942 2927 25943 2953
rect 25969 2927 25970 2953
rect 25942 2674 25970 2927
rect 25942 2225 25970 2646
rect 25942 2199 25943 2225
rect 25969 2199 25970 2225
rect 25942 2170 25970 2199
rect 25382 2169 25970 2170
rect 25382 2143 25943 2169
rect 25969 2143 25970 2169
rect 25382 2142 25970 2143
rect 24766 1834 24794 2142
rect 24766 1801 24794 1806
rect 24430 1751 24431 1777
rect 24457 1751 24458 1777
rect 24430 1745 24458 1751
rect 25606 1777 25634 2142
rect 25942 2137 25970 2142
rect 25998 3346 26026 3351
rect 25606 1751 25607 1777
rect 25633 1751 25634 1777
rect 25606 1721 25634 1751
rect 25606 1695 25607 1721
rect 25633 1695 25634 1721
rect 25606 1689 25634 1695
rect 25998 1694 26026 3318
rect 26222 2953 26250 3711
rect 26838 3738 26866 4102
rect 26894 3906 26922 4214
rect 26894 3873 26922 3878
rect 26838 3710 26922 3738
rect 26894 3345 26922 3710
rect 26894 3319 26895 3345
rect 26921 3319 26922 3345
rect 26894 3313 26922 3319
rect 26222 2927 26223 2953
rect 26249 2927 26250 2953
rect 26222 2562 26250 2927
rect 26222 2170 26250 2534
rect 26726 2562 26754 2567
rect 26726 2515 26754 2534
rect 26222 2123 26250 2142
rect 26390 2506 26418 2511
rect 25886 1666 26026 1694
rect 26390 1777 26418 2478
rect 26390 1751 26391 1777
rect 26417 1751 26418 1777
rect 26390 1722 26418 1751
rect 26390 1689 26418 1694
rect 26726 2282 26754 2287
rect 24573 1582 25035 1587
rect 24573 1581 24582 1582
rect 24573 1555 24574 1581
rect 24573 1554 24582 1555
rect 24610 1554 24634 1582
rect 24662 1554 24686 1582
rect 24714 1581 24738 1582
rect 24766 1581 24790 1582
rect 24724 1555 24738 1581
rect 24786 1555 24790 1581
rect 24714 1554 24738 1555
rect 24766 1554 24790 1555
rect 24818 1581 24842 1582
rect 24870 1581 24894 1582
rect 24818 1555 24822 1581
rect 24870 1555 24884 1581
rect 24818 1554 24842 1555
rect 24870 1554 24894 1555
rect 24922 1554 24946 1582
rect 24974 1554 24998 1582
rect 25026 1581 25035 1582
rect 25034 1555 25035 1581
rect 25026 1554 25035 1555
rect 24573 1549 25035 1554
rect 25494 462 25690 490
rect 25494 400 25522 462
rect 12782 350 13034 378
rect 13160 0 13216 400
rect 14392 0 14448 400
rect 15624 0 15680 400
rect 16856 0 16912 400
rect 18088 0 18144 400
rect 19320 0 19376 400
rect 20552 0 20608 400
rect 21784 0 21840 400
rect 23016 0 23072 400
rect 24248 0 24304 400
rect 25480 0 25536 400
rect 25662 378 25690 462
rect 25886 378 25914 1666
rect 26726 400 26754 2254
rect 26950 2282 26978 9199
rect 27622 9225 27650 9254
rect 27622 9199 27623 9225
rect 27649 9199 27650 9225
rect 27622 9193 27650 9199
rect 27073 9030 27535 9035
rect 27073 9029 27082 9030
rect 27073 9003 27074 9029
rect 27073 9002 27082 9003
rect 27110 9002 27134 9030
rect 27162 9002 27186 9030
rect 27214 9029 27238 9030
rect 27266 9029 27290 9030
rect 27224 9003 27238 9029
rect 27286 9003 27290 9029
rect 27214 9002 27238 9003
rect 27266 9002 27290 9003
rect 27318 9029 27342 9030
rect 27370 9029 27394 9030
rect 27318 9003 27322 9029
rect 27370 9003 27384 9029
rect 27318 9002 27342 9003
rect 27370 9002 27394 9003
rect 27422 9002 27446 9030
rect 27474 9002 27498 9030
rect 27526 9029 27535 9030
rect 27534 9003 27535 9029
rect 27526 9002 27535 9003
rect 27073 8997 27535 9002
rect 27566 8890 27594 8895
rect 27398 8497 27426 8503
rect 27398 8471 27399 8497
rect 27425 8471 27426 8497
rect 27398 8441 27426 8471
rect 27398 8415 27399 8441
rect 27425 8415 27426 8441
rect 27398 8386 27426 8415
rect 27398 8353 27426 8358
rect 27073 8246 27535 8251
rect 27073 8245 27082 8246
rect 27073 8219 27074 8245
rect 27073 8218 27082 8219
rect 27110 8218 27134 8246
rect 27162 8218 27186 8246
rect 27214 8245 27238 8246
rect 27266 8245 27290 8246
rect 27224 8219 27238 8245
rect 27286 8219 27290 8245
rect 27214 8218 27238 8219
rect 27266 8218 27290 8219
rect 27318 8245 27342 8246
rect 27370 8245 27394 8246
rect 27318 8219 27322 8245
rect 27370 8219 27384 8245
rect 27318 8218 27342 8219
rect 27370 8218 27394 8219
rect 27422 8218 27446 8246
rect 27474 8218 27498 8246
rect 27526 8245 27535 8246
rect 27534 8219 27535 8245
rect 27526 8218 27535 8219
rect 27073 8213 27535 8218
rect 27566 8162 27594 8862
rect 27734 8833 27762 9254
rect 27734 8807 27735 8833
rect 27761 8807 27762 8833
rect 27734 8778 27762 8807
rect 27398 8134 27594 8162
rect 27622 8777 27762 8778
rect 27622 8751 27735 8777
rect 27761 8751 27762 8777
rect 27622 8750 27762 8751
rect 27398 7713 27426 8134
rect 27398 7687 27399 7713
rect 27425 7687 27426 7713
rect 27398 7657 27426 7687
rect 27398 7631 27399 7657
rect 27425 7631 27426 7657
rect 27398 7625 27426 7631
rect 27073 7462 27535 7467
rect 27073 7461 27082 7462
rect 27073 7435 27074 7461
rect 27073 7434 27082 7435
rect 27110 7434 27134 7462
rect 27162 7434 27186 7462
rect 27214 7461 27238 7462
rect 27266 7461 27290 7462
rect 27224 7435 27238 7461
rect 27286 7435 27290 7461
rect 27214 7434 27238 7435
rect 27266 7434 27290 7435
rect 27318 7461 27342 7462
rect 27370 7461 27394 7462
rect 27318 7435 27322 7461
rect 27370 7435 27384 7461
rect 27318 7434 27342 7435
rect 27370 7434 27394 7435
rect 27422 7434 27446 7462
rect 27474 7434 27498 7462
rect 27526 7461 27535 7462
rect 27534 7435 27535 7461
rect 27526 7434 27535 7435
rect 27073 7429 27535 7434
rect 27622 7266 27650 8750
rect 27734 8745 27762 8750
rect 27678 8386 27706 8391
rect 27678 8049 27706 8358
rect 27678 8023 27679 8049
rect 27705 8023 27706 8049
rect 27678 7993 27706 8023
rect 27678 7967 27679 7993
rect 27705 7967 27706 7993
rect 27678 7961 27706 7967
rect 27902 7574 27930 9983
rect 27846 7546 27930 7574
rect 27958 10010 27986 10015
rect 27958 9170 27986 9982
rect 28350 10010 28378 10015
rect 28350 9963 28378 9982
rect 28182 9618 28210 9623
rect 28406 9618 28434 10038
rect 28182 9617 28434 9618
rect 28182 9591 28183 9617
rect 28209 9591 28407 9617
rect 28433 9591 28434 9617
rect 28182 9590 28434 9591
rect 28182 9585 28210 9590
rect 28406 9585 28434 9590
rect 28798 10010 28826 10374
rect 29470 10066 29498 11550
rect 29526 11545 29554 11550
rect 29974 11185 30002 11191
rect 29974 11159 29975 11185
rect 30001 11159 30002 11185
rect 29974 11130 30002 11159
rect 30086 11130 30114 11830
rect 30590 11578 30618 11583
rect 30702 11578 30730 11943
rect 31430 11969 31682 11970
rect 31430 11943 31599 11969
rect 31625 11943 31682 11969
rect 31430 11942 31682 11943
rect 30590 11577 30786 11578
rect 30590 11551 30591 11577
rect 30617 11551 30786 11577
rect 30590 11550 30786 11551
rect 30590 11545 30618 11550
rect 29974 11129 30114 11130
rect 29974 11103 29975 11129
rect 30001 11103 30114 11129
rect 29974 11102 30114 11103
rect 29974 11097 30002 11102
rect 29573 10990 30035 10995
rect 29573 10989 29582 10990
rect 29573 10963 29574 10989
rect 29573 10962 29582 10963
rect 29610 10962 29634 10990
rect 29662 10962 29686 10990
rect 29714 10989 29738 10990
rect 29766 10989 29790 10990
rect 29724 10963 29738 10989
rect 29786 10963 29790 10989
rect 29714 10962 29738 10963
rect 29766 10962 29790 10963
rect 29818 10989 29842 10990
rect 29870 10989 29894 10990
rect 29818 10963 29822 10989
rect 29870 10963 29884 10989
rect 29818 10962 29842 10963
rect 29870 10962 29894 10963
rect 29922 10962 29946 10990
rect 29974 10962 29998 10990
rect 30026 10989 30035 10990
rect 30034 10963 30035 10989
rect 30026 10962 30035 10963
rect 29573 10957 30035 10962
rect 29974 10850 30002 10855
rect 30086 10850 30114 11102
rect 29974 10849 30114 10850
rect 29974 10823 29975 10849
rect 30001 10823 30114 10849
rect 29974 10822 30114 10823
rect 30758 11185 30786 11550
rect 30758 11159 30759 11185
rect 30785 11159 30786 11185
rect 29974 10793 30002 10822
rect 29974 10767 29975 10793
rect 30001 10767 30002 10793
rect 29974 10401 30002 10767
rect 29974 10375 29975 10401
rect 30001 10375 30002 10401
rect 29974 10345 30002 10375
rect 29974 10319 29975 10345
rect 30001 10319 30002 10345
rect 29974 10290 30002 10319
rect 30310 10793 30338 10799
rect 30310 10767 30311 10793
rect 30337 10767 30338 10793
rect 29974 10262 30226 10290
rect 29573 10206 30035 10211
rect 29573 10205 29582 10206
rect 29573 10179 29574 10205
rect 29573 10178 29582 10179
rect 29610 10178 29634 10206
rect 29662 10178 29686 10206
rect 29714 10205 29738 10206
rect 29766 10205 29790 10206
rect 29724 10179 29738 10205
rect 29786 10179 29790 10205
rect 29714 10178 29738 10179
rect 29766 10178 29790 10179
rect 29818 10205 29842 10206
rect 29870 10205 29894 10206
rect 29818 10179 29822 10205
rect 29870 10179 29884 10205
rect 29818 10178 29842 10179
rect 29870 10178 29894 10179
rect 29922 10178 29946 10206
rect 29974 10178 29998 10206
rect 30026 10205 30035 10206
rect 30034 10179 30035 10205
rect 30026 10178 30035 10179
rect 29573 10173 30035 10178
rect 29470 10033 29498 10038
rect 29806 10066 29834 10071
rect 28798 9617 28826 9982
rect 28798 9591 28799 9617
rect 28825 9591 28826 9617
rect 27678 7266 27706 7271
rect 27622 7265 27706 7266
rect 27622 7239 27679 7265
rect 27705 7239 27706 7265
rect 27622 7238 27706 7239
rect 27678 7209 27706 7238
rect 27678 7183 27679 7209
rect 27705 7183 27706 7209
rect 27566 6874 27594 6879
rect 27073 6678 27535 6683
rect 27073 6677 27082 6678
rect 27073 6651 27074 6677
rect 27073 6650 27082 6651
rect 27110 6650 27134 6678
rect 27162 6650 27186 6678
rect 27214 6677 27238 6678
rect 27266 6677 27290 6678
rect 27224 6651 27238 6677
rect 27286 6651 27290 6677
rect 27214 6650 27238 6651
rect 27266 6650 27290 6651
rect 27318 6677 27342 6678
rect 27370 6677 27394 6678
rect 27318 6651 27322 6677
rect 27370 6651 27384 6677
rect 27318 6650 27342 6651
rect 27370 6650 27394 6651
rect 27422 6650 27446 6678
rect 27474 6650 27498 6678
rect 27526 6677 27535 6678
rect 27534 6651 27535 6677
rect 27526 6650 27535 6651
rect 27073 6645 27535 6650
rect 27398 6146 27426 6151
rect 27566 6146 27594 6846
rect 27678 6874 27706 7183
rect 27678 6841 27706 6846
rect 27790 6874 27818 6879
rect 27790 6827 27818 6846
rect 27846 6481 27874 7546
rect 27846 6455 27847 6481
rect 27873 6455 27874 6481
rect 27846 6425 27874 6455
rect 27846 6399 27847 6425
rect 27873 6399 27874 6425
rect 27846 6393 27874 6399
rect 27398 6145 27594 6146
rect 27398 6119 27399 6145
rect 27425 6119 27594 6145
rect 27398 6118 27594 6119
rect 27398 6089 27426 6118
rect 27398 6063 27399 6089
rect 27425 6063 27426 6089
rect 27398 6057 27426 6063
rect 27073 5894 27535 5899
rect 27073 5893 27082 5894
rect 27073 5867 27074 5893
rect 27073 5866 27082 5867
rect 27110 5866 27134 5894
rect 27162 5866 27186 5894
rect 27214 5893 27238 5894
rect 27266 5893 27290 5894
rect 27224 5867 27238 5893
rect 27286 5867 27290 5893
rect 27214 5866 27238 5867
rect 27266 5866 27290 5867
rect 27318 5893 27342 5894
rect 27370 5893 27394 5894
rect 27318 5867 27322 5893
rect 27370 5867 27384 5893
rect 27318 5866 27342 5867
rect 27370 5866 27394 5867
rect 27422 5866 27446 5894
rect 27474 5866 27498 5894
rect 27526 5893 27535 5894
rect 27534 5867 27535 5893
rect 27526 5866 27535 5867
rect 27073 5861 27535 5866
rect 27622 5697 27650 5703
rect 27622 5671 27623 5697
rect 27649 5671 27650 5697
rect 27622 5642 27650 5671
rect 27678 5642 27706 5647
rect 27622 5641 27706 5642
rect 27622 5615 27679 5641
rect 27705 5615 27706 5641
rect 27622 5614 27706 5615
rect 27006 5586 27034 5591
rect 27006 4914 27034 5558
rect 27073 5110 27535 5115
rect 27073 5109 27082 5110
rect 27073 5083 27074 5109
rect 27073 5082 27082 5083
rect 27110 5082 27134 5110
rect 27162 5082 27186 5110
rect 27214 5109 27238 5110
rect 27266 5109 27290 5110
rect 27224 5083 27238 5109
rect 27286 5083 27290 5109
rect 27214 5082 27238 5083
rect 27266 5082 27290 5083
rect 27318 5109 27342 5110
rect 27370 5109 27394 5110
rect 27318 5083 27322 5109
rect 27370 5083 27384 5109
rect 27318 5082 27342 5083
rect 27370 5082 27394 5083
rect 27422 5082 27446 5110
rect 27474 5082 27498 5110
rect 27526 5109 27535 5110
rect 27534 5083 27535 5109
rect 27526 5082 27535 5083
rect 27073 5077 27535 5082
rect 27006 4881 27034 4886
rect 27174 5026 27202 5031
rect 27174 4914 27202 4998
rect 27398 4914 27426 4919
rect 27174 4913 27426 4914
rect 27174 4887 27175 4913
rect 27201 4887 27399 4913
rect 27425 4887 27426 4913
rect 27174 4886 27426 4887
rect 27174 4577 27202 4886
rect 27398 4881 27426 4886
rect 27174 4551 27175 4577
rect 27201 4551 27202 4577
rect 27174 4522 27202 4551
rect 27174 4489 27202 4494
rect 27073 4326 27535 4331
rect 27073 4325 27082 4326
rect 27073 4299 27074 4325
rect 27073 4298 27082 4299
rect 27110 4298 27134 4326
rect 27162 4298 27186 4326
rect 27214 4325 27238 4326
rect 27266 4325 27290 4326
rect 27224 4299 27238 4325
rect 27286 4299 27290 4325
rect 27214 4298 27238 4299
rect 27266 4298 27290 4299
rect 27318 4325 27342 4326
rect 27370 4325 27394 4326
rect 27318 4299 27322 4325
rect 27370 4299 27384 4325
rect 27318 4298 27342 4299
rect 27370 4298 27394 4299
rect 27422 4298 27446 4326
rect 27474 4298 27498 4326
rect 27526 4325 27535 4326
rect 27534 4299 27535 4325
rect 27526 4298 27535 4299
rect 27073 4293 27535 4298
rect 27510 4242 27538 4247
rect 27510 4129 27538 4214
rect 27510 4103 27511 4129
rect 27537 4103 27538 4129
rect 27510 4097 27538 4103
rect 27174 3906 27202 3911
rect 27174 3793 27202 3878
rect 27174 3767 27175 3793
rect 27201 3767 27202 3793
rect 27174 3737 27202 3767
rect 27174 3711 27175 3737
rect 27201 3711 27202 3737
rect 27174 3705 27202 3711
rect 27073 3542 27535 3547
rect 27073 3541 27082 3542
rect 27073 3515 27074 3541
rect 27073 3514 27082 3515
rect 27110 3514 27134 3542
rect 27162 3514 27186 3542
rect 27214 3541 27238 3542
rect 27266 3541 27290 3542
rect 27224 3515 27238 3541
rect 27286 3515 27290 3541
rect 27214 3514 27238 3515
rect 27266 3514 27290 3515
rect 27318 3541 27342 3542
rect 27370 3541 27394 3542
rect 27318 3515 27322 3541
rect 27370 3515 27384 3541
rect 27318 3514 27342 3515
rect 27370 3514 27394 3515
rect 27422 3514 27446 3542
rect 27474 3514 27498 3542
rect 27526 3541 27535 3542
rect 27534 3515 27535 3541
rect 27526 3514 27535 3515
rect 27073 3509 27535 3514
rect 27622 3066 27650 5614
rect 27678 5609 27706 5614
rect 27398 3038 27650 3066
rect 27398 3009 27426 3038
rect 27398 2983 27399 3009
rect 27425 2983 27426 3009
rect 27398 2953 27426 2983
rect 27398 2927 27399 2953
rect 27425 2927 27426 2953
rect 27398 2921 27426 2927
rect 27073 2758 27535 2763
rect 27073 2757 27082 2758
rect 27073 2731 27074 2757
rect 27073 2730 27082 2731
rect 27110 2730 27134 2758
rect 27162 2730 27186 2758
rect 27214 2757 27238 2758
rect 27266 2757 27290 2758
rect 27224 2731 27238 2757
rect 27286 2731 27290 2757
rect 27214 2730 27238 2731
rect 27266 2730 27290 2731
rect 27318 2757 27342 2758
rect 27370 2757 27394 2758
rect 27318 2731 27322 2757
rect 27370 2731 27384 2757
rect 27318 2730 27342 2731
rect 27370 2730 27394 2731
rect 27422 2730 27446 2758
rect 27474 2730 27498 2758
rect 27526 2757 27535 2758
rect 27534 2731 27535 2757
rect 27526 2730 27535 2731
rect 27073 2725 27535 2730
rect 26950 2249 26978 2254
rect 27622 2674 27650 3038
rect 27398 2226 27426 2231
rect 27398 2169 27426 2198
rect 27398 2143 27399 2169
rect 27425 2143 27426 2169
rect 27398 2137 27426 2143
rect 27073 1974 27535 1979
rect 27073 1973 27082 1974
rect 27073 1947 27074 1973
rect 27073 1946 27082 1947
rect 27110 1946 27134 1974
rect 27162 1946 27186 1974
rect 27214 1973 27238 1974
rect 27266 1973 27290 1974
rect 27224 1947 27238 1973
rect 27286 1947 27290 1973
rect 27214 1946 27238 1947
rect 27266 1946 27290 1947
rect 27318 1973 27342 1974
rect 27370 1973 27394 1974
rect 27318 1947 27322 1973
rect 27370 1947 27384 1973
rect 27318 1946 27342 1947
rect 27370 1946 27394 1947
rect 27422 1946 27446 1974
rect 27474 1946 27498 1974
rect 27526 1973 27535 1974
rect 27534 1947 27535 1973
rect 27526 1946 27535 1947
rect 27073 1941 27535 1946
rect 27566 1778 27594 1783
rect 27622 1778 27650 2646
rect 27678 4242 27706 4247
rect 27678 4073 27706 4214
rect 27678 4047 27679 4073
rect 27705 4047 27706 4073
rect 27678 3345 27706 4047
rect 27678 3319 27679 3345
rect 27705 3319 27706 3345
rect 27678 3289 27706 3319
rect 27678 3263 27679 3289
rect 27705 3263 27706 3289
rect 27678 2561 27706 3263
rect 27678 2535 27679 2561
rect 27705 2535 27706 2561
rect 27678 2505 27706 2535
rect 27678 2479 27679 2505
rect 27705 2479 27706 2505
rect 27678 2226 27706 2479
rect 27678 2193 27706 2198
rect 27566 1777 27650 1778
rect 27566 1751 27567 1777
rect 27593 1751 27650 1777
rect 27566 1750 27650 1751
rect 27566 1721 27594 1750
rect 27566 1695 27567 1721
rect 27593 1695 27594 1721
rect 27566 1689 27594 1695
rect 27958 400 27986 9142
rect 28350 6873 28378 6879
rect 28350 6847 28351 6873
rect 28377 6847 28378 6873
rect 28350 6762 28378 6847
rect 28350 6729 28378 6734
rect 28238 5026 28266 5031
rect 28182 4746 28210 4751
rect 28070 4578 28098 4583
rect 28070 4466 28098 4550
rect 28070 4214 28098 4438
rect 28014 4186 28098 4214
rect 28182 4214 28210 4718
rect 28238 4578 28266 4998
rect 28462 4914 28490 4919
rect 28238 4512 28266 4550
rect 28294 4858 28322 4863
rect 28182 4186 28266 4214
rect 28014 3738 28042 4186
rect 28238 4153 28266 4158
rect 28182 3738 28210 3743
rect 28014 3737 28210 3738
rect 28014 3711 28015 3737
rect 28041 3711 28183 3737
rect 28209 3711 28210 3737
rect 28014 3710 28210 3711
rect 28014 3705 28042 3710
rect 28070 3009 28098 3710
rect 28182 3705 28210 3710
rect 28294 3737 28322 4830
rect 28350 4521 28378 4527
rect 28350 4495 28351 4521
rect 28377 4495 28378 4521
rect 28350 4214 28378 4495
rect 28462 4522 28490 4886
rect 28462 4489 28490 4494
rect 28742 4522 28770 4527
rect 28742 4475 28770 4494
rect 28686 4242 28714 4247
rect 28350 4186 28546 4214
rect 28294 3711 28295 3737
rect 28321 3711 28322 3737
rect 28294 3705 28322 3711
rect 28462 4130 28490 4135
rect 28462 3345 28490 4102
rect 28462 3319 28463 3345
rect 28489 3319 28490 3345
rect 28070 2983 28071 3009
rect 28097 2983 28098 3009
rect 28070 2954 28098 2983
rect 28350 3010 28378 3015
rect 28350 2963 28378 2982
rect 28182 2954 28210 2959
rect 28070 2953 28210 2954
rect 28070 2927 28183 2953
rect 28209 2927 28210 2953
rect 28070 2926 28210 2927
rect 28182 2921 28210 2926
rect 28070 2618 28098 2623
rect 28070 2225 28098 2590
rect 28462 2562 28490 3319
rect 28518 3010 28546 4186
rect 28686 4129 28714 4214
rect 28686 4103 28687 4129
rect 28713 4103 28714 4129
rect 28686 4097 28714 4103
rect 28518 2977 28546 2982
rect 28462 2515 28490 2534
rect 28742 2953 28770 2959
rect 28742 2927 28743 2953
rect 28769 2927 28770 2953
rect 28742 2562 28770 2927
rect 28070 2199 28071 2225
rect 28097 2199 28098 2225
rect 28070 2170 28098 2199
rect 28182 2170 28210 2175
rect 28070 2169 28210 2170
rect 28070 2143 28183 2169
rect 28209 2143 28210 2169
rect 28070 2142 28210 2143
rect 28182 2137 28210 2142
rect 28350 2169 28378 2175
rect 28350 2143 28351 2169
rect 28377 2143 28378 2169
rect 28350 2114 28378 2143
rect 28742 2169 28770 2534
rect 28742 2143 28743 2169
rect 28769 2143 28770 2169
rect 28742 2137 28770 2143
rect 28350 2081 28378 2086
rect 28518 1778 28546 1783
rect 28518 1731 28546 1750
rect 25662 350 25914 378
rect 26712 0 26768 400
rect 27944 0 28000 400
rect 28798 378 28826 9591
rect 29414 10009 29442 10015
rect 29414 9983 29415 10009
rect 29441 9983 29442 10009
rect 29414 9617 29442 9983
rect 29806 10009 29834 10038
rect 29806 9983 29807 10009
rect 29833 9983 29834 10009
rect 29414 9591 29415 9617
rect 29441 9591 29442 9617
rect 29414 9226 29442 9591
rect 29694 9618 29722 9623
rect 29806 9618 29834 9983
rect 30030 10066 30058 10071
rect 30030 10010 30058 10038
rect 30030 10009 30114 10010
rect 30030 9983 30031 10009
rect 30057 9983 30114 10009
rect 30030 9982 30114 9983
rect 30030 9977 30058 9982
rect 29694 9617 29834 9618
rect 29694 9591 29695 9617
rect 29721 9591 29807 9617
rect 29833 9591 29834 9617
rect 29694 9590 29834 9591
rect 29694 9585 29722 9590
rect 29806 9585 29834 9590
rect 30086 9898 30114 9982
rect 29573 9422 30035 9427
rect 29573 9421 29582 9422
rect 29573 9395 29574 9421
rect 29573 9394 29582 9395
rect 29610 9394 29634 9422
rect 29662 9394 29686 9422
rect 29714 9421 29738 9422
rect 29766 9421 29790 9422
rect 29724 9395 29738 9421
rect 29786 9395 29790 9421
rect 29714 9394 29738 9395
rect 29766 9394 29790 9395
rect 29818 9421 29842 9422
rect 29870 9421 29894 9422
rect 29818 9395 29822 9421
rect 29870 9395 29884 9421
rect 29818 9394 29842 9395
rect 29870 9394 29894 9395
rect 29922 9394 29946 9422
rect 29974 9394 29998 9422
rect 30026 9421 30035 9422
rect 30034 9395 30035 9421
rect 30026 9394 30035 9395
rect 29573 9389 30035 9394
rect 29414 9193 29442 9198
rect 29526 9226 29554 9231
rect 28854 8834 28882 8839
rect 28854 8787 28882 8806
rect 29414 8834 29442 8839
rect 29526 8834 29554 9198
rect 29442 8806 29554 8834
rect 29414 8768 29442 8806
rect 29573 8638 30035 8643
rect 29573 8637 29582 8638
rect 29573 8611 29574 8637
rect 29573 8610 29582 8611
rect 29610 8610 29634 8638
rect 29662 8610 29686 8638
rect 29714 8637 29738 8638
rect 29766 8637 29790 8638
rect 29724 8611 29738 8637
rect 29786 8611 29790 8637
rect 29714 8610 29738 8611
rect 29766 8610 29790 8611
rect 29818 8637 29842 8638
rect 29870 8637 29894 8638
rect 29818 8611 29822 8637
rect 29870 8611 29884 8637
rect 29818 8610 29842 8611
rect 29870 8610 29894 8611
rect 29922 8610 29946 8638
rect 29974 8610 29998 8638
rect 30026 8637 30035 8638
rect 30034 8611 30035 8637
rect 30026 8610 30035 8611
rect 29573 8605 30035 8610
rect 29414 8441 29442 8447
rect 29414 8415 29415 8441
rect 29441 8415 29442 8441
rect 29358 8050 29386 8055
rect 29414 8050 29442 8415
rect 29358 8049 29442 8050
rect 29358 8023 29359 8049
rect 29385 8023 29442 8049
rect 29358 8022 29442 8023
rect 29862 8442 29890 8447
rect 30086 8442 30114 9870
rect 29862 8441 30114 8442
rect 29862 8415 29863 8441
rect 29889 8415 30087 8441
rect 30113 8415 30114 8441
rect 29862 8414 30114 8415
rect 29862 8049 29890 8414
rect 29862 8023 29863 8049
rect 29889 8023 29890 8049
rect 29358 7657 29386 8022
rect 29862 8017 29890 8023
rect 30086 7993 30114 8414
rect 30086 7967 30087 7993
rect 30113 7967 30114 7993
rect 30086 7961 30114 7967
rect 30198 9281 30226 10262
rect 30198 9255 30199 9281
rect 30225 9255 30226 9281
rect 30198 9225 30226 9255
rect 30198 9199 30199 9225
rect 30225 9199 30226 9225
rect 30198 8834 30226 9199
rect 30198 8777 30226 8806
rect 30198 8751 30199 8777
rect 30225 8751 30226 8777
rect 29573 7854 30035 7859
rect 29573 7853 29582 7854
rect 29573 7827 29574 7853
rect 29573 7826 29582 7827
rect 29610 7826 29634 7854
rect 29662 7826 29686 7854
rect 29714 7853 29738 7854
rect 29766 7853 29790 7854
rect 29724 7827 29738 7853
rect 29786 7827 29790 7853
rect 29714 7826 29738 7827
rect 29766 7826 29790 7827
rect 29818 7853 29842 7854
rect 29870 7853 29894 7854
rect 29818 7827 29822 7853
rect 29870 7827 29884 7853
rect 29818 7826 29842 7827
rect 29870 7826 29894 7827
rect 29922 7826 29946 7854
rect 29974 7826 29998 7854
rect 30026 7853 30035 7854
rect 30034 7827 30035 7853
rect 30026 7826 30035 7827
rect 29573 7821 30035 7826
rect 29358 7631 29359 7657
rect 29385 7631 29386 7657
rect 28854 7265 28882 7271
rect 28854 7239 28855 7265
rect 28881 7239 28882 7265
rect 28854 6762 28882 7239
rect 28854 6481 28882 6734
rect 28854 6455 28855 6481
rect 28881 6455 28882 6481
rect 28854 6449 28882 6455
rect 29358 7265 29386 7631
rect 29358 7239 29359 7265
rect 29385 7239 29386 7265
rect 29358 6873 29386 7239
rect 30198 7713 30226 8751
rect 30198 7687 30199 7713
rect 30225 7687 30226 7713
rect 30198 7657 30226 7687
rect 30198 7631 30199 7657
rect 30225 7631 30226 7657
rect 30198 7265 30226 7631
rect 30198 7239 30199 7265
rect 30225 7239 30226 7265
rect 30198 7209 30226 7239
rect 30198 7183 30199 7209
rect 30225 7183 30226 7209
rect 29573 7070 30035 7075
rect 29573 7069 29582 7070
rect 29573 7043 29574 7069
rect 29573 7042 29582 7043
rect 29610 7042 29634 7070
rect 29662 7042 29686 7070
rect 29714 7069 29738 7070
rect 29766 7069 29790 7070
rect 29724 7043 29738 7069
rect 29786 7043 29790 7069
rect 29714 7042 29738 7043
rect 29766 7042 29790 7043
rect 29818 7069 29842 7070
rect 29870 7069 29894 7070
rect 29818 7043 29822 7069
rect 29870 7043 29884 7069
rect 29818 7042 29842 7043
rect 29870 7042 29894 7043
rect 29922 7042 29946 7070
rect 29974 7042 29998 7070
rect 30026 7069 30035 7070
rect 30034 7043 30035 7069
rect 30026 7042 30035 7043
rect 29573 7037 30035 7042
rect 29358 6847 29359 6873
rect 29385 6847 29386 6873
rect 29358 6762 29386 6847
rect 29358 6481 29386 6734
rect 29358 6455 29359 6481
rect 29385 6455 29386 6481
rect 29358 6089 29386 6455
rect 30198 6929 30226 7183
rect 30198 6903 30199 6929
rect 30225 6903 30226 6929
rect 30198 6873 30226 6903
rect 30198 6847 30199 6873
rect 30225 6847 30226 6873
rect 30198 6481 30226 6847
rect 30198 6455 30199 6481
rect 30225 6455 30226 6481
rect 30198 6425 30226 6455
rect 30198 6399 30199 6425
rect 30225 6399 30226 6425
rect 29573 6286 30035 6291
rect 29573 6285 29582 6286
rect 29573 6259 29574 6285
rect 29573 6258 29582 6259
rect 29610 6258 29634 6286
rect 29662 6258 29686 6286
rect 29714 6285 29738 6286
rect 29766 6285 29790 6286
rect 29724 6259 29738 6285
rect 29786 6259 29790 6285
rect 29714 6258 29738 6259
rect 29766 6258 29790 6259
rect 29818 6285 29842 6286
rect 29870 6285 29894 6286
rect 29818 6259 29822 6285
rect 29870 6259 29884 6285
rect 29818 6258 29842 6259
rect 29870 6258 29894 6259
rect 29922 6258 29946 6286
rect 29974 6258 29998 6286
rect 30026 6285 30035 6286
rect 30034 6259 30035 6285
rect 30026 6258 30035 6259
rect 29573 6253 30035 6258
rect 29358 6063 29359 6089
rect 29385 6063 29386 6089
rect 29358 5697 29386 6063
rect 29358 5671 29359 5697
rect 29385 5671 29386 5697
rect 29358 5306 29386 5671
rect 30198 6145 30226 6399
rect 30198 6119 30199 6145
rect 30225 6119 30226 6145
rect 30198 6089 30226 6119
rect 30198 6063 30199 6089
rect 30225 6063 30226 6089
rect 30198 5866 30226 6063
rect 30198 5697 30226 5838
rect 30198 5671 30199 5697
rect 30225 5671 30226 5697
rect 30198 5641 30226 5671
rect 30198 5615 30199 5641
rect 30225 5615 30226 5641
rect 29573 5502 30035 5507
rect 29573 5501 29582 5502
rect 29573 5475 29574 5501
rect 29573 5474 29582 5475
rect 29610 5474 29634 5502
rect 29662 5474 29686 5502
rect 29714 5501 29738 5502
rect 29766 5501 29790 5502
rect 29724 5475 29738 5501
rect 29786 5475 29790 5501
rect 29714 5474 29738 5475
rect 29766 5474 29790 5475
rect 29818 5501 29842 5502
rect 29870 5501 29894 5502
rect 29818 5475 29822 5501
rect 29870 5475 29884 5501
rect 29818 5474 29842 5475
rect 29870 5474 29894 5475
rect 29922 5474 29946 5502
rect 29974 5474 29998 5502
rect 30026 5501 30035 5502
rect 30034 5475 30035 5501
rect 30026 5474 30035 5475
rect 29573 5469 30035 5474
rect 29358 5259 29386 5278
rect 30198 5361 30226 5615
rect 30198 5335 30199 5361
rect 30225 5335 30226 5361
rect 30198 5305 30226 5335
rect 30198 5279 30199 5305
rect 30225 5279 30226 5305
rect 30198 5273 30226 5279
rect 30254 10066 30282 10071
rect 30142 5026 30170 5031
rect 29302 4913 29330 4919
rect 29302 4887 29303 4913
rect 29329 4887 29330 4913
rect 29302 4857 29330 4887
rect 30142 4913 30170 4998
rect 30142 4887 30143 4913
rect 30169 4887 30170 4913
rect 30142 4881 30170 4887
rect 29302 4831 29303 4857
rect 29329 4831 29330 4857
rect 29302 4522 29330 4831
rect 30030 4858 30058 4863
rect 30030 4811 30058 4830
rect 29573 4718 30035 4723
rect 29573 4717 29582 4718
rect 29573 4691 29574 4717
rect 29573 4690 29582 4691
rect 29610 4690 29634 4718
rect 29662 4690 29686 4718
rect 29714 4717 29738 4718
rect 29766 4717 29790 4718
rect 29724 4691 29738 4717
rect 29786 4691 29790 4717
rect 29714 4690 29738 4691
rect 29766 4690 29790 4691
rect 29818 4717 29842 4718
rect 29870 4717 29894 4718
rect 29818 4691 29822 4717
rect 29870 4691 29884 4717
rect 29818 4690 29842 4691
rect 29870 4690 29894 4691
rect 29922 4690 29946 4718
rect 29974 4690 29998 4718
rect 30026 4717 30035 4718
rect 30034 4691 30035 4717
rect 30026 4690 30035 4691
rect 29573 4685 30035 4690
rect 29414 4522 29442 4527
rect 29302 4521 29442 4522
rect 29302 4495 29303 4521
rect 29329 4495 29415 4521
rect 29441 4495 29442 4521
rect 29302 4494 29442 4495
rect 29302 4489 29330 4494
rect 28910 4242 28938 4247
rect 28910 4129 28938 4214
rect 28910 4103 28911 4129
rect 28937 4103 28938 4129
rect 28910 4097 28938 4103
rect 29414 4242 29442 4494
rect 28966 3737 28994 3743
rect 28966 3711 28967 3737
rect 28993 3711 28994 3737
rect 28966 2450 28994 3711
rect 28966 1778 28994 2422
rect 28966 1745 28994 1750
rect 29358 3345 29386 3351
rect 29358 3319 29359 3345
rect 29385 3319 29386 3345
rect 29358 3289 29386 3319
rect 29358 3263 29359 3289
rect 29385 3263 29386 3289
rect 29358 2954 29386 3263
rect 29358 2674 29386 2926
rect 29358 2561 29386 2646
rect 29358 2535 29359 2561
rect 29385 2535 29386 2561
rect 29358 2505 29386 2535
rect 29358 2479 29359 2505
rect 29385 2479 29386 2505
rect 29358 1777 29386 2479
rect 29414 2170 29442 4214
rect 30086 4129 30114 4135
rect 30086 4103 30087 4129
rect 30113 4103 30114 4129
rect 29573 3934 30035 3939
rect 29573 3933 29582 3934
rect 29573 3907 29574 3933
rect 29573 3906 29582 3907
rect 29610 3906 29634 3934
rect 29662 3906 29686 3934
rect 29714 3933 29738 3934
rect 29766 3933 29790 3934
rect 29724 3907 29738 3933
rect 29786 3907 29790 3933
rect 29714 3906 29738 3907
rect 29766 3906 29790 3907
rect 29818 3933 29842 3934
rect 29870 3933 29894 3934
rect 29818 3907 29822 3933
rect 29870 3907 29884 3933
rect 29818 3906 29842 3907
rect 29870 3906 29894 3907
rect 29922 3906 29946 3934
rect 29974 3906 29998 3934
rect 30026 3933 30035 3934
rect 30034 3907 30035 3933
rect 30026 3906 30035 3907
rect 29573 3901 30035 3906
rect 29694 3793 29722 3799
rect 29694 3767 29695 3793
rect 29721 3767 29722 3793
rect 29470 3738 29498 3743
rect 29694 3738 29722 3767
rect 29470 3737 29722 3738
rect 29470 3711 29471 3737
rect 29497 3711 29722 3737
rect 29470 3710 29722 3711
rect 29470 2954 29498 3710
rect 30030 3290 30058 3295
rect 30086 3290 30114 4103
rect 30058 3262 30114 3290
rect 30030 3243 30058 3262
rect 29573 3150 30035 3155
rect 29573 3149 29582 3150
rect 29573 3123 29574 3149
rect 29573 3122 29582 3123
rect 29610 3122 29634 3150
rect 29662 3122 29686 3150
rect 29714 3149 29738 3150
rect 29766 3149 29790 3150
rect 29724 3123 29738 3149
rect 29786 3123 29790 3149
rect 29714 3122 29738 3123
rect 29766 3122 29790 3123
rect 29818 3149 29842 3150
rect 29870 3149 29894 3150
rect 29818 3123 29822 3149
rect 29870 3123 29884 3149
rect 29818 3122 29842 3123
rect 29870 3122 29894 3123
rect 29922 3122 29946 3150
rect 29974 3122 29998 3150
rect 30026 3149 30035 3150
rect 30034 3123 30035 3149
rect 30026 3122 30035 3123
rect 29573 3117 30035 3122
rect 29470 2921 29498 2926
rect 29918 3009 29946 3015
rect 29918 2983 29919 3009
rect 29945 2983 29946 3009
rect 29918 2954 29946 2983
rect 29918 2907 29946 2926
rect 30086 3010 30114 3262
rect 30086 2561 30114 2982
rect 30086 2535 30087 2561
rect 30113 2535 30114 2561
rect 30086 2529 30114 2535
rect 30142 4074 30170 4079
rect 30142 3289 30170 4046
rect 30142 3263 30143 3289
rect 30169 3263 30170 3289
rect 30142 2618 30170 3263
rect 30142 2561 30170 2590
rect 30142 2535 30143 2561
rect 30169 2535 30170 2561
rect 30142 2529 30170 2535
rect 29573 2366 30035 2371
rect 29573 2365 29582 2366
rect 29573 2339 29574 2365
rect 29573 2338 29582 2339
rect 29610 2338 29634 2366
rect 29662 2338 29686 2366
rect 29714 2365 29738 2366
rect 29766 2365 29790 2366
rect 29724 2339 29738 2365
rect 29786 2339 29790 2365
rect 29714 2338 29738 2339
rect 29766 2338 29790 2339
rect 29818 2365 29842 2366
rect 29870 2365 29894 2366
rect 29818 2339 29822 2365
rect 29870 2339 29884 2365
rect 29818 2338 29842 2339
rect 29870 2338 29894 2339
rect 29922 2338 29946 2366
rect 29974 2338 29998 2366
rect 30026 2365 30035 2366
rect 30034 2339 30035 2365
rect 30026 2338 30035 2339
rect 29573 2333 30035 2338
rect 29414 2137 29442 2142
rect 29918 2225 29946 2231
rect 29918 2199 29919 2225
rect 29945 2199 29946 2225
rect 29918 2170 29946 2199
rect 29918 2123 29946 2142
rect 29358 1751 29359 1777
rect 29385 1751 29386 1777
rect 29358 1721 29386 1751
rect 29358 1695 29359 1721
rect 29385 1695 29386 1721
rect 29358 1689 29386 1695
rect 29573 1582 30035 1587
rect 29573 1581 29582 1582
rect 29573 1555 29574 1581
rect 29573 1554 29582 1555
rect 29610 1554 29634 1582
rect 29662 1554 29686 1582
rect 29714 1581 29738 1582
rect 29766 1581 29790 1582
rect 29724 1555 29738 1581
rect 29786 1555 29790 1581
rect 29714 1554 29738 1555
rect 29766 1554 29790 1555
rect 29818 1581 29842 1582
rect 29870 1581 29894 1582
rect 29818 1555 29822 1581
rect 29870 1555 29884 1581
rect 29818 1554 29842 1555
rect 29870 1554 29894 1555
rect 29922 1554 29946 1582
rect 29974 1554 29998 1582
rect 30026 1581 30035 1582
rect 30034 1555 30035 1581
rect 30026 1554 30035 1555
rect 29573 1549 30035 1554
rect 30254 882 30282 10038
rect 30310 10010 30338 10767
rect 30310 9977 30338 9982
rect 30702 10401 30730 10407
rect 30702 10375 30703 10401
rect 30729 10375 30730 10401
rect 30702 10010 30730 10375
rect 30758 10066 30786 11159
rect 31430 10849 31458 11942
rect 31598 11937 31626 11942
rect 31654 11913 31682 11942
rect 31654 11887 31655 11913
rect 31681 11887 31682 11913
rect 31654 11881 31682 11887
rect 31486 11634 31514 11639
rect 31486 11577 31514 11606
rect 31934 11634 31962 19614
rect 32270 19530 32298 19614
rect 32424 19600 32480 20000
rect 36974 19614 37282 19642
rect 32438 19530 32466 19600
rect 32270 19502 32466 19530
rect 32073 18438 32535 18443
rect 32073 18437 32082 18438
rect 32073 18411 32074 18437
rect 32073 18410 32082 18411
rect 32110 18410 32134 18438
rect 32162 18410 32186 18438
rect 32214 18437 32238 18438
rect 32266 18437 32290 18438
rect 32224 18411 32238 18437
rect 32286 18411 32290 18437
rect 32214 18410 32238 18411
rect 32266 18410 32290 18411
rect 32318 18437 32342 18438
rect 32370 18437 32394 18438
rect 32318 18411 32322 18437
rect 32370 18411 32384 18437
rect 32318 18410 32342 18411
rect 32370 18410 32394 18411
rect 32422 18410 32446 18438
rect 32474 18410 32498 18438
rect 32526 18437 32535 18438
rect 32534 18411 32535 18437
rect 32526 18410 32535 18411
rect 32073 18405 32535 18410
rect 34573 18046 35035 18051
rect 34573 18045 34582 18046
rect 34573 18019 34574 18045
rect 34573 18018 34582 18019
rect 34610 18018 34634 18046
rect 34662 18018 34686 18046
rect 34714 18045 34738 18046
rect 34766 18045 34790 18046
rect 34724 18019 34738 18045
rect 34786 18019 34790 18045
rect 34714 18018 34738 18019
rect 34766 18018 34790 18019
rect 34818 18045 34842 18046
rect 34870 18045 34894 18046
rect 34818 18019 34822 18045
rect 34870 18019 34884 18045
rect 34818 18018 34842 18019
rect 34870 18018 34894 18019
rect 34922 18018 34946 18046
rect 34974 18018 34998 18046
rect 35026 18045 35035 18046
rect 35034 18019 35035 18045
rect 35026 18018 35035 18019
rect 34573 18013 35035 18018
rect 32073 17654 32535 17659
rect 32073 17653 32082 17654
rect 32073 17627 32074 17653
rect 32073 17626 32082 17627
rect 32110 17626 32134 17654
rect 32162 17626 32186 17654
rect 32214 17653 32238 17654
rect 32266 17653 32290 17654
rect 32224 17627 32238 17653
rect 32286 17627 32290 17653
rect 32214 17626 32238 17627
rect 32266 17626 32290 17627
rect 32318 17653 32342 17654
rect 32370 17653 32394 17654
rect 32318 17627 32322 17653
rect 32370 17627 32384 17653
rect 32318 17626 32342 17627
rect 32370 17626 32394 17627
rect 32422 17626 32446 17654
rect 32474 17626 32498 17654
rect 32526 17653 32535 17654
rect 32534 17627 32535 17653
rect 32526 17626 32535 17627
rect 32073 17621 32535 17626
rect 34573 17262 35035 17267
rect 34573 17261 34582 17262
rect 34573 17235 34574 17261
rect 34573 17234 34582 17235
rect 34610 17234 34634 17262
rect 34662 17234 34686 17262
rect 34714 17261 34738 17262
rect 34766 17261 34790 17262
rect 34724 17235 34738 17261
rect 34786 17235 34790 17261
rect 34714 17234 34738 17235
rect 34766 17234 34790 17235
rect 34818 17261 34842 17262
rect 34870 17261 34894 17262
rect 34818 17235 34822 17261
rect 34870 17235 34884 17261
rect 34818 17234 34842 17235
rect 34870 17234 34894 17235
rect 34922 17234 34946 17262
rect 34974 17234 34998 17262
rect 35026 17261 35035 17262
rect 35034 17235 35035 17261
rect 35026 17234 35035 17235
rect 34573 17229 35035 17234
rect 32073 16870 32535 16875
rect 32073 16869 32082 16870
rect 32073 16843 32074 16869
rect 32073 16842 32082 16843
rect 32110 16842 32134 16870
rect 32162 16842 32186 16870
rect 32214 16869 32238 16870
rect 32266 16869 32290 16870
rect 32224 16843 32238 16869
rect 32286 16843 32290 16869
rect 32214 16842 32238 16843
rect 32266 16842 32290 16843
rect 32318 16869 32342 16870
rect 32370 16869 32394 16870
rect 32318 16843 32322 16869
rect 32370 16843 32384 16869
rect 32318 16842 32342 16843
rect 32370 16842 32394 16843
rect 32422 16842 32446 16870
rect 32474 16842 32498 16870
rect 32526 16869 32535 16870
rect 32534 16843 32535 16869
rect 32526 16842 32535 16843
rect 32073 16837 32535 16842
rect 34573 16478 35035 16483
rect 34573 16477 34582 16478
rect 34573 16451 34574 16477
rect 34573 16450 34582 16451
rect 34610 16450 34634 16478
rect 34662 16450 34686 16478
rect 34714 16477 34738 16478
rect 34766 16477 34790 16478
rect 34724 16451 34738 16477
rect 34786 16451 34790 16477
rect 34714 16450 34738 16451
rect 34766 16450 34790 16451
rect 34818 16477 34842 16478
rect 34870 16477 34894 16478
rect 34818 16451 34822 16477
rect 34870 16451 34884 16477
rect 34818 16450 34842 16451
rect 34870 16450 34894 16451
rect 34922 16450 34946 16478
rect 34974 16450 34998 16478
rect 35026 16477 35035 16478
rect 35034 16451 35035 16477
rect 35026 16450 35035 16451
rect 34573 16445 35035 16450
rect 32073 16086 32535 16091
rect 32073 16085 32082 16086
rect 32073 16059 32074 16085
rect 32073 16058 32082 16059
rect 32110 16058 32134 16086
rect 32162 16058 32186 16086
rect 32214 16085 32238 16086
rect 32266 16085 32290 16086
rect 32224 16059 32238 16085
rect 32286 16059 32290 16085
rect 32214 16058 32238 16059
rect 32266 16058 32290 16059
rect 32318 16085 32342 16086
rect 32370 16085 32394 16086
rect 32318 16059 32322 16085
rect 32370 16059 32384 16085
rect 32318 16058 32342 16059
rect 32370 16058 32394 16059
rect 32422 16058 32446 16086
rect 32474 16058 32498 16086
rect 32526 16085 32535 16086
rect 32534 16059 32535 16085
rect 32526 16058 32535 16059
rect 32073 16053 32535 16058
rect 34573 15694 35035 15699
rect 34573 15693 34582 15694
rect 34573 15667 34574 15693
rect 34573 15666 34582 15667
rect 34610 15666 34634 15694
rect 34662 15666 34686 15694
rect 34714 15693 34738 15694
rect 34766 15693 34790 15694
rect 34724 15667 34738 15693
rect 34786 15667 34790 15693
rect 34714 15666 34738 15667
rect 34766 15666 34790 15667
rect 34818 15693 34842 15694
rect 34870 15693 34894 15694
rect 34818 15667 34822 15693
rect 34870 15667 34884 15693
rect 34818 15666 34842 15667
rect 34870 15666 34894 15667
rect 34922 15666 34946 15694
rect 34974 15666 34998 15694
rect 35026 15693 35035 15694
rect 35034 15667 35035 15693
rect 35026 15666 35035 15667
rect 34573 15661 35035 15666
rect 32073 15302 32535 15307
rect 32073 15301 32082 15302
rect 32073 15275 32074 15301
rect 32073 15274 32082 15275
rect 32110 15274 32134 15302
rect 32162 15274 32186 15302
rect 32214 15301 32238 15302
rect 32266 15301 32290 15302
rect 32224 15275 32238 15301
rect 32286 15275 32290 15301
rect 32214 15274 32238 15275
rect 32266 15274 32290 15275
rect 32318 15301 32342 15302
rect 32370 15301 32394 15302
rect 32318 15275 32322 15301
rect 32370 15275 32384 15301
rect 32318 15274 32342 15275
rect 32370 15274 32394 15275
rect 32422 15274 32446 15302
rect 32474 15274 32498 15302
rect 32526 15301 32535 15302
rect 32534 15275 32535 15301
rect 32526 15274 32535 15275
rect 32073 15269 32535 15274
rect 34573 14910 35035 14915
rect 34573 14909 34582 14910
rect 34573 14883 34574 14909
rect 34573 14882 34582 14883
rect 34610 14882 34634 14910
rect 34662 14882 34686 14910
rect 34714 14909 34738 14910
rect 34766 14909 34790 14910
rect 34724 14883 34738 14909
rect 34786 14883 34790 14909
rect 34714 14882 34738 14883
rect 34766 14882 34790 14883
rect 34818 14909 34842 14910
rect 34870 14909 34894 14910
rect 34818 14883 34822 14909
rect 34870 14883 34884 14909
rect 34818 14882 34842 14883
rect 34870 14882 34894 14883
rect 34922 14882 34946 14910
rect 34974 14882 34998 14910
rect 35026 14909 35035 14910
rect 35034 14883 35035 14909
rect 35026 14882 35035 14883
rect 34573 14877 35035 14882
rect 32073 14518 32535 14523
rect 32073 14517 32082 14518
rect 32073 14491 32074 14517
rect 32073 14490 32082 14491
rect 32110 14490 32134 14518
rect 32162 14490 32186 14518
rect 32214 14517 32238 14518
rect 32266 14517 32290 14518
rect 32224 14491 32238 14517
rect 32286 14491 32290 14517
rect 32214 14490 32238 14491
rect 32266 14490 32290 14491
rect 32318 14517 32342 14518
rect 32370 14517 32394 14518
rect 32318 14491 32322 14517
rect 32370 14491 32384 14517
rect 32318 14490 32342 14491
rect 32370 14490 32394 14491
rect 32422 14490 32446 14518
rect 32474 14490 32498 14518
rect 32526 14517 32535 14518
rect 32534 14491 32535 14517
rect 32526 14490 32535 14491
rect 32073 14485 32535 14490
rect 34573 14126 35035 14131
rect 34573 14125 34582 14126
rect 34573 14099 34574 14125
rect 34573 14098 34582 14099
rect 34610 14098 34634 14126
rect 34662 14098 34686 14126
rect 34714 14125 34738 14126
rect 34766 14125 34790 14126
rect 34724 14099 34738 14125
rect 34786 14099 34790 14125
rect 34714 14098 34738 14099
rect 34766 14098 34790 14099
rect 34818 14125 34842 14126
rect 34870 14125 34894 14126
rect 34818 14099 34822 14125
rect 34870 14099 34884 14125
rect 34818 14098 34842 14099
rect 34870 14098 34894 14099
rect 34922 14098 34946 14126
rect 34974 14098 34998 14126
rect 35026 14125 35035 14126
rect 35034 14099 35035 14125
rect 35026 14098 35035 14099
rect 34573 14093 35035 14098
rect 32073 13734 32535 13739
rect 32073 13733 32082 13734
rect 32073 13707 32074 13733
rect 32073 13706 32082 13707
rect 32110 13706 32134 13734
rect 32162 13706 32186 13734
rect 32214 13733 32238 13734
rect 32266 13733 32290 13734
rect 32224 13707 32238 13733
rect 32286 13707 32290 13733
rect 32214 13706 32238 13707
rect 32266 13706 32290 13707
rect 32318 13733 32342 13734
rect 32370 13733 32394 13734
rect 32318 13707 32322 13733
rect 32370 13707 32384 13733
rect 32318 13706 32342 13707
rect 32370 13706 32394 13707
rect 32422 13706 32446 13734
rect 32474 13706 32498 13734
rect 32526 13733 32535 13734
rect 32534 13707 32535 13733
rect 32526 13706 32535 13707
rect 32073 13701 32535 13706
rect 34573 13342 35035 13347
rect 34573 13341 34582 13342
rect 34573 13315 34574 13341
rect 34573 13314 34582 13315
rect 34610 13314 34634 13342
rect 34662 13314 34686 13342
rect 34714 13341 34738 13342
rect 34766 13341 34790 13342
rect 34724 13315 34738 13341
rect 34786 13315 34790 13341
rect 34714 13314 34738 13315
rect 34766 13314 34790 13315
rect 34818 13341 34842 13342
rect 34870 13341 34894 13342
rect 34818 13315 34822 13341
rect 34870 13315 34884 13341
rect 34818 13314 34842 13315
rect 34870 13314 34894 13315
rect 34922 13314 34946 13342
rect 34974 13314 34998 13342
rect 35026 13341 35035 13342
rect 35034 13315 35035 13341
rect 35026 13314 35035 13315
rect 34573 13309 35035 13314
rect 32073 12950 32535 12955
rect 32073 12949 32082 12950
rect 32073 12923 32074 12949
rect 32073 12922 32082 12923
rect 32110 12922 32134 12950
rect 32162 12922 32186 12950
rect 32214 12949 32238 12950
rect 32266 12949 32290 12950
rect 32224 12923 32238 12949
rect 32286 12923 32290 12949
rect 32214 12922 32238 12923
rect 32266 12922 32290 12923
rect 32318 12949 32342 12950
rect 32370 12949 32394 12950
rect 32318 12923 32322 12949
rect 32370 12923 32384 12949
rect 32318 12922 32342 12923
rect 32370 12922 32394 12923
rect 32422 12922 32446 12950
rect 32474 12922 32498 12950
rect 32526 12949 32535 12950
rect 32534 12923 32535 12949
rect 32526 12922 32535 12923
rect 32073 12917 32535 12922
rect 34573 12558 35035 12563
rect 34573 12557 34582 12558
rect 34573 12531 34574 12557
rect 34573 12530 34582 12531
rect 34610 12530 34634 12558
rect 34662 12530 34686 12558
rect 34714 12557 34738 12558
rect 34766 12557 34790 12558
rect 34724 12531 34738 12557
rect 34786 12531 34790 12557
rect 34714 12530 34738 12531
rect 34766 12530 34790 12531
rect 34818 12557 34842 12558
rect 34870 12557 34894 12558
rect 34818 12531 34822 12557
rect 34870 12531 34884 12557
rect 34818 12530 34842 12531
rect 34870 12530 34894 12531
rect 34922 12530 34946 12558
rect 34974 12530 34998 12558
rect 35026 12557 35035 12558
rect 35034 12531 35035 12557
rect 35026 12530 35035 12531
rect 34573 12525 35035 12530
rect 32073 12166 32535 12171
rect 32073 12165 32082 12166
rect 32073 12139 32074 12165
rect 32073 12138 32082 12139
rect 32110 12138 32134 12166
rect 32162 12138 32186 12166
rect 32214 12165 32238 12166
rect 32266 12165 32290 12166
rect 32224 12139 32238 12165
rect 32286 12139 32290 12165
rect 32214 12138 32238 12139
rect 32266 12138 32290 12139
rect 32318 12165 32342 12166
rect 32370 12165 32394 12166
rect 32318 12139 32322 12165
rect 32370 12139 32384 12165
rect 32318 12138 32342 12139
rect 32370 12138 32394 12139
rect 32422 12138 32446 12166
rect 32474 12138 32498 12166
rect 32526 12165 32535 12166
rect 32534 12139 32535 12165
rect 32526 12138 32535 12139
rect 32073 12133 32535 12138
rect 31934 11601 31962 11606
rect 32438 11969 32466 11975
rect 32438 11943 32439 11969
rect 32465 11943 32466 11969
rect 31486 11551 31487 11577
rect 31513 11551 31514 11577
rect 31486 11186 31514 11551
rect 32438 11578 32466 11943
rect 32830 11970 32858 11975
rect 32830 11923 32858 11942
rect 33110 11970 33138 11975
rect 33110 11914 33138 11942
rect 33110 11913 33194 11914
rect 33110 11887 33111 11913
rect 33137 11887 33194 11913
rect 33110 11886 33194 11887
rect 33110 11881 33138 11886
rect 32438 11545 32466 11550
rect 32774 11578 32802 11583
rect 32073 11382 32535 11387
rect 32073 11381 32082 11382
rect 32073 11355 32074 11381
rect 32073 11354 32082 11355
rect 32110 11354 32134 11382
rect 32162 11354 32186 11382
rect 32214 11381 32238 11382
rect 32266 11381 32290 11382
rect 32224 11355 32238 11381
rect 32286 11355 32290 11381
rect 32214 11354 32238 11355
rect 32266 11354 32290 11355
rect 32318 11381 32342 11382
rect 32370 11381 32394 11382
rect 32318 11355 32322 11381
rect 32370 11355 32384 11381
rect 32318 11354 32342 11355
rect 32370 11354 32394 11355
rect 32422 11354 32446 11382
rect 32474 11354 32498 11382
rect 32526 11381 32535 11382
rect 32534 11355 32535 11381
rect 32526 11354 32535 11355
rect 32073 11349 32535 11354
rect 32438 11186 32466 11191
rect 31486 11185 31682 11186
rect 31486 11159 31487 11185
rect 31513 11159 31682 11185
rect 31486 11158 31682 11159
rect 31486 11153 31514 11158
rect 31430 10823 31431 10849
rect 31457 10823 31458 10849
rect 31430 10793 31458 10823
rect 31430 10767 31431 10793
rect 31457 10767 31458 10793
rect 31262 10402 31290 10407
rect 31430 10402 31458 10767
rect 30758 10033 30786 10038
rect 31094 10401 31458 10402
rect 31094 10375 31263 10401
rect 31289 10375 31431 10401
rect 31457 10375 31458 10401
rect 31094 10374 31458 10375
rect 30702 9977 30730 9982
rect 30814 10010 30842 10015
rect 30814 9730 30842 9982
rect 30814 9697 30842 9702
rect 31094 9898 31122 10374
rect 31262 10369 31290 10374
rect 31430 10369 31458 10374
rect 31654 11129 31682 11158
rect 32438 11139 32466 11158
rect 32774 11186 32802 11550
rect 33166 11578 33194 11886
rect 34573 11774 35035 11779
rect 34573 11773 34582 11774
rect 34573 11747 34574 11773
rect 34573 11746 34582 11747
rect 34610 11746 34634 11774
rect 34662 11746 34686 11774
rect 34714 11773 34738 11774
rect 34766 11773 34790 11774
rect 34724 11747 34738 11773
rect 34786 11747 34790 11773
rect 34714 11746 34738 11747
rect 34766 11746 34790 11747
rect 34818 11773 34842 11774
rect 34870 11773 34894 11774
rect 34818 11747 34822 11773
rect 34870 11747 34884 11773
rect 34818 11746 34842 11747
rect 34870 11746 34894 11747
rect 34922 11746 34946 11774
rect 34974 11746 34998 11774
rect 35026 11773 35035 11774
rect 35034 11747 35035 11773
rect 35026 11746 35035 11747
rect 34573 11741 35035 11746
rect 33166 11512 33194 11550
rect 33614 11578 33642 11583
rect 33614 11531 33642 11550
rect 34510 11578 34538 11583
rect 34510 11242 34538 11550
rect 31654 11103 31655 11129
rect 31681 11103 31682 11129
rect 31654 10094 31682 11103
rect 32774 10793 32802 11158
rect 33110 11185 33138 11191
rect 33110 11159 33111 11185
rect 33137 11159 33138 11185
rect 33110 11129 33138 11159
rect 33110 11103 33111 11129
rect 33137 11103 33138 11129
rect 33110 10794 33138 11103
rect 33166 10794 33194 10799
rect 33390 10794 33418 10799
rect 32774 10767 32775 10793
rect 32801 10767 32802 10793
rect 32073 10598 32535 10603
rect 32073 10597 32082 10598
rect 32073 10571 32074 10597
rect 32073 10570 32082 10571
rect 32110 10570 32134 10598
rect 32162 10570 32186 10598
rect 32214 10597 32238 10598
rect 32266 10597 32290 10598
rect 32224 10571 32238 10597
rect 32286 10571 32290 10597
rect 32214 10570 32238 10571
rect 32266 10570 32290 10571
rect 32318 10597 32342 10598
rect 32370 10597 32394 10598
rect 32318 10571 32322 10597
rect 32370 10571 32384 10597
rect 32318 10570 32342 10571
rect 32370 10570 32394 10571
rect 32422 10570 32446 10598
rect 32474 10570 32498 10598
rect 32526 10597 32535 10598
rect 32534 10571 32535 10597
rect 32526 10570 32535 10571
rect 32073 10565 32535 10570
rect 31486 10066 31682 10094
rect 32158 10401 32186 10407
rect 32158 10375 32159 10401
rect 32185 10375 32186 10401
rect 32158 10066 32186 10375
rect 31374 10010 31402 10015
rect 31486 10010 31514 10066
rect 32158 10033 32186 10038
rect 31374 10009 31514 10010
rect 31374 9983 31375 10009
rect 31401 9983 31487 10009
rect 31513 9983 31514 10009
rect 31374 9982 31514 9983
rect 31374 9977 31402 9982
rect 30982 9617 31010 9623
rect 30982 9591 30983 9617
rect 31009 9591 31010 9617
rect 30982 9226 31010 9591
rect 30982 8834 31010 9198
rect 31094 9618 31122 9870
rect 31150 9618 31178 9623
rect 31094 9617 31178 9618
rect 31094 9591 31151 9617
rect 31177 9591 31178 9617
rect 31094 9590 31178 9591
rect 31094 9226 31122 9590
rect 31150 9585 31178 9590
rect 31374 9618 31402 9623
rect 31150 9226 31178 9231
rect 31374 9226 31402 9590
rect 31094 9225 31402 9226
rect 31094 9199 31151 9225
rect 31177 9199 31375 9225
rect 31401 9199 31402 9225
rect 31094 9198 31402 9199
rect 30982 8833 31066 8834
rect 30982 8807 30983 8833
rect 31009 8807 31066 8833
rect 30982 8806 31066 8807
rect 30982 8801 31010 8806
rect 31038 8442 31066 8806
rect 31038 8395 31066 8414
rect 30758 8049 30786 8055
rect 30758 8023 30759 8049
rect 30785 8023 30786 8049
rect 30758 7657 30786 8023
rect 31094 8050 31122 9198
rect 31150 9193 31178 9198
rect 31374 9193 31402 9198
rect 31150 8834 31178 8839
rect 31150 8787 31178 8806
rect 31374 8834 31402 8839
rect 31430 8834 31458 9982
rect 31486 9977 31514 9982
rect 32774 9898 32802 10767
rect 32886 10793 33418 10794
rect 32886 10767 33167 10793
rect 33193 10767 33391 10793
rect 33417 10767 33418 10793
rect 32886 10766 33418 10767
rect 32830 10066 32858 10071
rect 32830 10009 32858 10038
rect 32830 9983 32831 10009
rect 32857 9983 32858 10009
rect 32830 9977 32858 9983
rect 32886 10010 32914 10766
rect 33166 10761 33194 10766
rect 33390 10761 33418 10766
rect 34454 10793 34482 10799
rect 34454 10767 34455 10793
rect 34481 10767 34482 10793
rect 33110 10401 33138 10407
rect 33110 10375 33111 10401
rect 33137 10375 33138 10401
rect 33110 10345 33138 10375
rect 33110 10319 33111 10345
rect 33137 10319 33138 10345
rect 33110 10094 33138 10319
rect 32073 9814 32535 9819
rect 32073 9813 32082 9814
rect 32073 9787 32074 9813
rect 32073 9786 32082 9787
rect 32110 9786 32134 9814
rect 32162 9786 32186 9814
rect 32214 9813 32238 9814
rect 32266 9813 32290 9814
rect 32224 9787 32238 9813
rect 32286 9787 32290 9813
rect 32214 9786 32238 9787
rect 32266 9786 32290 9787
rect 32318 9813 32342 9814
rect 32370 9813 32394 9814
rect 32318 9787 32322 9813
rect 32370 9787 32384 9813
rect 32318 9786 32342 9787
rect 32370 9786 32394 9787
rect 32422 9786 32446 9814
rect 32474 9786 32498 9814
rect 32526 9813 32535 9814
rect 32534 9787 32535 9813
rect 32526 9786 32535 9787
rect 32073 9781 32535 9786
rect 31402 8806 31458 8834
rect 31990 9730 32018 9735
rect 31990 8834 32018 9702
rect 32158 9730 32186 9735
rect 32158 9617 32186 9702
rect 32158 9591 32159 9617
rect 32185 9591 32186 9617
rect 32158 9585 32186 9591
rect 32073 9030 32535 9035
rect 32073 9029 32082 9030
rect 32073 9003 32074 9029
rect 32073 9002 32082 9003
rect 32110 9002 32134 9030
rect 32162 9002 32186 9030
rect 32214 9029 32238 9030
rect 32266 9029 32290 9030
rect 32224 9003 32238 9029
rect 32286 9003 32290 9029
rect 32214 9002 32238 9003
rect 32266 9002 32290 9003
rect 32318 9029 32342 9030
rect 32370 9029 32394 9030
rect 32318 9003 32322 9029
rect 32370 9003 32384 9029
rect 32318 9002 32342 9003
rect 32370 9002 32394 9003
rect 32422 9002 32446 9030
rect 32474 9002 32498 9030
rect 32526 9029 32535 9030
rect 32534 9003 32535 9029
rect 32526 9002 32535 9003
rect 32073 8997 32535 9002
rect 32158 8834 32186 8839
rect 31990 8833 32186 8834
rect 31990 8807 32159 8833
rect 32185 8807 32186 8833
rect 31990 8806 32186 8807
rect 31374 8787 31402 8806
rect 31430 8498 31458 8806
rect 31318 8442 31346 8447
rect 31430 8442 31458 8470
rect 31318 8441 31458 8442
rect 31318 8415 31319 8441
rect 31345 8415 31431 8441
rect 31457 8415 31458 8441
rect 31318 8414 31458 8415
rect 31318 8409 31346 8414
rect 31430 8409 31458 8414
rect 31934 8442 31962 8447
rect 31150 8050 31178 8055
rect 31374 8050 31402 8055
rect 31094 8049 31402 8050
rect 31094 8023 31151 8049
rect 31177 8023 31375 8049
rect 31401 8023 31402 8049
rect 31094 8022 31402 8023
rect 31150 8017 31178 8022
rect 30758 7631 30759 7657
rect 30785 7631 30786 7657
rect 30758 7574 30786 7631
rect 31206 7657 31234 8022
rect 31206 7631 31207 7657
rect 31233 7631 31234 7657
rect 31206 7625 31234 7631
rect 31374 7657 31402 8022
rect 31934 8050 31962 8414
rect 32158 8442 32186 8806
rect 32158 8409 32186 8414
rect 32718 8442 32746 8447
rect 32718 8395 32746 8414
rect 32073 8246 32535 8251
rect 32073 8245 32082 8246
rect 32073 8219 32074 8245
rect 32073 8218 32082 8219
rect 32110 8218 32134 8246
rect 32162 8218 32186 8246
rect 32214 8245 32238 8246
rect 32266 8245 32290 8246
rect 32224 8219 32238 8245
rect 32286 8219 32290 8245
rect 32214 8218 32238 8219
rect 32266 8218 32290 8219
rect 32318 8245 32342 8246
rect 32370 8245 32394 8246
rect 32318 8219 32322 8245
rect 32370 8219 32384 8245
rect 32318 8218 32342 8219
rect 32370 8218 32394 8219
rect 32422 8218 32446 8246
rect 32474 8218 32498 8246
rect 32526 8245 32535 8246
rect 32534 8219 32535 8245
rect 32526 8218 32535 8219
rect 32073 8213 32535 8218
rect 31934 8017 31962 8022
rect 32438 8050 32466 8055
rect 31374 7631 31375 7657
rect 31401 7631 31402 7657
rect 31374 7574 31402 7631
rect 32438 7602 32466 8022
rect 32774 7994 32802 9870
rect 32830 9618 32858 9623
rect 32830 9571 32858 9590
rect 32830 9225 32858 9231
rect 32830 9199 32831 9225
rect 32857 9199 32858 9225
rect 32830 9170 32858 9199
rect 32830 9137 32858 9142
rect 32886 8890 32914 9982
rect 32942 10066 32970 10071
rect 32942 9450 32970 10038
rect 32942 9417 32970 9422
rect 33054 10066 33138 10094
rect 34454 10402 34482 10767
rect 34510 10794 34538 11214
rect 35126 11242 35154 11247
rect 34958 11186 34986 11191
rect 34958 11139 34986 11158
rect 35126 11185 35154 11214
rect 35126 11159 35127 11185
rect 35153 11159 35154 11185
rect 35126 11153 35154 11159
rect 35350 11242 35378 11247
rect 35350 11185 35378 11214
rect 35350 11159 35351 11185
rect 35377 11159 35378 11185
rect 34573 10990 35035 10995
rect 34573 10989 34582 10990
rect 34573 10963 34574 10989
rect 34573 10962 34582 10963
rect 34610 10962 34634 10990
rect 34662 10962 34686 10990
rect 34714 10989 34738 10990
rect 34766 10989 34790 10990
rect 34724 10963 34738 10989
rect 34786 10963 34790 10989
rect 34714 10962 34738 10963
rect 34766 10962 34790 10963
rect 34818 10989 34842 10990
rect 34870 10989 34894 10990
rect 34818 10963 34822 10989
rect 34870 10963 34884 10989
rect 34818 10962 34842 10963
rect 34870 10962 34894 10963
rect 34922 10962 34946 10990
rect 34974 10962 34998 10990
rect 35026 10989 35035 10990
rect 35034 10963 35035 10989
rect 35026 10962 35035 10963
rect 34573 10957 35035 10962
rect 34622 10794 34650 10799
rect 34846 10794 34874 10799
rect 34510 10793 34874 10794
rect 34510 10767 34623 10793
rect 34649 10767 34847 10793
rect 34873 10767 34874 10793
rect 34510 10766 34874 10767
rect 34622 10761 34650 10766
rect 34846 10761 34874 10766
rect 34454 10122 34482 10374
rect 34958 10402 34986 10407
rect 34958 10355 34986 10374
rect 35238 10402 35266 10407
rect 35350 10402 35378 11159
rect 35238 10401 35378 10402
rect 35238 10375 35239 10401
rect 35265 10375 35351 10401
rect 35377 10375 35378 10401
rect 35238 10374 35378 10375
rect 35238 10369 35266 10374
rect 35350 10346 35378 10374
rect 36134 11186 36162 11191
rect 36134 10514 36162 11158
rect 36694 10793 36722 10799
rect 36694 10767 36695 10793
rect 36721 10767 36722 10793
rect 36694 10738 36722 10767
rect 36694 10705 36722 10710
rect 36134 10486 36442 10514
rect 36134 10401 36162 10486
rect 36134 10375 36135 10401
rect 36161 10375 36162 10401
rect 36134 10369 36162 10375
rect 36246 10402 36274 10407
rect 35350 10313 35378 10318
rect 34573 10206 35035 10211
rect 34573 10205 34582 10206
rect 34573 10179 34574 10205
rect 34573 10178 34582 10179
rect 34610 10178 34634 10206
rect 34662 10178 34686 10206
rect 34714 10205 34738 10206
rect 34766 10205 34790 10206
rect 34724 10179 34738 10205
rect 34786 10179 34790 10205
rect 34714 10178 34738 10179
rect 34766 10178 34790 10179
rect 34818 10205 34842 10206
rect 34870 10205 34894 10206
rect 34818 10179 34822 10205
rect 34870 10179 34884 10205
rect 34818 10178 34842 10179
rect 34870 10178 34894 10179
rect 34922 10178 34946 10206
rect 34974 10178 34998 10206
rect 35026 10205 35035 10206
rect 35034 10179 35035 10205
rect 35026 10178 35035 10179
rect 34573 10173 35035 10178
rect 34454 10089 34482 10094
rect 32886 8857 32914 8862
rect 32774 7961 32802 7966
rect 32830 8833 32858 8839
rect 32830 8807 32831 8833
rect 32857 8807 32858 8833
rect 32830 8778 32858 8807
rect 33054 8778 33082 10066
rect 33166 10009 33194 10015
rect 33166 9983 33167 10009
rect 33193 9983 33194 10009
rect 33110 9618 33138 9623
rect 33110 9562 33138 9590
rect 33166 9562 33194 9983
rect 33110 9561 33194 9562
rect 33110 9535 33111 9561
rect 33137 9535 33194 9561
rect 33110 9534 33194 9535
rect 33110 9529 33138 9534
rect 33166 9225 33194 9534
rect 33166 9199 33167 9225
rect 33193 9199 33194 9225
rect 33110 8778 33138 8783
rect 33054 8750 33110 8778
rect 32830 8498 32858 8750
rect 33110 8731 33138 8750
rect 30758 7546 30954 7574
rect 31374 7546 31626 7574
rect 32438 7569 32466 7574
rect 32606 7602 32634 7607
rect 30926 7265 30954 7546
rect 30926 7239 30927 7265
rect 30953 7239 30954 7265
rect 30926 6874 30954 7239
rect 31598 7265 31626 7546
rect 32073 7462 32535 7467
rect 32073 7461 32082 7462
rect 32073 7435 32074 7461
rect 32073 7434 32082 7435
rect 32110 7434 32134 7462
rect 32162 7434 32186 7462
rect 32214 7461 32238 7462
rect 32266 7461 32290 7462
rect 32224 7435 32238 7461
rect 32286 7435 32290 7461
rect 32214 7434 32238 7435
rect 32266 7434 32290 7435
rect 32318 7461 32342 7462
rect 32370 7461 32394 7462
rect 32318 7435 32322 7461
rect 32370 7435 32384 7461
rect 32318 7434 32342 7435
rect 32370 7434 32394 7435
rect 32422 7434 32446 7462
rect 32474 7434 32498 7462
rect 32526 7461 32535 7462
rect 32534 7435 32535 7461
rect 32526 7434 32535 7435
rect 32073 7429 32535 7434
rect 31598 7239 31599 7265
rect 31625 7239 31626 7265
rect 31598 7210 31626 7239
rect 32438 7266 32466 7271
rect 32606 7266 32634 7574
rect 32438 7265 32634 7266
rect 32438 7239 32439 7265
rect 32465 7239 32634 7265
rect 32438 7238 32634 7239
rect 32830 7266 32858 8470
rect 33166 8441 33194 9199
rect 33166 8415 33167 8441
rect 33193 8415 33194 8441
rect 33166 8386 33194 8415
rect 33166 8049 33194 8358
rect 33614 10009 33642 10015
rect 33614 9983 33615 10009
rect 33641 9983 33642 10009
rect 33614 9225 33642 9983
rect 34454 10009 34482 10015
rect 34454 9983 34455 10009
rect 34481 9983 34482 10009
rect 34454 9898 34482 9983
rect 34622 10010 34650 10015
rect 34622 9963 34650 9982
rect 34846 10010 34874 10015
rect 34846 9963 34874 9982
rect 35126 10010 35154 10015
rect 34454 9506 34482 9870
rect 34454 9473 34482 9478
rect 34958 9617 34986 9623
rect 34958 9591 34959 9617
rect 34985 9591 34986 9617
rect 34958 9506 34986 9591
rect 35126 9618 35154 9982
rect 35350 9618 35378 9623
rect 35126 9617 35350 9618
rect 35126 9591 35127 9617
rect 35153 9591 35350 9617
rect 35126 9590 35350 9591
rect 36246 9618 36274 10374
rect 36414 9954 36442 10486
rect 36414 9921 36442 9926
rect 36694 10009 36722 10015
rect 36694 9983 36695 10009
rect 36721 9983 36722 10009
rect 36694 9954 36722 9983
rect 36694 9921 36722 9926
rect 36414 9618 36442 9623
rect 36246 9617 36722 9618
rect 36246 9591 36415 9617
rect 36441 9591 36722 9617
rect 36246 9590 36722 9591
rect 35126 9585 35154 9590
rect 35350 9552 35378 9590
rect 36414 9585 36442 9590
rect 34958 9473 34986 9478
rect 36414 9506 36442 9511
rect 33614 9199 33615 9225
rect 33641 9199 33642 9225
rect 33614 8441 33642 9199
rect 33614 8415 33615 8441
rect 33641 8415 33642 8441
rect 33614 8386 33642 8415
rect 34174 9450 34202 9455
rect 34174 9282 34202 9422
rect 34573 9422 35035 9427
rect 34573 9421 34582 9422
rect 34573 9395 34574 9421
rect 34573 9394 34582 9395
rect 34610 9394 34634 9422
rect 34662 9394 34686 9422
rect 34714 9421 34738 9422
rect 34766 9421 34790 9422
rect 34724 9395 34738 9421
rect 34786 9395 34790 9421
rect 34714 9394 34738 9395
rect 34766 9394 34790 9395
rect 34818 9421 34842 9422
rect 34870 9421 34894 9422
rect 34818 9395 34822 9421
rect 34870 9395 34884 9421
rect 34818 9394 34842 9395
rect 34870 9394 34894 9395
rect 34922 9394 34946 9422
rect 34974 9394 34998 9422
rect 35026 9421 35035 9422
rect 35034 9395 35035 9421
rect 35026 9394 35035 9395
rect 34573 9389 35035 9394
rect 34174 9225 34202 9254
rect 34174 9199 34175 9225
rect 34201 9199 34202 9225
rect 34174 8441 34202 9199
rect 34678 9282 34706 9287
rect 34678 8834 34706 9254
rect 34510 8833 34706 8834
rect 34510 8807 34679 8833
rect 34705 8807 34706 8833
rect 34510 8806 34706 8807
rect 34174 8415 34175 8441
rect 34201 8415 34202 8441
rect 34174 8409 34202 8415
rect 34398 8442 34426 8447
rect 33614 8353 33642 8358
rect 33166 8023 33167 8049
rect 33193 8023 33194 8049
rect 33166 7993 33194 8023
rect 33614 8050 33642 8055
rect 33726 8050 33754 8055
rect 33614 8049 33754 8050
rect 33614 8023 33615 8049
rect 33641 8023 33727 8049
rect 33753 8023 33754 8049
rect 33614 8022 33754 8023
rect 33614 8017 33642 8022
rect 33166 7967 33167 7993
rect 33193 7967 33194 7993
rect 32438 7233 32466 7238
rect 32830 7233 32858 7238
rect 32998 7657 33026 7663
rect 32998 7631 32999 7657
rect 33025 7631 33026 7657
rect 32998 7602 33026 7631
rect 31654 7210 31682 7215
rect 31598 7209 31682 7210
rect 31598 7183 31655 7209
rect 31681 7183 31682 7209
rect 31598 7182 31682 7183
rect 31598 6929 31626 7182
rect 31654 7177 31682 7182
rect 31598 6903 31599 6929
rect 31625 6903 31626 6929
rect 30926 6873 31010 6874
rect 30926 6847 30927 6873
rect 30953 6847 31010 6873
rect 30926 6846 31010 6847
rect 30926 6841 30954 6846
rect 30982 6481 31010 6846
rect 31598 6873 31626 6903
rect 31598 6847 31599 6873
rect 31625 6847 31626 6873
rect 31598 6841 31626 6847
rect 32998 6873 33026 7574
rect 32998 6847 32999 6873
rect 33025 6847 33026 6873
rect 32998 6762 33026 6847
rect 32998 6729 33026 6734
rect 33166 7658 33194 7967
rect 33390 7658 33418 7663
rect 33166 7657 33390 7658
rect 33166 7631 33167 7657
rect 33193 7631 33390 7657
rect 33166 7630 33390 7631
rect 32073 6678 32535 6683
rect 32073 6677 32082 6678
rect 32073 6651 32074 6677
rect 32073 6650 32082 6651
rect 32110 6650 32134 6678
rect 32162 6650 32186 6678
rect 32214 6677 32238 6678
rect 32266 6677 32290 6678
rect 32224 6651 32238 6677
rect 32286 6651 32290 6677
rect 32214 6650 32238 6651
rect 32266 6650 32290 6651
rect 32318 6677 32342 6678
rect 32370 6677 32394 6678
rect 32318 6651 32322 6677
rect 32370 6651 32384 6677
rect 32318 6650 32342 6651
rect 32370 6650 32394 6651
rect 32422 6650 32446 6678
rect 32474 6650 32498 6678
rect 32526 6677 32535 6678
rect 32534 6651 32535 6677
rect 32526 6650 32535 6651
rect 32073 6645 32535 6650
rect 30982 6455 30983 6481
rect 31009 6455 31010 6481
rect 30926 6090 30954 6095
rect 30982 6090 31010 6455
rect 30926 6089 31010 6090
rect 30926 6063 30927 6089
rect 30953 6063 31010 6089
rect 30926 6062 31010 6063
rect 30926 6057 30954 6062
rect 30982 5697 31010 6062
rect 30982 5671 30983 5697
rect 31009 5671 31010 5697
rect 30926 5306 30954 5311
rect 30982 5306 31010 5671
rect 31822 6481 31850 6487
rect 31822 6455 31823 6481
rect 31849 6455 31850 6481
rect 31822 6425 31850 6455
rect 32438 6482 32466 6487
rect 33166 6482 33194 7630
rect 33390 7592 33418 7630
rect 33726 7574 33754 8022
rect 33894 7994 33922 7999
rect 33894 7993 33978 7994
rect 33894 7967 33895 7993
rect 33921 7967 33978 7993
rect 33894 7966 33978 7967
rect 33894 7961 33922 7966
rect 33726 7546 33810 7574
rect 33334 7266 33362 7271
rect 33334 7209 33362 7238
rect 33782 7265 33810 7546
rect 33782 7239 33783 7265
rect 33809 7239 33810 7265
rect 33334 7183 33335 7209
rect 33361 7183 33362 7209
rect 33334 6762 33362 7183
rect 33334 6729 33362 6734
rect 33614 7209 33642 7215
rect 33614 7183 33615 7209
rect 33641 7183 33642 7209
rect 33334 6482 33362 6487
rect 32438 6481 32746 6482
rect 32438 6455 32439 6481
rect 32465 6455 32746 6481
rect 32438 6454 32746 6455
rect 33166 6481 33362 6482
rect 33166 6455 33335 6481
rect 33361 6455 33362 6481
rect 33166 6454 33362 6455
rect 32438 6449 32466 6454
rect 31822 6399 31823 6425
rect 31849 6399 31850 6425
rect 31822 6145 31850 6399
rect 31822 6119 31823 6145
rect 31849 6119 31850 6145
rect 31822 6089 31850 6119
rect 31822 6063 31823 6089
rect 31849 6063 31850 6089
rect 31822 5866 31850 6063
rect 32718 6089 32746 6454
rect 33334 6425 33362 6454
rect 33334 6399 33335 6425
rect 33361 6399 33362 6425
rect 32718 6063 32719 6089
rect 32745 6063 32746 6089
rect 32073 5894 32535 5899
rect 32073 5893 32082 5894
rect 32073 5867 32074 5893
rect 32073 5866 32082 5867
rect 32110 5866 32134 5894
rect 32162 5866 32186 5894
rect 32214 5893 32238 5894
rect 32266 5893 32290 5894
rect 32224 5867 32238 5893
rect 32286 5867 32290 5893
rect 32214 5866 32238 5867
rect 32266 5866 32290 5867
rect 32318 5893 32342 5894
rect 32370 5893 32394 5894
rect 32318 5867 32322 5893
rect 32370 5867 32384 5893
rect 32318 5866 32342 5867
rect 32370 5866 32394 5867
rect 32422 5866 32446 5894
rect 32474 5866 32498 5894
rect 32526 5893 32535 5894
rect 32534 5867 32535 5893
rect 32526 5866 32535 5867
rect 32073 5861 32535 5866
rect 31822 5698 31850 5838
rect 31878 5698 31906 5703
rect 31822 5697 31906 5698
rect 31822 5671 31879 5697
rect 31905 5671 31906 5697
rect 31822 5670 31906 5671
rect 31878 5641 31906 5670
rect 32438 5698 32466 5703
rect 32438 5651 32466 5670
rect 32718 5698 32746 6063
rect 33278 6090 33306 6095
rect 33334 6090 33362 6399
rect 33390 6090 33418 6095
rect 33278 6089 33418 6090
rect 33278 6063 33279 6089
rect 33305 6063 33391 6089
rect 33417 6063 33418 6089
rect 33278 6062 33418 6063
rect 33278 6057 33306 6062
rect 31878 5615 31879 5641
rect 31905 5615 31906 5641
rect 30954 5278 31010 5306
rect 30926 5240 30954 5278
rect 30366 5026 30394 5031
rect 30366 4913 30394 4998
rect 30366 4887 30367 4913
rect 30393 4887 30394 4913
rect 30366 4881 30394 4887
rect 30982 4913 31010 5278
rect 31822 5361 31850 5367
rect 31822 5335 31823 5361
rect 31849 5335 31850 5361
rect 31822 5306 31850 5335
rect 31878 5306 31906 5615
rect 31822 5305 31906 5306
rect 31822 5279 31823 5305
rect 31849 5279 31906 5305
rect 31822 5278 31906 5279
rect 31822 5273 31850 5278
rect 30982 4887 30983 4913
rect 31009 4887 31010 4913
rect 30478 4521 30506 4527
rect 30478 4495 30479 4521
rect 30505 4495 30506 4521
rect 30310 4074 30338 4079
rect 30310 4027 30338 4046
rect 30478 3737 30506 4495
rect 30982 4242 31010 4887
rect 31878 4913 31906 5278
rect 32718 5306 32746 5670
rect 33334 5697 33362 6062
rect 33390 6057 33418 6062
rect 33334 5671 33335 5697
rect 33361 5671 33362 5697
rect 33334 5641 33362 5671
rect 33334 5615 33335 5641
rect 33361 5615 33362 5641
rect 32073 5110 32535 5115
rect 32073 5109 32082 5110
rect 32073 5083 32074 5109
rect 32073 5082 32082 5083
rect 32110 5082 32134 5110
rect 32162 5082 32186 5110
rect 32214 5109 32238 5110
rect 32266 5109 32290 5110
rect 32224 5083 32238 5109
rect 32286 5083 32290 5109
rect 32214 5082 32238 5083
rect 32266 5082 32290 5083
rect 32318 5109 32342 5110
rect 32370 5109 32394 5110
rect 32318 5083 32322 5109
rect 32370 5083 32384 5109
rect 32318 5082 32342 5083
rect 32370 5082 32394 5083
rect 32422 5082 32446 5110
rect 32474 5082 32498 5110
rect 32526 5109 32535 5110
rect 32534 5083 32535 5109
rect 32526 5082 32535 5083
rect 32073 5077 32535 5082
rect 32158 4914 32186 4919
rect 31878 4887 31879 4913
rect 31905 4887 31906 4913
rect 31878 4857 31906 4887
rect 31990 4913 32186 4914
rect 31990 4887 32159 4913
rect 32185 4887 32186 4913
rect 31990 4886 32186 4887
rect 31878 4831 31879 4857
rect 31905 4831 31906 4857
rect 30982 4129 31010 4214
rect 30982 4103 30983 4129
rect 31009 4103 31010 4129
rect 30478 3711 30479 3737
rect 30505 3711 30506 3737
rect 30478 3402 30506 3711
rect 30478 3369 30506 3374
rect 30814 3850 30842 3855
rect 30702 3346 30730 3351
rect 30310 3289 30338 3295
rect 30310 3263 30311 3289
rect 30337 3263 30338 3289
rect 30310 3010 30338 3263
rect 30310 2618 30338 2982
rect 30310 2561 30338 2590
rect 30310 2535 30311 2561
rect 30337 2535 30338 2561
rect 30310 2529 30338 2535
rect 30366 2953 30394 2959
rect 30366 2927 30367 2953
rect 30393 2927 30394 2953
rect 30310 2170 30338 2175
rect 30366 2170 30394 2927
rect 30702 2562 30730 3318
rect 30702 2529 30730 2534
rect 30814 2561 30842 3822
rect 30982 3402 31010 4103
rect 31374 4577 31402 4583
rect 31374 4551 31375 4577
rect 31401 4551 31402 4577
rect 31374 4521 31402 4551
rect 31374 4495 31375 4521
rect 31401 4495 31402 4521
rect 31374 3793 31402 4495
rect 31374 3767 31375 3793
rect 31401 3767 31402 3793
rect 31374 3738 31402 3767
rect 31878 4129 31906 4831
rect 31878 4103 31879 4129
rect 31905 4103 31906 4129
rect 31878 4073 31906 4103
rect 31878 4047 31879 4073
rect 31905 4047 31906 4073
rect 31878 3738 31906 4047
rect 31374 3737 31906 3738
rect 31374 3711 31375 3737
rect 31401 3711 31906 3737
rect 31374 3710 31906 3711
rect 31934 4858 31962 4863
rect 31934 4522 31962 4830
rect 31934 3738 31962 4494
rect 31990 4242 32018 4886
rect 32158 4881 32186 4886
rect 32046 4522 32074 4527
rect 32046 4475 32074 4494
rect 32158 4521 32186 4527
rect 32158 4495 32159 4521
rect 32185 4495 32186 4521
rect 32158 4466 32186 4495
rect 32158 4433 32186 4438
rect 32326 4521 32354 4527
rect 32326 4495 32327 4521
rect 32353 4495 32354 4521
rect 32326 4466 32354 4495
rect 32326 4433 32354 4438
rect 32718 4521 32746 5278
rect 33278 5306 33306 5311
rect 33334 5306 33362 5615
rect 33390 5306 33418 5311
rect 33278 5305 33418 5306
rect 33278 5279 33279 5305
rect 33305 5279 33391 5305
rect 33417 5279 33418 5305
rect 33278 5278 33418 5279
rect 33278 5273 33306 5278
rect 33390 5250 33418 5278
rect 33334 4914 33362 4919
rect 33390 4914 33418 5222
rect 33614 5082 33642 7183
rect 33782 7210 33810 7239
rect 33894 7210 33922 7215
rect 33782 7209 33922 7210
rect 33782 7183 33895 7209
rect 33921 7183 33922 7209
rect 33782 7182 33922 7183
rect 33670 6481 33698 6487
rect 33670 6455 33671 6481
rect 33697 6455 33698 6481
rect 33670 5922 33698 6455
rect 33670 5697 33698 5894
rect 33670 5671 33671 5697
rect 33697 5671 33698 5697
rect 33670 5665 33698 5671
rect 33726 6482 33754 6487
rect 33726 5641 33754 6454
rect 33726 5615 33727 5641
rect 33753 5615 33754 5641
rect 33670 5082 33698 5087
rect 33614 5054 33670 5082
rect 33334 4913 33418 4914
rect 33334 4887 33335 4913
rect 33361 4887 33418 4913
rect 33334 4886 33418 4887
rect 33670 4913 33698 5054
rect 33670 4887 33671 4913
rect 33697 4887 33698 4913
rect 33334 4857 33362 4886
rect 33334 4831 33335 4857
rect 33361 4831 33362 4857
rect 32718 4495 32719 4521
rect 32745 4495 32746 4521
rect 32073 4326 32535 4331
rect 32073 4325 32082 4326
rect 32073 4299 32074 4325
rect 32073 4298 32082 4299
rect 32110 4298 32134 4326
rect 32162 4298 32186 4326
rect 32214 4325 32238 4326
rect 32266 4325 32290 4326
rect 32224 4299 32238 4325
rect 32286 4299 32290 4325
rect 32214 4298 32238 4299
rect 32266 4298 32290 4299
rect 32318 4325 32342 4326
rect 32370 4325 32394 4326
rect 32318 4299 32322 4325
rect 32370 4299 32384 4325
rect 32318 4298 32342 4299
rect 32370 4298 32394 4299
rect 32422 4298 32446 4326
rect 32474 4298 32498 4326
rect 32526 4325 32535 4326
rect 32534 4299 32535 4325
rect 32526 4298 32535 4299
rect 32073 4293 32535 4298
rect 31990 4209 32018 4214
rect 32158 4242 32186 4247
rect 32158 4129 32186 4214
rect 32718 4242 32746 4495
rect 33278 4522 33306 4527
rect 33334 4522 33362 4831
rect 33390 4522 33418 4527
rect 33278 4521 33418 4522
rect 33278 4495 33279 4521
rect 33305 4495 33391 4521
rect 33417 4495 33418 4521
rect 33278 4494 33418 4495
rect 33278 4489 33306 4494
rect 32718 4209 32746 4214
rect 32158 4103 32159 4129
rect 32185 4103 32186 4129
rect 32158 4097 32186 4103
rect 33334 4129 33362 4494
rect 33390 4489 33418 4494
rect 33334 4103 33335 4129
rect 33361 4103 33362 4129
rect 33334 4073 33362 4103
rect 33334 4047 33335 4073
rect 33361 4047 33362 4073
rect 32046 3738 32074 3743
rect 31934 3737 32074 3738
rect 31934 3711 32047 3737
rect 32073 3711 32074 3737
rect 31934 3710 32074 3711
rect 31374 3705 31402 3710
rect 30982 3369 31010 3374
rect 31598 3346 31626 3351
rect 30814 2535 30815 2561
rect 30841 2535 30842 2561
rect 30814 2529 30842 2535
rect 31262 3009 31290 3015
rect 31262 2983 31263 3009
rect 31289 2983 31290 3009
rect 31262 2953 31290 2983
rect 31262 2927 31263 2953
rect 31289 2927 31290 2953
rect 30310 2169 30394 2170
rect 30310 2143 30311 2169
rect 30337 2143 30394 2169
rect 30310 2142 30394 2143
rect 31262 2170 31290 2927
rect 31318 2954 31346 2959
rect 31318 2226 31346 2926
rect 31374 2226 31402 2231
rect 31318 2225 31402 2226
rect 31318 2199 31375 2225
rect 31401 2199 31402 2225
rect 31318 2198 31402 2199
rect 30310 1778 30338 2142
rect 31262 2137 31290 2142
rect 31374 2169 31402 2198
rect 31374 2143 31375 2169
rect 31401 2143 31402 2169
rect 31374 2137 31402 2143
rect 31486 2170 31514 2175
rect 30310 1712 30338 1750
rect 31486 1777 31514 2142
rect 31486 1751 31487 1777
rect 31513 1751 31514 1777
rect 31486 1722 31514 1751
rect 31486 1689 31514 1694
rect 31598 1694 31626 3318
rect 31878 3345 31906 3710
rect 31878 3319 31879 3345
rect 31905 3319 31906 3345
rect 31878 3289 31906 3319
rect 31878 3263 31879 3289
rect 31905 3263 31906 3289
rect 31878 2561 31906 3263
rect 31878 2535 31879 2561
rect 31905 2535 31906 2561
rect 31878 2505 31906 2535
rect 31878 2479 31879 2505
rect 31905 2479 31906 2505
rect 31878 1778 31906 2479
rect 31990 2954 32018 3710
rect 32046 3705 32074 3710
rect 32158 3738 32186 3743
rect 32158 3691 32186 3710
rect 32326 3738 32354 3743
rect 32326 3691 32354 3710
rect 32886 3737 32914 3743
rect 32886 3711 32887 3737
rect 32913 3711 32914 3737
rect 32073 3542 32535 3547
rect 32073 3541 32082 3542
rect 32073 3515 32074 3541
rect 32073 3514 32082 3515
rect 32110 3514 32134 3542
rect 32162 3514 32186 3542
rect 32214 3541 32238 3542
rect 32266 3541 32290 3542
rect 32224 3515 32238 3541
rect 32286 3515 32290 3541
rect 32214 3514 32238 3515
rect 32266 3514 32290 3515
rect 32318 3541 32342 3542
rect 32370 3541 32394 3542
rect 32318 3515 32322 3541
rect 32370 3515 32384 3541
rect 32318 3514 32342 3515
rect 32370 3514 32394 3515
rect 32422 3514 32446 3542
rect 32474 3514 32498 3542
rect 32526 3541 32535 3542
rect 32534 3515 32535 3541
rect 32526 3514 32535 3515
rect 32073 3509 32535 3514
rect 32438 3345 32466 3351
rect 32438 3319 32439 3345
rect 32465 3319 32466 3345
rect 32158 3010 32186 3015
rect 32158 2963 32186 2982
rect 32326 3010 32354 3015
rect 32326 2963 32354 2982
rect 32046 2954 32074 2959
rect 31990 2953 32074 2954
rect 31990 2927 32047 2953
rect 32073 2927 32074 2953
rect 31990 2926 32074 2927
rect 31990 2170 32018 2926
rect 32046 2921 32074 2926
rect 32438 2898 32466 3319
rect 32718 3346 32746 3351
rect 32830 3346 32858 3351
rect 32718 3345 32858 3346
rect 32718 3319 32719 3345
rect 32745 3319 32831 3345
rect 32857 3319 32858 3345
rect 32718 3318 32858 3319
rect 32718 3313 32746 3318
rect 32830 2954 32858 3318
rect 32830 2921 32858 2926
rect 32886 3010 32914 3711
rect 32438 2865 32466 2870
rect 32073 2758 32535 2763
rect 32073 2757 32082 2758
rect 32073 2731 32074 2757
rect 32073 2730 32082 2731
rect 32110 2730 32134 2758
rect 32162 2730 32186 2758
rect 32214 2757 32238 2758
rect 32266 2757 32290 2758
rect 32224 2731 32238 2757
rect 32286 2731 32290 2757
rect 32214 2730 32238 2731
rect 32266 2730 32290 2731
rect 32318 2757 32342 2758
rect 32370 2757 32394 2758
rect 32318 2731 32322 2757
rect 32370 2731 32384 2757
rect 32318 2730 32342 2731
rect 32370 2730 32394 2731
rect 32422 2730 32446 2758
rect 32474 2730 32498 2758
rect 32526 2757 32535 2758
rect 32534 2731 32535 2757
rect 32526 2730 32535 2731
rect 32073 2725 32535 2730
rect 32158 2562 32186 2567
rect 32158 2515 32186 2534
rect 32606 2562 32634 2567
rect 32158 2226 32186 2231
rect 32158 2179 32186 2198
rect 32326 2226 32354 2231
rect 32326 2179 32354 2198
rect 32102 2170 32130 2175
rect 31990 2142 32102 2170
rect 32102 2123 32130 2142
rect 32606 2170 32634 2534
rect 32718 2170 32746 2175
rect 32606 2169 32746 2170
rect 32606 2143 32719 2169
rect 32745 2143 32746 2169
rect 32606 2142 32746 2143
rect 32073 1974 32535 1979
rect 32073 1973 32082 1974
rect 32073 1947 32074 1973
rect 32073 1946 32082 1947
rect 32110 1946 32134 1974
rect 32162 1946 32186 1974
rect 32214 1973 32238 1974
rect 32266 1973 32290 1974
rect 32224 1947 32238 1973
rect 32286 1947 32290 1973
rect 32214 1946 32238 1947
rect 32266 1946 32290 1947
rect 32318 1973 32342 1974
rect 32370 1973 32394 1974
rect 32318 1947 32322 1973
rect 32370 1947 32384 1973
rect 32318 1946 32342 1947
rect 32370 1946 32394 1947
rect 32422 1946 32446 1974
rect 32474 1946 32498 1974
rect 32526 1973 32535 1974
rect 32534 1947 32535 1973
rect 32526 1946 32535 1947
rect 32073 1941 32535 1946
rect 31878 1745 31906 1750
rect 32550 1778 32578 1783
rect 32606 1778 32634 2142
rect 32718 2137 32746 2142
rect 32550 1777 32634 1778
rect 32550 1751 32551 1777
rect 32577 1751 32634 1777
rect 32550 1750 32634 1751
rect 32550 1745 32578 1750
rect 31598 1666 31682 1694
rect 30254 854 30450 882
rect 29022 462 29218 490
rect 29022 378 29050 462
rect 29190 400 29218 462
rect 30422 400 30450 854
rect 31654 400 31682 1666
rect 32886 400 32914 2982
rect 32998 2953 33026 2959
rect 32998 2927 32999 2953
rect 33025 2927 33026 2953
rect 32998 2898 33026 2927
rect 33166 2954 33194 2959
rect 33166 2907 33194 2926
rect 32998 2865 33026 2870
rect 33334 2561 33362 4047
rect 33670 4129 33698 4887
rect 33670 4103 33671 4129
rect 33697 4103 33698 4129
rect 33670 3345 33698 4103
rect 33670 3319 33671 3345
rect 33697 3319 33698 3345
rect 33390 2954 33418 2959
rect 33390 2907 33418 2926
rect 33334 2535 33335 2561
rect 33361 2535 33362 2561
rect 33334 2506 33362 2535
rect 33334 2459 33362 2478
rect 33670 2561 33698 3319
rect 33670 2535 33671 2561
rect 33697 2535 33698 2561
rect 33670 2170 33698 2535
rect 33726 4858 33754 5615
rect 33782 5026 33810 7182
rect 33894 7177 33922 7182
rect 33894 6929 33922 6935
rect 33894 6903 33895 6929
rect 33921 6903 33922 6929
rect 33894 6873 33922 6903
rect 33894 6847 33895 6873
rect 33921 6847 33922 6873
rect 33894 6762 33922 6847
rect 33894 6729 33922 6734
rect 33894 6482 33922 6487
rect 33894 5697 33922 6454
rect 33894 5671 33895 5697
rect 33921 5671 33922 5697
rect 33894 5665 33922 5671
rect 33782 4993 33810 4998
rect 33894 4858 33922 4863
rect 33726 4857 33922 4858
rect 33726 4831 33727 4857
rect 33753 4831 33895 4857
rect 33921 4831 33922 4857
rect 33726 4830 33922 4831
rect 33726 4074 33754 4830
rect 33894 4825 33922 4830
rect 33894 4074 33922 4079
rect 33726 4073 33922 4074
rect 33726 4047 33727 4073
rect 33753 4047 33895 4073
rect 33921 4047 33922 4073
rect 33726 4046 33922 4047
rect 33726 3346 33754 4046
rect 33894 4041 33922 4046
rect 33894 3793 33922 3799
rect 33894 3767 33895 3793
rect 33921 3767 33922 3793
rect 33894 3738 33922 3767
rect 33894 3691 33922 3710
rect 33894 3346 33922 3351
rect 33726 3345 33922 3346
rect 33726 3319 33895 3345
rect 33921 3319 33922 3345
rect 33726 3318 33922 3319
rect 33726 3289 33754 3318
rect 33894 3313 33922 3318
rect 33726 3263 33727 3289
rect 33753 3263 33754 3289
rect 33726 2618 33754 3263
rect 33726 2590 33922 2618
rect 33726 2505 33754 2590
rect 33894 2561 33922 2590
rect 33894 2535 33895 2561
rect 33921 2535 33922 2561
rect 33894 2529 33922 2535
rect 33726 2479 33727 2505
rect 33753 2479 33754 2505
rect 33726 2226 33754 2479
rect 33726 2193 33754 2198
rect 33838 2506 33866 2511
rect 33838 2225 33866 2478
rect 33950 2450 33978 7966
rect 34398 7657 34426 8414
rect 34510 8050 34538 8806
rect 34678 8801 34706 8806
rect 35238 9281 35266 9287
rect 35238 9255 35239 9281
rect 35265 9255 35266 9281
rect 35238 9225 35266 9255
rect 35238 9199 35239 9225
rect 35265 9199 35266 9225
rect 34573 8638 35035 8643
rect 34573 8637 34582 8638
rect 34573 8611 34574 8637
rect 34573 8610 34582 8611
rect 34610 8610 34634 8638
rect 34662 8610 34686 8638
rect 34714 8637 34738 8638
rect 34766 8637 34790 8638
rect 34724 8611 34738 8637
rect 34786 8611 34790 8637
rect 34714 8610 34738 8611
rect 34766 8610 34790 8611
rect 34818 8637 34842 8638
rect 34870 8637 34894 8638
rect 34818 8611 34822 8637
rect 34870 8611 34884 8637
rect 34818 8610 34842 8611
rect 34870 8610 34894 8611
rect 34922 8610 34946 8638
rect 34974 8610 34998 8638
rect 35026 8637 35035 8638
rect 35034 8611 35035 8637
rect 35026 8610 35035 8611
rect 34573 8605 35035 8610
rect 34678 8050 34706 8055
rect 34510 8022 34678 8050
rect 34678 7984 34706 8022
rect 34573 7854 35035 7859
rect 34573 7853 34582 7854
rect 34573 7827 34574 7853
rect 34573 7826 34582 7827
rect 34610 7826 34634 7854
rect 34662 7826 34686 7854
rect 34714 7853 34738 7854
rect 34766 7853 34790 7854
rect 34724 7827 34738 7853
rect 34786 7827 34790 7853
rect 34714 7826 34738 7827
rect 34766 7826 34790 7827
rect 34818 7853 34842 7854
rect 34870 7853 34894 7854
rect 34818 7827 34822 7853
rect 34870 7827 34884 7853
rect 34818 7826 34842 7827
rect 34870 7826 34894 7827
rect 34922 7826 34946 7854
rect 34974 7826 34998 7854
rect 35026 7853 35035 7854
rect 35034 7827 35035 7853
rect 35026 7826 35035 7827
rect 34573 7821 35035 7826
rect 34398 7631 34399 7657
rect 34425 7631 34426 7657
rect 34398 7266 34426 7631
rect 35238 7713 35266 9199
rect 36190 9170 36218 9175
rect 35854 8833 35882 8839
rect 35854 8807 35855 8833
rect 35881 8807 35882 8833
rect 35854 8778 35882 8807
rect 35798 8750 35854 8778
rect 35238 7687 35239 7713
rect 35265 7687 35266 7713
rect 35238 7658 35266 7687
rect 35238 7574 35266 7630
rect 35182 7546 35266 7574
rect 35350 8497 35378 8503
rect 35350 8471 35351 8497
rect 35377 8471 35378 8497
rect 35350 8441 35378 8471
rect 35350 8415 35351 8441
rect 35377 8415 35378 8441
rect 35350 7546 35378 8415
rect 35798 7658 35826 8750
rect 35854 8731 35882 8750
rect 34398 7233 34426 7238
rect 34958 7266 34986 7271
rect 34958 7219 34986 7238
rect 34573 7070 35035 7075
rect 34573 7069 34582 7070
rect 34573 7043 34574 7069
rect 34573 7042 34582 7043
rect 34610 7042 34634 7070
rect 34662 7042 34686 7070
rect 34714 7069 34738 7070
rect 34766 7069 34790 7070
rect 34724 7043 34738 7069
rect 34786 7043 34790 7069
rect 34714 7042 34738 7043
rect 34766 7042 34790 7043
rect 34818 7069 34842 7070
rect 34870 7069 34894 7070
rect 34818 7043 34822 7069
rect 34870 7043 34884 7069
rect 34818 7042 34842 7043
rect 34870 7042 34894 7043
rect 34922 7042 34946 7070
rect 34974 7042 34998 7070
rect 35026 7069 35035 7070
rect 35034 7043 35035 7069
rect 35026 7042 35035 7043
rect 34573 7037 35035 7042
rect 35182 6930 35210 7546
rect 35350 7513 35378 7518
rect 35518 7546 35546 7551
rect 35182 6897 35210 6902
rect 35294 6929 35322 6935
rect 35294 6903 35295 6929
rect 35321 6903 35322 6929
rect 34398 6873 34426 6879
rect 34398 6847 34399 6873
rect 34425 6847 34426 6873
rect 34398 6706 34426 6847
rect 35294 6874 35322 6903
rect 35294 6827 35322 6846
rect 34398 6482 34426 6678
rect 35350 6762 35378 6767
rect 35518 6762 35546 7518
rect 35798 7265 35826 7630
rect 35798 7239 35799 7265
rect 35825 7239 35826 7265
rect 35798 7209 35826 7239
rect 35798 7183 35799 7209
rect 35825 7183 35826 7209
rect 35798 7177 35826 7183
rect 35854 8049 35882 8055
rect 35854 8023 35855 8049
rect 35881 8023 35882 8049
rect 35854 7993 35882 8023
rect 35854 7967 35855 7993
rect 35881 7967 35882 7993
rect 35854 7546 35882 7967
rect 35854 7210 35882 7518
rect 36134 8050 36162 8055
rect 36134 7658 36162 8022
rect 36134 7265 36162 7630
rect 36190 7574 36218 9142
rect 36414 8834 36442 9478
rect 36694 9225 36722 9590
rect 36694 9199 36695 9225
rect 36721 9199 36722 9225
rect 36694 9193 36722 9199
rect 36414 8833 36722 8834
rect 36414 8807 36415 8833
rect 36441 8807 36722 8833
rect 36414 8806 36722 8807
rect 36414 8801 36442 8806
rect 36694 8441 36722 8806
rect 36694 8415 36695 8441
rect 36721 8415 36722 8441
rect 36694 8409 36722 8415
rect 36974 8778 37002 19614
rect 37254 19530 37282 19614
rect 37408 19600 37464 20000
rect 37422 19530 37450 19600
rect 37254 19502 37450 19530
rect 37073 18438 37535 18443
rect 37073 18437 37082 18438
rect 37073 18411 37074 18437
rect 37073 18410 37082 18411
rect 37110 18410 37134 18438
rect 37162 18410 37186 18438
rect 37214 18437 37238 18438
rect 37266 18437 37290 18438
rect 37224 18411 37238 18437
rect 37286 18411 37290 18437
rect 37214 18410 37238 18411
rect 37266 18410 37290 18411
rect 37318 18437 37342 18438
rect 37370 18437 37394 18438
rect 37318 18411 37322 18437
rect 37370 18411 37384 18437
rect 37318 18410 37342 18411
rect 37370 18410 37394 18411
rect 37422 18410 37446 18438
rect 37474 18410 37498 18438
rect 37526 18437 37535 18438
rect 37534 18411 37535 18437
rect 37526 18410 37535 18411
rect 37073 18405 37535 18410
rect 37073 17654 37535 17659
rect 37073 17653 37082 17654
rect 37073 17627 37074 17653
rect 37073 17626 37082 17627
rect 37110 17626 37134 17654
rect 37162 17626 37186 17654
rect 37214 17653 37238 17654
rect 37266 17653 37290 17654
rect 37224 17627 37238 17653
rect 37286 17627 37290 17653
rect 37214 17626 37238 17627
rect 37266 17626 37290 17627
rect 37318 17653 37342 17654
rect 37370 17653 37394 17654
rect 37318 17627 37322 17653
rect 37370 17627 37384 17653
rect 37318 17626 37342 17627
rect 37370 17626 37394 17627
rect 37422 17626 37446 17654
rect 37474 17626 37498 17654
rect 37526 17653 37535 17654
rect 37534 17627 37535 17653
rect 37526 17626 37535 17627
rect 37073 17621 37535 17626
rect 37073 16870 37535 16875
rect 37073 16869 37082 16870
rect 37073 16843 37074 16869
rect 37073 16842 37082 16843
rect 37110 16842 37134 16870
rect 37162 16842 37186 16870
rect 37214 16869 37238 16870
rect 37266 16869 37290 16870
rect 37224 16843 37238 16869
rect 37286 16843 37290 16869
rect 37214 16842 37238 16843
rect 37266 16842 37290 16843
rect 37318 16869 37342 16870
rect 37370 16869 37394 16870
rect 37318 16843 37322 16869
rect 37370 16843 37384 16869
rect 37318 16842 37342 16843
rect 37370 16842 37394 16843
rect 37422 16842 37446 16870
rect 37474 16842 37498 16870
rect 37526 16869 37535 16870
rect 37534 16843 37535 16869
rect 37526 16842 37535 16843
rect 37073 16837 37535 16842
rect 37073 16086 37535 16091
rect 37073 16085 37082 16086
rect 37073 16059 37074 16085
rect 37073 16058 37082 16059
rect 37110 16058 37134 16086
rect 37162 16058 37186 16086
rect 37214 16085 37238 16086
rect 37266 16085 37290 16086
rect 37224 16059 37238 16085
rect 37286 16059 37290 16085
rect 37214 16058 37238 16059
rect 37266 16058 37290 16059
rect 37318 16085 37342 16086
rect 37370 16085 37394 16086
rect 37318 16059 37322 16085
rect 37370 16059 37384 16085
rect 37318 16058 37342 16059
rect 37370 16058 37394 16059
rect 37422 16058 37446 16086
rect 37474 16058 37498 16086
rect 37526 16085 37535 16086
rect 37534 16059 37535 16085
rect 37526 16058 37535 16059
rect 37073 16053 37535 16058
rect 37073 15302 37535 15307
rect 37073 15301 37082 15302
rect 37073 15275 37074 15301
rect 37073 15274 37082 15275
rect 37110 15274 37134 15302
rect 37162 15274 37186 15302
rect 37214 15301 37238 15302
rect 37266 15301 37290 15302
rect 37224 15275 37238 15301
rect 37286 15275 37290 15301
rect 37214 15274 37238 15275
rect 37266 15274 37290 15275
rect 37318 15301 37342 15302
rect 37370 15301 37394 15302
rect 37318 15275 37322 15301
rect 37370 15275 37384 15301
rect 37318 15274 37342 15275
rect 37370 15274 37394 15275
rect 37422 15274 37446 15302
rect 37474 15274 37498 15302
rect 37526 15301 37535 15302
rect 37534 15275 37535 15301
rect 37526 15274 37535 15275
rect 37073 15269 37535 15274
rect 37073 14518 37535 14523
rect 37073 14517 37082 14518
rect 37073 14491 37074 14517
rect 37073 14490 37082 14491
rect 37110 14490 37134 14518
rect 37162 14490 37186 14518
rect 37214 14517 37238 14518
rect 37266 14517 37290 14518
rect 37224 14491 37238 14517
rect 37286 14491 37290 14517
rect 37214 14490 37238 14491
rect 37266 14490 37290 14491
rect 37318 14517 37342 14518
rect 37370 14517 37394 14518
rect 37318 14491 37322 14517
rect 37370 14491 37384 14517
rect 37318 14490 37342 14491
rect 37370 14490 37394 14491
rect 37422 14490 37446 14518
rect 37474 14490 37498 14518
rect 37526 14517 37535 14518
rect 37534 14491 37535 14517
rect 37526 14490 37535 14491
rect 37073 14485 37535 14490
rect 37073 13734 37535 13739
rect 37073 13733 37082 13734
rect 37073 13707 37074 13733
rect 37073 13706 37082 13707
rect 37110 13706 37134 13734
rect 37162 13706 37186 13734
rect 37214 13733 37238 13734
rect 37266 13733 37290 13734
rect 37224 13707 37238 13733
rect 37286 13707 37290 13733
rect 37214 13706 37238 13707
rect 37266 13706 37290 13707
rect 37318 13733 37342 13734
rect 37370 13733 37394 13734
rect 37318 13707 37322 13733
rect 37370 13707 37384 13733
rect 37318 13706 37342 13707
rect 37370 13706 37394 13707
rect 37422 13706 37446 13734
rect 37474 13706 37498 13734
rect 37526 13733 37535 13734
rect 37534 13707 37535 13733
rect 37526 13706 37535 13707
rect 37073 13701 37535 13706
rect 37073 12950 37535 12955
rect 37073 12949 37082 12950
rect 37073 12923 37074 12949
rect 37073 12922 37082 12923
rect 37110 12922 37134 12950
rect 37162 12922 37186 12950
rect 37214 12949 37238 12950
rect 37266 12949 37290 12950
rect 37224 12923 37238 12949
rect 37286 12923 37290 12949
rect 37214 12922 37238 12923
rect 37266 12922 37290 12923
rect 37318 12949 37342 12950
rect 37370 12949 37394 12950
rect 37318 12923 37322 12949
rect 37370 12923 37384 12949
rect 37318 12922 37342 12923
rect 37370 12922 37394 12923
rect 37422 12922 37446 12950
rect 37474 12922 37498 12950
rect 37526 12949 37535 12950
rect 37534 12923 37535 12949
rect 37526 12922 37535 12923
rect 37073 12917 37535 12922
rect 37073 12166 37535 12171
rect 37073 12165 37082 12166
rect 37073 12139 37074 12165
rect 37073 12138 37082 12139
rect 37110 12138 37134 12166
rect 37162 12138 37186 12166
rect 37214 12165 37238 12166
rect 37266 12165 37290 12166
rect 37224 12139 37238 12165
rect 37286 12139 37290 12165
rect 37214 12138 37238 12139
rect 37266 12138 37290 12139
rect 37318 12165 37342 12166
rect 37370 12165 37394 12166
rect 37318 12139 37322 12165
rect 37370 12139 37384 12165
rect 37318 12138 37342 12139
rect 37370 12138 37394 12139
rect 37422 12138 37446 12166
rect 37474 12138 37498 12166
rect 37526 12165 37535 12166
rect 37534 12139 37535 12165
rect 37526 12138 37535 12139
rect 37073 12133 37535 12138
rect 37073 11382 37535 11387
rect 37073 11381 37082 11382
rect 37073 11355 37074 11381
rect 37073 11354 37082 11355
rect 37110 11354 37134 11382
rect 37162 11354 37186 11382
rect 37214 11381 37238 11382
rect 37266 11381 37290 11382
rect 37224 11355 37238 11381
rect 37286 11355 37290 11381
rect 37214 11354 37238 11355
rect 37266 11354 37290 11355
rect 37318 11381 37342 11382
rect 37370 11381 37394 11382
rect 37318 11355 37322 11381
rect 37370 11355 37384 11381
rect 37318 11354 37342 11355
rect 37370 11354 37394 11355
rect 37422 11354 37446 11382
rect 37474 11354 37498 11382
rect 37526 11381 37535 11382
rect 37534 11355 37535 11381
rect 37526 11354 37535 11355
rect 37073 11349 37535 11354
rect 37310 11185 37338 11191
rect 37310 11159 37311 11185
rect 37337 11159 37338 11185
rect 37310 11130 37338 11159
rect 37310 11129 37674 11130
rect 37310 11103 37311 11129
rect 37337 11103 37674 11129
rect 37310 11102 37674 11103
rect 37310 11097 37338 11102
rect 37646 10849 37674 11102
rect 37646 10823 37647 10849
rect 37673 10823 37674 10849
rect 37646 10793 37674 10823
rect 37646 10767 37647 10793
rect 37673 10767 37674 10793
rect 37073 10598 37535 10603
rect 37073 10597 37082 10598
rect 37073 10571 37074 10597
rect 37073 10570 37082 10571
rect 37110 10570 37134 10598
rect 37162 10570 37186 10598
rect 37214 10597 37238 10598
rect 37266 10597 37290 10598
rect 37224 10571 37238 10597
rect 37286 10571 37290 10597
rect 37214 10570 37238 10571
rect 37266 10570 37290 10571
rect 37318 10597 37342 10598
rect 37370 10597 37394 10598
rect 37318 10571 37322 10597
rect 37370 10571 37384 10597
rect 37318 10570 37342 10571
rect 37370 10570 37394 10571
rect 37422 10570 37446 10598
rect 37474 10570 37498 10598
rect 37526 10597 37535 10598
rect 37534 10571 37535 10597
rect 37526 10570 37535 10571
rect 37073 10565 37535 10570
rect 37310 10401 37338 10407
rect 37310 10375 37311 10401
rect 37337 10375 37338 10401
rect 37310 10346 37338 10375
rect 37310 10299 37338 10318
rect 37590 10346 37618 10351
rect 37073 9814 37535 9819
rect 37073 9813 37082 9814
rect 37073 9787 37074 9813
rect 37073 9786 37082 9787
rect 37110 9786 37134 9814
rect 37162 9786 37186 9814
rect 37214 9813 37238 9814
rect 37266 9813 37290 9814
rect 37224 9787 37238 9813
rect 37286 9787 37290 9813
rect 37214 9786 37238 9787
rect 37266 9786 37290 9787
rect 37318 9813 37342 9814
rect 37370 9813 37394 9814
rect 37318 9787 37322 9813
rect 37370 9787 37384 9813
rect 37318 9786 37342 9787
rect 37370 9786 37394 9787
rect 37422 9786 37446 9814
rect 37474 9786 37498 9814
rect 37526 9813 37535 9814
rect 37534 9787 37535 9813
rect 37526 9786 37535 9787
rect 37073 9781 37535 9786
rect 37310 9617 37338 9623
rect 37310 9591 37311 9617
rect 37337 9591 37338 9617
rect 37310 9562 37338 9591
rect 37310 9515 37338 9534
rect 37073 9030 37535 9035
rect 37073 9029 37082 9030
rect 37073 9003 37074 9029
rect 37073 9002 37082 9003
rect 37110 9002 37134 9030
rect 37162 9002 37186 9030
rect 37214 9029 37238 9030
rect 37266 9029 37290 9030
rect 37224 9003 37238 9029
rect 37286 9003 37290 9029
rect 37214 9002 37238 9003
rect 37266 9002 37290 9003
rect 37318 9029 37342 9030
rect 37370 9029 37394 9030
rect 37318 9003 37322 9029
rect 37370 9003 37384 9029
rect 37318 9002 37342 9003
rect 37370 9002 37394 9003
rect 37422 9002 37446 9030
rect 37474 9002 37498 9030
rect 37526 9029 37535 9030
rect 37534 9003 37535 9029
rect 37526 9002 37535 9003
rect 37073 8997 37535 9002
rect 36974 8050 37002 8750
rect 37310 8833 37338 8839
rect 37310 8807 37311 8833
rect 37337 8807 37338 8833
rect 37310 8778 37338 8807
rect 37590 8778 37618 10318
rect 37646 10065 37674 10767
rect 37646 10039 37647 10065
rect 37673 10039 37674 10065
rect 37646 10009 37674 10039
rect 37646 9983 37647 10009
rect 37673 9983 37674 10009
rect 37646 9562 37674 9983
rect 37646 9281 37674 9534
rect 37646 9255 37647 9281
rect 37673 9255 37674 9281
rect 37646 9225 37674 9255
rect 37646 9199 37647 9225
rect 37673 9199 37674 9225
rect 37646 9193 37674 9199
rect 37310 8777 37674 8778
rect 37310 8751 37311 8777
rect 37337 8751 37674 8777
rect 37310 8750 37674 8751
rect 37310 8745 37338 8750
rect 37646 8497 37674 8750
rect 37646 8471 37647 8497
rect 37673 8471 37674 8497
rect 37646 8441 37674 8471
rect 37646 8415 37647 8441
rect 37673 8415 37674 8441
rect 37646 8409 37674 8415
rect 37073 8246 37535 8251
rect 37073 8245 37082 8246
rect 37073 8219 37074 8245
rect 37073 8218 37082 8219
rect 37110 8218 37134 8246
rect 37162 8218 37186 8246
rect 37214 8245 37238 8246
rect 37266 8245 37290 8246
rect 37224 8219 37238 8245
rect 37286 8219 37290 8245
rect 37214 8218 37238 8219
rect 37266 8218 37290 8219
rect 37318 8245 37342 8246
rect 37370 8245 37394 8246
rect 37318 8219 37322 8245
rect 37370 8219 37384 8245
rect 37318 8218 37342 8219
rect 37370 8218 37394 8219
rect 37422 8218 37446 8246
rect 37474 8218 37498 8246
rect 37526 8245 37535 8246
rect 37534 8219 37535 8245
rect 37526 8218 37535 8219
rect 37073 8213 37535 8218
rect 36974 8049 37114 8050
rect 36974 8023 36975 8049
rect 37001 8023 37114 8049
rect 36974 8022 37114 8023
rect 36974 8017 37002 8022
rect 37086 7994 37114 8022
rect 37086 7993 37170 7994
rect 37086 7967 37087 7993
rect 37113 7967 37170 7993
rect 37086 7966 37170 7967
rect 37086 7961 37114 7966
rect 36694 7658 36722 7663
rect 36190 7546 36442 7574
rect 36134 7239 36135 7265
rect 36161 7239 36162 7265
rect 36134 7233 36162 7239
rect 35854 7177 35882 7182
rect 35378 6734 35546 6762
rect 35630 6874 35658 6879
rect 34678 6482 34706 6487
rect 34398 6481 34706 6482
rect 34398 6455 34679 6481
rect 34705 6455 34706 6481
rect 34398 6454 34706 6455
rect 34454 6090 34482 6095
rect 34510 6090 34538 6454
rect 34678 6449 34706 6454
rect 34573 6286 35035 6291
rect 34573 6285 34582 6286
rect 34573 6259 34574 6285
rect 34573 6258 34582 6259
rect 34610 6258 34634 6286
rect 34662 6258 34686 6286
rect 34714 6285 34738 6286
rect 34766 6285 34790 6286
rect 34724 6259 34738 6285
rect 34786 6259 34790 6285
rect 34714 6258 34738 6259
rect 34766 6258 34790 6259
rect 34818 6285 34842 6286
rect 34870 6285 34894 6286
rect 34818 6259 34822 6285
rect 34870 6259 34884 6285
rect 34818 6258 34842 6259
rect 34870 6258 34894 6259
rect 34922 6258 34946 6286
rect 34974 6258 34998 6286
rect 35026 6285 35035 6286
rect 35034 6259 35035 6285
rect 35026 6258 35035 6259
rect 34573 6253 35035 6258
rect 34454 6089 34538 6090
rect 34454 6063 34455 6089
rect 34481 6063 34538 6089
rect 34454 6062 34538 6063
rect 34454 6057 34482 6062
rect 34510 5698 34538 6062
rect 35350 6145 35378 6734
rect 35630 6481 35658 6846
rect 35630 6455 35631 6481
rect 35657 6455 35658 6481
rect 35630 6425 35658 6455
rect 35630 6399 35631 6425
rect 35657 6399 35658 6425
rect 35630 6393 35658 6399
rect 35686 6873 35714 6879
rect 35686 6847 35687 6873
rect 35713 6847 35714 6873
rect 35350 6119 35351 6145
rect 35377 6119 35378 6145
rect 35350 6089 35378 6119
rect 35630 6090 35658 6095
rect 35350 6063 35351 6089
rect 35377 6063 35378 6089
rect 35350 6057 35378 6063
rect 35574 6089 35658 6090
rect 35574 6063 35631 6089
rect 35657 6063 35658 6089
rect 35574 6062 35658 6063
rect 35574 5922 35602 6062
rect 35630 6057 35658 6062
rect 34678 5698 34706 5703
rect 34510 5697 34706 5698
rect 34510 5671 34679 5697
rect 34705 5671 34706 5697
rect 34510 5670 34706 5671
rect 34174 5306 34202 5311
rect 34174 5259 34202 5278
rect 34510 4914 34538 5670
rect 34678 5665 34706 5670
rect 35238 5698 35266 5703
rect 35350 5698 35378 5703
rect 35238 5697 35378 5698
rect 35238 5671 35239 5697
rect 35265 5671 35351 5697
rect 35377 5671 35378 5697
rect 35238 5670 35378 5671
rect 35238 5665 35266 5670
rect 34573 5502 35035 5507
rect 34573 5501 34582 5502
rect 34573 5475 34574 5501
rect 34573 5474 34582 5475
rect 34610 5474 34634 5502
rect 34662 5474 34686 5502
rect 34714 5501 34738 5502
rect 34766 5501 34790 5502
rect 34724 5475 34738 5501
rect 34786 5475 34790 5501
rect 34714 5474 34738 5475
rect 34766 5474 34790 5475
rect 34818 5501 34842 5502
rect 34870 5501 34894 5502
rect 34818 5475 34822 5501
rect 34870 5475 34884 5501
rect 34818 5474 34842 5475
rect 34870 5474 34894 5475
rect 34922 5474 34946 5502
rect 34974 5474 34998 5502
rect 35026 5501 35035 5502
rect 35034 5475 35035 5501
rect 35026 5474 35035 5475
rect 34573 5469 35035 5474
rect 34622 5305 34650 5311
rect 34622 5279 34623 5305
rect 34649 5279 34650 5305
rect 34622 5250 34650 5279
rect 34622 5217 34650 5222
rect 34846 5305 34874 5311
rect 34846 5279 34847 5305
rect 34873 5279 34874 5305
rect 34846 5250 34874 5279
rect 34846 5217 34874 5222
rect 34678 4914 34706 4919
rect 34510 4913 34706 4914
rect 34510 4887 34679 4913
rect 34705 4887 34706 4913
rect 34510 4886 34706 4887
rect 34454 4522 34482 4527
rect 34510 4522 34538 4886
rect 34678 4881 34706 4886
rect 35238 4914 35266 4919
rect 35350 4914 35378 5670
rect 35238 4913 35378 4914
rect 35238 4887 35239 4913
rect 35265 4887 35351 4913
rect 35377 4887 35378 4913
rect 35238 4886 35378 4887
rect 35238 4881 35266 4886
rect 34573 4718 35035 4723
rect 34573 4717 34582 4718
rect 34573 4691 34574 4717
rect 34573 4690 34582 4691
rect 34610 4690 34634 4718
rect 34662 4690 34686 4718
rect 34714 4717 34738 4718
rect 34766 4717 34790 4718
rect 34724 4691 34738 4717
rect 34786 4691 34790 4717
rect 34714 4690 34738 4691
rect 34766 4690 34790 4691
rect 34818 4717 34842 4718
rect 34870 4717 34894 4718
rect 34818 4691 34822 4717
rect 34870 4691 34884 4717
rect 34818 4690 34842 4691
rect 34870 4690 34894 4691
rect 34922 4690 34946 4718
rect 34974 4690 34998 4718
rect 35026 4717 35035 4718
rect 35034 4691 35035 4717
rect 35026 4690 35035 4691
rect 34573 4685 35035 4690
rect 34454 4521 34538 4522
rect 34454 4495 34455 4521
rect 34481 4495 34538 4521
rect 34454 4494 34538 4495
rect 34454 4489 34482 4494
rect 34510 4130 34538 4494
rect 35350 4577 35378 4886
rect 35350 4551 35351 4577
rect 35377 4551 35378 4577
rect 35350 4521 35378 4551
rect 35350 4495 35351 4521
rect 35377 4495 35378 4521
rect 34678 4130 34706 4135
rect 34510 4129 34706 4130
rect 34510 4103 34679 4129
rect 34705 4103 34706 4129
rect 34510 4102 34706 4103
rect 34174 3737 34202 3743
rect 34174 3711 34175 3737
rect 34201 3711 34202 3737
rect 34174 3346 34202 3711
rect 34174 3010 34202 3318
rect 34174 2953 34202 2982
rect 34174 2927 34175 2953
rect 34201 2927 34202 2953
rect 34174 2921 34202 2927
rect 34454 3738 34482 3743
rect 33950 2417 33978 2422
rect 34230 2898 34258 2903
rect 33838 2199 33839 2225
rect 33865 2199 33866 2225
rect 33670 2137 33698 2142
rect 33838 2169 33866 2199
rect 33838 2143 33839 2169
rect 33865 2143 33866 2169
rect 33838 2137 33866 2143
rect 34230 2169 34258 2870
rect 34230 2143 34231 2169
rect 34257 2143 34258 2169
rect 34118 2114 34146 2119
rect 33446 1778 33474 1783
rect 33446 1721 33474 1750
rect 33446 1695 33447 1721
rect 33473 1695 33474 1721
rect 33446 1689 33474 1695
rect 34118 400 34146 2086
rect 34230 1777 34258 2143
rect 34230 1751 34231 1777
rect 34257 1751 34258 1777
rect 34230 1745 34258 1751
rect 34454 1778 34482 3710
rect 34510 3346 34538 4102
rect 34678 4097 34706 4102
rect 34573 3934 35035 3939
rect 34573 3933 34582 3934
rect 34573 3907 34574 3933
rect 34573 3906 34582 3907
rect 34610 3906 34634 3934
rect 34662 3906 34686 3934
rect 34714 3933 34738 3934
rect 34766 3933 34790 3934
rect 34724 3907 34738 3933
rect 34786 3907 34790 3933
rect 34714 3906 34738 3907
rect 34766 3906 34790 3907
rect 34818 3933 34842 3934
rect 34870 3933 34894 3934
rect 34818 3907 34822 3933
rect 34870 3907 34884 3933
rect 34818 3906 34842 3907
rect 34870 3906 34894 3907
rect 34922 3906 34946 3934
rect 34974 3906 34998 3934
rect 35026 3933 35035 3934
rect 35034 3907 35035 3933
rect 35026 3906 35035 3907
rect 34573 3901 35035 3906
rect 35350 3793 35378 4495
rect 35574 4914 35602 5894
rect 35686 5754 35714 6847
rect 35798 6874 35826 6879
rect 35910 6874 35938 6879
rect 35798 6873 35938 6874
rect 35798 6847 35799 6873
rect 35825 6847 35911 6873
rect 35937 6847 35938 6873
rect 35798 6846 35938 6847
rect 35798 6482 35826 6846
rect 35910 6841 35938 6846
rect 36414 6482 36442 7546
rect 36694 6873 36722 7630
rect 37142 7658 37170 7966
rect 37366 7658 37394 7663
rect 37142 7657 37394 7658
rect 37142 7631 37143 7657
rect 37169 7631 37367 7657
rect 37393 7631 37394 7657
rect 37142 7630 37394 7631
rect 37142 7625 37170 7630
rect 37366 7625 37394 7630
rect 37073 7462 37535 7467
rect 37073 7461 37082 7462
rect 37073 7435 37074 7461
rect 37073 7434 37082 7435
rect 37110 7434 37134 7462
rect 37162 7434 37186 7462
rect 37214 7461 37238 7462
rect 37266 7461 37290 7462
rect 37224 7435 37238 7461
rect 37286 7435 37290 7461
rect 37214 7434 37238 7435
rect 37266 7434 37290 7435
rect 37318 7461 37342 7462
rect 37370 7461 37394 7462
rect 37318 7435 37322 7461
rect 37370 7435 37384 7461
rect 37318 7434 37342 7435
rect 37370 7434 37394 7435
rect 37422 7434 37446 7462
rect 37474 7434 37498 7462
rect 37526 7461 37535 7462
rect 37534 7435 37535 7461
rect 37526 7434 37535 7435
rect 37073 7429 37535 7434
rect 36694 6847 36695 6873
rect 36721 6847 36722 6873
rect 36694 6841 36722 6847
rect 36750 7266 36778 7271
rect 35826 6454 35994 6482
rect 35798 6449 35826 6454
rect 35686 5721 35714 5726
rect 35742 6090 35770 6095
rect 35910 6090 35938 6095
rect 35742 6089 35938 6090
rect 35742 6063 35743 6089
rect 35769 6063 35911 6089
rect 35937 6063 35938 6089
rect 35742 6062 35938 6063
rect 35742 5362 35770 6062
rect 35910 6057 35938 6062
rect 35910 5362 35938 5367
rect 35742 5361 35938 5362
rect 35742 5335 35911 5361
rect 35937 5335 35938 5361
rect 35742 5334 35938 5335
rect 35630 5305 35658 5311
rect 35630 5279 35631 5305
rect 35657 5279 35658 5305
rect 35630 5082 35658 5279
rect 35630 5049 35658 5054
rect 35742 5305 35770 5334
rect 35910 5329 35938 5334
rect 35742 5279 35743 5305
rect 35769 5279 35770 5305
rect 35742 5026 35770 5279
rect 35742 4993 35770 4998
rect 35574 4522 35602 4886
rect 35686 4522 35714 4527
rect 35798 4522 35826 4527
rect 35966 4522 35994 6454
rect 36414 6481 36722 6482
rect 36414 6455 36415 6481
rect 36441 6455 36722 6481
rect 36414 6454 36722 6455
rect 36414 6449 36442 6454
rect 36694 6089 36722 6454
rect 36694 6063 36695 6089
rect 36721 6063 36722 6089
rect 36694 6057 36722 6063
rect 35574 4521 35714 4522
rect 35574 4495 35687 4521
rect 35713 4495 35714 4521
rect 35574 4494 35714 4495
rect 35350 3767 35351 3793
rect 35377 3767 35378 3793
rect 35350 3738 35378 3767
rect 34510 3313 34538 3318
rect 34678 3346 34706 3351
rect 34678 3299 34706 3318
rect 34573 3150 35035 3155
rect 34573 3149 34582 3150
rect 34573 3123 34574 3149
rect 34573 3122 34582 3123
rect 34610 3122 34634 3150
rect 34662 3122 34686 3150
rect 34714 3149 34738 3150
rect 34766 3149 34790 3150
rect 34724 3123 34738 3149
rect 34786 3123 34790 3149
rect 34714 3122 34738 3123
rect 34766 3122 34790 3123
rect 34818 3149 34842 3150
rect 34870 3149 34894 3150
rect 34818 3123 34822 3149
rect 34870 3123 34884 3149
rect 34818 3122 34842 3123
rect 34870 3122 34894 3123
rect 34922 3122 34946 3150
rect 34974 3122 34998 3150
rect 35026 3149 35035 3150
rect 35034 3123 35035 3149
rect 35026 3122 35035 3123
rect 34573 3117 35035 3122
rect 34678 3010 34706 3015
rect 34678 2561 34706 2982
rect 35350 3009 35378 3710
rect 35630 4186 35658 4191
rect 35630 3738 35658 4158
rect 35630 3345 35658 3710
rect 35630 3319 35631 3345
rect 35657 3319 35658 3345
rect 35630 3289 35658 3319
rect 35630 3263 35631 3289
rect 35657 3263 35658 3289
rect 35630 3257 35658 3263
rect 35686 3737 35714 4494
rect 35686 3711 35687 3737
rect 35713 3711 35714 3737
rect 35686 3290 35714 3711
rect 35350 2983 35351 3009
rect 35377 2983 35378 3009
rect 35350 2953 35378 2983
rect 35350 2927 35351 2953
rect 35377 2927 35378 2953
rect 35350 2921 35378 2927
rect 35686 2953 35714 3262
rect 35742 4521 35994 4522
rect 35742 4495 35799 4521
rect 35825 4495 35967 4521
rect 35993 4495 35994 4521
rect 35742 4494 35994 4495
rect 35742 3793 35770 4494
rect 35798 4489 35826 4494
rect 35966 4489 35994 4494
rect 36134 5697 36162 5703
rect 36134 5671 36135 5697
rect 36161 5671 36162 5697
rect 36134 4913 36162 5671
rect 36134 4887 36135 4913
rect 36161 4887 36162 4913
rect 35854 4186 35882 4191
rect 35854 4129 35882 4158
rect 35854 4103 35855 4129
rect 35881 4103 35882 4129
rect 35854 4073 35882 4103
rect 35854 4047 35855 4073
rect 35881 4047 35882 4073
rect 35854 4041 35882 4047
rect 36134 4129 36162 4887
rect 36134 4103 36135 4129
rect 36161 4103 36162 4129
rect 35742 3767 35743 3793
rect 35769 3767 35770 3793
rect 35742 3682 35770 3767
rect 35910 3737 35938 3743
rect 35910 3711 35911 3737
rect 35937 3711 35938 3737
rect 35910 3682 35938 3711
rect 35742 3654 35938 3682
rect 35742 3010 35770 3654
rect 36134 3346 36162 4103
rect 36134 3299 36162 3318
rect 36694 5305 36722 5311
rect 36694 5279 36695 5305
rect 36721 5279 36722 5305
rect 36694 4521 36722 5279
rect 36694 4495 36695 4521
rect 36721 4495 36722 4521
rect 36694 3737 36722 4495
rect 36694 3711 36695 3737
rect 36721 3711 36722 3737
rect 36694 3346 36722 3711
rect 36694 3313 36722 3318
rect 35910 3010 35938 3015
rect 35742 3009 35938 3010
rect 35742 2983 35743 3009
rect 35769 2983 35911 3009
rect 35937 2983 35938 3009
rect 35742 2982 35938 2983
rect 35742 2977 35770 2982
rect 35686 2927 35687 2953
rect 35713 2927 35714 2953
rect 35686 2921 35714 2927
rect 35910 2898 35938 2982
rect 36750 2953 36778 7238
rect 37310 7265 37338 7271
rect 37310 7239 37311 7265
rect 37337 7239 37338 7265
rect 37310 7210 37338 7239
rect 37310 7163 37338 7182
rect 37646 7210 37674 7215
rect 37646 6929 37674 7182
rect 37646 6903 37647 6929
rect 37673 6903 37674 6929
rect 37646 6873 37674 6903
rect 37646 6847 37647 6873
rect 37673 6847 37674 6873
rect 37646 6841 37674 6847
rect 37073 6678 37535 6683
rect 37073 6677 37082 6678
rect 37073 6651 37074 6677
rect 37073 6650 37082 6651
rect 37110 6650 37134 6678
rect 37162 6650 37186 6678
rect 37214 6677 37238 6678
rect 37266 6677 37290 6678
rect 37224 6651 37238 6677
rect 37286 6651 37290 6677
rect 37214 6650 37238 6651
rect 37266 6650 37290 6651
rect 37318 6677 37342 6678
rect 37370 6677 37394 6678
rect 37318 6651 37322 6677
rect 37370 6651 37384 6677
rect 37318 6650 37342 6651
rect 37370 6650 37394 6651
rect 37422 6650 37446 6678
rect 37474 6650 37498 6678
rect 37526 6677 37535 6678
rect 37534 6651 37535 6677
rect 37526 6650 37535 6651
rect 37073 6645 37535 6650
rect 37254 6481 37282 6487
rect 37254 6455 37255 6481
rect 37281 6455 37282 6481
rect 37254 6425 37282 6455
rect 37254 6399 37255 6425
rect 37281 6399 37282 6425
rect 37254 6090 37282 6399
rect 37366 6090 37394 6095
rect 37254 6089 37366 6090
rect 37254 6063 37255 6089
rect 37281 6063 37366 6089
rect 37254 6062 37366 6063
rect 37254 6057 37282 6062
rect 37366 6024 37394 6062
rect 37646 6090 37674 6095
rect 37073 5894 37535 5899
rect 37073 5893 37082 5894
rect 37073 5867 37074 5893
rect 37073 5866 37082 5867
rect 37110 5866 37134 5894
rect 37162 5866 37186 5894
rect 37214 5893 37238 5894
rect 37266 5893 37290 5894
rect 37224 5867 37238 5893
rect 37286 5867 37290 5893
rect 37214 5866 37238 5867
rect 37266 5866 37290 5867
rect 37318 5893 37342 5894
rect 37370 5893 37394 5894
rect 37318 5867 37322 5893
rect 37370 5867 37384 5893
rect 37318 5866 37342 5867
rect 37370 5866 37394 5867
rect 37422 5866 37446 5894
rect 37474 5866 37498 5894
rect 37526 5893 37535 5894
rect 37534 5867 37535 5893
rect 37526 5866 37535 5867
rect 37073 5861 37535 5866
rect 37310 5697 37338 5703
rect 37310 5671 37311 5697
rect 37337 5671 37338 5697
rect 37310 5641 37338 5671
rect 37310 5615 37311 5641
rect 37337 5615 37338 5641
rect 37310 5362 37338 5615
rect 37590 5642 37618 5647
rect 37590 5595 37618 5614
rect 37646 5362 37674 6062
rect 37310 5361 37674 5362
rect 37310 5335 37647 5361
rect 37673 5335 37674 5361
rect 37310 5334 37674 5335
rect 37646 5305 37674 5334
rect 37646 5279 37647 5305
rect 37673 5279 37674 5305
rect 37073 5110 37535 5115
rect 37073 5109 37082 5110
rect 37073 5083 37074 5109
rect 37073 5082 37082 5083
rect 37110 5082 37134 5110
rect 37162 5082 37186 5110
rect 37214 5109 37238 5110
rect 37266 5109 37290 5110
rect 37224 5083 37238 5109
rect 37286 5083 37290 5109
rect 37214 5082 37238 5083
rect 37266 5082 37290 5083
rect 37318 5109 37342 5110
rect 37370 5109 37394 5110
rect 37318 5083 37322 5109
rect 37370 5083 37384 5109
rect 37318 5082 37342 5083
rect 37370 5082 37394 5083
rect 37422 5082 37446 5110
rect 37474 5082 37498 5110
rect 37526 5109 37535 5110
rect 37534 5083 37535 5109
rect 37526 5082 37535 5083
rect 37073 5077 37535 5082
rect 37310 4913 37338 4919
rect 37310 4887 37311 4913
rect 37337 4887 37338 4913
rect 37310 4857 37338 4887
rect 37310 4831 37311 4857
rect 37337 4831 37338 4857
rect 37310 4578 37338 4831
rect 37590 4858 37618 4863
rect 37590 4811 37618 4830
rect 37646 4578 37674 5279
rect 37310 4577 37674 4578
rect 37310 4551 37647 4577
rect 37673 4551 37674 4577
rect 37310 4550 37674 4551
rect 37646 4521 37674 4550
rect 37646 4495 37647 4521
rect 37673 4495 37674 4521
rect 37073 4326 37535 4331
rect 37073 4325 37082 4326
rect 37073 4299 37074 4325
rect 37073 4298 37082 4299
rect 37110 4298 37134 4326
rect 37162 4298 37186 4326
rect 37214 4325 37238 4326
rect 37266 4325 37290 4326
rect 37224 4299 37238 4325
rect 37286 4299 37290 4325
rect 37214 4298 37238 4299
rect 37266 4298 37290 4299
rect 37318 4325 37342 4326
rect 37370 4325 37394 4326
rect 37318 4299 37322 4325
rect 37370 4299 37384 4325
rect 37318 4298 37342 4299
rect 37370 4298 37394 4299
rect 37422 4298 37446 4326
rect 37474 4298 37498 4326
rect 37526 4325 37535 4326
rect 37534 4299 37535 4325
rect 37526 4298 37535 4299
rect 37073 4293 37535 4298
rect 37086 4130 37114 4135
rect 37086 4073 37114 4102
rect 37086 4047 37087 4073
rect 37113 4047 37114 4073
rect 37086 4041 37114 4047
rect 37590 4073 37618 4079
rect 37590 4047 37591 4073
rect 37617 4047 37618 4073
rect 37590 3738 37618 4047
rect 37073 3542 37535 3547
rect 37073 3541 37082 3542
rect 37073 3515 37074 3541
rect 37073 3514 37082 3515
rect 37110 3514 37134 3542
rect 37162 3514 37186 3542
rect 37214 3541 37238 3542
rect 37266 3541 37290 3542
rect 37224 3515 37238 3541
rect 37286 3515 37290 3541
rect 37214 3514 37238 3515
rect 37266 3514 37290 3515
rect 37318 3541 37342 3542
rect 37370 3541 37394 3542
rect 37318 3515 37322 3541
rect 37370 3515 37384 3541
rect 37318 3514 37342 3515
rect 37370 3514 37394 3515
rect 37422 3514 37446 3542
rect 37474 3514 37498 3542
rect 37526 3541 37535 3542
rect 37534 3515 37535 3541
rect 37526 3514 37535 3515
rect 37073 3509 37535 3514
rect 37142 3402 37170 3407
rect 37142 2954 37170 3374
rect 37310 3345 37338 3351
rect 37310 3319 37311 3345
rect 37337 3319 37338 3345
rect 37310 3289 37338 3319
rect 37310 3263 37311 3289
rect 37337 3263 37338 3289
rect 37310 3066 37338 3263
rect 37310 3033 37338 3038
rect 37590 3289 37618 3710
rect 37590 3263 37591 3289
rect 37617 3263 37618 3289
rect 37366 2954 37394 2959
rect 36750 2927 36751 2953
rect 36777 2927 36778 2953
rect 36750 2921 36778 2927
rect 36974 2953 37394 2954
rect 36974 2927 37143 2953
rect 37169 2927 37367 2953
rect 37393 2927 37394 2953
rect 36974 2926 37394 2927
rect 35910 2865 35938 2870
rect 34678 2535 34679 2561
rect 34705 2535 34706 2561
rect 34678 2529 34706 2535
rect 35854 2561 35882 2567
rect 35854 2535 35855 2561
rect 35881 2535 35882 2561
rect 35854 2506 35882 2535
rect 35854 2459 35882 2478
rect 36134 2561 36162 2567
rect 36134 2535 36135 2561
rect 36161 2535 36162 2561
rect 34573 2366 35035 2371
rect 34573 2365 34582 2366
rect 34573 2339 34574 2365
rect 34573 2338 34582 2339
rect 34610 2338 34634 2366
rect 34662 2338 34686 2366
rect 34714 2365 34738 2366
rect 34766 2365 34790 2366
rect 34724 2339 34738 2365
rect 34786 2339 34790 2365
rect 34714 2338 34738 2339
rect 34766 2338 34790 2339
rect 34818 2365 34842 2366
rect 34870 2365 34894 2366
rect 34818 2339 34822 2365
rect 34870 2339 34884 2365
rect 34818 2338 34842 2339
rect 34870 2338 34894 2339
rect 34922 2338 34946 2366
rect 34974 2338 34998 2366
rect 35026 2365 35035 2366
rect 35034 2339 35035 2365
rect 35026 2338 35035 2339
rect 34573 2333 35035 2338
rect 36134 2282 36162 2535
rect 36974 2561 37002 2926
rect 37142 2921 37170 2926
rect 37366 2921 37394 2926
rect 37073 2758 37535 2763
rect 37073 2757 37082 2758
rect 37073 2731 37074 2757
rect 37073 2730 37082 2731
rect 37110 2730 37134 2758
rect 37162 2730 37186 2758
rect 37214 2757 37238 2758
rect 37266 2757 37290 2758
rect 37224 2731 37238 2757
rect 37286 2731 37290 2757
rect 37214 2730 37238 2731
rect 37266 2730 37290 2731
rect 37318 2757 37342 2758
rect 37370 2757 37394 2758
rect 37318 2731 37322 2757
rect 37370 2731 37384 2757
rect 37318 2730 37342 2731
rect 37370 2730 37394 2731
rect 37422 2730 37446 2758
rect 37474 2730 37498 2758
rect 37526 2757 37535 2758
rect 37534 2731 37535 2757
rect 37526 2730 37535 2731
rect 37073 2725 37535 2730
rect 37590 2674 37618 3263
rect 36974 2535 36975 2561
rect 37001 2535 37002 2561
rect 36974 2506 37002 2535
rect 37534 2646 37618 2674
rect 37646 3793 37674 4495
rect 37646 3767 37647 3793
rect 37673 3767 37674 3793
rect 37646 3737 37674 3767
rect 37646 3711 37647 3737
rect 37673 3711 37674 3737
rect 37646 3066 37674 3711
rect 37086 2506 37114 2511
rect 36974 2505 37114 2506
rect 36974 2479 37087 2505
rect 37113 2479 37114 2505
rect 36974 2478 37114 2479
rect 34454 1745 34482 1750
rect 35182 2225 35210 2231
rect 35182 2199 35183 2225
rect 35209 2199 35210 2225
rect 35182 2169 35210 2199
rect 35742 2226 35770 2231
rect 35742 2179 35770 2198
rect 35910 2226 35938 2231
rect 35910 2179 35938 2198
rect 35182 2143 35183 2169
rect 35209 2143 35210 2169
rect 35182 1777 35210 2143
rect 35686 2170 35714 2175
rect 35686 2123 35714 2142
rect 35182 1751 35183 1777
rect 35209 1751 35210 1777
rect 35182 1722 35210 1751
rect 35182 1689 35210 1694
rect 35350 1778 35378 1783
rect 36134 1778 36162 2254
rect 36582 2450 36610 2455
rect 36190 1778 36218 1783
rect 36134 1777 36218 1778
rect 36134 1751 36191 1777
rect 36217 1751 36218 1777
rect 36134 1750 36218 1751
rect 34573 1582 35035 1587
rect 34573 1581 34582 1582
rect 34573 1555 34574 1581
rect 34573 1554 34582 1555
rect 34610 1554 34634 1582
rect 34662 1554 34686 1582
rect 34714 1581 34738 1582
rect 34766 1581 34790 1582
rect 34724 1555 34738 1581
rect 34786 1555 34790 1581
rect 34714 1554 34738 1555
rect 34766 1554 34790 1555
rect 34818 1581 34842 1582
rect 34870 1581 34894 1582
rect 34818 1555 34822 1581
rect 34870 1555 34884 1581
rect 34818 1554 34842 1555
rect 34870 1554 34894 1555
rect 34922 1554 34946 1582
rect 34974 1554 34998 1582
rect 35026 1581 35035 1582
rect 35034 1555 35035 1581
rect 35026 1554 35035 1555
rect 34573 1549 35035 1554
rect 35350 400 35378 1750
rect 36190 1745 36218 1750
rect 36582 400 36610 2422
rect 36694 2282 36722 2287
rect 36694 2169 36722 2254
rect 36694 2143 36695 2169
rect 36721 2143 36722 2169
rect 36694 2137 36722 2143
rect 36974 1778 37002 2478
rect 37086 2473 37114 2478
rect 37534 2170 37562 2646
rect 37590 2505 37618 2511
rect 37590 2479 37591 2505
rect 37617 2479 37618 2505
rect 37590 2394 37618 2479
rect 37590 2361 37618 2366
rect 37646 2506 37674 3038
rect 37534 2137 37562 2142
rect 37646 2225 37674 2478
rect 37646 2199 37647 2225
rect 37673 2199 37674 2225
rect 37646 2169 37674 2199
rect 37702 5642 37730 5647
rect 37870 5642 37898 5647
rect 37702 5641 37898 5642
rect 37702 5615 37703 5641
rect 37729 5615 37871 5641
rect 37897 5615 37898 5641
rect 37702 5614 37898 5615
rect 37702 5026 37730 5614
rect 37870 5609 37898 5614
rect 38990 5642 39018 5647
rect 37702 4858 37730 4998
rect 37870 4858 37898 4863
rect 37702 4857 37898 4858
rect 37702 4831 37703 4857
rect 37729 4831 37871 4857
rect 37897 4831 37898 4857
rect 37702 4830 37898 4831
rect 37702 4074 37730 4830
rect 37870 4825 37898 4830
rect 38206 4858 38234 4863
rect 38206 4521 38234 4830
rect 38654 4857 38682 4863
rect 38654 4831 38655 4857
rect 38681 4831 38682 4857
rect 38206 4495 38207 4521
rect 38233 4495 38234 4521
rect 37870 4074 37898 4079
rect 37702 4073 37898 4074
rect 37702 4047 37703 4073
rect 37729 4047 37871 4073
rect 37897 4047 37898 4073
rect 37702 4046 37898 4047
rect 37702 3290 37730 4046
rect 37870 4041 37898 4046
rect 38150 3738 38178 3743
rect 38150 3691 38178 3710
rect 37870 3290 37898 3295
rect 37702 3289 37898 3290
rect 37702 3263 37703 3289
rect 37729 3263 37871 3289
rect 37897 3263 37898 3289
rect 37702 3262 37898 3263
rect 37702 2506 37730 3262
rect 37870 3257 37898 3262
rect 38206 2953 38234 4495
rect 38206 2927 38207 2953
rect 38233 2927 38234 2953
rect 37870 2506 37898 2511
rect 37702 2505 37898 2506
rect 37702 2479 37703 2505
rect 37729 2479 37871 2505
rect 37897 2479 37898 2505
rect 37702 2478 37898 2479
rect 37702 2226 37730 2478
rect 37870 2473 37898 2478
rect 38206 2506 38234 2927
rect 37702 2193 37730 2198
rect 38150 2450 38178 2455
rect 38150 2225 38178 2422
rect 38206 2394 38234 2478
rect 38206 2361 38234 2366
rect 38262 4522 38290 4527
rect 38430 4522 38458 4527
rect 38262 4521 38458 4522
rect 38262 4495 38263 4521
rect 38289 4495 38431 4521
rect 38457 4495 38458 4521
rect 38262 4494 38458 4495
rect 38262 3738 38290 4494
rect 38430 4489 38458 4494
rect 38598 4242 38626 4247
rect 38430 3738 38458 3743
rect 38598 3738 38626 4214
rect 38654 4186 38682 4831
rect 38766 4858 38794 4863
rect 38934 4858 38962 4863
rect 38766 4857 38962 4858
rect 38766 4831 38767 4857
rect 38793 4831 38935 4857
rect 38961 4831 38962 4857
rect 38766 4830 38962 4831
rect 38710 4522 38738 4527
rect 38766 4522 38794 4830
rect 38934 4825 38962 4830
rect 38822 4522 38850 4527
rect 38710 4521 38850 4522
rect 38710 4495 38711 4521
rect 38737 4495 38823 4521
rect 38849 4495 38850 4521
rect 38710 4494 38850 4495
rect 38710 4489 38738 4494
rect 38822 4242 38850 4494
rect 38990 4522 39018 5614
rect 38990 4521 39130 4522
rect 38990 4495 38991 4521
rect 39017 4495 39130 4521
rect 38990 4494 39130 4495
rect 38990 4489 39018 4494
rect 38654 4158 38738 4186
rect 38654 4073 38682 4079
rect 38654 4047 38655 4073
rect 38681 4047 38682 4073
rect 38654 3962 38682 4047
rect 38654 3929 38682 3934
rect 38654 3738 38682 3743
rect 38262 3737 38654 3738
rect 38262 3711 38263 3737
rect 38289 3711 38431 3737
rect 38457 3711 38654 3737
rect 38262 3710 38654 3711
rect 38262 3010 38290 3710
rect 38430 3705 38458 3710
rect 38654 3672 38682 3710
rect 38654 3289 38682 3295
rect 38654 3263 38655 3289
rect 38681 3263 38682 3289
rect 38430 3010 38458 3015
rect 38262 3009 38458 3010
rect 38262 2983 38431 3009
rect 38457 2983 38458 3009
rect 38262 2982 38458 2983
rect 38262 2953 38290 2982
rect 38430 2977 38458 2982
rect 38262 2927 38263 2953
rect 38289 2927 38290 2953
rect 38150 2199 38151 2225
rect 38177 2199 38178 2225
rect 37646 2143 37647 2169
rect 37673 2143 37674 2169
rect 37646 2137 37674 2143
rect 37814 2170 37842 2175
rect 37073 1974 37535 1979
rect 37073 1973 37082 1974
rect 37073 1947 37074 1973
rect 37073 1946 37082 1947
rect 37110 1946 37134 1974
rect 37162 1946 37186 1974
rect 37214 1973 37238 1974
rect 37266 1973 37290 1974
rect 37224 1947 37238 1973
rect 37286 1947 37290 1973
rect 37214 1946 37238 1947
rect 37266 1946 37290 1947
rect 37318 1973 37342 1974
rect 37370 1973 37394 1974
rect 37318 1947 37322 1973
rect 37370 1947 37384 1973
rect 37318 1946 37342 1947
rect 37370 1946 37394 1947
rect 37422 1946 37446 1974
rect 37474 1946 37498 1974
rect 37526 1973 37535 1974
rect 37534 1947 37535 1973
rect 37526 1946 37535 1947
rect 37073 1941 37535 1946
rect 36974 1777 37170 1778
rect 36974 1751 36975 1777
rect 37001 1751 37170 1777
rect 36974 1750 37170 1751
rect 36974 1745 37002 1750
rect 37142 1721 37170 1750
rect 37142 1695 37143 1721
rect 37169 1695 37170 1721
rect 37142 1689 37170 1695
rect 37814 400 37842 2142
rect 38150 2170 38178 2199
rect 38150 1777 38178 2142
rect 38150 1751 38151 1777
rect 38177 1751 38178 1777
rect 38150 1745 38178 1751
rect 38262 2226 38290 2927
rect 38654 2953 38682 3263
rect 38654 2927 38655 2953
rect 38681 2927 38682 2953
rect 38262 1778 38290 2198
rect 38318 2898 38346 2903
rect 38318 2226 38346 2870
rect 38654 2898 38682 2927
rect 38654 2562 38682 2870
rect 38710 2674 38738 4158
rect 38822 4130 38850 4214
rect 38934 4130 38962 4135
rect 38822 4129 38962 4130
rect 38822 4103 38823 4129
rect 38849 4103 38935 4129
rect 38961 4103 38962 4129
rect 38822 4102 38962 4103
rect 38822 4097 38850 4102
rect 38934 4097 38962 4102
rect 38934 3962 38962 3967
rect 38822 3738 38850 3743
rect 38822 3691 38850 3710
rect 38822 3289 38850 3295
rect 38822 3263 38823 3289
rect 38849 3263 38850 3289
rect 38822 2953 38850 3263
rect 38822 2927 38823 2953
rect 38849 2927 38850 2953
rect 38822 2898 38850 2927
rect 38822 2865 38850 2870
rect 38934 3289 38962 3934
rect 38990 3738 39018 3743
rect 38990 3737 39074 3738
rect 38990 3711 38991 3737
rect 39017 3711 39074 3737
rect 38990 3710 39074 3711
rect 38990 3705 39018 3710
rect 38934 3263 38935 3289
rect 38961 3263 38962 3289
rect 38934 2953 38962 3263
rect 38934 2927 38935 2953
rect 38961 2927 38962 2953
rect 38710 2646 38850 2674
rect 38766 2562 38794 2567
rect 38654 2561 38794 2562
rect 38654 2535 38655 2561
rect 38681 2535 38767 2561
rect 38793 2535 38794 2561
rect 38654 2534 38794 2535
rect 38430 2226 38458 2231
rect 38318 2225 38458 2226
rect 38318 2199 38431 2225
rect 38457 2199 38458 2225
rect 38318 2198 38458 2199
rect 38318 2169 38346 2198
rect 38430 2193 38458 2198
rect 38318 2143 38319 2169
rect 38345 2143 38346 2169
rect 38318 2137 38346 2143
rect 38430 1778 38458 1783
rect 38262 1777 38458 1778
rect 38262 1751 38263 1777
rect 38289 1751 38431 1777
rect 38457 1751 38458 1777
rect 38262 1750 38458 1751
rect 38262 1745 38290 1750
rect 38430 1745 38458 1750
rect 38654 1778 38682 2534
rect 38766 2529 38794 2534
rect 38710 2226 38738 2231
rect 38710 2179 38738 2198
rect 38822 2114 38850 2646
rect 38934 2505 38962 2927
rect 38934 2479 38935 2505
rect 38961 2479 38962 2505
rect 38878 2226 38906 2231
rect 38878 2179 38906 2198
rect 38934 2170 38962 2479
rect 38934 2123 38962 2142
rect 39046 2506 39074 3710
rect 38822 2081 38850 2086
rect 38822 1778 38850 1783
rect 38654 1777 38850 1778
rect 38654 1751 38655 1777
rect 38681 1751 38823 1777
rect 38849 1751 38850 1777
rect 38654 1750 38850 1751
rect 38654 1745 38682 1750
rect 38822 1745 38850 1750
rect 38934 1778 38962 1783
rect 38934 1731 38962 1750
rect 39046 400 39074 2478
rect 39102 1778 39130 4494
rect 39102 1745 39130 1750
rect 28798 350 29050 378
rect 29176 0 29232 400
rect 30408 0 30464 400
rect 31640 0 31696 400
rect 32872 0 32928 400
rect 34104 0 34160 400
rect 35336 0 35392 400
rect 36568 0 36624 400
rect 37800 0 37856 400
rect 39032 0 39088 400
<< via2 >>
rect 2082 18437 2110 18438
rect 2082 18411 2100 18437
rect 2100 18411 2110 18437
rect 2082 18410 2110 18411
rect 2134 18437 2162 18438
rect 2134 18411 2136 18437
rect 2136 18411 2162 18437
rect 2134 18410 2162 18411
rect 2186 18437 2214 18438
rect 2238 18437 2266 18438
rect 2186 18411 2198 18437
rect 2198 18411 2214 18437
rect 2238 18411 2260 18437
rect 2260 18411 2266 18437
rect 2186 18410 2214 18411
rect 2238 18410 2266 18411
rect 2290 18410 2318 18438
rect 2342 18437 2370 18438
rect 2394 18437 2422 18438
rect 2342 18411 2348 18437
rect 2348 18411 2370 18437
rect 2394 18411 2410 18437
rect 2410 18411 2422 18437
rect 2342 18410 2370 18411
rect 2394 18410 2422 18411
rect 2446 18437 2474 18438
rect 2446 18411 2472 18437
rect 2472 18411 2474 18437
rect 2446 18410 2474 18411
rect 2498 18437 2526 18438
rect 2498 18411 2508 18437
rect 2508 18411 2526 18437
rect 2498 18410 2526 18411
rect 2082 17653 2110 17654
rect 2082 17627 2100 17653
rect 2100 17627 2110 17653
rect 2082 17626 2110 17627
rect 2134 17653 2162 17654
rect 2134 17627 2136 17653
rect 2136 17627 2162 17653
rect 2134 17626 2162 17627
rect 2186 17653 2214 17654
rect 2238 17653 2266 17654
rect 2186 17627 2198 17653
rect 2198 17627 2214 17653
rect 2238 17627 2260 17653
rect 2260 17627 2266 17653
rect 2186 17626 2214 17627
rect 2238 17626 2266 17627
rect 2290 17626 2318 17654
rect 2342 17653 2370 17654
rect 2394 17653 2422 17654
rect 2342 17627 2348 17653
rect 2348 17627 2370 17653
rect 2394 17627 2410 17653
rect 2410 17627 2422 17653
rect 2342 17626 2370 17627
rect 2394 17626 2422 17627
rect 2446 17653 2474 17654
rect 2446 17627 2472 17653
rect 2472 17627 2474 17653
rect 2446 17626 2474 17627
rect 2498 17653 2526 17654
rect 2498 17627 2508 17653
rect 2508 17627 2526 17653
rect 2498 17626 2526 17627
rect 2082 16869 2110 16870
rect 2082 16843 2100 16869
rect 2100 16843 2110 16869
rect 2082 16842 2110 16843
rect 2134 16869 2162 16870
rect 2134 16843 2136 16869
rect 2136 16843 2162 16869
rect 2134 16842 2162 16843
rect 2186 16869 2214 16870
rect 2238 16869 2266 16870
rect 2186 16843 2198 16869
rect 2198 16843 2214 16869
rect 2238 16843 2260 16869
rect 2260 16843 2266 16869
rect 2186 16842 2214 16843
rect 2238 16842 2266 16843
rect 2290 16842 2318 16870
rect 2342 16869 2370 16870
rect 2394 16869 2422 16870
rect 2342 16843 2348 16869
rect 2348 16843 2370 16869
rect 2394 16843 2410 16869
rect 2410 16843 2422 16869
rect 2342 16842 2370 16843
rect 2394 16842 2422 16843
rect 2446 16869 2474 16870
rect 2446 16843 2472 16869
rect 2472 16843 2474 16869
rect 2446 16842 2474 16843
rect 2498 16869 2526 16870
rect 2498 16843 2508 16869
rect 2508 16843 2526 16869
rect 2498 16842 2526 16843
rect 2082 16085 2110 16086
rect 2082 16059 2100 16085
rect 2100 16059 2110 16085
rect 2082 16058 2110 16059
rect 2134 16085 2162 16086
rect 2134 16059 2136 16085
rect 2136 16059 2162 16085
rect 2134 16058 2162 16059
rect 2186 16085 2214 16086
rect 2238 16085 2266 16086
rect 2186 16059 2198 16085
rect 2198 16059 2214 16085
rect 2238 16059 2260 16085
rect 2260 16059 2266 16085
rect 2186 16058 2214 16059
rect 2238 16058 2266 16059
rect 2290 16058 2318 16086
rect 2342 16085 2370 16086
rect 2394 16085 2422 16086
rect 2342 16059 2348 16085
rect 2348 16059 2370 16085
rect 2394 16059 2410 16085
rect 2410 16059 2422 16085
rect 2342 16058 2370 16059
rect 2394 16058 2422 16059
rect 2446 16085 2474 16086
rect 2446 16059 2472 16085
rect 2472 16059 2474 16085
rect 2446 16058 2474 16059
rect 2498 16085 2526 16086
rect 2498 16059 2508 16085
rect 2508 16059 2526 16085
rect 2498 16058 2526 16059
rect 2082 15301 2110 15302
rect 2082 15275 2100 15301
rect 2100 15275 2110 15301
rect 2082 15274 2110 15275
rect 2134 15301 2162 15302
rect 2134 15275 2136 15301
rect 2136 15275 2162 15301
rect 2134 15274 2162 15275
rect 2186 15301 2214 15302
rect 2238 15301 2266 15302
rect 2186 15275 2198 15301
rect 2198 15275 2214 15301
rect 2238 15275 2260 15301
rect 2260 15275 2266 15301
rect 2186 15274 2214 15275
rect 2238 15274 2266 15275
rect 2290 15274 2318 15302
rect 2342 15301 2370 15302
rect 2394 15301 2422 15302
rect 2342 15275 2348 15301
rect 2348 15275 2370 15301
rect 2394 15275 2410 15301
rect 2410 15275 2422 15301
rect 2342 15274 2370 15275
rect 2394 15274 2422 15275
rect 2446 15301 2474 15302
rect 2446 15275 2472 15301
rect 2472 15275 2474 15301
rect 2446 15274 2474 15275
rect 2498 15301 2526 15302
rect 2498 15275 2508 15301
rect 2508 15275 2526 15301
rect 2498 15274 2526 15275
rect 2422 14686 2450 14714
rect 2590 14686 2618 14714
rect 2082 14517 2110 14518
rect 2082 14491 2100 14517
rect 2100 14491 2110 14517
rect 2082 14490 2110 14491
rect 2134 14517 2162 14518
rect 2134 14491 2136 14517
rect 2136 14491 2162 14517
rect 2134 14490 2162 14491
rect 2186 14517 2214 14518
rect 2238 14517 2266 14518
rect 2186 14491 2198 14517
rect 2198 14491 2214 14517
rect 2238 14491 2260 14517
rect 2260 14491 2266 14517
rect 2186 14490 2214 14491
rect 2238 14490 2266 14491
rect 2290 14490 2318 14518
rect 2342 14517 2370 14518
rect 2394 14517 2422 14518
rect 2342 14491 2348 14517
rect 2348 14491 2370 14517
rect 2394 14491 2410 14517
rect 2410 14491 2422 14517
rect 2342 14490 2370 14491
rect 2394 14490 2422 14491
rect 2446 14517 2474 14518
rect 2446 14491 2472 14517
rect 2472 14491 2474 14517
rect 2446 14490 2474 14491
rect 2498 14517 2526 14518
rect 2498 14491 2508 14517
rect 2508 14491 2526 14517
rect 2498 14490 2526 14491
rect 2478 14350 2506 14378
rect 2422 14321 2450 14322
rect 2422 14295 2423 14321
rect 2423 14295 2449 14321
rect 2449 14295 2450 14321
rect 2422 14294 2450 14295
rect 2590 14294 2618 14322
rect 2082 13733 2110 13734
rect 2082 13707 2100 13733
rect 2100 13707 2110 13733
rect 2082 13706 2110 13707
rect 2134 13733 2162 13734
rect 2134 13707 2136 13733
rect 2136 13707 2162 13733
rect 2134 13706 2162 13707
rect 2186 13733 2214 13734
rect 2238 13733 2266 13734
rect 2186 13707 2198 13733
rect 2198 13707 2214 13733
rect 2238 13707 2260 13733
rect 2260 13707 2266 13733
rect 2186 13706 2214 13707
rect 2238 13706 2266 13707
rect 2290 13706 2318 13734
rect 2342 13733 2370 13734
rect 2394 13733 2422 13734
rect 2342 13707 2348 13733
rect 2348 13707 2370 13733
rect 2394 13707 2410 13733
rect 2410 13707 2422 13733
rect 2342 13706 2370 13707
rect 2394 13706 2422 13707
rect 2446 13733 2474 13734
rect 2446 13707 2472 13733
rect 2472 13707 2474 13733
rect 2446 13706 2474 13707
rect 2498 13733 2526 13734
rect 2498 13707 2508 13733
rect 2508 13707 2526 13733
rect 2498 13706 2526 13707
rect 1974 13118 2002 13146
rect 4582 18045 4610 18046
rect 4582 18019 4600 18045
rect 4600 18019 4610 18045
rect 4582 18018 4610 18019
rect 4634 18045 4662 18046
rect 4634 18019 4636 18045
rect 4636 18019 4662 18045
rect 4634 18018 4662 18019
rect 4686 18045 4714 18046
rect 4738 18045 4766 18046
rect 4686 18019 4698 18045
rect 4698 18019 4714 18045
rect 4738 18019 4760 18045
rect 4760 18019 4766 18045
rect 4686 18018 4714 18019
rect 4738 18018 4766 18019
rect 4790 18018 4818 18046
rect 4842 18045 4870 18046
rect 4894 18045 4922 18046
rect 4842 18019 4848 18045
rect 4848 18019 4870 18045
rect 4894 18019 4910 18045
rect 4910 18019 4922 18045
rect 4842 18018 4870 18019
rect 4894 18018 4922 18019
rect 4946 18045 4974 18046
rect 4946 18019 4972 18045
rect 4972 18019 4974 18045
rect 4946 18018 4974 18019
rect 4998 18045 5026 18046
rect 4998 18019 5008 18045
rect 5008 18019 5026 18045
rect 4998 18018 5026 18019
rect 4582 17261 4610 17262
rect 4582 17235 4600 17261
rect 4600 17235 4610 17261
rect 4582 17234 4610 17235
rect 4634 17261 4662 17262
rect 4634 17235 4636 17261
rect 4636 17235 4662 17261
rect 4634 17234 4662 17235
rect 4686 17261 4714 17262
rect 4738 17261 4766 17262
rect 4686 17235 4698 17261
rect 4698 17235 4714 17261
rect 4738 17235 4760 17261
rect 4760 17235 4766 17261
rect 4686 17234 4714 17235
rect 4738 17234 4766 17235
rect 4790 17234 4818 17262
rect 4842 17261 4870 17262
rect 4894 17261 4922 17262
rect 4842 17235 4848 17261
rect 4848 17235 4870 17261
rect 4894 17235 4910 17261
rect 4910 17235 4922 17261
rect 4842 17234 4870 17235
rect 4894 17234 4922 17235
rect 4946 17261 4974 17262
rect 4946 17235 4972 17261
rect 4972 17235 4974 17261
rect 4946 17234 4974 17235
rect 4998 17261 5026 17262
rect 4998 17235 5008 17261
rect 5008 17235 5026 17261
rect 4998 17234 5026 17235
rect 4582 16477 4610 16478
rect 4582 16451 4600 16477
rect 4600 16451 4610 16477
rect 4582 16450 4610 16451
rect 4634 16477 4662 16478
rect 4634 16451 4636 16477
rect 4636 16451 4662 16477
rect 4634 16450 4662 16451
rect 4686 16477 4714 16478
rect 4738 16477 4766 16478
rect 4686 16451 4698 16477
rect 4698 16451 4714 16477
rect 4738 16451 4760 16477
rect 4760 16451 4766 16477
rect 4686 16450 4714 16451
rect 4738 16450 4766 16451
rect 4790 16450 4818 16478
rect 4842 16477 4870 16478
rect 4894 16477 4922 16478
rect 4842 16451 4848 16477
rect 4848 16451 4870 16477
rect 4894 16451 4910 16477
rect 4910 16451 4922 16477
rect 4842 16450 4870 16451
rect 4894 16450 4922 16451
rect 4946 16477 4974 16478
rect 4946 16451 4972 16477
rect 4972 16451 4974 16477
rect 4946 16450 4974 16451
rect 4998 16477 5026 16478
rect 4998 16451 5008 16477
rect 5008 16451 5026 16477
rect 4998 16450 5026 16451
rect 7082 18437 7110 18438
rect 7082 18411 7100 18437
rect 7100 18411 7110 18437
rect 7082 18410 7110 18411
rect 7134 18437 7162 18438
rect 7134 18411 7136 18437
rect 7136 18411 7162 18437
rect 7134 18410 7162 18411
rect 7186 18437 7214 18438
rect 7238 18437 7266 18438
rect 7186 18411 7198 18437
rect 7198 18411 7214 18437
rect 7238 18411 7260 18437
rect 7260 18411 7266 18437
rect 7186 18410 7214 18411
rect 7238 18410 7266 18411
rect 7290 18410 7318 18438
rect 7342 18437 7370 18438
rect 7394 18437 7422 18438
rect 7342 18411 7348 18437
rect 7348 18411 7370 18437
rect 7394 18411 7410 18437
rect 7410 18411 7422 18437
rect 7342 18410 7370 18411
rect 7394 18410 7422 18411
rect 7446 18437 7474 18438
rect 7446 18411 7472 18437
rect 7472 18411 7474 18437
rect 7446 18410 7474 18411
rect 7498 18437 7526 18438
rect 7498 18411 7508 18437
rect 7508 18411 7526 18437
rect 7498 18410 7526 18411
rect 12082 18437 12110 18438
rect 12082 18411 12100 18437
rect 12100 18411 12110 18437
rect 12082 18410 12110 18411
rect 12134 18437 12162 18438
rect 12134 18411 12136 18437
rect 12136 18411 12162 18437
rect 12134 18410 12162 18411
rect 12186 18437 12214 18438
rect 12238 18437 12266 18438
rect 12186 18411 12198 18437
rect 12198 18411 12214 18437
rect 12238 18411 12260 18437
rect 12260 18411 12266 18437
rect 12186 18410 12214 18411
rect 12238 18410 12266 18411
rect 12290 18410 12318 18438
rect 12342 18437 12370 18438
rect 12394 18437 12422 18438
rect 12342 18411 12348 18437
rect 12348 18411 12370 18437
rect 12394 18411 12410 18437
rect 12410 18411 12422 18437
rect 12342 18410 12370 18411
rect 12394 18410 12422 18411
rect 12446 18437 12474 18438
rect 12446 18411 12472 18437
rect 12472 18411 12474 18437
rect 12446 18410 12474 18411
rect 12498 18437 12526 18438
rect 12498 18411 12508 18437
rect 12508 18411 12526 18437
rect 12498 18410 12526 18411
rect 9582 18045 9610 18046
rect 9582 18019 9600 18045
rect 9600 18019 9610 18045
rect 9582 18018 9610 18019
rect 9634 18045 9662 18046
rect 9634 18019 9636 18045
rect 9636 18019 9662 18045
rect 9634 18018 9662 18019
rect 9686 18045 9714 18046
rect 9738 18045 9766 18046
rect 9686 18019 9698 18045
rect 9698 18019 9714 18045
rect 9738 18019 9760 18045
rect 9760 18019 9766 18045
rect 9686 18018 9714 18019
rect 9738 18018 9766 18019
rect 9790 18018 9818 18046
rect 9842 18045 9870 18046
rect 9894 18045 9922 18046
rect 9842 18019 9848 18045
rect 9848 18019 9870 18045
rect 9894 18019 9910 18045
rect 9910 18019 9922 18045
rect 9842 18018 9870 18019
rect 9894 18018 9922 18019
rect 9946 18045 9974 18046
rect 9946 18019 9972 18045
rect 9972 18019 9974 18045
rect 9946 18018 9974 18019
rect 9998 18045 10026 18046
rect 9998 18019 10008 18045
rect 10008 18019 10026 18045
rect 9998 18018 10026 18019
rect 14582 18045 14610 18046
rect 14582 18019 14600 18045
rect 14600 18019 14610 18045
rect 14582 18018 14610 18019
rect 14634 18045 14662 18046
rect 14634 18019 14636 18045
rect 14636 18019 14662 18045
rect 14634 18018 14662 18019
rect 14686 18045 14714 18046
rect 14738 18045 14766 18046
rect 14686 18019 14698 18045
rect 14698 18019 14714 18045
rect 14738 18019 14760 18045
rect 14760 18019 14766 18045
rect 14686 18018 14714 18019
rect 14738 18018 14766 18019
rect 14790 18018 14818 18046
rect 14842 18045 14870 18046
rect 14894 18045 14922 18046
rect 14842 18019 14848 18045
rect 14848 18019 14870 18045
rect 14894 18019 14910 18045
rect 14910 18019 14922 18045
rect 14842 18018 14870 18019
rect 14894 18018 14922 18019
rect 14946 18045 14974 18046
rect 14946 18019 14972 18045
rect 14972 18019 14974 18045
rect 14946 18018 14974 18019
rect 14998 18045 15026 18046
rect 14998 18019 15008 18045
rect 15008 18019 15026 18045
rect 14998 18018 15026 18019
rect 7082 17653 7110 17654
rect 7082 17627 7100 17653
rect 7100 17627 7110 17653
rect 7082 17626 7110 17627
rect 7134 17653 7162 17654
rect 7134 17627 7136 17653
rect 7136 17627 7162 17653
rect 7134 17626 7162 17627
rect 7186 17653 7214 17654
rect 7238 17653 7266 17654
rect 7186 17627 7198 17653
rect 7198 17627 7214 17653
rect 7238 17627 7260 17653
rect 7260 17627 7266 17653
rect 7186 17626 7214 17627
rect 7238 17626 7266 17627
rect 7290 17626 7318 17654
rect 7342 17653 7370 17654
rect 7394 17653 7422 17654
rect 7342 17627 7348 17653
rect 7348 17627 7370 17653
rect 7394 17627 7410 17653
rect 7410 17627 7422 17653
rect 7342 17626 7370 17627
rect 7394 17626 7422 17627
rect 7446 17653 7474 17654
rect 7446 17627 7472 17653
rect 7472 17627 7474 17653
rect 7446 17626 7474 17627
rect 7498 17653 7526 17654
rect 7498 17627 7508 17653
rect 7508 17627 7526 17653
rect 7498 17626 7526 17627
rect 12082 17653 12110 17654
rect 12082 17627 12100 17653
rect 12100 17627 12110 17653
rect 12082 17626 12110 17627
rect 12134 17653 12162 17654
rect 12134 17627 12136 17653
rect 12136 17627 12162 17653
rect 12134 17626 12162 17627
rect 12186 17653 12214 17654
rect 12238 17653 12266 17654
rect 12186 17627 12198 17653
rect 12198 17627 12214 17653
rect 12238 17627 12260 17653
rect 12260 17627 12266 17653
rect 12186 17626 12214 17627
rect 12238 17626 12266 17627
rect 12290 17626 12318 17654
rect 12342 17653 12370 17654
rect 12394 17653 12422 17654
rect 12342 17627 12348 17653
rect 12348 17627 12370 17653
rect 12394 17627 12410 17653
rect 12410 17627 12422 17653
rect 12342 17626 12370 17627
rect 12394 17626 12422 17627
rect 12446 17653 12474 17654
rect 12446 17627 12472 17653
rect 12472 17627 12474 17653
rect 12446 17626 12474 17627
rect 12498 17653 12526 17654
rect 12498 17627 12508 17653
rect 12508 17627 12526 17653
rect 12498 17626 12526 17627
rect 9582 17261 9610 17262
rect 9582 17235 9600 17261
rect 9600 17235 9610 17261
rect 9582 17234 9610 17235
rect 9634 17261 9662 17262
rect 9634 17235 9636 17261
rect 9636 17235 9662 17261
rect 9634 17234 9662 17235
rect 9686 17261 9714 17262
rect 9738 17261 9766 17262
rect 9686 17235 9698 17261
rect 9698 17235 9714 17261
rect 9738 17235 9760 17261
rect 9760 17235 9766 17261
rect 9686 17234 9714 17235
rect 9738 17234 9766 17235
rect 9790 17234 9818 17262
rect 9842 17261 9870 17262
rect 9894 17261 9922 17262
rect 9842 17235 9848 17261
rect 9848 17235 9870 17261
rect 9894 17235 9910 17261
rect 9910 17235 9922 17261
rect 9842 17234 9870 17235
rect 9894 17234 9922 17235
rect 9946 17261 9974 17262
rect 9946 17235 9972 17261
rect 9972 17235 9974 17261
rect 9946 17234 9974 17235
rect 9998 17261 10026 17262
rect 9998 17235 10008 17261
rect 10008 17235 10026 17261
rect 9998 17234 10026 17235
rect 7082 16869 7110 16870
rect 7082 16843 7100 16869
rect 7100 16843 7110 16869
rect 7082 16842 7110 16843
rect 7134 16869 7162 16870
rect 7134 16843 7136 16869
rect 7136 16843 7162 16869
rect 7134 16842 7162 16843
rect 7186 16869 7214 16870
rect 7238 16869 7266 16870
rect 7186 16843 7198 16869
rect 7198 16843 7214 16869
rect 7238 16843 7260 16869
rect 7260 16843 7266 16869
rect 7186 16842 7214 16843
rect 7238 16842 7266 16843
rect 7290 16842 7318 16870
rect 7342 16869 7370 16870
rect 7394 16869 7422 16870
rect 7342 16843 7348 16869
rect 7348 16843 7370 16869
rect 7394 16843 7410 16869
rect 7410 16843 7422 16869
rect 7342 16842 7370 16843
rect 7394 16842 7422 16843
rect 7446 16869 7474 16870
rect 7446 16843 7472 16869
rect 7472 16843 7474 16869
rect 7446 16842 7474 16843
rect 7498 16869 7526 16870
rect 7498 16843 7508 16869
rect 7508 16843 7526 16869
rect 7498 16842 7526 16843
rect 5894 16254 5922 16282
rect 6118 16281 6146 16282
rect 6118 16255 6119 16281
rect 6119 16255 6145 16281
rect 6145 16255 6146 16281
rect 6118 16254 6146 16255
rect 7518 16281 7546 16282
rect 7518 16255 7519 16281
rect 7519 16255 7545 16281
rect 7545 16255 7546 16281
rect 7518 16254 7546 16255
rect 7082 16085 7110 16086
rect 7082 16059 7100 16085
rect 7100 16059 7110 16085
rect 7082 16058 7110 16059
rect 7134 16085 7162 16086
rect 7134 16059 7136 16085
rect 7136 16059 7162 16085
rect 7134 16058 7162 16059
rect 7186 16085 7214 16086
rect 7238 16085 7266 16086
rect 7186 16059 7198 16085
rect 7198 16059 7214 16085
rect 7238 16059 7260 16085
rect 7260 16059 7266 16085
rect 7186 16058 7214 16059
rect 7238 16058 7266 16059
rect 7290 16058 7318 16086
rect 7342 16085 7370 16086
rect 7394 16085 7422 16086
rect 7342 16059 7348 16085
rect 7348 16059 7370 16085
rect 7394 16059 7410 16085
rect 7410 16059 7422 16085
rect 7342 16058 7370 16059
rect 7394 16058 7422 16059
rect 7446 16085 7474 16086
rect 7446 16059 7472 16085
rect 7472 16059 7474 16085
rect 7446 16058 7474 16059
rect 7498 16085 7526 16086
rect 7498 16059 7508 16085
rect 7508 16059 7526 16085
rect 7498 16058 7526 16059
rect 4582 15693 4610 15694
rect 4582 15667 4600 15693
rect 4600 15667 4610 15693
rect 4582 15666 4610 15667
rect 4634 15693 4662 15694
rect 4634 15667 4636 15693
rect 4636 15667 4662 15693
rect 4634 15666 4662 15667
rect 4686 15693 4714 15694
rect 4738 15693 4766 15694
rect 4686 15667 4698 15693
rect 4698 15667 4714 15693
rect 4738 15667 4760 15693
rect 4760 15667 4766 15693
rect 4686 15666 4714 15667
rect 4738 15666 4766 15667
rect 4790 15666 4818 15694
rect 4842 15693 4870 15694
rect 4894 15693 4922 15694
rect 4842 15667 4848 15693
rect 4848 15667 4870 15693
rect 4894 15667 4910 15693
rect 4910 15667 4922 15693
rect 4842 15666 4870 15667
rect 4894 15666 4922 15667
rect 4946 15693 4974 15694
rect 4946 15667 4972 15693
rect 4972 15667 4974 15693
rect 4946 15666 4974 15667
rect 4998 15693 5026 15694
rect 4998 15667 5008 15693
rect 5008 15667 5026 15693
rect 4998 15666 5026 15667
rect 3038 14713 3066 14714
rect 3038 14687 3039 14713
rect 3039 14687 3065 14713
rect 3065 14687 3066 14713
rect 3038 14686 3066 14687
rect 3598 14713 3626 14714
rect 3598 14687 3599 14713
rect 3599 14687 3625 14713
rect 3625 14687 3626 14713
rect 3598 14686 3626 14687
rect 3822 14630 3850 14658
rect 4582 14909 4610 14910
rect 4582 14883 4600 14909
rect 4600 14883 4610 14909
rect 4582 14882 4610 14883
rect 4634 14909 4662 14910
rect 4634 14883 4636 14909
rect 4636 14883 4662 14909
rect 4634 14882 4662 14883
rect 4686 14909 4714 14910
rect 4738 14909 4766 14910
rect 4686 14883 4698 14909
rect 4698 14883 4714 14909
rect 4738 14883 4760 14909
rect 4760 14883 4766 14909
rect 4686 14882 4714 14883
rect 4738 14882 4766 14883
rect 4790 14882 4818 14910
rect 4842 14909 4870 14910
rect 4894 14909 4922 14910
rect 4842 14883 4848 14909
rect 4848 14883 4870 14909
rect 4894 14883 4910 14909
rect 4910 14883 4922 14909
rect 4842 14882 4870 14883
rect 4894 14882 4922 14883
rect 4946 14909 4974 14910
rect 4946 14883 4972 14909
rect 4972 14883 4974 14909
rect 4946 14882 4974 14883
rect 4998 14909 5026 14910
rect 4998 14883 5008 14909
rect 5008 14883 5026 14909
rect 4998 14882 5026 14883
rect 5278 14686 5306 14714
rect 4494 14350 4522 14378
rect 3822 14321 3850 14322
rect 3822 14295 3823 14321
rect 3823 14295 3849 14321
rect 3849 14295 3850 14321
rect 3822 14294 3850 14295
rect 3374 13398 3402 13426
rect 2366 13145 2394 13146
rect 2366 13119 2367 13145
rect 2367 13119 2393 13145
rect 2393 13119 2394 13145
rect 2366 13118 2394 13119
rect 2082 12949 2110 12950
rect 2082 12923 2100 12949
rect 2100 12923 2110 12949
rect 2082 12922 2110 12923
rect 2134 12949 2162 12950
rect 2134 12923 2136 12949
rect 2136 12923 2162 12949
rect 2134 12922 2162 12923
rect 2186 12949 2214 12950
rect 2238 12949 2266 12950
rect 2186 12923 2198 12949
rect 2198 12923 2214 12949
rect 2238 12923 2260 12949
rect 2260 12923 2266 12949
rect 2186 12922 2214 12923
rect 2238 12922 2266 12923
rect 2290 12922 2318 12950
rect 2342 12949 2370 12950
rect 2394 12949 2422 12950
rect 2342 12923 2348 12949
rect 2348 12923 2370 12949
rect 2394 12923 2410 12949
rect 2410 12923 2422 12949
rect 2342 12922 2370 12923
rect 2394 12922 2422 12923
rect 2446 12949 2474 12950
rect 2446 12923 2472 12949
rect 2472 12923 2474 12949
rect 2446 12922 2474 12923
rect 2498 12949 2526 12950
rect 2498 12923 2508 12949
rect 2508 12923 2526 12949
rect 2498 12922 2526 12923
rect 2198 12670 2226 12698
rect 2646 12614 2674 12642
rect 2758 13145 2786 13146
rect 2758 13119 2759 13145
rect 2759 13119 2785 13145
rect 2785 13119 2786 13145
rect 2758 13118 2786 13119
rect 4998 14350 5026 14378
rect 5838 14713 5866 14714
rect 5838 14687 5839 14713
rect 5839 14687 5865 14713
rect 5865 14687 5866 14713
rect 5838 14686 5866 14687
rect 6006 14742 6034 14770
rect 5278 14321 5306 14322
rect 5278 14295 5279 14321
rect 5279 14295 5305 14321
rect 5305 14295 5306 14321
rect 5278 14294 5306 14295
rect 4582 14125 4610 14126
rect 4582 14099 4600 14125
rect 4600 14099 4610 14125
rect 4582 14098 4610 14099
rect 4634 14125 4662 14126
rect 4634 14099 4636 14125
rect 4636 14099 4662 14125
rect 4634 14098 4662 14099
rect 4686 14125 4714 14126
rect 4738 14125 4766 14126
rect 4686 14099 4698 14125
rect 4698 14099 4714 14125
rect 4738 14099 4760 14125
rect 4760 14099 4766 14125
rect 4686 14098 4714 14099
rect 4738 14098 4766 14099
rect 4790 14098 4818 14126
rect 4842 14125 4870 14126
rect 4894 14125 4922 14126
rect 4842 14099 4848 14125
rect 4848 14099 4870 14125
rect 4894 14099 4910 14125
rect 4910 14099 4922 14125
rect 4842 14098 4870 14099
rect 4894 14098 4922 14099
rect 4946 14125 4974 14126
rect 4946 14099 4972 14125
rect 4972 14099 4974 14125
rect 4946 14098 4974 14099
rect 4998 14125 5026 14126
rect 4998 14099 5008 14125
rect 5008 14099 5026 14125
rect 4998 14098 5026 14099
rect 3822 13398 3850 13426
rect 4102 13510 4130 13538
rect 3318 13145 3346 13146
rect 3318 13119 3319 13145
rect 3319 13119 3345 13145
rect 3345 13119 3346 13145
rect 3318 13118 3346 13119
rect 2758 12670 2786 12698
rect 5838 13929 5866 13930
rect 5838 13903 5839 13929
rect 5839 13903 5865 13929
rect 5865 13903 5866 13929
rect 5838 13902 5866 13903
rect 5278 13537 5306 13538
rect 5278 13511 5279 13537
rect 5279 13511 5305 13537
rect 5305 13511 5306 13537
rect 5278 13510 5306 13511
rect 5838 13510 5866 13538
rect 4582 13341 4610 13342
rect 4582 13315 4600 13341
rect 4600 13315 4610 13341
rect 4582 13314 4610 13315
rect 4634 13341 4662 13342
rect 4634 13315 4636 13341
rect 4636 13315 4662 13341
rect 4634 13314 4662 13315
rect 4686 13341 4714 13342
rect 4738 13341 4766 13342
rect 4686 13315 4698 13341
rect 4698 13315 4714 13341
rect 4738 13315 4760 13341
rect 4760 13315 4766 13341
rect 4686 13314 4714 13315
rect 4738 13314 4766 13315
rect 4790 13314 4818 13342
rect 4842 13341 4870 13342
rect 4894 13341 4922 13342
rect 4842 13315 4848 13341
rect 4848 13315 4870 13341
rect 4894 13315 4910 13341
rect 4910 13315 4922 13341
rect 4842 13314 4870 13315
rect 4894 13314 4922 13315
rect 4946 13341 4974 13342
rect 4946 13315 4972 13341
rect 4972 13315 4974 13341
rect 4946 13314 4974 13315
rect 4998 13341 5026 13342
rect 4998 13315 5008 13341
rect 5008 13315 5026 13341
rect 4998 13314 5026 13315
rect 3038 12334 3066 12362
rect 2082 12165 2110 12166
rect 2082 12139 2100 12165
rect 2100 12139 2110 12165
rect 2082 12138 2110 12139
rect 2134 12165 2162 12166
rect 2134 12139 2136 12165
rect 2136 12139 2162 12165
rect 2134 12138 2162 12139
rect 2186 12165 2214 12166
rect 2238 12165 2266 12166
rect 2186 12139 2198 12165
rect 2198 12139 2214 12165
rect 2238 12139 2260 12165
rect 2260 12139 2266 12165
rect 2186 12138 2214 12139
rect 2238 12138 2266 12139
rect 2290 12138 2318 12166
rect 2342 12165 2370 12166
rect 2394 12165 2422 12166
rect 2342 12139 2348 12165
rect 2348 12139 2370 12165
rect 2394 12139 2410 12165
rect 2410 12139 2422 12165
rect 2342 12138 2370 12139
rect 2394 12138 2422 12139
rect 2446 12165 2474 12166
rect 2446 12139 2472 12165
rect 2472 12139 2474 12165
rect 2446 12138 2474 12139
rect 2498 12165 2526 12166
rect 2498 12139 2508 12165
rect 2508 12139 2526 12165
rect 2498 12138 2526 12139
rect 1862 10766 1890 10794
rect 1638 9198 1666 9226
rect 1414 8414 1442 8442
rect 1918 9310 1946 9338
rect 1862 9225 1890 9226
rect 1862 9199 1863 9225
rect 1863 9199 1889 9225
rect 1889 9199 1890 9225
rect 1862 9198 1890 9199
rect 1862 8441 1890 8442
rect 1862 8415 1863 8441
rect 1863 8415 1889 8441
rect 1889 8415 1890 8441
rect 1862 8414 1890 8415
rect 1918 6454 1946 6482
rect 1806 4129 1834 4130
rect 1806 4103 1807 4129
rect 1807 4103 1833 4129
rect 1833 4103 1834 4129
rect 1806 4102 1834 4103
rect 1918 4102 1946 4130
rect 1918 3598 1946 3626
rect 1190 2646 1218 2674
rect 1638 2198 1666 2226
rect 3598 12361 3626 12362
rect 3598 12335 3599 12361
rect 3599 12335 3625 12361
rect 3625 12335 3626 12361
rect 3598 12334 3626 12335
rect 4102 12334 4130 12362
rect 4326 12558 4354 12586
rect 4102 11969 4130 11970
rect 4102 11943 4103 11969
rect 4103 11943 4129 11969
rect 4129 11943 4130 11969
rect 4102 11942 4130 11943
rect 4582 12557 4610 12558
rect 4582 12531 4600 12557
rect 4600 12531 4610 12557
rect 4582 12530 4610 12531
rect 4634 12557 4662 12558
rect 4634 12531 4636 12557
rect 4636 12531 4662 12557
rect 4634 12530 4662 12531
rect 4686 12557 4714 12558
rect 4738 12557 4766 12558
rect 4686 12531 4698 12557
rect 4698 12531 4714 12557
rect 4738 12531 4760 12557
rect 4760 12531 4766 12557
rect 4686 12530 4714 12531
rect 4738 12530 4766 12531
rect 4790 12530 4818 12558
rect 4842 12557 4870 12558
rect 4894 12557 4922 12558
rect 4842 12531 4848 12557
rect 4848 12531 4870 12557
rect 4894 12531 4910 12557
rect 4910 12531 4922 12557
rect 4842 12530 4870 12531
rect 4894 12530 4922 12531
rect 4946 12557 4974 12558
rect 4946 12531 4972 12557
rect 4972 12531 4974 12557
rect 4946 12530 4974 12531
rect 4998 12557 5026 12558
rect 4998 12531 5008 12557
rect 5008 12531 5026 12557
rect 4998 12530 5026 12531
rect 5278 11969 5306 11970
rect 5278 11943 5279 11969
rect 5279 11943 5305 11969
rect 5305 11943 5306 11969
rect 5278 11942 5306 11943
rect 4582 11773 4610 11774
rect 4582 11747 4600 11773
rect 4600 11747 4610 11773
rect 4582 11746 4610 11747
rect 4634 11773 4662 11774
rect 4634 11747 4636 11773
rect 4636 11747 4662 11773
rect 4634 11746 4662 11747
rect 4686 11773 4714 11774
rect 4738 11773 4766 11774
rect 4686 11747 4698 11773
rect 4698 11747 4714 11773
rect 4738 11747 4760 11773
rect 4760 11747 4766 11773
rect 4686 11746 4714 11747
rect 4738 11746 4766 11747
rect 4790 11746 4818 11774
rect 4842 11773 4870 11774
rect 4894 11773 4922 11774
rect 4842 11747 4848 11773
rect 4848 11747 4870 11773
rect 4894 11747 4910 11773
rect 4910 11747 4922 11773
rect 4842 11746 4870 11747
rect 4894 11746 4922 11747
rect 4946 11773 4974 11774
rect 4946 11747 4972 11773
rect 4972 11747 4974 11773
rect 4946 11746 4974 11747
rect 4998 11773 5026 11774
rect 4998 11747 5008 11773
rect 5008 11747 5026 11773
rect 4998 11746 5026 11747
rect 2082 11381 2110 11382
rect 2082 11355 2100 11381
rect 2100 11355 2110 11381
rect 2082 11354 2110 11355
rect 2134 11381 2162 11382
rect 2134 11355 2136 11381
rect 2136 11355 2162 11381
rect 2134 11354 2162 11355
rect 2186 11381 2214 11382
rect 2238 11381 2266 11382
rect 2186 11355 2198 11381
rect 2198 11355 2214 11381
rect 2238 11355 2260 11381
rect 2260 11355 2266 11381
rect 2186 11354 2214 11355
rect 2238 11354 2266 11355
rect 2290 11354 2318 11382
rect 2342 11381 2370 11382
rect 2394 11381 2422 11382
rect 2342 11355 2348 11381
rect 2348 11355 2370 11381
rect 2394 11355 2410 11381
rect 2410 11355 2422 11381
rect 2342 11354 2370 11355
rect 2394 11354 2422 11355
rect 2446 11381 2474 11382
rect 2446 11355 2472 11381
rect 2472 11355 2474 11381
rect 2446 11354 2474 11355
rect 2498 11381 2526 11382
rect 2498 11355 2508 11381
rect 2508 11355 2526 11381
rect 2498 11354 2526 11355
rect 2478 10878 2506 10906
rect 2590 10878 2618 10906
rect 2086 10793 2114 10794
rect 2086 10767 2087 10793
rect 2087 10767 2113 10793
rect 2113 10767 2114 10793
rect 2086 10766 2114 10767
rect 2082 10597 2110 10598
rect 2082 10571 2100 10597
rect 2100 10571 2110 10597
rect 2082 10570 2110 10571
rect 2134 10597 2162 10598
rect 2134 10571 2136 10597
rect 2136 10571 2162 10597
rect 2134 10570 2162 10571
rect 2186 10597 2214 10598
rect 2238 10597 2266 10598
rect 2186 10571 2198 10597
rect 2198 10571 2214 10597
rect 2238 10571 2260 10597
rect 2260 10571 2266 10597
rect 2186 10570 2214 10571
rect 2238 10570 2266 10571
rect 2290 10570 2318 10598
rect 2342 10597 2370 10598
rect 2394 10597 2422 10598
rect 2342 10571 2348 10597
rect 2348 10571 2370 10597
rect 2394 10571 2410 10597
rect 2410 10571 2422 10597
rect 2342 10570 2370 10571
rect 2394 10570 2422 10571
rect 2446 10597 2474 10598
rect 2446 10571 2472 10597
rect 2472 10571 2474 10597
rect 2446 10570 2474 10571
rect 2498 10597 2526 10598
rect 2498 10571 2508 10597
rect 2508 10571 2526 10597
rect 2498 10570 2526 10571
rect 3038 10878 3066 10906
rect 2082 9813 2110 9814
rect 2082 9787 2100 9813
rect 2100 9787 2110 9813
rect 2082 9786 2110 9787
rect 2134 9813 2162 9814
rect 2134 9787 2136 9813
rect 2136 9787 2162 9813
rect 2134 9786 2162 9787
rect 2186 9813 2214 9814
rect 2238 9813 2266 9814
rect 2186 9787 2198 9813
rect 2198 9787 2214 9813
rect 2238 9787 2260 9813
rect 2260 9787 2266 9813
rect 2186 9786 2214 9787
rect 2238 9786 2266 9787
rect 2290 9786 2318 9814
rect 2342 9813 2370 9814
rect 2394 9813 2422 9814
rect 2342 9787 2348 9813
rect 2348 9787 2370 9813
rect 2394 9787 2410 9813
rect 2410 9787 2422 9813
rect 2342 9786 2370 9787
rect 2394 9786 2422 9787
rect 2446 9813 2474 9814
rect 2446 9787 2472 9813
rect 2472 9787 2474 9813
rect 2446 9786 2474 9787
rect 2498 9813 2526 9814
rect 2498 9787 2508 9813
rect 2508 9787 2526 9813
rect 2498 9786 2526 9787
rect 4582 10989 4610 10990
rect 4582 10963 4600 10989
rect 4600 10963 4610 10989
rect 4582 10962 4610 10963
rect 4634 10989 4662 10990
rect 4634 10963 4636 10989
rect 4636 10963 4662 10989
rect 4634 10962 4662 10963
rect 4686 10989 4714 10990
rect 4738 10989 4766 10990
rect 4686 10963 4698 10989
rect 4698 10963 4714 10989
rect 4738 10963 4760 10989
rect 4760 10963 4766 10989
rect 4686 10962 4714 10963
rect 4738 10962 4766 10963
rect 4790 10962 4818 10990
rect 4842 10989 4870 10990
rect 4894 10989 4922 10990
rect 4842 10963 4848 10989
rect 4848 10963 4870 10989
rect 4894 10963 4910 10989
rect 4910 10963 4922 10989
rect 4842 10962 4870 10963
rect 4894 10962 4922 10963
rect 4946 10989 4974 10990
rect 4946 10963 4972 10989
rect 4972 10963 4974 10989
rect 4946 10962 4974 10963
rect 4998 10989 5026 10990
rect 4998 10963 5008 10989
rect 5008 10963 5026 10989
rect 4998 10962 5026 10963
rect 5278 10766 5306 10794
rect 3822 10401 3850 10402
rect 3822 10375 3823 10401
rect 3823 10375 3849 10401
rect 3849 10375 3850 10401
rect 3822 10374 3850 10375
rect 5838 10934 5866 10962
rect 5838 10793 5866 10794
rect 5838 10767 5839 10793
rect 5839 10767 5865 10793
rect 5865 10767 5866 10793
rect 5838 10766 5866 10767
rect 5278 10401 5306 10402
rect 5278 10375 5279 10401
rect 5279 10375 5305 10401
rect 5305 10375 5306 10401
rect 5278 10374 5306 10375
rect 4582 10205 4610 10206
rect 4582 10179 4600 10205
rect 4600 10179 4610 10205
rect 4582 10178 4610 10179
rect 4634 10205 4662 10206
rect 4634 10179 4636 10205
rect 4636 10179 4662 10205
rect 4634 10178 4662 10179
rect 4686 10205 4714 10206
rect 4738 10205 4766 10206
rect 4686 10179 4698 10205
rect 4698 10179 4714 10205
rect 4738 10179 4760 10205
rect 4760 10179 4766 10205
rect 4686 10178 4714 10179
rect 4738 10178 4766 10179
rect 4790 10178 4818 10206
rect 4842 10205 4870 10206
rect 4894 10205 4922 10206
rect 4842 10179 4848 10205
rect 4848 10179 4870 10205
rect 4894 10179 4910 10205
rect 4910 10179 4922 10205
rect 4842 10178 4870 10179
rect 4894 10178 4922 10179
rect 4946 10205 4974 10206
rect 4946 10179 4972 10205
rect 4972 10179 4974 10205
rect 4946 10178 4974 10179
rect 4998 10205 5026 10206
rect 4998 10179 5008 10205
rect 5008 10179 5026 10205
rect 4998 10178 5026 10179
rect 3822 9617 3850 9618
rect 3822 9591 3823 9617
rect 3823 9591 3849 9617
rect 3849 9591 3850 9617
rect 3822 9590 3850 9591
rect 2478 9310 2506 9338
rect 2030 9254 2058 9282
rect 3374 9281 3402 9282
rect 3374 9255 3375 9281
rect 3375 9255 3401 9281
rect 3401 9255 3402 9281
rect 3374 9254 3402 9255
rect 2082 9029 2110 9030
rect 2082 9003 2100 9029
rect 2100 9003 2110 9029
rect 2082 9002 2110 9003
rect 2134 9029 2162 9030
rect 2134 9003 2136 9029
rect 2136 9003 2162 9029
rect 2134 9002 2162 9003
rect 2186 9029 2214 9030
rect 2238 9029 2266 9030
rect 2186 9003 2198 9029
rect 2198 9003 2214 9029
rect 2238 9003 2260 9029
rect 2260 9003 2266 9029
rect 2186 9002 2214 9003
rect 2238 9002 2266 9003
rect 2290 9002 2318 9030
rect 2342 9029 2370 9030
rect 2394 9029 2422 9030
rect 2342 9003 2348 9029
rect 2348 9003 2370 9029
rect 2394 9003 2410 9029
rect 2410 9003 2422 9029
rect 2342 9002 2370 9003
rect 2394 9002 2422 9003
rect 2446 9029 2474 9030
rect 2446 9003 2472 9029
rect 2472 9003 2474 9029
rect 2446 9002 2474 9003
rect 2498 9029 2526 9030
rect 2498 9003 2508 9029
rect 2508 9003 2526 9029
rect 2498 9002 2526 9003
rect 2082 8245 2110 8246
rect 2082 8219 2100 8245
rect 2100 8219 2110 8245
rect 2082 8218 2110 8219
rect 2134 8245 2162 8246
rect 2134 8219 2136 8245
rect 2136 8219 2162 8245
rect 2134 8218 2162 8219
rect 2186 8245 2214 8246
rect 2238 8245 2266 8246
rect 2186 8219 2198 8245
rect 2198 8219 2214 8245
rect 2238 8219 2260 8245
rect 2260 8219 2266 8245
rect 2186 8218 2214 8219
rect 2238 8218 2266 8219
rect 2290 8218 2318 8246
rect 2342 8245 2370 8246
rect 2394 8245 2422 8246
rect 2342 8219 2348 8245
rect 2348 8219 2370 8245
rect 2394 8219 2410 8245
rect 2410 8219 2422 8245
rect 2342 8218 2370 8219
rect 2394 8218 2422 8219
rect 2446 8245 2474 8246
rect 2446 8219 2472 8245
rect 2472 8219 2474 8245
rect 2446 8218 2474 8219
rect 2498 8245 2526 8246
rect 2498 8219 2508 8245
rect 2508 8219 2526 8245
rect 2498 8218 2526 8219
rect 2082 7461 2110 7462
rect 2082 7435 2100 7461
rect 2100 7435 2110 7461
rect 2082 7434 2110 7435
rect 2134 7461 2162 7462
rect 2134 7435 2136 7461
rect 2136 7435 2162 7461
rect 2134 7434 2162 7435
rect 2186 7461 2214 7462
rect 2238 7461 2266 7462
rect 2186 7435 2198 7461
rect 2198 7435 2214 7461
rect 2238 7435 2260 7461
rect 2260 7435 2266 7461
rect 2186 7434 2214 7435
rect 2238 7434 2266 7435
rect 2290 7434 2318 7462
rect 2342 7461 2370 7462
rect 2394 7461 2422 7462
rect 2342 7435 2348 7461
rect 2348 7435 2370 7461
rect 2394 7435 2410 7461
rect 2410 7435 2422 7461
rect 2342 7434 2370 7435
rect 2394 7434 2422 7435
rect 2446 7461 2474 7462
rect 2446 7435 2472 7461
rect 2472 7435 2474 7461
rect 2446 7434 2474 7435
rect 2498 7461 2526 7462
rect 2498 7435 2508 7461
rect 2508 7435 2526 7461
rect 2498 7434 2526 7435
rect 2478 7265 2506 7266
rect 2478 7239 2479 7265
rect 2479 7239 2505 7265
rect 2505 7239 2506 7265
rect 2478 7238 2506 7239
rect 2590 7238 2618 7266
rect 3822 9254 3850 9282
rect 3038 7238 3066 7266
rect 3038 6873 3066 6874
rect 3038 6847 3039 6873
rect 3039 6847 3065 6873
rect 3065 6847 3066 6873
rect 3038 6846 3066 6847
rect 3598 6873 3626 6874
rect 3598 6847 3599 6873
rect 3599 6847 3625 6873
rect 3625 6847 3626 6873
rect 3598 6846 3626 6847
rect 2082 6677 2110 6678
rect 2082 6651 2100 6677
rect 2100 6651 2110 6677
rect 2082 6650 2110 6651
rect 2134 6677 2162 6678
rect 2134 6651 2136 6677
rect 2136 6651 2162 6677
rect 2134 6650 2162 6651
rect 2186 6677 2214 6678
rect 2238 6677 2266 6678
rect 2186 6651 2198 6677
rect 2198 6651 2214 6677
rect 2238 6651 2260 6677
rect 2260 6651 2266 6677
rect 2186 6650 2214 6651
rect 2238 6650 2266 6651
rect 2290 6650 2318 6678
rect 2342 6677 2370 6678
rect 2394 6677 2422 6678
rect 2342 6651 2348 6677
rect 2348 6651 2370 6677
rect 2394 6651 2410 6677
rect 2410 6651 2422 6677
rect 2342 6650 2370 6651
rect 2394 6650 2422 6651
rect 2446 6677 2474 6678
rect 2446 6651 2472 6677
rect 2472 6651 2474 6677
rect 2446 6650 2474 6651
rect 2498 6677 2526 6678
rect 2498 6651 2508 6677
rect 2508 6651 2526 6677
rect 2498 6650 2526 6651
rect 2198 6481 2226 6482
rect 2198 6455 2199 6481
rect 2199 6455 2225 6481
rect 2225 6455 2226 6481
rect 2198 6454 2226 6455
rect 2758 6454 2786 6482
rect 2082 5893 2110 5894
rect 2082 5867 2100 5893
rect 2100 5867 2110 5893
rect 2082 5866 2110 5867
rect 2134 5893 2162 5894
rect 2134 5867 2136 5893
rect 2136 5867 2162 5893
rect 2134 5866 2162 5867
rect 2186 5893 2214 5894
rect 2238 5893 2266 5894
rect 2186 5867 2198 5893
rect 2198 5867 2214 5893
rect 2238 5867 2260 5893
rect 2260 5867 2266 5893
rect 2186 5866 2214 5867
rect 2238 5866 2266 5867
rect 2290 5866 2318 5894
rect 2342 5893 2370 5894
rect 2394 5893 2422 5894
rect 2342 5867 2348 5893
rect 2348 5867 2370 5893
rect 2394 5867 2410 5893
rect 2410 5867 2422 5893
rect 2342 5866 2370 5867
rect 2394 5866 2422 5867
rect 2446 5893 2474 5894
rect 2446 5867 2472 5893
rect 2472 5867 2474 5893
rect 2446 5866 2474 5867
rect 2498 5893 2526 5894
rect 2498 5867 2508 5893
rect 2508 5867 2526 5893
rect 2498 5866 2526 5867
rect 2082 5109 2110 5110
rect 2082 5083 2100 5109
rect 2100 5083 2110 5109
rect 2082 5082 2110 5083
rect 2134 5109 2162 5110
rect 2134 5083 2136 5109
rect 2136 5083 2162 5109
rect 2134 5082 2162 5083
rect 2186 5109 2214 5110
rect 2238 5109 2266 5110
rect 2186 5083 2198 5109
rect 2198 5083 2214 5109
rect 2238 5083 2260 5109
rect 2260 5083 2266 5109
rect 2186 5082 2214 5083
rect 2238 5082 2266 5083
rect 2290 5082 2318 5110
rect 2342 5109 2370 5110
rect 2394 5109 2422 5110
rect 2342 5083 2348 5109
rect 2348 5083 2370 5109
rect 2394 5083 2410 5109
rect 2410 5083 2422 5109
rect 2342 5082 2370 5083
rect 2394 5082 2422 5083
rect 2446 5109 2474 5110
rect 2446 5083 2472 5109
rect 2472 5083 2474 5109
rect 2446 5082 2474 5083
rect 2498 5109 2526 5110
rect 2498 5083 2508 5109
rect 2508 5083 2526 5109
rect 2498 5082 2526 5083
rect 2082 4325 2110 4326
rect 2082 4299 2100 4325
rect 2100 4299 2110 4325
rect 2082 4298 2110 4299
rect 2134 4325 2162 4326
rect 2134 4299 2136 4325
rect 2136 4299 2162 4325
rect 2134 4298 2162 4299
rect 2186 4325 2214 4326
rect 2238 4325 2266 4326
rect 2186 4299 2198 4325
rect 2198 4299 2214 4325
rect 2238 4299 2260 4325
rect 2260 4299 2266 4325
rect 2186 4298 2214 4299
rect 2238 4298 2266 4299
rect 2290 4298 2318 4326
rect 2342 4325 2370 4326
rect 2394 4325 2422 4326
rect 2342 4299 2348 4325
rect 2348 4299 2370 4325
rect 2394 4299 2410 4325
rect 2410 4299 2422 4325
rect 2342 4298 2370 4299
rect 2394 4298 2422 4299
rect 2446 4325 2474 4326
rect 2446 4299 2472 4325
rect 2472 4299 2474 4325
rect 2446 4298 2474 4299
rect 2498 4325 2526 4326
rect 2498 4299 2508 4325
rect 2508 4299 2526 4325
rect 2498 4298 2526 4299
rect 4046 9926 4074 9954
rect 3990 6510 4018 6538
rect 3598 5305 3626 5306
rect 3598 5279 3599 5305
rect 3599 5279 3625 5305
rect 3625 5279 3626 5305
rect 3598 5278 3626 5279
rect 2758 4521 2786 4522
rect 2758 4495 2759 4521
rect 2759 4495 2785 4521
rect 2785 4495 2786 4521
rect 2758 4494 2786 4495
rect 2982 4494 3010 4522
rect 2030 4129 2058 4130
rect 2030 4103 2031 4129
rect 2031 4103 2057 4129
rect 2057 4103 2058 4129
rect 2030 4102 2058 4103
rect 2030 3598 2058 3626
rect 3318 4521 3346 4522
rect 3318 4495 3319 4521
rect 3319 4495 3345 4521
rect 3345 4495 3346 4521
rect 3318 4494 3346 4495
rect 3598 4494 3626 4522
rect 3262 3766 3290 3794
rect 2478 3598 2506 3626
rect 2082 3541 2110 3542
rect 2082 3515 2100 3541
rect 2100 3515 2110 3541
rect 2082 3514 2110 3515
rect 2134 3541 2162 3542
rect 2134 3515 2136 3541
rect 2136 3515 2162 3541
rect 2134 3514 2162 3515
rect 2186 3541 2214 3542
rect 2238 3541 2266 3542
rect 2186 3515 2198 3541
rect 2198 3515 2214 3541
rect 2238 3515 2260 3541
rect 2260 3515 2266 3541
rect 2186 3514 2214 3515
rect 2238 3514 2266 3515
rect 2290 3514 2318 3542
rect 2342 3541 2370 3542
rect 2394 3541 2422 3542
rect 2342 3515 2348 3541
rect 2348 3515 2370 3541
rect 2394 3515 2410 3541
rect 2410 3515 2422 3541
rect 2342 3514 2370 3515
rect 2394 3514 2422 3515
rect 2446 3541 2474 3542
rect 2446 3515 2472 3541
rect 2472 3515 2474 3541
rect 2446 3514 2474 3515
rect 2498 3541 2526 3542
rect 2498 3515 2508 3541
rect 2508 3515 2526 3541
rect 2498 3514 2526 3515
rect 2082 2757 2110 2758
rect 2082 2731 2100 2757
rect 2100 2731 2110 2757
rect 2082 2730 2110 2731
rect 2134 2757 2162 2758
rect 2134 2731 2136 2757
rect 2136 2731 2162 2757
rect 2134 2730 2162 2731
rect 2186 2757 2214 2758
rect 2238 2757 2266 2758
rect 2186 2731 2198 2757
rect 2198 2731 2214 2757
rect 2238 2731 2260 2757
rect 2260 2731 2266 2757
rect 2186 2730 2214 2731
rect 2238 2730 2266 2731
rect 2290 2730 2318 2758
rect 2342 2757 2370 2758
rect 2394 2757 2422 2758
rect 2342 2731 2348 2757
rect 2348 2731 2370 2757
rect 2394 2731 2410 2757
rect 2410 2731 2422 2757
rect 2342 2730 2370 2731
rect 2394 2730 2422 2731
rect 2446 2757 2474 2758
rect 2446 2731 2472 2757
rect 2472 2731 2474 2757
rect 2446 2730 2474 2731
rect 2498 2757 2526 2758
rect 2498 2731 2508 2757
rect 2508 2731 2526 2757
rect 2498 2730 2526 2731
rect 2478 2590 2506 2618
rect 1974 2534 2002 2562
rect 2366 2534 2394 2562
rect 3038 2590 3066 2618
rect 2590 2254 2618 2282
rect 3038 2169 3066 2170
rect 3038 2143 3039 2169
rect 3039 2143 3065 2169
rect 3065 2143 3066 2169
rect 3038 2142 3066 2143
rect 2082 1973 2110 1974
rect 2082 1947 2100 1973
rect 2100 1947 2110 1973
rect 2082 1946 2110 1947
rect 2134 1973 2162 1974
rect 2134 1947 2136 1973
rect 2136 1947 2162 1973
rect 2134 1946 2162 1947
rect 2186 1973 2214 1974
rect 2238 1973 2266 1974
rect 2186 1947 2198 1973
rect 2198 1947 2214 1973
rect 2238 1947 2260 1973
rect 2260 1947 2266 1973
rect 2186 1946 2214 1947
rect 2238 1946 2266 1947
rect 2290 1946 2318 1974
rect 2342 1973 2370 1974
rect 2394 1973 2422 1974
rect 2342 1947 2348 1973
rect 2348 1947 2370 1973
rect 2394 1947 2410 1973
rect 2410 1947 2422 1973
rect 2342 1946 2370 1947
rect 2394 1946 2422 1947
rect 2446 1973 2474 1974
rect 2446 1947 2472 1973
rect 2472 1947 2474 1973
rect 2446 1946 2474 1947
rect 2498 1973 2526 1974
rect 2498 1947 2508 1973
rect 2508 1947 2526 1973
rect 2498 1946 2526 1947
rect 2086 1862 2114 1890
rect 5446 10710 5474 10738
rect 4582 9421 4610 9422
rect 4582 9395 4600 9421
rect 4600 9395 4610 9421
rect 4582 9394 4610 9395
rect 4634 9421 4662 9422
rect 4634 9395 4636 9421
rect 4636 9395 4662 9421
rect 4634 9394 4662 9395
rect 4686 9421 4714 9422
rect 4738 9421 4766 9422
rect 4686 9395 4698 9421
rect 4698 9395 4714 9421
rect 4738 9395 4760 9421
rect 4760 9395 4766 9421
rect 4686 9394 4714 9395
rect 4738 9394 4766 9395
rect 4790 9394 4818 9422
rect 4842 9421 4870 9422
rect 4894 9421 4922 9422
rect 4842 9395 4848 9421
rect 4848 9395 4870 9421
rect 4894 9395 4910 9421
rect 4910 9395 4922 9421
rect 4842 9394 4870 9395
rect 4894 9394 4922 9395
rect 4946 9421 4974 9422
rect 4946 9395 4972 9421
rect 4972 9395 4974 9421
rect 4946 9394 4974 9395
rect 4998 9421 5026 9422
rect 4998 9395 5008 9421
rect 5008 9395 5026 9421
rect 4998 9394 5026 9395
rect 4494 9225 4522 9226
rect 4494 9199 4495 9225
rect 4495 9199 4521 9225
rect 4521 9199 4522 9225
rect 4494 9198 4522 9199
rect 5110 9198 5138 9226
rect 4998 8833 5026 8834
rect 4998 8807 4999 8833
rect 4999 8807 5025 8833
rect 5025 8807 5026 8833
rect 4998 8806 5026 8807
rect 5110 8806 5138 8834
rect 4582 8637 4610 8638
rect 4582 8611 4600 8637
rect 4600 8611 4610 8637
rect 4582 8610 4610 8611
rect 4634 8637 4662 8638
rect 4634 8611 4636 8637
rect 4636 8611 4662 8637
rect 4634 8610 4662 8611
rect 4686 8637 4714 8638
rect 4738 8637 4766 8638
rect 4686 8611 4698 8637
rect 4698 8611 4714 8637
rect 4738 8611 4760 8637
rect 4760 8611 4766 8637
rect 4686 8610 4714 8611
rect 4738 8610 4766 8611
rect 4790 8610 4818 8638
rect 4842 8637 4870 8638
rect 4894 8637 4922 8638
rect 4842 8611 4848 8637
rect 4848 8611 4870 8637
rect 4894 8611 4910 8637
rect 4910 8611 4922 8637
rect 4842 8610 4870 8611
rect 4894 8610 4922 8611
rect 4946 8637 4974 8638
rect 4946 8611 4972 8637
rect 4972 8611 4974 8637
rect 4946 8610 4974 8611
rect 4998 8637 5026 8638
rect 4998 8611 5008 8637
rect 5008 8611 5026 8637
rect 4998 8610 5026 8611
rect 4494 8441 4522 8442
rect 4494 8415 4495 8441
rect 4495 8415 4521 8441
rect 4521 8415 4522 8441
rect 4494 8414 4522 8415
rect 4582 7853 4610 7854
rect 4582 7827 4600 7853
rect 4600 7827 4610 7853
rect 4582 7826 4610 7827
rect 4634 7853 4662 7854
rect 4634 7827 4636 7853
rect 4636 7827 4662 7853
rect 4634 7826 4662 7827
rect 4686 7853 4714 7854
rect 4738 7853 4766 7854
rect 4686 7827 4698 7853
rect 4698 7827 4714 7853
rect 4738 7827 4760 7853
rect 4760 7827 4766 7853
rect 4686 7826 4714 7827
rect 4738 7826 4766 7827
rect 4790 7826 4818 7854
rect 4842 7853 4870 7854
rect 4894 7853 4922 7854
rect 4842 7827 4848 7853
rect 4848 7827 4870 7853
rect 4894 7827 4910 7853
rect 4910 7827 4922 7853
rect 4842 7826 4870 7827
rect 4894 7826 4922 7827
rect 4946 7853 4974 7854
rect 4946 7827 4972 7853
rect 4972 7827 4974 7853
rect 4946 7826 4974 7827
rect 4998 7853 5026 7854
rect 4998 7827 5008 7853
rect 5008 7827 5026 7853
rect 4998 7826 5026 7827
rect 4494 7182 4522 7210
rect 4998 7209 5026 7210
rect 4998 7183 4999 7209
rect 4999 7183 5025 7209
rect 5025 7183 5026 7209
rect 4998 7182 5026 7183
rect 4582 7069 4610 7070
rect 4582 7043 4600 7069
rect 4600 7043 4610 7069
rect 4582 7042 4610 7043
rect 4634 7069 4662 7070
rect 4634 7043 4636 7069
rect 4636 7043 4662 7069
rect 4634 7042 4662 7043
rect 4686 7069 4714 7070
rect 4738 7069 4766 7070
rect 4686 7043 4698 7069
rect 4698 7043 4714 7069
rect 4738 7043 4760 7069
rect 4760 7043 4766 7069
rect 4686 7042 4714 7043
rect 4738 7042 4766 7043
rect 4790 7042 4818 7070
rect 4842 7069 4870 7070
rect 4894 7069 4922 7070
rect 4842 7043 4848 7069
rect 4848 7043 4870 7069
rect 4894 7043 4910 7069
rect 4910 7043 4922 7069
rect 4842 7042 4870 7043
rect 4894 7042 4922 7043
rect 4946 7069 4974 7070
rect 4946 7043 4972 7069
rect 4972 7043 4974 7069
rect 4946 7042 4974 7043
rect 4998 7069 5026 7070
rect 4998 7043 5008 7069
rect 5008 7043 5026 7069
rect 4998 7042 5026 7043
rect 4102 6846 4130 6874
rect 4102 6481 4130 6482
rect 4102 6455 4103 6481
rect 4103 6455 4129 6481
rect 4129 6455 4130 6481
rect 4102 6454 4130 6455
rect 4270 6510 4298 6538
rect 4582 6285 4610 6286
rect 4582 6259 4600 6285
rect 4600 6259 4610 6285
rect 4582 6258 4610 6259
rect 4634 6285 4662 6286
rect 4634 6259 4636 6285
rect 4636 6259 4662 6285
rect 4634 6258 4662 6259
rect 4686 6285 4714 6286
rect 4738 6285 4766 6286
rect 4686 6259 4698 6285
rect 4698 6259 4714 6285
rect 4738 6259 4760 6285
rect 4760 6259 4766 6285
rect 4686 6258 4714 6259
rect 4738 6258 4766 6259
rect 4790 6258 4818 6286
rect 4842 6285 4870 6286
rect 4894 6285 4922 6286
rect 4842 6259 4848 6285
rect 4848 6259 4870 6285
rect 4894 6259 4910 6285
rect 4910 6259 4922 6285
rect 4842 6258 4870 6259
rect 4894 6258 4922 6259
rect 4946 6285 4974 6286
rect 4946 6259 4972 6285
rect 4972 6259 4974 6285
rect 4946 6258 4974 6259
rect 4998 6285 5026 6286
rect 4998 6259 5008 6285
rect 5008 6259 5026 6285
rect 4998 6258 5026 6259
rect 4102 5278 4130 5306
rect 4102 5054 4130 5082
rect 4582 5501 4610 5502
rect 4582 5475 4600 5501
rect 4600 5475 4610 5501
rect 4582 5474 4610 5475
rect 4634 5501 4662 5502
rect 4634 5475 4636 5501
rect 4636 5475 4662 5501
rect 4634 5474 4662 5475
rect 4686 5501 4714 5502
rect 4738 5501 4766 5502
rect 4686 5475 4698 5501
rect 4698 5475 4714 5501
rect 4738 5475 4760 5501
rect 4760 5475 4766 5501
rect 4686 5474 4714 5475
rect 4738 5474 4766 5475
rect 4790 5474 4818 5502
rect 4842 5501 4870 5502
rect 4894 5501 4922 5502
rect 4842 5475 4848 5501
rect 4848 5475 4870 5501
rect 4894 5475 4910 5501
rect 4910 5475 4922 5501
rect 4842 5474 4870 5475
rect 4894 5474 4922 5475
rect 4946 5501 4974 5502
rect 4946 5475 4972 5501
rect 4972 5475 4974 5501
rect 4946 5474 4974 5475
rect 4998 5501 5026 5502
rect 4998 5475 5008 5501
rect 5008 5475 5026 5501
rect 4998 5474 5026 5475
rect 4582 4717 4610 4718
rect 4582 4691 4600 4717
rect 4600 4691 4610 4717
rect 4582 4690 4610 4691
rect 4634 4717 4662 4718
rect 4634 4691 4636 4717
rect 4636 4691 4662 4717
rect 4634 4690 4662 4691
rect 4686 4717 4714 4718
rect 4738 4717 4766 4718
rect 4686 4691 4698 4717
rect 4698 4691 4714 4717
rect 4738 4691 4760 4717
rect 4760 4691 4766 4717
rect 4686 4690 4714 4691
rect 4738 4690 4766 4691
rect 4790 4690 4818 4718
rect 4842 4717 4870 4718
rect 4894 4717 4922 4718
rect 4842 4691 4848 4717
rect 4848 4691 4870 4717
rect 4894 4691 4910 4717
rect 4910 4691 4922 4717
rect 4842 4690 4870 4691
rect 4894 4690 4922 4691
rect 4946 4717 4974 4718
rect 4946 4691 4972 4717
rect 4972 4691 4974 4717
rect 4946 4690 4974 4691
rect 4998 4717 5026 4718
rect 4998 4691 5008 4717
rect 5008 4691 5026 4717
rect 4998 4690 5026 4691
rect 3542 2590 3570 2618
rect 3598 2422 3626 2450
rect 5278 4214 5306 4242
rect 4270 4158 4298 4186
rect 4494 4158 4522 4186
rect 4998 4158 5026 4186
rect 4582 3933 4610 3934
rect 4582 3907 4600 3933
rect 4600 3907 4610 3933
rect 4582 3906 4610 3907
rect 4634 3933 4662 3934
rect 4634 3907 4636 3933
rect 4636 3907 4662 3933
rect 4634 3906 4662 3907
rect 4686 3933 4714 3934
rect 4738 3933 4766 3934
rect 4686 3907 4698 3933
rect 4698 3907 4714 3933
rect 4738 3907 4760 3933
rect 4760 3907 4766 3933
rect 4686 3906 4714 3907
rect 4738 3906 4766 3907
rect 4790 3906 4818 3934
rect 4842 3933 4870 3934
rect 4894 3933 4922 3934
rect 4842 3907 4848 3933
rect 4848 3907 4870 3933
rect 4894 3907 4910 3933
rect 4910 3907 4922 3933
rect 4842 3906 4870 3907
rect 4894 3906 4922 3907
rect 4946 3933 4974 3934
rect 4946 3907 4972 3933
rect 4972 3907 4974 3933
rect 4946 3906 4974 3907
rect 4998 3933 5026 3934
rect 4998 3907 5008 3933
rect 5008 3907 5026 3933
rect 4998 3906 5026 3907
rect 4494 3598 4522 3626
rect 4046 2590 4074 2618
rect 4582 3149 4610 3150
rect 4582 3123 4600 3149
rect 4600 3123 4610 3149
rect 4582 3122 4610 3123
rect 4634 3149 4662 3150
rect 4634 3123 4636 3149
rect 4636 3123 4662 3149
rect 4634 3122 4662 3123
rect 4686 3149 4714 3150
rect 4738 3149 4766 3150
rect 4686 3123 4698 3149
rect 4698 3123 4714 3149
rect 4738 3123 4760 3149
rect 4760 3123 4766 3149
rect 4686 3122 4714 3123
rect 4738 3122 4766 3123
rect 4790 3122 4818 3150
rect 4842 3149 4870 3150
rect 4894 3149 4922 3150
rect 4842 3123 4848 3149
rect 4848 3123 4870 3149
rect 4894 3123 4910 3149
rect 4910 3123 4922 3149
rect 4842 3122 4870 3123
rect 4894 3122 4922 3123
rect 4946 3149 4974 3150
rect 4946 3123 4972 3149
rect 4972 3123 4974 3149
rect 4946 3122 4974 3123
rect 4998 3149 5026 3150
rect 4998 3123 5008 3149
rect 5008 3123 5026 3149
rect 4998 3122 5026 3123
rect 5558 8833 5586 8834
rect 5558 8807 5559 8833
rect 5559 8807 5585 8833
rect 5585 8807 5586 8833
rect 5558 8806 5586 8807
rect 5950 9617 5978 9618
rect 5950 9591 5951 9617
rect 5951 9591 5977 9617
rect 5977 9591 5978 9617
rect 5950 9590 5978 9591
rect 5894 8806 5922 8834
rect 5558 7630 5586 7658
rect 6398 14350 6426 14378
rect 6398 13537 6426 13538
rect 6398 13511 6399 13537
rect 6399 13511 6425 13537
rect 6425 13511 6426 13537
rect 6398 13510 6426 13511
rect 6454 13454 6482 13482
rect 6398 11774 6426 11802
rect 6230 9590 6258 9618
rect 6846 14630 6874 14658
rect 7014 15470 7042 15498
rect 7294 15497 7322 15498
rect 7294 15471 7295 15497
rect 7295 15471 7321 15497
rect 7321 15471 7322 15497
rect 7294 15470 7322 15471
rect 7082 15301 7110 15302
rect 7082 15275 7100 15301
rect 7100 15275 7110 15301
rect 7082 15274 7110 15275
rect 7134 15301 7162 15302
rect 7134 15275 7136 15301
rect 7136 15275 7162 15301
rect 7134 15274 7162 15275
rect 7186 15301 7214 15302
rect 7238 15301 7266 15302
rect 7186 15275 7198 15301
rect 7198 15275 7214 15301
rect 7238 15275 7260 15301
rect 7260 15275 7266 15301
rect 7186 15274 7214 15275
rect 7238 15274 7266 15275
rect 7290 15274 7318 15302
rect 7342 15301 7370 15302
rect 7394 15301 7422 15302
rect 7342 15275 7348 15301
rect 7348 15275 7370 15301
rect 7394 15275 7410 15301
rect 7410 15275 7422 15301
rect 7342 15274 7370 15275
rect 7394 15274 7422 15275
rect 7446 15301 7474 15302
rect 7446 15275 7472 15301
rect 7472 15275 7474 15301
rect 7446 15274 7474 15275
rect 7498 15301 7526 15302
rect 7498 15275 7508 15301
rect 7508 15275 7526 15301
rect 7498 15274 7526 15275
rect 7798 15889 7826 15890
rect 7798 15863 7799 15889
rect 7799 15863 7825 15889
rect 7825 15863 7826 15889
rect 7798 15862 7826 15863
rect 7798 15470 7826 15498
rect 7574 15022 7602 15050
rect 6902 13510 6930 13538
rect 6958 13958 6986 13986
rect 7082 14517 7110 14518
rect 7082 14491 7100 14517
rect 7100 14491 7110 14517
rect 7082 14490 7110 14491
rect 7134 14517 7162 14518
rect 7134 14491 7136 14517
rect 7136 14491 7162 14517
rect 7134 14490 7162 14491
rect 7186 14517 7214 14518
rect 7238 14517 7266 14518
rect 7186 14491 7198 14517
rect 7198 14491 7214 14517
rect 7238 14491 7260 14517
rect 7260 14491 7266 14517
rect 7186 14490 7214 14491
rect 7238 14490 7266 14491
rect 7290 14490 7318 14518
rect 7342 14517 7370 14518
rect 7394 14517 7422 14518
rect 7342 14491 7348 14517
rect 7348 14491 7370 14517
rect 7394 14491 7410 14517
rect 7410 14491 7422 14517
rect 7342 14490 7370 14491
rect 7394 14490 7422 14491
rect 7446 14517 7474 14518
rect 7446 14491 7472 14517
rect 7472 14491 7474 14517
rect 7446 14490 7474 14491
rect 7498 14517 7526 14518
rect 7498 14491 7508 14517
rect 7508 14491 7526 14517
rect 7498 14490 7526 14491
rect 9582 16477 9610 16478
rect 9582 16451 9600 16477
rect 9600 16451 9610 16477
rect 9582 16450 9610 16451
rect 9634 16477 9662 16478
rect 9634 16451 9636 16477
rect 9636 16451 9662 16477
rect 9634 16450 9662 16451
rect 9686 16477 9714 16478
rect 9738 16477 9766 16478
rect 9686 16451 9698 16477
rect 9698 16451 9714 16477
rect 9738 16451 9760 16477
rect 9760 16451 9766 16477
rect 9686 16450 9714 16451
rect 9738 16450 9766 16451
rect 9790 16450 9818 16478
rect 9842 16477 9870 16478
rect 9894 16477 9922 16478
rect 9842 16451 9848 16477
rect 9848 16451 9870 16477
rect 9894 16451 9910 16477
rect 9910 16451 9922 16477
rect 9842 16450 9870 16451
rect 9894 16450 9922 16451
rect 9946 16477 9974 16478
rect 9946 16451 9972 16477
rect 9972 16451 9974 16477
rect 9946 16450 9974 16451
rect 9998 16477 10026 16478
rect 9998 16451 10008 16477
rect 10008 16451 10026 16477
rect 9998 16450 10026 16451
rect 10150 16310 10178 16338
rect 9310 15862 9338 15890
rect 9478 16254 9506 16282
rect 9982 16281 10010 16282
rect 9982 16255 9983 16281
rect 9983 16255 10009 16281
rect 10009 16255 10010 16281
rect 9982 16254 10010 16255
rect 10822 16337 10850 16338
rect 10822 16311 10823 16337
rect 10823 16311 10849 16337
rect 10849 16311 10850 16337
rect 10822 16310 10850 16311
rect 9582 15693 9610 15694
rect 9582 15667 9600 15693
rect 9600 15667 9610 15693
rect 9582 15666 9610 15667
rect 9634 15693 9662 15694
rect 9634 15667 9636 15693
rect 9636 15667 9662 15693
rect 9634 15666 9662 15667
rect 9686 15693 9714 15694
rect 9738 15693 9766 15694
rect 9686 15667 9698 15693
rect 9698 15667 9714 15693
rect 9738 15667 9760 15693
rect 9760 15667 9766 15693
rect 9686 15666 9714 15667
rect 9738 15666 9766 15667
rect 9790 15666 9818 15694
rect 9842 15693 9870 15694
rect 9894 15693 9922 15694
rect 9842 15667 9848 15693
rect 9848 15667 9870 15693
rect 9894 15667 9910 15693
rect 9910 15667 9922 15693
rect 9842 15666 9870 15667
rect 9894 15666 9922 15667
rect 9946 15693 9974 15694
rect 9946 15667 9972 15693
rect 9972 15667 9974 15693
rect 9946 15666 9974 15667
rect 9998 15693 10026 15694
rect 9998 15667 10008 15693
rect 10008 15667 10026 15693
rect 9998 15666 10026 15667
rect 8974 15105 9002 15106
rect 8974 15079 8975 15105
rect 8975 15079 9001 15105
rect 9001 15079 9002 15105
rect 8974 15078 9002 15079
rect 7014 13902 7042 13930
rect 7082 13733 7110 13734
rect 7082 13707 7100 13733
rect 7100 13707 7110 13733
rect 7082 13706 7110 13707
rect 7134 13733 7162 13734
rect 7134 13707 7136 13733
rect 7136 13707 7162 13733
rect 7134 13706 7162 13707
rect 7186 13733 7214 13734
rect 7238 13733 7266 13734
rect 7186 13707 7198 13733
rect 7198 13707 7214 13733
rect 7238 13707 7260 13733
rect 7260 13707 7266 13733
rect 7186 13706 7214 13707
rect 7238 13706 7266 13707
rect 7290 13706 7318 13734
rect 7342 13733 7370 13734
rect 7394 13733 7422 13734
rect 7342 13707 7348 13733
rect 7348 13707 7370 13733
rect 7394 13707 7410 13733
rect 7410 13707 7422 13733
rect 7342 13706 7370 13707
rect 7394 13706 7422 13707
rect 7446 13733 7474 13734
rect 7446 13707 7472 13733
rect 7472 13707 7474 13733
rect 7446 13706 7474 13707
rect 7498 13733 7526 13734
rect 7498 13707 7508 13733
rect 7508 13707 7526 13733
rect 7498 13706 7526 13707
rect 6958 13454 6986 13482
rect 7082 12949 7110 12950
rect 7082 12923 7100 12949
rect 7100 12923 7110 12949
rect 7082 12922 7110 12923
rect 7134 12949 7162 12950
rect 7134 12923 7136 12949
rect 7136 12923 7162 12949
rect 7134 12922 7162 12923
rect 7186 12949 7214 12950
rect 7238 12949 7266 12950
rect 7186 12923 7198 12949
rect 7198 12923 7214 12949
rect 7238 12923 7260 12949
rect 7260 12923 7266 12949
rect 7186 12922 7214 12923
rect 7238 12922 7266 12923
rect 7290 12922 7318 12950
rect 7342 12949 7370 12950
rect 7394 12949 7422 12950
rect 7342 12923 7348 12949
rect 7348 12923 7370 12949
rect 7394 12923 7410 12949
rect 7410 12923 7422 12949
rect 7342 12922 7370 12923
rect 7394 12922 7422 12923
rect 7446 12949 7474 12950
rect 7446 12923 7472 12949
rect 7472 12923 7474 12949
rect 7446 12922 7474 12923
rect 7498 12949 7526 12950
rect 7498 12923 7508 12949
rect 7508 12923 7526 12949
rect 7498 12922 7526 12923
rect 8470 13985 8498 13986
rect 8470 13959 8471 13985
rect 8471 13959 8497 13985
rect 8497 13959 8498 13985
rect 8470 13958 8498 13959
rect 8974 13958 9002 13986
rect 10150 15134 10178 15162
rect 10934 16254 10962 16282
rect 12614 17318 12642 17346
rect 12082 16869 12110 16870
rect 12082 16843 12100 16869
rect 12100 16843 12110 16869
rect 12082 16842 12110 16843
rect 12134 16869 12162 16870
rect 12134 16843 12136 16869
rect 12136 16843 12162 16869
rect 12134 16842 12162 16843
rect 12186 16869 12214 16870
rect 12238 16869 12266 16870
rect 12186 16843 12198 16869
rect 12198 16843 12214 16869
rect 12238 16843 12260 16869
rect 12260 16843 12266 16869
rect 12186 16842 12214 16843
rect 12238 16842 12266 16843
rect 12290 16842 12318 16870
rect 12342 16869 12370 16870
rect 12394 16869 12422 16870
rect 12342 16843 12348 16869
rect 12348 16843 12370 16869
rect 12394 16843 12410 16869
rect 12410 16843 12422 16869
rect 12342 16842 12370 16843
rect 12394 16842 12422 16843
rect 12446 16869 12474 16870
rect 12446 16843 12472 16869
rect 12472 16843 12474 16869
rect 12446 16842 12474 16843
rect 12498 16869 12526 16870
rect 12498 16843 12508 16869
rect 12508 16843 12526 16869
rect 12498 16842 12526 16843
rect 11998 16590 12026 16618
rect 12334 16590 12362 16618
rect 11382 16310 11410 16338
rect 11158 16281 11186 16282
rect 11158 16255 11159 16281
rect 11159 16255 11185 16281
rect 11185 16255 11186 16281
rect 11158 16254 11186 16255
rect 12614 16534 12642 16562
rect 12082 16085 12110 16086
rect 12082 16059 12100 16085
rect 12100 16059 12110 16085
rect 12082 16058 12110 16059
rect 12134 16085 12162 16086
rect 12134 16059 12136 16085
rect 12136 16059 12162 16085
rect 12134 16058 12162 16059
rect 12186 16085 12214 16086
rect 12238 16085 12266 16086
rect 12186 16059 12198 16085
rect 12198 16059 12214 16085
rect 12238 16059 12260 16085
rect 12260 16059 12266 16085
rect 12186 16058 12214 16059
rect 12238 16058 12266 16059
rect 12290 16058 12318 16086
rect 12342 16085 12370 16086
rect 12394 16085 12422 16086
rect 12342 16059 12348 16085
rect 12348 16059 12370 16085
rect 12394 16059 12410 16085
rect 12410 16059 12422 16085
rect 12342 16058 12370 16059
rect 12394 16058 12422 16059
rect 12446 16085 12474 16086
rect 12446 16059 12472 16085
rect 12472 16059 12474 16085
rect 12446 16058 12474 16059
rect 12498 16085 12526 16086
rect 12498 16059 12508 16085
rect 12508 16059 12526 16085
rect 12498 16058 12526 16059
rect 14582 17261 14610 17262
rect 14582 17235 14600 17261
rect 14600 17235 14610 17261
rect 14582 17234 14610 17235
rect 14634 17261 14662 17262
rect 14634 17235 14636 17261
rect 14636 17235 14662 17261
rect 14634 17234 14662 17235
rect 14686 17261 14714 17262
rect 14738 17261 14766 17262
rect 14686 17235 14698 17261
rect 14698 17235 14714 17261
rect 14738 17235 14760 17261
rect 14760 17235 14766 17261
rect 14686 17234 14714 17235
rect 14738 17234 14766 17235
rect 14790 17234 14818 17262
rect 14842 17261 14870 17262
rect 14894 17261 14922 17262
rect 14842 17235 14848 17261
rect 14848 17235 14870 17261
rect 14894 17235 14910 17261
rect 14910 17235 14922 17261
rect 14842 17234 14870 17235
rect 14894 17234 14922 17235
rect 14946 17261 14974 17262
rect 14946 17235 14972 17261
rect 14972 17235 14974 17261
rect 14946 17234 14974 17235
rect 14998 17261 15026 17262
rect 14998 17235 15008 17261
rect 15008 17235 15026 17261
rect 14998 17234 15026 17235
rect 12950 16142 12978 16170
rect 11102 15862 11130 15890
rect 9582 14909 9610 14910
rect 9582 14883 9600 14909
rect 9600 14883 9610 14909
rect 9582 14882 9610 14883
rect 9634 14909 9662 14910
rect 9634 14883 9636 14909
rect 9636 14883 9662 14909
rect 9634 14882 9662 14883
rect 9686 14909 9714 14910
rect 9738 14909 9766 14910
rect 9686 14883 9698 14909
rect 9698 14883 9714 14909
rect 9738 14883 9760 14909
rect 9760 14883 9766 14909
rect 9686 14882 9714 14883
rect 9738 14882 9766 14883
rect 9790 14882 9818 14910
rect 9842 14909 9870 14910
rect 9894 14909 9922 14910
rect 9842 14883 9848 14909
rect 9848 14883 9870 14909
rect 9894 14883 9910 14909
rect 9910 14883 9922 14909
rect 9842 14882 9870 14883
rect 9894 14882 9922 14883
rect 9946 14909 9974 14910
rect 9946 14883 9972 14909
rect 9972 14883 9974 14909
rect 9946 14882 9974 14883
rect 9998 14909 10026 14910
rect 9998 14883 10008 14909
rect 10008 14883 10026 14909
rect 9998 14882 10026 14883
rect 9582 14125 9610 14126
rect 9582 14099 9600 14125
rect 9600 14099 9610 14125
rect 9582 14098 9610 14099
rect 9634 14125 9662 14126
rect 9634 14099 9636 14125
rect 9636 14099 9662 14125
rect 9634 14098 9662 14099
rect 9686 14125 9714 14126
rect 9738 14125 9766 14126
rect 9686 14099 9698 14125
rect 9698 14099 9714 14125
rect 9738 14099 9760 14125
rect 9760 14099 9766 14125
rect 9686 14098 9714 14099
rect 9738 14098 9766 14099
rect 9790 14098 9818 14126
rect 9842 14125 9870 14126
rect 9894 14125 9922 14126
rect 9842 14099 9848 14125
rect 9848 14099 9870 14125
rect 9894 14099 9910 14125
rect 9910 14099 9922 14125
rect 9842 14098 9870 14099
rect 9894 14098 9922 14099
rect 9946 14125 9974 14126
rect 9946 14099 9972 14125
rect 9972 14099 9974 14125
rect 9946 14098 9974 14099
rect 9998 14125 10026 14126
rect 9998 14099 10008 14125
rect 10008 14099 10026 14125
rect 9998 14098 10026 14099
rect 9582 13341 9610 13342
rect 9582 13315 9600 13341
rect 9600 13315 9610 13341
rect 9582 13314 9610 13315
rect 9634 13341 9662 13342
rect 9634 13315 9636 13341
rect 9636 13315 9662 13341
rect 9634 13314 9662 13315
rect 9686 13341 9714 13342
rect 9738 13341 9766 13342
rect 9686 13315 9698 13341
rect 9698 13315 9714 13341
rect 9738 13315 9760 13341
rect 9760 13315 9766 13341
rect 9686 13314 9714 13315
rect 9738 13314 9766 13315
rect 9790 13314 9818 13342
rect 9842 13341 9870 13342
rect 9894 13341 9922 13342
rect 9842 13315 9848 13341
rect 9848 13315 9870 13341
rect 9894 13315 9910 13341
rect 9910 13315 9922 13341
rect 9842 13314 9870 13315
rect 9894 13314 9922 13315
rect 9946 13341 9974 13342
rect 9946 13315 9972 13341
rect 9972 13315 9974 13341
rect 9946 13314 9974 13315
rect 9998 13341 10026 13342
rect 9998 13315 10008 13341
rect 10008 13315 10026 13341
rect 9998 13314 10026 13315
rect 7082 12165 7110 12166
rect 7082 12139 7100 12165
rect 7100 12139 7110 12165
rect 7082 12138 7110 12139
rect 7134 12165 7162 12166
rect 7134 12139 7136 12165
rect 7136 12139 7162 12165
rect 7134 12138 7162 12139
rect 7186 12165 7214 12166
rect 7238 12165 7266 12166
rect 7186 12139 7198 12165
rect 7198 12139 7214 12165
rect 7238 12139 7260 12165
rect 7260 12139 7266 12165
rect 7186 12138 7214 12139
rect 7238 12138 7266 12139
rect 7290 12138 7318 12166
rect 7342 12165 7370 12166
rect 7394 12165 7422 12166
rect 7342 12139 7348 12165
rect 7348 12139 7370 12165
rect 7394 12139 7410 12165
rect 7410 12139 7422 12165
rect 7342 12138 7370 12139
rect 7394 12138 7422 12139
rect 7446 12165 7474 12166
rect 7446 12139 7472 12165
rect 7472 12139 7474 12165
rect 7446 12138 7474 12139
rect 7498 12165 7526 12166
rect 7498 12139 7508 12165
rect 7508 12139 7526 12165
rect 7498 12138 7526 12139
rect 7014 11774 7042 11802
rect 9582 12557 9610 12558
rect 9582 12531 9600 12557
rect 9600 12531 9610 12557
rect 9582 12530 9610 12531
rect 9634 12557 9662 12558
rect 9634 12531 9636 12557
rect 9636 12531 9662 12557
rect 9634 12530 9662 12531
rect 9686 12557 9714 12558
rect 9738 12557 9766 12558
rect 9686 12531 9698 12557
rect 9698 12531 9714 12557
rect 9738 12531 9760 12557
rect 9760 12531 9766 12557
rect 9686 12530 9714 12531
rect 9738 12530 9766 12531
rect 9790 12530 9818 12558
rect 9842 12557 9870 12558
rect 9894 12557 9922 12558
rect 9842 12531 9848 12557
rect 9848 12531 9870 12557
rect 9894 12531 9910 12557
rect 9910 12531 9922 12557
rect 9842 12530 9870 12531
rect 9894 12530 9922 12531
rect 9946 12557 9974 12558
rect 9946 12531 9972 12557
rect 9972 12531 9974 12557
rect 9946 12530 9974 12531
rect 9998 12557 10026 12558
rect 9998 12531 10008 12557
rect 10008 12531 10026 12557
rect 9998 12530 10026 12531
rect 8470 11969 8498 11970
rect 8470 11943 8471 11969
rect 8471 11943 8497 11969
rect 8497 11943 8498 11969
rect 8470 11942 8498 11943
rect 7082 11381 7110 11382
rect 7082 11355 7100 11381
rect 7100 11355 7110 11381
rect 7082 11354 7110 11355
rect 7134 11381 7162 11382
rect 7134 11355 7136 11381
rect 7136 11355 7162 11381
rect 7134 11354 7162 11355
rect 7186 11381 7214 11382
rect 7238 11381 7266 11382
rect 7186 11355 7198 11381
rect 7198 11355 7214 11381
rect 7238 11355 7260 11381
rect 7260 11355 7266 11381
rect 7186 11354 7214 11355
rect 7238 11354 7266 11355
rect 7290 11354 7318 11382
rect 7342 11381 7370 11382
rect 7394 11381 7422 11382
rect 7342 11355 7348 11381
rect 7348 11355 7370 11381
rect 7394 11355 7410 11381
rect 7410 11355 7422 11381
rect 7342 11354 7370 11355
rect 7394 11354 7422 11355
rect 7446 11381 7474 11382
rect 7446 11355 7472 11381
rect 7472 11355 7474 11381
rect 7446 11354 7474 11355
rect 7498 11381 7526 11382
rect 7498 11355 7508 11381
rect 7508 11355 7526 11381
rect 7498 11354 7526 11355
rect 10878 14294 10906 14322
rect 12082 15301 12110 15302
rect 12082 15275 12100 15301
rect 12100 15275 12110 15301
rect 12082 15274 12110 15275
rect 12134 15301 12162 15302
rect 12134 15275 12136 15301
rect 12136 15275 12162 15301
rect 12134 15274 12162 15275
rect 12186 15301 12214 15302
rect 12238 15301 12266 15302
rect 12186 15275 12198 15301
rect 12198 15275 12214 15301
rect 12238 15275 12260 15301
rect 12260 15275 12266 15301
rect 12186 15274 12214 15275
rect 12238 15274 12266 15275
rect 12290 15274 12318 15302
rect 12342 15301 12370 15302
rect 12394 15301 12422 15302
rect 12342 15275 12348 15301
rect 12348 15275 12370 15301
rect 12394 15275 12410 15301
rect 12410 15275 12422 15301
rect 12342 15274 12370 15275
rect 12394 15274 12422 15275
rect 12446 15301 12474 15302
rect 12446 15275 12472 15301
rect 12472 15275 12474 15301
rect 12446 15274 12474 15275
rect 12498 15301 12526 15302
rect 12498 15275 12508 15301
rect 12508 15275 12526 15301
rect 12498 15274 12526 15275
rect 11214 13398 11242 13426
rect 11550 13398 11578 13426
rect 8358 11774 8386 11802
rect 6118 8441 6146 8442
rect 6118 8415 6119 8441
rect 6119 8415 6145 8441
rect 6145 8415 6146 8441
rect 6118 8414 6146 8415
rect 6118 7657 6146 7658
rect 6118 7631 6119 7657
rect 6119 7631 6145 7657
rect 6145 7631 6146 7657
rect 6118 7630 6146 7631
rect 6510 7686 6538 7714
rect 5558 6481 5586 6482
rect 5558 6455 5559 6481
rect 5559 6455 5585 6481
rect 5585 6455 5586 6481
rect 5558 6454 5586 6455
rect 5558 5054 5586 5082
rect 6454 7209 6482 7210
rect 6454 7183 6455 7209
rect 6455 7183 6481 7209
rect 6481 7183 6482 7209
rect 6454 7182 6482 7183
rect 5782 4606 5810 4634
rect 5446 2646 5474 2674
rect 5726 3345 5754 3346
rect 5726 3319 5727 3345
rect 5727 3319 5753 3345
rect 5753 3319 5754 3345
rect 5726 3318 5754 3319
rect 4998 2561 5026 2562
rect 4998 2535 4999 2561
rect 4999 2535 5025 2561
rect 5025 2535 5026 2561
rect 4998 2534 5026 2535
rect 5726 2561 5754 2562
rect 5726 2535 5727 2561
rect 5727 2535 5753 2561
rect 5753 2535 5754 2561
rect 5726 2534 5754 2535
rect 4102 2422 4130 2450
rect 4582 2365 4610 2366
rect 4582 2339 4600 2365
rect 4600 2339 4610 2365
rect 4582 2338 4610 2339
rect 4634 2365 4662 2366
rect 4634 2339 4636 2365
rect 4636 2339 4662 2365
rect 4634 2338 4662 2339
rect 4686 2365 4714 2366
rect 4738 2365 4766 2366
rect 4686 2339 4698 2365
rect 4698 2339 4714 2365
rect 4738 2339 4760 2365
rect 4760 2339 4766 2365
rect 4686 2338 4714 2339
rect 4738 2338 4766 2339
rect 4790 2338 4818 2366
rect 4842 2365 4870 2366
rect 4894 2365 4922 2366
rect 4842 2339 4848 2365
rect 4848 2339 4870 2365
rect 4894 2339 4910 2365
rect 4910 2339 4922 2365
rect 4842 2338 4870 2339
rect 4894 2338 4922 2339
rect 4946 2365 4974 2366
rect 4946 2339 4972 2365
rect 4972 2339 4974 2365
rect 4946 2338 4974 2339
rect 4998 2365 5026 2366
rect 4998 2339 5008 2365
rect 5008 2339 5026 2365
rect 4998 2338 5026 2339
rect 3934 1862 3962 1890
rect 4494 2225 4522 2226
rect 4494 2199 4495 2225
rect 4495 2199 4521 2225
rect 4521 2199 4522 2225
rect 4494 2198 4522 2199
rect 5502 2142 5530 2170
rect 4494 2086 4522 2114
rect 5502 1638 5530 1666
rect 4582 1581 4610 1582
rect 4582 1555 4600 1581
rect 4600 1555 4610 1581
rect 4582 1554 4610 1555
rect 4634 1581 4662 1582
rect 4634 1555 4636 1581
rect 4636 1555 4662 1581
rect 4634 1554 4662 1555
rect 4686 1581 4714 1582
rect 4738 1581 4766 1582
rect 4686 1555 4698 1581
rect 4698 1555 4714 1581
rect 4738 1555 4760 1581
rect 4760 1555 4766 1581
rect 4686 1554 4714 1555
rect 4738 1554 4766 1555
rect 4790 1554 4818 1582
rect 4842 1581 4870 1582
rect 4894 1581 4922 1582
rect 4842 1555 4848 1581
rect 4848 1555 4870 1581
rect 4894 1555 4910 1581
rect 4910 1555 4922 1581
rect 4842 1554 4870 1555
rect 4894 1554 4922 1555
rect 4946 1581 4974 1582
rect 4946 1555 4972 1581
rect 4972 1555 4974 1581
rect 4946 1554 4974 1555
rect 4998 1581 5026 1582
rect 4998 1555 5008 1581
rect 5008 1555 5026 1581
rect 4998 1554 5026 1555
rect 6510 5305 6538 5306
rect 6510 5279 6511 5305
rect 6511 5279 6537 5305
rect 6537 5279 6538 5305
rect 6510 5278 6538 5279
rect 6006 4521 6034 4522
rect 6006 4495 6007 4521
rect 6007 4495 6033 4521
rect 6033 4495 6034 4521
rect 6006 4494 6034 4495
rect 6006 4214 6034 4242
rect 6454 4158 6482 4186
rect 6006 3345 6034 3346
rect 6006 3319 6007 3345
rect 6007 3319 6033 3345
rect 6033 3319 6034 3345
rect 6006 3318 6034 3319
rect 5838 2534 5866 2562
rect 6454 2561 6482 2562
rect 6454 2535 6455 2561
rect 6455 2535 6481 2561
rect 6481 2535 6482 2561
rect 6454 2534 6482 2535
rect 6342 2198 6370 2226
rect 6398 1721 6426 1722
rect 6398 1695 6399 1721
rect 6399 1695 6425 1721
rect 6425 1695 6426 1721
rect 6398 1694 6426 1695
rect 7294 10934 7322 10962
rect 7574 10934 7602 10962
rect 7082 10597 7110 10598
rect 7082 10571 7100 10597
rect 7100 10571 7110 10597
rect 7082 10570 7110 10571
rect 7134 10597 7162 10598
rect 7134 10571 7136 10597
rect 7136 10571 7162 10597
rect 7134 10570 7162 10571
rect 7186 10597 7214 10598
rect 7238 10597 7266 10598
rect 7186 10571 7198 10597
rect 7198 10571 7214 10597
rect 7238 10571 7260 10597
rect 7260 10571 7266 10597
rect 7186 10570 7214 10571
rect 7238 10570 7266 10571
rect 7290 10570 7318 10598
rect 7342 10597 7370 10598
rect 7394 10597 7422 10598
rect 7342 10571 7348 10597
rect 7348 10571 7370 10597
rect 7394 10571 7410 10597
rect 7410 10571 7422 10597
rect 7342 10570 7370 10571
rect 7394 10570 7422 10571
rect 7446 10597 7474 10598
rect 7446 10571 7472 10597
rect 7472 10571 7474 10597
rect 7446 10570 7474 10571
rect 7498 10597 7526 10598
rect 7498 10571 7508 10597
rect 7508 10571 7526 10597
rect 7498 10570 7526 10571
rect 7014 10009 7042 10010
rect 7014 9983 7015 10009
rect 7015 9983 7041 10009
rect 7041 9983 7042 10009
rect 7014 9982 7042 9983
rect 7082 9813 7110 9814
rect 7082 9787 7100 9813
rect 7100 9787 7110 9813
rect 7082 9786 7110 9787
rect 7134 9813 7162 9814
rect 7134 9787 7136 9813
rect 7136 9787 7162 9813
rect 7134 9786 7162 9787
rect 7186 9813 7214 9814
rect 7238 9813 7266 9814
rect 7186 9787 7198 9813
rect 7198 9787 7214 9813
rect 7238 9787 7260 9813
rect 7260 9787 7266 9813
rect 7186 9786 7214 9787
rect 7238 9786 7266 9787
rect 7290 9786 7318 9814
rect 7342 9813 7370 9814
rect 7394 9813 7422 9814
rect 7342 9787 7348 9813
rect 7348 9787 7370 9813
rect 7394 9787 7410 9813
rect 7410 9787 7422 9813
rect 7342 9786 7370 9787
rect 7394 9786 7422 9787
rect 7446 9813 7474 9814
rect 7446 9787 7472 9813
rect 7472 9787 7474 9813
rect 7446 9786 7474 9787
rect 7498 9813 7526 9814
rect 7498 9787 7508 9813
rect 7508 9787 7526 9813
rect 7498 9786 7526 9787
rect 10430 11969 10458 11970
rect 10430 11943 10431 11969
rect 10431 11943 10457 11969
rect 10457 11943 10458 11969
rect 10430 11942 10458 11943
rect 9582 11773 9610 11774
rect 9582 11747 9600 11773
rect 9600 11747 9610 11773
rect 9582 11746 9610 11747
rect 9634 11773 9662 11774
rect 9634 11747 9636 11773
rect 9636 11747 9662 11773
rect 9634 11746 9662 11747
rect 9686 11773 9714 11774
rect 9738 11773 9766 11774
rect 9686 11747 9698 11773
rect 9698 11747 9714 11773
rect 9738 11747 9760 11773
rect 9760 11747 9766 11773
rect 9686 11746 9714 11747
rect 9738 11746 9766 11747
rect 9790 11746 9818 11774
rect 9842 11773 9870 11774
rect 9894 11773 9922 11774
rect 9842 11747 9848 11773
rect 9848 11747 9870 11773
rect 9894 11747 9910 11773
rect 9910 11747 9922 11773
rect 9842 11746 9870 11747
rect 9894 11746 9922 11747
rect 9946 11773 9974 11774
rect 9946 11747 9972 11773
rect 9972 11747 9974 11773
rect 9946 11746 9974 11747
rect 9998 11773 10026 11774
rect 9998 11747 10008 11773
rect 10008 11747 10026 11773
rect 9998 11746 10026 11747
rect 9254 10934 9282 10962
rect 9582 10989 9610 10990
rect 9582 10963 9600 10989
rect 9600 10963 9610 10989
rect 9582 10962 9610 10963
rect 9634 10989 9662 10990
rect 9634 10963 9636 10989
rect 9636 10963 9662 10989
rect 9634 10962 9662 10963
rect 9686 10989 9714 10990
rect 9738 10989 9766 10990
rect 9686 10963 9698 10989
rect 9698 10963 9714 10989
rect 9738 10963 9760 10989
rect 9760 10963 9766 10989
rect 9686 10962 9714 10963
rect 9738 10962 9766 10963
rect 9790 10962 9818 10990
rect 9842 10989 9870 10990
rect 9894 10989 9922 10990
rect 9842 10963 9848 10989
rect 9848 10963 9870 10989
rect 9894 10963 9910 10989
rect 9910 10963 9922 10989
rect 9842 10962 9870 10963
rect 9894 10962 9922 10963
rect 9946 10989 9974 10990
rect 9946 10963 9972 10989
rect 9972 10963 9974 10989
rect 9946 10962 9974 10963
rect 9998 10989 10026 10990
rect 9998 10963 10008 10989
rect 10008 10963 10026 10989
rect 9998 10962 10026 10963
rect 8806 10094 8834 10122
rect 8750 9982 8778 10010
rect 7082 9029 7110 9030
rect 7082 9003 7100 9029
rect 7100 9003 7110 9029
rect 7082 9002 7110 9003
rect 7134 9029 7162 9030
rect 7134 9003 7136 9029
rect 7136 9003 7162 9029
rect 7134 9002 7162 9003
rect 7186 9029 7214 9030
rect 7238 9029 7266 9030
rect 7186 9003 7198 9029
rect 7198 9003 7214 9029
rect 7238 9003 7260 9029
rect 7260 9003 7266 9029
rect 7186 9002 7214 9003
rect 7238 9002 7266 9003
rect 7290 9002 7318 9030
rect 7342 9029 7370 9030
rect 7394 9029 7422 9030
rect 7342 9003 7348 9029
rect 7348 9003 7370 9029
rect 7394 9003 7410 9029
rect 7410 9003 7422 9029
rect 7342 9002 7370 9003
rect 7394 9002 7422 9003
rect 7446 9029 7474 9030
rect 7446 9003 7472 9029
rect 7472 9003 7474 9029
rect 7446 9002 7474 9003
rect 7498 9029 7526 9030
rect 7498 9003 7508 9029
rect 7508 9003 7526 9029
rect 7498 9002 7526 9003
rect 7014 8414 7042 8442
rect 7082 8245 7110 8246
rect 7082 8219 7100 8245
rect 7100 8219 7110 8245
rect 7082 8218 7110 8219
rect 7134 8245 7162 8246
rect 7134 8219 7136 8245
rect 7136 8219 7162 8245
rect 7134 8218 7162 8219
rect 7186 8245 7214 8246
rect 7238 8245 7266 8246
rect 7186 8219 7198 8245
rect 7198 8219 7214 8245
rect 7238 8219 7260 8245
rect 7260 8219 7266 8245
rect 7186 8218 7214 8219
rect 7238 8218 7266 8219
rect 7290 8218 7318 8246
rect 7342 8245 7370 8246
rect 7394 8245 7422 8246
rect 7342 8219 7348 8245
rect 7348 8219 7370 8245
rect 7394 8219 7410 8245
rect 7410 8219 7422 8245
rect 7342 8218 7370 8219
rect 7394 8218 7422 8219
rect 7446 8245 7474 8246
rect 7446 8219 7472 8245
rect 7472 8219 7474 8245
rect 7446 8218 7474 8219
rect 7498 8245 7526 8246
rect 7498 8219 7508 8245
rect 7508 8219 7526 8245
rect 7498 8218 7526 8219
rect 7294 7518 7322 7546
rect 8750 8049 8778 8050
rect 8750 8023 8751 8049
rect 8751 8023 8777 8049
rect 8777 8023 8778 8049
rect 8750 8022 8778 8023
rect 7574 7630 7602 7658
rect 7082 7461 7110 7462
rect 7082 7435 7100 7461
rect 7100 7435 7110 7461
rect 7082 7434 7110 7435
rect 7134 7461 7162 7462
rect 7134 7435 7136 7461
rect 7136 7435 7162 7461
rect 7134 7434 7162 7435
rect 7186 7461 7214 7462
rect 7238 7461 7266 7462
rect 7186 7435 7198 7461
rect 7198 7435 7214 7461
rect 7238 7435 7260 7461
rect 7260 7435 7266 7461
rect 7186 7434 7214 7435
rect 7238 7434 7266 7435
rect 7290 7434 7318 7462
rect 7342 7461 7370 7462
rect 7394 7461 7422 7462
rect 7342 7435 7348 7461
rect 7348 7435 7370 7461
rect 7394 7435 7410 7461
rect 7410 7435 7422 7461
rect 7342 7434 7370 7435
rect 7394 7434 7422 7435
rect 7446 7461 7474 7462
rect 7446 7435 7472 7461
rect 7472 7435 7474 7461
rect 7446 7434 7474 7435
rect 7498 7461 7526 7462
rect 7498 7435 7508 7461
rect 7508 7435 7526 7461
rect 7498 7434 7526 7435
rect 7742 7686 7770 7714
rect 6958 7182 6986 7210
rect 7798 7518 7826 7546
rect 8470 7462 8498 7490
rect 7082 6677 7110 6678
rect 7082 6651 7100 6677
rect 7100 6651 7110 6677
rect 7082 6650 7110 6651
rect 7134 6677 7162 6678
rect 7134 6651 7136 6677
rect 7136 6651 7162 6677
rect 7134 6650 7162 6651
rect 7186 6677 7214 6678
rect 7238 6677 7266 6678
rect 7186 6651 7198 6677
rect 7198 6651 7214 6677
rect 7238 6651 7260 6677
rect 7260 6651 7266 6677
rect 7186 6650 7214 6651
rect 7238 6650 7266 6651
rect 7290 6650 7318 6678
rect 7342 6677 7370 6678
rect 7394 6677 7422 6678
rect 7342 6651 7348 6677
rect 7348 6651 7370 6677
rect 7394 6651 7410 6677
rect 7410 6651 7422 6677
rect 7342 6650 7370 6651
rect 7394 6650 7422 6651
rect 7446 6677 7474 6678
rect 7446 6651 7472 6677
rect 7472 6651 7474 6677
rect 7446 6650 7474 6651
rect 7498 6677 7526 6678
rect 7498 6651 7508 6677
rect 7508 6651 7526 6677
rect 7498 6650 7526 6651
rect 7574 6089 7602 6090
rect 7574 6063 7575 6089
rect 7575 6063 7601 6089
rect 7601 6063 7602 6089
rect 7574 6062 7602 6063
rect 8078 6062 8106 6090
rect 7082 5893 7110 5894
rect 7082 5867 7100 5893
rect 7100 5867 7110 5893
rect 7082 5866 7110 5867
rect 7134 5893 7162 5894
rect 7134 5867 7136 5893
rect 7136 5867 7162 5893
rect 7134 5866 7162 5867
rect 7186 5893 7214 5894
rect 7238 5893 7266 5894
rect 7186 5867 7198 5893
rect 7198 5867 7214 5893
rect 7238 5867 7260 5893
rect 7260 5867 7266 5893
rect 7186 5866 7214 5867
rect 7238 5866 7266 5867
rect 7290 5866 7318 5894
rect 7342 5893 7370 5894
rect 7394 5893 7422 5894
rect 7342 5867 7348 5893
rect 7348 5867 7370 5893
rect 7394 5867 7410 5893
rect 7410 5867 7422 5893
rect 7342 5866 7370 5867
rect 7394 5866 7422 5867
rect 7446 5893 7474 5894
rect 7446 5867 7472 5893
rect 7472 5867 7474 5893
rect 7446 5866 7474 5867
rect 7498 5893 7526 5894
rect 7498 5867 7508 5893
rect 7508 5867 7526 5893
rect 7498 5866 7526 5867
rect 8078 5838 8106 5866
rect 7742 5305 7770 5306
rect 7742 5279 7743 5305
rect 7743 5279 7769 5305
rect 7769 5279 7770 5305
rect 7742 5278 7770 5279
rect 7966 5305 7994 5306
rect 7966 5279 7967 5305
rect 7967 5279 7993 5305
rect 7993 5279 7994 5305
rect 7966 5278 7994 5279
rect 8246 5278 8274 5306
rect 7082 5109 7110 5110
rect 7082 5083 7100 5109
rect 7100 5083 7110 5109
rect 7082 5082 7110 5083
rect 7134 5109 7162 5110
rect 7134 5083 7136 5109
rect 7136 5083 7162 5109
rect 7134 5082 7162 5083
rect 7186 5109 7214 5110
rect 7238 5109 7266 5110
rect 7186 5083 7198 5109
rect 7198 5083 7214 5109
rect 7238 5083 7260 5109
rect 7260 5083 7266 5109
rect 7186 5082 7214 5083
rect 7238 5082 7266 5083
rect 7290 5082 7318 5110
rect 7342 5109 7370 5110
rect 7394 5109 7422 5110
rect 7342 5083 7348 5109
rect 7348 5083 7370 5109
rect 7394 5083 7410 5109
rect 7410 5083 7422 5109
rect 7342 5082 7370 5083
rect 7394 5082 7422 5083
rect 7446 5109 7474 5110
rect 7446 5083 7472 5109
rect 7472 5083 7474 5109
rect 7446 5082 7474 5083
rect 7498 5109 7526 5110
rect 7498 5083 7508 5109
rect 7508 5083 7526 5109
rect 7498 5082 7526 5083
rect 7294 4521 7322 4522
rect 7294 4495 7295 4521
rect 7295 4495 7321 4521
rect 7321 4495 7322 4521
rect 7294 4494 7322 4495
rect 7574 4494 7602 4522
rect 7082 4325 7110 4326
rect 7082 4299 7100 4325
rect 7100 4299 7110 4325
rect 7082 4298 7110 4299
rect 7134 4325 7162 4326
rect 7134 4299 7136 4325
rect 7136 4299 7162 4325
rect 7134 4298 7162 4299
rect 7186 4325 7214 4326
rect 7238 4325 7266 4326
rect 7186 4299 7198 4325
rect 7198 4299 7214 4325
rect 7238 4299 7260 4325
rect 7260 4299 7266 4325
rect 7186 4298 7214 4299
rect 7238 4298 7266 4299
rect 7290 4298 7318 4326
rect 7342 4325 7370 4326
rect 7394 4325 7422 4326
rect 7342 4299 7348 4325
rect 7348 4299 7370 4325
rect 7394 4299 7410 4325
rect 7410 4299 7422 4325
rect 7342 4298 7370 4299
rect 7394 4298 7422 4299
rect 7446 4325 7474 4326
rect 7446 4299 7472 4325
rect 7472 4299 7474 4325
rect 7446 4298 7474 4299
rect 7498 4325 7526 4326
rect 7498 4299 7508 4325
rect 7508 4299 7526 4325
rect 7498 4298 7526 4299
rect 7014 4158 7042 4186
rect 7082 3541 7110 3542
rect 7082 3515 7100 3541
rect 7100 3515 7110 3541
rect 7082 3514 7110 3515
rect 7134 3541 7162 3542
rect 7134 3515 7136 3541
rect 7136 3515 7162 3541
rect 7134 3514 7162 3515
rect 7186 3541 7214 3542
rect 7238 3541 7266 3542
rect 7186 3515 7198 3541
rect 7198 3515 7214 3541
rect 7238 3515 7260 3541
rect 7260 3515 7266 3541
rect 7186 3514 7214 3515
rect 7238 3514 7266 3515
rect 7290 3514 7318 3542
rect 7342 3541 7370 3542
rect 7394 3541 7422 3542
rect 7342 3515 7348 3541
rect 7348 3515 7370 3541
rect 7394 3515 7410 3541
rect 7410 3515 7422 3541
rect 7342 3514 7370 3515
rect 7394 3514 7422 3515
rect 7446 3541 7474 3542
rect 7446 3515 7472 3541
rect 7472 3515 7474 3541
rect 7446 3514 7474 3515
rect 7498 3541 7526 3542
rect 7498 3515 7508 3541
rect 7508 3515 7526 3541
rect 7498 3514 7526 3515
rect 12446 14713 12474 14714
rect 12446 14687 12447 14713
rect 12447 14687 12473 14713
rect 12473 14687 12474 14713
rect 12446 14686 12474 14687
rect 12838 14686 12866 14714
rect 12082 14517 12110 14518
rect 12082 14491 12100 14517
rect 12100 14491 12110 14517
rect 12082 14490 12110 14491
rect 12134 14517 12162 14518
rect 12134 14491 12136 14517
rect 12136 14491 12162 14517
rect 12134 14490 12162 14491
rect 12186 14517 12214 14518
rect 12238 14517 12266 14518
rect 12186 14491 12198 14517
rect 12198 14491 12214 14517
rect 12238 14491 12260 14517
rect 12260 14491 12266 14517
rect 12186 14490 12214 14491
rect 12238 14490 12266 14491
rect 12290 14490 12318 14518
rect 12342 14517 12370 14518
rect 12394 14517 12422 14518
rect 12342 14491 12348 14517
rect 12348 14491 12370 14517
rect 12394 14491 12410 14517
rect 12410 14491 12422 14517
rect 12342 14490 12370 14491
rect 12394 14490 12422 14491
rect 12446 14517 12474 14518
rect 12446 14491 12472 14517
rect 12472 14491 12474 14517
rect 12446 14490 12474 14491
rect 12498 14517 12526 14518
rect 12498 14491 12508 14517
rect 12508 14491 12526 14517
rect 12498 14490 12526 14491
rect 12446 14294 12474 14322
rect 12894 14321 12922 14322
rect 12894 14295 12895 14321
rect 12895 14295 12921 14321
rect 12921 14295 12922 14321
rect 12894 14294 12922 14295
rect 12082 13733 12110 13734
rect 12082 13707 12100 13733
rect 12100 13707 12110 13733
rect 12082 13706 12110 13707
rect 12134 13733 12162 13734
rect 12134 13707 12136 13733
rect 12136 13707 12162 13733
rect 12134 13706 12162 13707
rect 12186 13733 12214 13734
rect 12238 13733 12266 13734
rect 12186 13707 12198 13733
rect 12198 13707 12214 13733
rect 12238 13707 12260 13733
rect 12260 13707 12266 13733
rect 12186 13706 12214 13707
rect 12238 13706 12266 13707
rect 12290 13706 12318 13734
rect 12342 13733 12370 13734
rect 12394 13733 12422 13734
rect 12342 13707 12348 13733
rect 12348 13707 12370 13733
rect 12394 13707 12410 13733
rect 12410 13707 12422 13733
rect 12342 13706 12370 13707
rect 12394 13706 12422 13707
rect 12446 13733 12474 13734
rect 12446 13707 12472 13733
rect 12472 13707 12474 13733
rect 12446 13706 12474 13707
rect 12498 13733 12526 13734
rect 12498 13707 12508 13733
rect 12508 13707 12526 13733
rect 12498 13706 12526 13707
rect 12670 13398 12698 13426
rect 13454 16617 13482 16618
rect 13454 16591 13455 16617
rect 13455 16591 13481 16617
rect 13481 16591 13482 16617
rect 13454 16590 13482 16591
rect 13790 16590 13818 16618
rect 14582 16477 14610 16478
rect 14582 16451 14600 16477
rect 14600 16451 14610 16477
rect 14582 16450 14610 16451
rect 14634 16477 14662 16478
rect 14634 16451 14636 16477
rect 14636 16451 14662 16477
rect 14634 16450 14662 16451
rect 14686 16477 14714 16478
rect 14738 16477 14766 16478
rect 14686 16451 14698 16477
rect 14698 16451 14714 16477
rect 14738 16451 14760 16477
rect 14760 16451 14766 16477
rect 14686 16450 14714 16451
rect 14738 16450 14766 16451
rect 14790 16450 14818 16478
rect 14842 16477 14870 16478
rect 14894 16477 14922 16478
rect 14842 16451 14848 16477
rect 14848 16451 14870 16477
rect 14894 16451 14910 16477
rect 14910 16451 14922 16477
rect 14842 16450 14870 16451
rect 14894 16450 14922 16451
rect 14946 16477 14974 16478
rect 14946 16451 14972 16477
rect 14972 16451 14974 16477
rect 14946 16450 14974 16451
rect 14998 16477 15026 16478
rect 14998 16451 15008 16477
rect 15008 16451 15026 16477
rect 14998 16450 15026 16451
rect 13286 16142 13314 16170
rect 13062 15078 13090 15106
rect 13062 14742 13090 14770
rect 15414 15918 15442 15946
rect 15078 15889 15106 15890
rect 15078 15863 15079 15889
rect 15079 15863 15105 15889
rect 15105 15863 15106 15889
rect 15078 15862 15106 15863
rect 14582 15693 14610 15694
rect 14582 15667 14600 15693
rect 14600 15667 14610 15693
rect 14582 15666 14610 15667
rect 14634 15693 14662 15694
rect 14634 15667 14636 15693
rect 14636 15667 14662 15693
rect 14634 15666 14662 15667
rect 14686 15693 14714 15694
rect 14738 15693 14766 15694
rect 14686 15667 14698 15693
rect 14698 15667 14714 15693
rect 14738 15667 14760 15693
rect 14760 15667 14766 15693
rect 14686 15666 14714 15667
rect 14738 15666 14766 15667
rect 14790 15666 14818 15694
rect 14842 15693 14870 15694
rect 14894 15693 14922 15694
rect 14842 15667 14848 15693
rect 14848 15667 14870 15693
rect 14894 15667 14910 15693
rect 14910 15667 14922 15693
rect 14842 15666 14870 15667
rect 14894 15666 14922 15667
rect 14946 15693 14974 15694
rect 14946 15667 14972 15693
rect 14972 15667 14974 15693
rect 14946 15666 14974 15667
rect 14998 15693 15026 15694
rect 14998 15667 15008 15693
rect 15008 15667 15026 15693
rect 14998 15666 15026 15667
rect 14294 15078 14322 15106
rect 14798 15105 14826 15106
rect 14798 15079 14799 15105
rect 14799 15079 14825 15105
rect 14825 15079 14826 15105
rect 14798 15078 14826 15079
rect 14582 14909 14610 14910
rect 14582 14883 14600 14909
rect 14600 14883 14610 14909
rect 14582 14882 14610 14883
rect 14634 14909 14662 14910
rect 14634 14883 14636 14909
rect 14636 14883 14662 14909
rect 14634 14882 14662 14883
rect 14686 14909 14714 14910
rect 14738 14909 14766 14910
rect 14686 14883 14698 14909
rect 14698 14883 14714 14909
rect 14738 14883 14760 14909
rect 14760 14883 14766 14909
rect 14686 14882 14714 14883
rect 14738 14882 14766 14883
rect 14790 14882 14818 14910
rect 14842 14909 14870 14910
rect 14894 14909 14922 14910
rect 14842 14883 14848 14909
rect 14848 14883 14870 14909
rect 14894 14883 14910 14909
rect 14910 14883 14922 14909
rect 14842 14882 14870 14883
rect 14894 14882 14922 14883
rect 14946 14909 14974 14910
rect 14946 14883 14972 14909
rect 14972 14883 14974 14909
rect 14946 14882 14974 14883
rect 14998 14909 15026 14910
rect 14998 14883 15008 14909
rect 15008 14883 15026 14909
rect 14998 14882 15026 14883
rect 16814 15918 16842 15946
rect 12950 13118 12978 13146
rect 12082 12949 12110 12950
rect 12082 12923 12100 12949
rect 12100 12923 12110 12949
rect 12082 12922 12110 12923
rect 12134 12949 12162 12950
rect 12134 12923 12136 12949
rect 12136 12923 12162 12949
rect 12134 12922 12162 12923
rect 12186 12949 12214 12950
rect 12238 12949 12266 12950
rect 12186 12923 12198 12949
rect 12198 12923 12214 12949
rect 12238 12923 12260 12949
rect 12260 12923 12266 12949
rect 12186 12922 12214 12923
rect 12238 12922 12266 12923
rect 12290 12922 12318 12950
rect 12342 12949 12370 12950
rect 12394 12949 12422 12950
rect 12342 12923 12348 12949
rect 12348 12923 12370 12949
rect 12394 12923 12410 12949
rect 12410 12923 12422 12949
rect 12342 12922 12370 12923
rect 12394 12922 12422 12923
rect 12446 12949 12474 12950
rect 12446 12923 12472 12949
rect 12472 12923 12474 12949
rect 12446 12922 12474 12923
rect 12498 12949 12526 12950
rect 12498 12923 12508 12949
rect 12508 12923 12526 12949
rect 12498 12922 12526 12923
rect 14014 14321 14042 14322
rect 14014 14295 14015 14321
rect 14015 14295 14041 14321
rect 14041 14295 14042 14321
rect 14014 14294 14042 14295
rect 13118 13398 13146 13426
rect 13398 13118 13426 13146
rect 14014 13145 14042 13146
rect 14014 13119 14015 13145
rect 14015 13119 14041 13145
rect 14041 13119 14042 13145
rect 14014 13118 14042 13119
rect 12082 12165 12110 12166
rect 12082 12139 12100 12165
rect 12100 12139 12110 12165
rect 12082 12138 12110 12139
rect 12134 12165 12162 12166
rect 12134 12139 12136 12165
rect 12136 12139 12162 12165
rect 12134 12138 12162 12139
rect 12186 12165 12214 12166
rect 12238 12165 12266 12166
rect 12186 12139 12198 12165
rect 12198 12139 12214 12165
rect 12238 12139 12260 12165
rect 12260 12139 12266 12165
rect 12186 12138 12214 12139
rect 12238 12138 12266 12139
rect 12290 12138 12318 12166
rect 12342 12165 12370 12166
rect 12394 12165 12422 12166
rect 12342 12139 12348 12165
rect 12348 12139 12370 12165
rect 12394 12139 12410 12165
rect 12410 12139 12422 12165
rect 12342 12138 12370 12139
rect 12394 12138 12422 12139
rect 12446 12165 12474 12166
rect 12446 12139 12472 12165
rect 12472 12139 12474 12165
rect 12446 12138 12474 12139
rect 12498 12165 12526 12166
rect 12498 12139 12508 12165
rect 12508 12139 12526 12165
rect 12498 12138 12526 12139
rect 11998 11774 12026 11802
rect 12082 11381 12110 11382
rect 12082 11355 12100 11381
rect 12100 11355 12110 11381
rect 12082 11354 12110 11355
rect 12134 11381 12162 11382
rect 12134 11355 12136 11381
rect 12136 11355 12162 11381
rect 12134 11354 12162 11355
rect 12186 11381 12214 11382
rect 12238 11381 12266 11382
rect 12186 11355 12198 11381
rect 12198 11355 12214 11381
rect 12238 11355 12260 11381
rect 12260 11355 12266 11381
rect 12186 11354 12214 11355
rect 12238 11354 12266 11355
rect 12290 11354 12318 11382
rect 12342 11381 12370 11382
rect 12394 11381 12422 11382
rect 12342 11355 12348 11381
rect 12348 11355 12370 11381
rect 12394 11355 12410 11381
rect 12410 11355 12422 11381
rect 12342 11354 12370 11355
rect 12394 11354 12422 11355
rect 12446 11381 12474 11382
rect 12446 11355 12472 11381
rect 12472 11355 12474 11381
rect 12446 11354 12474 11355
rect 12498 11381 12526 11382
rect 12498 11355 12508 11381
rect 12508 11355 12526 11381
rect 12498 11354 12526 11355
rect 9582 10205 9610 10206
rect 9582 10179 9600 10205
rect 9600 10179 9610 10205
rect 9582 10178 9610 10179
rect 9634 10205 9662 10206
rect 9634 10179 9636 10205
rect 9636 10179 9662 10205
rect 9634 10178 9662 10179
rect 9686 10205 9714 10206
rect 9738 10205 9766 10206
rect 9686 10179 9698 10205
rect 9698 10179 9714 10205
rect 9738 10179 9760 10205
rect 9760 10179 9766 10205
rect 9686 10178 9714 10179
rect 9738 10178 9766 10179
rect 9790 10178 9818 10206
rect 9842 10205 9870 10206
rect 9894 10205 9922 10206
rect 9842 10179 9848 10205
rect 9848 10179 9870 10205
rect 9894 10179 9910 10205
rect 9910 10179 9922 10205
rect 9842 10178 9870 10179
rect 9894 10178 9922 10179
rect 9946 10205 9974 10206
rect 9946 10179 9972 10205
rect 9972 10179 9974 10205
rect 9946 10178 9974 10179
rect 9998 10205 10026 10206
rect 9998 10179 10008 10205
rect 10008 10179 10026 10205
rect 9998 10178 10026 10179
rect 9582 9421 9610 9422
rect 9582 9395 9600 9421
rect 9600 9395 9610 9421
rect 9582 9394 9610 9395
rect 9634 9421 9662 9422
rect 9634 9395 9636 9421
rect 9636 9395 9662 9421
rect 9634 9394 9662 9395
rect 9686 9421 9714 9422
rect 9738 9421 9766 9422
rect 9686 9395 9698 9421
rect 9698 9395 9714 9421
rect 9738 9395 9760 9421
rect 9760 9395 9766 9421
rect 9686 9394 9714 9395
rect 9738 9394 9766 9395
rect 9790 9394 9818 9422
rect 9842 9421 9870 9422
rect 9894 9421 9922 9422
rect 9842 9395 9848 9421
rect 9848 9395 9870 9421
rect 9894 9395 9910 9421
rect 9910 9395 9922 9421
rect 9842 9394 9870 9395
rect 9894 9394 9922 9395
rect 9946 9421 9974 9422
rect 9946 9395 9972 9421
rect 9972 9395 9974 9421
rect 9946 9394 9974 9395
rect 9998 9421 10026 9422
rect 9998 9395 10008 9421
rect 10008 9395 10026 9421
rect 9998 9394 10026 9395
rect 12082 10597 12110 10598
rect 12082 10571 12100 10597
rect 12100 10571 12110 10597
rect 12082 10570 12110 10571
rect 12134 10597 12162 10598
rect 12134 10571 12136 10597
rect 12136 10571 12162 10597
rect 12134 10570 12162 10571
rect 12186 10597 12214 10598
rect 12238 10597 12266 10598
rect 12186 10571 12198 10597
rect 12198 10571 12214 10597
rect 12238 10571 12260 10597
rect 12260 10571 12266 10597
rect 12186 10570 12214 10571
rect 12238 10570 12266 10571
rect 12290 10570 12318 10598
rect 12342 10597 12370 10598
rect 12394 10597 12422 10598
rect 12342 10571 12348 10597
rect 12348 10571 12370 10597
rect 12394 10571 12410 10597
rect 12410 10571 12422 10597
rect 12342 10570 12370 10571
rect 12394 10570 12422 10571
rect 12446 10597 12474 10598
rect 12446 10571 12472 10597
rect 12472 10571 12474 10597
rect 12446 10570 12474 10571
rect 12498 10597 12526 10598
rect 12498 10571 12508 10597
rect 12508 10571 12526 10597
rect 12498 10570 12526 10571
rect 10542 9254 10570 9282
rect 10318 9225 10346 9226
rect 10318 9199 10319 9225
rect 10319 9199 10345 9225
rect 10345 9199 10346 9225
rect 10318 9198 10346 9199
rect 10486 9225 10514 9226
rect 10486 9199 10487 9225
rect 10487 9199 10513 9225
rect 10513 9199 10514 9225
rect 10486 9198 10514 9199
rect 9582 8637 9610 8638
rect 9582 8611 9600 8637
rect 9600 8611 9610 8637
rect 9582 8610 9610 8611
rect 9634 8637 9662 8638
rect 9634 8611 9636 8637
rect 9636 8611 9662 8637
rect 9634 8610 9662 8611
rect 9686 8637 9714 8638
rect 9738 8637 9766 8638
rect 9686 8611 9698 8637
rect 9698 8611 9714 8637
rect 9738 8611 9760 8637
rect 9760 8611 9766 8637
rect 9686 8610 9714 8611
rect 9738 8610 9766 8611
rect 9790 8610 9818 8638
rect 9842 8637 9870 8638
rect 9894 8637 9922 8638
rect 9842 8611 9848 8637
rect 9848 8611 9870 8637
rect 9894 8611 9910 8637
rect 9910 8611 9922 8637
rect 9842 8610 9870 8611
rect 9894 8610 9922 8611
rect 9946 8637 9974 8638
rect 9946 8611 9972 8637
rect 9972 8611 9974 8637
rect 9946 8610 9974 8611
rect 9998 8637 10026 8638
rect 9998 8611 10008 8637
rect 10008 8611 10026 8637
rect 9998 8610 10026 8611
rect 9814 8441 9842 8442
rect 9814 8415 9815 8441
rect 9815 8415 9841 8441
rect 9841 8415 9842 8441
rect 9814 8414 9842 8415
rect 10038 8414 10066 8442
rect 10150 8022 10178 8050
rect 9582 7853 9610 7854
rect 9582 7827 9600 7853
rect 9600 7827 9610 7853
rect 9582 7826 9610 7827
rect 9634 7853 9662 7854
rect 9634 7827 9636 7853
rect 9636 7827 9662 7853
rect 9634 7826 9662 7827
rect 9686 7853 9714 7854
rect 9738 7853 9766 7854
rect 9686 7827 9698 7853
rect 9698 7827 9714 7853
rect 9738 7827 9760 7853
rect 9760 7827 9766 7853
rect 9686 7826 9714 7827
rect 9738 7826 9766 7827
rect 9790 7826 9818 7854
rect 9842 7853 9870 7854
rect 9894 7853 9922 7854
rect 9842 7827 9848 7853
rect 9848 7827 9870 7853
rect 9894 7827 9910 7853
rect 9910 7827 9922 7853
rect 9842 7826 9870 7827
rect 9894 7826 9922 7827
rect 9946 7853 9974 7854
rect 9946 7827 9972 7853
rect 9972 7827 9974 7853
rect 9946 7826 9974 7827
rect 9998 7853 10026 7854
rect 9998 7827 10008 7853
rect 10008 7827 10026 7853
rect 9998 7826 10026 7827
rect 9254 7518 9282 7546
rect 10318 8022 10346 8050
rect 11998 10038 12026 10066
rect 12502 10038 12530 10066
rect 12950 10038 12978 10066
rect 14238 12390 14266 12418
rect 13342 11774 13370 11802
rect 14294 11046 14322 11074
rect 14582 14125 14610 14126
rect 14582 14099 14600 14125
rect 14600 14099 14610 14125
rect 14582 14098 14610 14099
rect 14634 14125 14662 14126
rect 14634 14099 14636 14125
rect 14636 14099 14662 14125
rect 14634 14098 14662 14099
rect 14686 14125 14714 14126
rect 14738 14125 14766 14126
rect 14686 14099 14698 14125
rect 14698 14099 14714 14125
rect 14738 14099 14760 14125
rect 14760 14099 14766 14125
rect 14686 14098 14714 14099
rect 14738 14098 14766 14099
rect 14790 14098 14818 14126
rect 14842 14125 14870 14126
rect 14894 14125 14922 14126
rect 14842 14099 14848 14125
rect 14848 14099 14870 14125
rect 14894 14099 14910 14125
rect 14910 14099 14922 14125
rect 14842 14098 14870 14099
rect 14894 14098 14922 14099
rect 14946 14125 14974 14126
rect 14946 14099 14972 14125
rect 14972 14099 14974 14125
rect 14946 14098 14974 14099
rect 14998 14125 15026 14126
rect 14998 14099 15008 14125
rect 15008 14099 15026 14125
rect 14998 14098 15026 14099
rect 14582 13341 14610 13342
rect 14582 13315 14600 13341
rect 14600 13315 14610 13341
rect 14582 13314 14610 13315
rect 14634 13341 14662 13342
rect 14634 13315 14636 13341
rect 14636 13315 14662 13341
rect 14634 13314 14662 13315
rect 14686 13341 14714 13342
rect 14738 13341 14766 13342
rect 14686 13315 14698 13341
rect 14698 13315 14714 13341
rect 14738 13315 14760 13341
rect 14760 13315 14766 13341
rect 14686 13314 14714 13315
rect 14738 13314 14766 13315
rect 14790 13314 14818 13342
rect 14842 13341 14870 13342
rect 14894 13341 14922 13342
rect 14842 13315 14848 13341
rect 14848 13315 14870 13341
rect 14894 13315 14910 13341
rect 14910 13315 14922 13341
rect 14842 13314 14870 13315
rect 14894 13314 14922 13315
rect 14946 13341 14974 13342
rect 14946 13315 14972 13341
rect 14972 13315 14974 13341
rect 14946 13314 14974 13315
rect 14998 13341 15026 13342
rect 14998 13315 15008 13341
rect 15008 13315 15026 13341
rect 14998 13314 15026 13315
rect 16478 15022 16506 15050
rect 16478 14686 16506 14714
rect 16534 15078 16562 15106
rect 16366 13902 16394 13930
rect 15470 13454 15498 13482
rect 15862 13481 15890 13482
rect 15862 13455 15863 13481
rect 15863 13455 15889 13481
rect 15889 13455 15890 13481
rect 15862 13454 15890 13455
rect 15302 13145 15330 13146
rect 15302 13119 15303 13145
rect 15303 13119 15329 13145
rect 15329 13119 15330 13145
rect 15302 13118 15330 13119
rect 14406 12417 14434 12418
rect 14406 12391 14407 12417
rect 14407 12391 14433 12417
rect 14433 12391 14434 12417
rect 14406 12390 14434 12391
rect 14582 12557 14610 12558
rect 14582 12531 14600 12557
rect 14600 12531 14610 12557
rect 14582 12530 14610 12531
rect 14634 12557 14662 12558
rect 14634 12531 14636 12557
rect 14636 12531 14662 12557
rect 14634 12530 14662 12531
rect 14686 12557 14714 12558
rect 14738 12557 14766 12558
rect 14686 12531 14698 12557
rect 14698 12531 14714 12557
rect 14738 12531 14760 12557
rect 14760 12531 14766 12557
rect 14686 12530 14714 12531
rect 14738 12530 14766 12531
rect 14790 12530 14818 12558
rect 14842 12557 14870 12558
rect 14894 12557 14922 12558
rect 14842 12531 14848 12557
rect 14848 12531 14870 12557
rect 14894 12531 14910 12557
rect 14910 12531 14922 12557
rect 14842 12530 14870 12531
rect 14894 12530 14922 12531
rect 14946 12557 14974 12558
rect 14946 12531 14972 12557
rect 14972 12531 14974 12557
rect 14946 12530 14974 12531
rect 14998 12557 15026 12558
rect 14998 12531 15008 12557
rect 15008 12531 15026 12557
rect 14998 12530 15026 12531
rect 14582 11773 14610 11774
rect 14582 11747 14600 11773
rect 14600 11747 14610 11773
rect 14582 11746 14610 11747
rect 14634 11773 14662 11774
rect 14634 11747 14636 11773
rect 14636 11747 14662 11773
rect 14634 11746 14662 11747
rect 14686 11773 14714 11774
rect 14738 11773 14766 11774
rect 14686 11747 14698 11773
rect 14698 11747 14714 11773
rect 14738 11747 14760 11773
rect 14760 11747 14766 11773
rect 14686 11746 14714 11747
rect 14738 11746 14766 11747
rect 14790 11746 14818 11774
rect 14842 11773 14870 11774
rect 14894 11773 14922 11774
rect 14842 11747 14848 11773
rect 14848 11747 14870 11773
rect 14894 11747 14910 11773
rect 14910 11747 14922 11773
rect 14842 11746 14870 11747
rect 14894 11746 14922 11747
rect 14946 11773 14974 11774
rect 14946 11747 14972 11773
rect 14972 11747 14974 11773
rect 14946 11746 14974 11747
rect 14998 11773 15026 11774
rect 14998 11747 15008 11773
rect 15008 11747 15026 11773
rect 14998 11746 15026 11747
rect 15078 11718 15106 11746
rect 14462 11046 14490 11074
rect 14582 10989 14610 10990
rect 14582 10963 14600 10989
rect 14600 10963 14610 10989
rect 14582 10962 14610 10963
rect 14634 10989 14662 10990
rect 14634 10963 14636 10989
rect 14636 10963 14662 10989
rect 14634 10962 14662 10963
rect 14686 10989 14714 10990
rect 14738 10989 14766 10990
rect 14686 10963 14698 10989
rect 14698 10963 14714 10989
rect 14738 10963 14760 10989
rect 14760 10963 14766 10989
rect 14686 10962 14714 10963
rect 14738 10962 14766 10963
rect 14790 10962 14818 10990
rect 14842 10989 14870 10990
rect 14894 10989 14922 10990
rect 14842 10963 14848 10989
rect 14848 10963 14870 10989
rect 14894 10963 14910 10989
rect 14910 10963 14922 10989
rect 14842 10962 14870 10963
rect 14894 10962 14922 10963
rect 14946 10989 14974 10990
rect 14946 10963 14972 10989
rect 14972 10963 14974 10989
rect 14946 10962 14974 10963
rect 14998 10989 15026 10990
rect 14998 10963 15008 10989
rect 15008 10963 15026 10989
rect 14998 10962 15026 10963
rect 14582 10205 14610 10206
rect 14582 10179 14600 10205
rect 14600 10179 14610 10205
rect 14582 10178 14610 10179
rect 14634 10205 14662 10206
rect 14634 10179 14636 10205
rect 14636 10179 14662 10205
rect 14634 10178 14662 10179
rect 14686 10205 14714 10206
rect 14738 10205 14766 10206
rect 14686 10179 14698 10205
rect 14698 10179 14714 10205
rect 14738 10179 14760 10205
rect 14760 10179 14766 10205
rect 14686 10178 14714 10179
rect 14738 10178 14766 10179
rect 14790 10178 14818 10206
rect 14842 10205 14870 10206
rect 14894 10205 14922 10206
rect 14842 10179 14848 10205
rect 14848 10179 14870 10205
rect 14894 10179 14910 10205
rect 14910 10179 14922 10205
rect 14842 10178 14870 10179
rect 14894 10178 14922 10179
rect 14946 10205 14974 10206
rect 14946 10179 14972 10205
rect 14972 10179 14974 10205
rect 14946 10178 14974 10179
rect 14998 10205 15026 10206
rect 14998 10179 15008 10205
rect 15008 10179 15026 10205
rect 14998 10178 15026 10179
rect 13342 9982 13370 10010
rect 12082 9813 12110 9814
rect 12082 9787 12100 9813
rect 12100 9787 12110 9813
rect 12082 9786 12110 9787
rect 12134 9813 12162 9814
rect 12134 9787 12136 9813
rect 12136 9787 12162 9813
rect 12134 9786 12162 9787
rect 12186 9813 12214 9814
rect 12238 9813 12266 9814
rect 12186 9787 12198 9813
rect 12198 9787 12214 9813
rect 12238 9787 12260 9813
rect 12260 9787 12266 9813
rect 12186 9786 12214 9787
rect 12238 9786 12266 9787
rect 12290 9786 12318 9814
rect 12342 9813 12370 9814
rect 12394 9813 12422 9814
rect 12342 9787 12348 9813
rect 12348 9787 12370 9813
rect 12394 9787 12410 9813
rect 12410 9787 12422 9813
rect 12342 9786 12370 9787
rect 12394 9786 12422 9787
rect 12446 9813 12474 9814
rect 12446 9787 12472 9813
rect 12472 9787 12474 9813
rect 12446 9786 12474 9787
rect 12498 9813 12526 9814
rect 12498 9787 12508 9813
rect 12508 9787 12526 9813
rect 12498 9786 12526 9787
rect 13622 10009 13650 10010
rect 13622 9983 13623 10009
rect 13623 9983 13649 10009
rect 13649 9983 13650 10009
rect 13622 9982 13650 9983
rect 11774 9254 11802 9282
rect 11942 9254 11970 9282
rect 13342 9254 13370 9282
rect 14014 9310 14042 9338
rect 12082 9029 12110 9030
rect 12082 9003 12100 9029
rect 12100 9003 12110 9029
rect 12082 9002 12110 9003
rect 12134 9029 12162 9030
rect 12134 9003 12136 9029
rect 12136 9003 12162 9029
rect 12134 9002 12162 9003
rect 12186 9029 12214 9030
rect 12238 9029 12266 9030
rect 12186 9003 12198 9029
rect 12198 9003 12214 9029
rect 12238 9003 12260 9029
rect 12260 9003 12266 9029
rect 12186 9002 12214 9003
rect 12238 9002 12266 9003
rect 12290 9002 12318 9030
rect 12342 9029 12370 9030
rect 12394 9029 12422 9030
rect 12342 9003 12348 9029
rect 12348 9003 12370 9029
rect 12394 9003 12410 9029
rect 12410 9003 12422 9029
rect 12342 9002 12370 9003
rect 12394 9002 12422 9003
rect 12446 9029 12474 9030
rect 12446 9003 12472 9029
rect 12472 9003 12474 9029
rect 12446 9002 12474 9003
rect 12498 9029 12526 9030
rect 12498 9003 12508 9029
rect 12508 9003 12526 9029
rect 12498 9002 12526 9003
rect 11438 8441 11466 8442
rect 11438 8415 11439 8441
rect 11439 8415 11465 8441
rect 11465 8415 11466 8441
rect 11438 8414 11466 8415
rect 10542 7966 10570 7994
rect 10206 7574 10234 7602
rect 9582 7069 9610 7070
rect 9582 7043 9600 7069
rect 9600 7043 9610 7069
rect 9582 7042 9610 7043
rect 9634 7069 9662 7070
rect 9634 7043 9636 7069
rect 9636 7043 9662 7069
rect 9634 7042 9662 7043
rect 9686 7069 9714 7070
rect 9738 7069 9766 7070
rect 9686 7043 9698 7069
rect 9698 7043 9714 7069
rect 9738 7043 9760 7069
rect 9760 7043 9766 7069
rect 9686 7042 9714 7043
rect 9738 7042 9766 7043
rect 9790 7042 9818 7070
rect 9842 7069 9870 7070
rect 9894 7069 9922 7070
rect 9842 7043 9848 7069
rect 9848 7043 9870 7069
rect 9894 7043 9910 7069
rect 9910 7043 9922 7069
rect 9842 7042 9870 7043
rect 9894 7042 9922 7043
rect 9946 7069 9974 7070
rect 9946 7043 9972 7069
rect 9972 7043 9974 7069
rect 9946 7042 9974 7043
rect 9998 7069 10026 7070
rect 9998 7043 10008 7069
rect 10008 7043 10026 7069
rect 9998 7042 10026 7043
rect 10374 6678 10402 6706
rect 9582 6285 9610 6286
rect 9582 6259 9600 6285
rect 9600 6259 9610 6285
rect 9582 6258 9610 6259
rect 9634 6285 9662 6286
rect 9634 6259 9636 6285
rect 9636 6259 9662 6285
rect 9634 6258 9662 6259
rect 9686 6285 9714 6286
rect 9738 6285 9766 6286
rect 9686 6259 9698 6285
rect 9698 6259 9714 6285
rect 9738 6259 9760 6285
rect 9760 6259 9766 6285
rect 9686 6258 9714 6259
rect 9738 6258 9766 6259
rect 9790 6258 9818 6286
rect 9842 6285 9870 6286
rect 9894 6285 9922 6286
rect 9842 6259 9848 6285
rect 9848 6259 9870 6285
rect 9894 6259 9910 6285
rect 9910 6259 9922 6285
rect 9842 6258 9870 6259
rect 9894 6258 9922 6259
rect 9946 6285 9974 6286
rect 9946 6259 9972 6285
rect 9972 6259 9974 6285
rect 9946 6258 9974 6259
rect 9998 6285 10026 6286
rect 9998 6259 10008 6285
rect 10008 6259 10026 6285
rect 9998 6258 10026 6259
rect 9534 5838 9562 5866
rect 10038 5838 10066 5866
rect 9582 5501 9610 5502
rect 9582 5475 9600 5501
rect 9600 5475 9610 5501
rect 9582 5474 9610 5475
rect 9634 5501 9662 5502
rect 9634 5475 9636 5501
rect 9636 5475 9662 5501
rect 9634 5474 9662 5475
rect 9686 5501 9714 5502
rect 9738 5501 9766 5502
rect 9686 5475 9698 5501
rect 9698 5475 9714 5501
rect 9738 5475 9760 5501
rect 9760 5475 9766 5501
rect 9686 5474 9714 5475
rect 9738 5474 9766 5475
rect 9790 5474 9818 5502
rect 9842 5501 9870 5502
rect 9894 5501 9922 5502
rect 9842 5475 9848 5501
rect 9848 5475 9870 5501
rect 9894 5475 9910 5501
rect 9910 5475 9922 5501
rect 9842 5474 9870 5475
rect 9894 5474 9922 5475
rect 9946 5501 9974 5502
rect 9946 5475 9972 5501
rect 9972 5475 9974 5501
rect 9946 5474 9974 5475
rect 9998 5501 10026 5502
rect 9998 5475 10008 5501
rect 10008 5475 10026 5501
rect 9998 5474 10026 5475
rect 9534 5278 9562 5306
rect 9814 5305 9842 5306
rect 9814 5279 9815 5305
rect 9815 5279 9841 5305
rect 9841 5279 9842 5305
rect 9814 5278 9842 5279
rect 10038 5222 10066 5250
rect 9582 4717 9610 4718
rect 9582 4691 9600 4717
rect 9600 4691 9610 4717
rect 9582 4690 9610 4691
rect 9634 4717 9662 4718
rect 9634 4691 9636 4717
rect 9636 4691 9662 4717
rect 9634 4690 9662 4691
rect 9686 4717 9714 4718
rect 9738 4717 9766 4718
rect 9686 4691 9698 4717
rect 9698 4691 9714 4717
rect 9738 4691 9760 4717
rect 9760 4691 9766 4717
rect 9686 4690 9714 4691
rect 9738 4690 9766 4691
rect 9790 4690 9818 4718
rect 9842 4717 9870 4718
rect 9894 4717 9922 4718
rect 9842 4691 9848 4717
rect 9848 4691 9870 4717
rect 9894 4691 9910 4717
rect 9910 4691 9922 4717
rect 9842 4690 9870 4691
rect 9894 4690 9922 4691
rect 9946 4717 9974 4718
rect 9946 4691 9972 4717
rect 9972 4691 9974 4717
rect 9946 4690 9974 4691
rect 9998 4717 10026 4718
rect 9998 4691 10008 4717
rect 10008 4691 10026 4717
rect 9998 4690 10026 4691
rect 9030 4494 9058 4522
rect 8806 3766 8834 3794
rect 8470 3737 8498 3738
rect 8470 3711 8471 3737
rect 8471 3711 8497 3737
rect 8497 3711 8498 3737
rect 8470 3710 8498 3711
rect 8974 3710 9002 3738
rect 8022 3430 8050 3458
rect 8302 3430 8330 3458
rect 8974 3374 9002 3402
rect 7082 2757 7110 2758
rect 7082 2731 7100 2757
rect 7100 2731 7110 2757
rect 7082 2730 7110 2731
rect 7134 2757 7162 2758
rect 7134 2731 7136 2757
rect 7136 2731 7162 2757
rect 7134 2730 7162 2731
rect 7186 2757 7214 2758
rect 7238 2757 7266 2758
rect 7186 2731 7198 2757
rect 7198 2731 7214 2757
rect 7238 2731 7260 2757
rect 7260 2731 7266 2757
rect 7186 2730 7214 2731
rect 7238 2730 7266 2731
rect 7290 2730 7318 2758
rect 7342 2757 7370 2758
rect 7394 2757 7422 2758
rect 7342 2731 7348 2757
rect 7348 2731 7370 2757
rect 7394 2731 7410 2757
rect 7410 2731 7422 2757
rect 7342 2730 7370 2731
rect 7394 2730 7422 2731
rect 7446 2757 7474 2758
rect 7446 2731 7472 2757
rect 7472 2731 7474 2757
rect 7446 2730 7474 2731
rect 7498 2757 7526 2758
rect 7498 2731 7508 2757
rect 7508 2731 7526 2757
rect 7498 2730 7526 2731
rect 7014 2534 7042 2562
rect 7574 2534 7602 2562
rect 8078 2561 8106 2562
rect 8078 2535 8079 2561
rect 8079 2535 8105 2561
rect 8105 2535 8106 2561
rect 8078 2534 8106 2535
rect 8470 2478 8498 2506
rect 10262 4521 10290 4522
rect 10262 4495 10263 4521
rect 10263 4495 10289 4521
rect 10289 4495 10290 4521
rect 10262 4494 10290 4495
rect 10486 4521 10514 4522
rect 10486 4495 10487 4521
rect 10487 4495 10513 4521
rect 10513 4495 10514 4521
rect 10486 4494 10514 4495
rect 9582 3933 9610 3934
rect 9582 3907 9600 3933
rect 9600 3907 9610 3933
rect 9582 3906 9610 3907
rect 9634 3933 9662 3934
rect 9634 3907 9636 3933
rect 9636 3907 9662 3933
rect 9634 3906 9662 3907
rect 9686 3933 9714 3934
rect 9738 3933 9766 3934
rect 9686 3907 9698 3933
rect 9698 3907 9714 3933
rect 9738 3907 9760 3933
rect 9760 3907 9766 3933
rect 9686 3906 9714 3907
rect 9738 3906 9766 3907
rect 9790 3906 9818 3934
rect 9842 3933 9870 3934
rect 9894 3933 9922 3934
rect 9842 3907 9848 3933
rect 9848 3907 9870 3933
rect 9894 3907 9910 3933
rect 9910 3907 9922 3933
rect 9842 3906 9870 3907
rect 9894 3906 9922 3907
rect 9946 3933 9974 3934
rect 9946 3907 9972 3933
rect 9972 3907 9974 3933
rect 9946 3906 9974 3907
rect 9998 3933 10026 3934
rect 9998 3907 10008 3933
rect 10008 3907 10026 3933
rect 9998 3906 10026 3907
rect 9478 3710 9506 3738
rect 9814 3737 9842 3738
rect 9814 3711 9815 3737
rect 9815 3711 9841 3737
rect 9841 3711 9842 3737
rect 9814 3710 9842 3711
rect 10486 3710 10514 3738
rect 9478 3374 9506 3402
rect 10486 3430 10514 3458
rect 9366 2534 9394 2562
rect 8974 2505 9002 2506
rect 8974 2479 8975 2505
rect 8975 2479 9001 2505
rect 9001 2479 9002 2505
rect 8974 2478 9002 2479
rect 8246 2254 8274 2282
rect 7014 2030 7042 2058
rect 7518 2030 7546 2058
rect 7082 1973 7110 1974
rect 7082 1947 7100 1973
rect 7100 1947 7110 1973
rect 7082 1946 7110 1947
rect 7134 1973 7162 1974
rect 7134 1947 7136 1973
rect 7136 1947 7162 1973
rect 7134 1946 7162 1947
rect 7186 1973 7214 1974
rect 7238 1973 7266 1974
rect 7186 1947 7198 1973
rect 7198 1947 7214 1973
rect 7238 1947 7260 1973
rect 7260 1947 7266 1973
rect 7186 1946 7214 1947
rect 7238 1946 7266 1947
rect 7290 1946 7318 1974
rect 7342 1973 7370 1974
rect 7394 1973 7422 1974
rect 7342 1947 7348 1973
rect 7348 1947 7370 1973
rect 7394 1947 7410 1973
rect 7410 1947 7422 1973
rect 7342 1946 7370 1947
rect 7394 1946 7422 1947
rect 7446 1973 7474 1974
rect 7446 1947 7472 1973
rect 7472 1947 7474 1973
rect 7446 1946 7474 1947
rect 7498 1973 7526 1974
rect 7498 1947 7508 1973
rect 7508 1947 7526 1973
rect 7498 1946 7526 1947
rect 7462 1862 7490 1890
rect 8974 1750 9002 1778
rect 9582 3149 9610 3150
rect 9582 3123 9600 3149
rect 9600 3123 9610 3149
rect 9582 3122 9610 3123
rect 9634 3149 9662 3150
rect 9634 3123 9636 3149
rect 9636 3123 9662 3149
rect 9634 3122 9662 3123
rect 9686 3149 9714 3150
rect 9738 3149 9766 3150
rect 9686 3123 9698 3149
rect 9698 3123 9714 3149
rect 9738 3123 9760 3149
rect 9760 3123 9766 3149
rect 9686 3122 9714 3123
rect 9738 3122 9766 3123
rect 9790 3122 9818 3150
rect 9842 3149 9870 3150
rect 9894 3149 9922 3150
rect 9842 3123 9848 3149
rect 9848 3123 9870 3149
rect 9894 3123 9910 3149
rect 9910 3123 9922 3149
rect 9842 3122 9870 3123
rect 9894 3122 9922 3123
rect 9946 3149 9974 3150
rect 9946 3123 9972 3149
rect 9972 3123 9974 3149
rect 9946 3122 9974 3123
rect 9998 3149 10026 3150
rect 9998 3123 10008 3149
rect 10008 3123 10026 3149
rect 9998 3122 10026 3123
rect 9366 1806 9394 1834
rect 9422 2422 9450 2450
rect 8358 1721 8386 1722
rect 8358 1695 8359 1721
rect 8359 1695 8385 1721
rect 8385 1695 8386 1721
rect 8358 1694 8386 1695
rect 9582 2365 9610 2366
rect 9582 2339 9600 2365
rect 9600 2339 9610 2365
rect 9582 2338 9610 2339
rect 9634 2365 9662 2366
rect 9634 2339 9636 2365
rect 9636 2339 9662 2365
rect 9634 2338 9662 2339
rect 9686 2365 9714 2366
rect 9738 2365 9766 2366
rect 9686 2339 9698 2365
rect 9698 2339 9714 2365
rect 9738 2339 9760 2365
rect 9760 2339 9766 2365
rect 9686 2338 9714 2339
rect 9738 2338 9766 2339
rect 9790 2338 9818 2366
rect 9842 2365 9870 2366
rect 9894 2365 9922 2366
rect 9842 2339 9848 2365
rect 9848 2339 9870 2365
rect 9894 2339 9910 2365
rect 9910 2339 9922 2365
rect 9842 2338 9870 2339
rect 9894 2338 9922 2339
rect 9946 2365 9974 2366
rect 9946 2339 9972 2365
rect 9972 2339 9974 2365
rect 9946 2338 9974 2339
rect 9998 2365 10026 2366
rect 9998 2339 10008 2365
rect 10008 2339 10026 2365
rect 9998 2338 10026 2339
rect 9478 2198 9506 2226
rect 10038 2198 10066 2226
rect 12082 8245 12110 8246
rect 12082 8219 12100 8245
rect 12100 8219 12110 8245
rect 12082 8218 12110 8219
rect 12134 8245 12162 8246
rect 12134 8219 12136 8245
rect 12136 8219 12162 8245
rect 12134 8218 12162 8219
rect 12186 8245 12214 8246
rect 12238 8245 12266 8246
rect 12186 8219 12198 8245
rect 12198 8219 12214 8245
rect 12238 8219 12260 8245
rect 12260 8219 12266 8245
rect 12186 8218 12214 8219
rect 12238 8218 12266 8219
rect 12290 8218 12318 8246
rect 12342 8245 12370 8246
rect 12394 8245 12422 8246
rect 12342 8219 12348 8245
rect 12348 8219 12370 8245
rect 12394 8219 12410 8245
rect 12410 8219 12422 8245
rect 12342 8218 12370 8219
rect 12394 8218 12422 8219
rect 12446 8245 12474 8246
rect 12446 8219 12472 8245
rect 12472 8219 12474 8245
rect 12446 8218 12474 8219
rect 12498 8245 12526 8246
rect 12498 8219 12508 8245
rect 12508 8219 12526 8245
rect 12498 8218 12526 8219
rect 15862 11046 15890 11074
rect 14406 8414 14434 8442
rect 12082 7461 12110 7462
rect 12082 7435 12100 7461
rect 12100 7435 12110 7461
rect 12082 7434 12110 7435
rect 12134 7461 12162 7462
rect 12134 7435 12136 7461
rect 12136 7435 12162 7461
rect 12134 7434 12162 7435
rect 12186 7461 12214 7462
rect 12238 7461 12266 7462
rect 12186 7435 12198 7461
rect 12198 7435 12214 7461
rect 12238 7435 12260 7461
rect 12260 7435 12266 7461
rect 12186 7434 12214 7435
rect 12238 7434 12266 7435
rect 12290 7434 12318 7462
rect 12342 7461 12370 7462
rect 12394 7461 12422 7462
rect 12342 7435 12348 7461
rect 12348 7435 12370 7461
rect 12394 7435 12410 7461
rect 12410 7435 12422 7461
rect 12342 7434 12370 7435
rect 12394 7434 12422 7435
rect 12446 7461 12474 7462
rect 12446 7435 12472 7461
rect 12472 7435 12474 7461
rect 12446 7434 12474 7435
rect 12498 7461 12526 7462
rect 12498 7435 12508 7461
rect 12508 7435 12526 7461
rect 12498 7434 12526 7435
rect 11998 7238 12026 7266
rect 11830 6678 11858 6706
rect 12082 6677 12110 6678
rect 12082 6651 12100 6677
rect 12100 6651 12110 6677
rect 12082 6650 12110 6651
rect 12134 6677 12162 6678
rect 12134 6651 12136 6677
rect 12136 6651 12162 6677
rect 12134 6650 12162 6651
rect 12186 6677 12214 6678
rect 12238 6677 12266 6678
rect 12186 6651 12198 6677
rect 12198 6651 12214 6677
rect 12238 6651 12260 6677
rect 12260 6651 12266 6677
rect 12186 6650 12214 6651
rect 12238 6650 12266 6651
rect 12290 6650 12318 6678
rect 12342 6677 12370 6678
rect 12394 6677 12422 6678
rect 12342 6651 12348 6677
rect 12348 6651 12370 6677
rect 12394 6651 12410 6677
rect 12410 6651 12422 6677
rect 12342 6650 12370 6651
rect 12394 6650 12422 6651
rect 12446 6677 12474 6678
rect 12446 6651 12472 6677
rect 12472 6651 12474 6677
rect 12446 6650 12474 6651
rect 12498 6677 12526 6678
rect 12498 6651 12508 6677
rect 12508 6651 12526 6677
rect 12498 6650 12526 6651
rect 11550 5838 11578 5866
rect 11550 5614 11578 5642
rect 11942 5670 11970 5698
rect 11550 5222 11578 5250
rect 11774 4521 11802 4522
rect 11774 4495 11775 4521
rect 11775 4495 11801 4521
rect 11801 4495 11802 4521
rect 11774 4494 11802 4495
rect 12082 5893 12110 5894
rect 12082 5867 12100 5893
rect 12100 5867 12110 5893
rect 12082 5866 12110 5867
rect 12134 5893 12162 5894
rect 12134 5867 12136 5893
rect 12136 5867 12162 5893
rect 12134 5866 12162 5867
rect 12186 5893 12214 5894
rect 12238 5893 12266 5894
rect 12186 5867 12198 5893
rect 12198 5867 12214 5893
rect 12238 5867 12260 5893
rect 12260 5867 12266 5893
rect 12186 5866 12214 5867
rect 12238 5866 12266 5867
rect 12290 5866 12318 5894
rect 12342 5893 12370 5894
rect 12394 5893 12422 5894
rect 12342 5867 12348 5893
rect 12348 5867 12370 5893
rect 12394 5867 12410 5893
rect 12410 5867 12422 5893
rect 12342 5866 12370 5867
rect 12394 5866 12422 5867
rect 12446 5893 12474 5894
rect 12446 5867 12472 5893
rect 12472 5867 12474 5893
rect 12446 5866 12474 5867
rect 12498 5893 12526 5894
rect 12498 5867 12508 5893
rect 12508 5867 12526 5893
rect 12498 5866 12526 5867
rect 12502 5697 12530 5698
rect 12502 5671 12503 5697
rect 12503 5671 12529 5697
rect 12529 5671 12530 5697
rect 12502 5670 12530 5671
rect 12726 5697 12754 5698
rect 12726 5671 12727 5697
rect 12727 5671 12753 5697
rect 12753 5671 12754 5697
rect 12726 5670 12754 5671
rect 12334 5614 12362 5642
rect 12614 5614 12642 5642
rect 12082 5109 12110 5110
rect 12082 5083 12100 5109
rect 12100 5083 12110 5109
rect 12082 5082 12110 5083
rect 12134 5109 12162 5110
rect 12134 5083 12136 5109
rect 12136 5083 12162 5109
rect 12134 5082 12162 5083
rect 12186 5109 12214 5110
rect 12238 5109 12266 5110
rect 12186 5083 12198 5109
rect 12198 5083 12214 5109
rect 12238 5083 12260 5109
rect 12260 5083 12266 5109
rect 12186 5082 12214 5083
rect 12238 5082 12266 5083
rect 12290 5082 12318 5110
rect 12342 5109 12370 5110
rect 12394 5109 12422 5110
rect 12342 5083 12348 5109
rect 12348 5083 12370 5109
rect 12394 5083 12410 5109
rect 12410 5083 12422 5109
rect 12342 5082 12370 5083
rect 12394 5082 12422 5083
rect 12446 5109 12474 5110
rect 12446 5083 12472 5109
rect 12472 5083 12474 5109
rect 12446 5082 12474 5083
rect 12498 5109 12526 5110
rect 12498 5083 12508 5109
rect 12508 5083 12526 5109
rect 12498 5082 12526 5083
rect 11942 4521 11970 4522
rect 11942 4495 11943 4521
rect 11943 4495 11969 4521
rect 11969 4495 11970 4521
rect 11942 4494 11970 4495
rect 12726 5278 12754 5306
rect 11382 4214 11410 4242
rect 10878 3737 10906 3738
rect 10878 3711 10879 3737
rect 10879 3711 10905 3737
rect 10905 3711 10906 3737
rect 10878 3710 10906 3711
rect 10542 2086 10570 2114
rect 11774 3710 11802 3738
rect 12082 4325 12110 4326
rect 12082 4299 12100 4325
rect 12100 4299 12110 4325
rect 12082 4298 12110 4299
rect 12134 4325 12162 4326
rect 12134 4299 12136 4325
rect 12136 4299 12162 4325
rect 12134 4298 12162 4299
rect 12186 4325 12214 4326
rect 12238 4325 12266 4326
rect 12186 4299 12198 4325
rect 12198 4299 12214 4325
rect 12238 4299 12260 4325
rect 12260 4299 12266 4325
rect 12186 4298 12214 4299
rect 12238 4298 12266 4299
rect 12290 4298 12318 4326
rect 12342 4325 12370 4326
rect 12394 4325 12422 4326
rect 12342 4299 12348 4325
rect 12348 4299 12370 4325
rect 12394 4299 12410 4325
rect 12410 4299 12422 4325
rect 12342 4298 12370 4299
rect 12394 4298 12422 4299
rect 12446 4325 12474 4326
rect 12446 4299 12472 4325
rect 12472 4299 12474 4325
rect 12446 4298 12474 4299
rect 12498 4325 12526 4326
rect 12498 4299 12508 4325
rect 12508 4299 12526 4325
rect 12498 4298 12526 4299
rect 11998 4214 12026 4242
rect 11942 3318 11970 3346
rect 12082 3541 12110 3542
rect 12082 3515 12100 3541
rect 12100 3515 12110 3541
rect 12082 3514 12110 3515
rect 12134 3541 12162 3542
rect 12134 3515 12136 3541
rect 12136 3515 12162 3541
rect 12134 3514 12162 3515
rect 12186 3541 12214 3542
rect 12238 3541 12266 3542
rect 12186 3515 12198 3541
rect 12198 3515 12214 3541
rect 12238 3515 12260 3541
rect 12260 3515 12266 3541
rect 12186 3514 12214 3515
rect 12238 3514 12266 3515
rect 12290 3514 12318 3542
rect 12342 3541 12370 3542
rect 12394 3541 12422 3542
rect 12342 3515 12348 3541
rect 12348 3515 12370 3541
rect 12394 3515 12410 3541
rect 12410 3515 12422 3541
rect 12342 3514 12370 3515
rect 12394 3514 12422 3515
rect 12446 3541 12474 3542
rect 12446 3515 12472 3541
rect 12472 3515 12474 3541
rect 12446 3514 12474 3515
rect 12498 3541 12526 3542
rect 12498 3515 12508 3541
rect 12508 3515 12526 3541
rect 12498 3514 12526 3515
rect 11774 3262 11802 3290
rect 10878 2142 10906 2170
rect 11382 2169 11410 2170
rect 11382 2143 11383 2169
rect 11383 2143 11409 2169
rect 11409 2143 11410 2169
rect 11382 2142 11410 2143
rect 10822 2086 10850 2114
rect 11382 1806 11410 1834
rect 9702 1777 9730 1778
rect 9702 1751 9703 1777
rect 9703 1751 9729 1777
rect 9729 1751 9730 1777
rect 9702 1750 9730 1751
rect 10710 1750 10738 1778
rect 9582 1581 9610 1582
rect 9582 1555 9600 1581
rect 9600 1555 9610 1581
rect 9582 1554 9610 1555
rect 9634 1581 9662 1582
rect 9634 1555 9636 1581
rect 9636 1555 9662 1581
rect 9634 1554 9662 1555
rect 9686 1581 9714 1582
rect 9738 1581 9766 1582
rect 9686 1555 9698 1581
rect 9698 1555 9714 1581
rect 9738 1555 9760 1581
rect 9760 1555 9766 1581
rect 9686 1554 9714 1555
rect 9738 1554 9766 1555
rect 9790 1554 9818 1582
rect 9842 1581 9870 1582
rect 9894 1581 9922 1582
rect 9842 1555 9848 1581
rect 9848 1555 9870 1581
rect 9894 1555 9910 1581
rect 9910 1555 9922 1581
rect 9842 1554 9870 1555
rect 9894 1554 9922 1555
rect 9946 1581 9974 1582
rect 9946 1555 9972 1581
rect 9972 1555 9974 1581
rect 9946 1554 9974 1555
rect 9998 1581 10026 1582
rect 9998 1555 10008 1581
rect 10008 1555 10026 1581
rect 9998 1554 10026 1555
rect 11774 2169 11802 2170
rect 11774 2143 11775 2169
rect 11775 2143 11801 2169
rect 11801 2143 11802 2169
rect 11774 2142 11802 2143
rect 11942 2169 11970 2170
rect 11942 2143 11943 2169
rect 11943 2143 11969 2169
rect 11969 2143 11970 2169
rect 11942 2142 11970 2143
rect 12334 3345 12362 3346
rect 12334 3319 12335 3345
rect 12335 3319 12361 3345
rect 12361 3319 12362 3345
rect 12334 3318 12362 3319
rect 12446 2953 12474 2954
rect 12446 2927 12447 2953
rect 12447 2927 12473 2953
rect 12473 2927 12474 2953
rect 12446 2926 12474 2927
rect 12082 2757 12110 2758
rect 12082 2731 12100 2757
rect 12100 2731 12110 2757
rect 12082 2730 12110 2731
rect 12134 2757 12162 2758
rect 12134 2731 12136 2757
rect 12136 2731 12162 2757
rect 12134 2730 12162 2731
rect 12186 2757 12214 2758
rect 12238 2757 12266 2758
rect 12186 2731 12198 2757
rect 12198 2731 12214 2757
rect 12238 2731 12260 2757
rect 12260 2731 12266 2757
rect 12186 2730 12214 2731
rect 12238 2730 12266 2731
rect 12290 2730 12318 2758
rect 12342 2757 12370 2758
rect 12394 2757 12422 2758
rect 12342 2731 12348 2757
rect 12348 2731 12370 2757
rect 12394 2731 12410 2757
rect 12410 2731 12422 2757
rect 12342 2730 12370 2731
rect 12394 2730 12422 2731
rect 12446 2757 12474 2758
rect 12446 2731 12472 2757
rect 12472 2731 12474 2757
rect 12446 2730 12474 2731
rect 12498 2757 12526 2758
rect 12498 2731 12508 2757
rect 12508 2731 12526 2757
rect 12498 2730 12526 2731
rect 12082 1973 12110 1974
rect 12082 1947 12100 1973
rect 12100 1947 12110 1973
rect 12082 1946 12110 1947
rect 12134 1973 12162 1974
rect 12134 1947 12136 1973
rect 12136 1947 12162 1973
rect 12134 1946 12162 1947
rect 12186 1973 12214 1974
rect 12238 1973 12266 1974
rect 12186 1947 12198 1973
rect 12198 1947 12214 1973
rect 12238 1947 12260 1973
rect 12260 1947 12266 1973
rect 12186 1946 12214 1947
rect 12238 1946 12266 1947
rect 12290 1946 12318 1974
rect 12342 1973 12370 1974
rect 12394 1973 12422 1974
rect 12342 1947 12348 1973
rect 12348 1947 12370 1973
rect 12394 1947 12410 1973
rect 12410 1947 12422 1973
rect 12342 1946 12370 1947
rect 12394 1946 12422 1947
rect 12446 1973 12474 1974
rect 12446 1947 12472 1973
rect 12472 1947 12474 1973
rect 12446 1946 12474 1947
rect 12498 1973 12526 1974
rect 12498 1947 12508 1973
rect 12508 1947 12526 1973
rect 12498 1946 12526 1947
rect 13118 7265 13146 7266
rect 13118 7239 13119 7265
rect 13119 7239 13145 7265
rect 13145 7239 13146 7265
rect 13118 7238 13146 7239
rect 14462 9590 14490 9618
rect 14798 9617 14826 9618
rect 14798 9591 14799 9617
rect 14799 9591 14825 9617
rect 14825 9591 14826 9617
rect 14798 9590 14826 9591
rect 15078 9590 15106 9618
rect 15750 10038 15778 10066
rect 14582 9421 14610 9422
rect 14582 9395 14600 9421
rect 14600 9395 14610 9421
rect 14582 9394 14610 9395
rect 14634 9421 14662 9422
rect 14634 9395 14636 9421
rect 14636 9395 14662 9421
rect 14634 9394 14662 9395
rect 14686 9421 14714 9422
rect 14738 9421 14766 9422
rect 14686 9395 14698 9421
rect 14698 9395 14714 9421
rect 14738 9395 14760 9421
rect 14760 9395 14766 9421
rect 14686 9394 14714 9395
rect 14738 9394 14766 9395
rect 14790 9394 14818 9422
rect 14842 9421 14870 9422
rect 14894 9421 14922 9422
rect 14842 9395 14848 9421
rect 14848 9395 14870 9421
rect 14894 9395 14910 9421
rect 14910 9395 14922 9421
rect 14842 9394 14870 9395
rect 14894 9394 14922 9395
rect 14946 9421 14974 9422
rect 14946 9395 14972 9421
rect 14972 9395 14974 9421
rect 14946 9394 14974 9395
rect 14998 9421 15026 9422
rect 14998 9395 15008 9421
rect 15008 9395 15026 9421
rect 14998 9394 15026 9395
rect 14462 9254 14490 9282
rect 15750 9590 15778 9618
rect 15134 9310 15162 9338
rect 15862 9590 15890 9618
rect 14582 8637 14610 8638
rect 14582 8611 14600 8637
rect 14600 8611 14610 8637
rect 14582 8610 14610 8611
rect 14634 8637 14662 8638
rect 14634 8611 14636 8637
rect 14636 8611 14662 8637
rect 14634 8610 14662 8611
rect 14686 8637 14714 8638
rect 14738 8637 14766 8638
rect 14686 8611 14698 8637
rect 14698 8611 14714 8637
rect 14738 8611 14760 8637
rect 14760 8611 14766 8637
rect 14686 8610 14714 8611
rect 14738 8610 14766 8611
rect 14790 8610 14818 8638
rect 14842 8637 14870 8638
rect 14894 8637 14922 8638
rect 14842 8611 14848 8637
rect 14848 8611 14870 8637
rect 14894 8611 14910 8637
rect 14910 8611 14922 8637
rect 14842 8610 14870 8611
rect 14894 8610 14922 8611
rect 14946 8637 14974 8638
rect 14946 8611 14972 8637
rect 14972 8611 14974 8637
rect 14946 8610 14974 8611
rect 14998 8637 15026 8638
rect 14998 8611 15008 8637
rect 15008 8611 15026 8637
rect 14998 8610 15026 8611
rect 14966 8414 14994 8442
rect 14582 7853 14610 7854
rect 14582 7827 14600 7853
rect 14600 7827 14610 7853
rect 14582 7826 14610 7827
rect 14634 7853 14662 7854
rect 14634 7827 14636 7853
rect 14636 7827 14662 7853
rect 14634 7826 14662 7827
rect 14686 7853 14714 7854
rect 14738 7853 14766 7854
rect 14686 7827 14698 7853
rect 14698 7827 14714 7853
rect 14738 7827 14760 7853
rect 14760 7827 14766 7853
rect 14686 7826 14714 7827
rect 14738 7826 14766 7827
rect 14790 7826 14818 7854
rect 14842 7853 14870 7854
rect 14894 7853 14922 7854
rect 14842 7827 14848 7853
rect 14848 7827 14870 7853
rect 14894 7827 14910 7853
rect 14910 7827 14922 7853
rect 14842 7826 14870 7827
rect 14894 7826 14922 7827
rect 14946 7853 14974 7854
rect 14946 7827 14972 7853
rect 14972 7827 14974 7853
rect 14946 7826 14974 7827
rect 14998 7853 15026 7854
rect 14998 7827 15008 7853
rect 15008 7827 15026 7853
rect 14998 7826 15026 7827
rect 13454 7265 13482 7266
rect 13454 7239 13455 7265
rect 13455 7239 13481 7265
rect 13481 7239 13482 7265
rect 13454 7238 13482 7239
rect 13118 6902 13146 6930
rect 16254 8414 16282 8442
rect 14582 7069 14610 7070
rect 14582 7043 14600 7069
rect 14600 7043 14610 7069
rect 14582 7042 14610 7043
rect 14634 7069 14662 7070
rect 14634 7043 14636 7069
rect 14636 7043 14662 7069
rect 14634 7042 14662 7043
rect 14686 7069 14714 7070
rect 14738 7069 14766 7070
rect 14686 7043 14698 7069
rect 14698 7043 14714 7069
rect 14738 7043 14760 7069
rect 14760 7043 14766 7069
rect 14686 7042 14714 7043
rect 14738 7042 14766 7043
rect 14790 7042 14818 7070
rect 14842 7069 14870 7070
rect 14894 7069 14922 7070
rect 14842 7043 14848 7069
rect 14848 7043 14870 7069
rect 14894 7043 14910 7069
rect 14910 7043 14922 7069
rect 14842 7042 14870 7043
rect 14894 7042 14922 7043
rect 14946 7069 14974 7070
rect 14946 7043 14972 7069
rect 14972 7043 14974 7069
rect 14946 7042 14974 7043
rect 14998 7069 15026 7070
rect 14998 7043 15008 7069
rect 15008 7043 15026 7069
rect 14998 7042 15026 7043
rect 14406 6902 14434 6930
rect 13510 6873 13538 6874
rect 13510 6847 13511 6873
rect 13511 6847 13537 6873
rect 13537 6847 13538 6873
rect 13510 6846 13538 6847
rect 15134 6873 15162 6874
rect 15134 6847 15135 6873
rect 15135 6847 15161 6873
rect 15161 6847 15162 6873
rect 15134 6846 15162 6847
rect 15246 6846 15274 6874
rect 13118 5614 13146 5642
rect 15750 6481 15778 6482
rect 15750 6455 15751 6481
rect 15751 6455 15777 6481
rect 15777 6455 15778 6481
rect 15750 6454 15778 6455
rect 14582 6285 14610 6286
rect 14582 6259 14600 6285
rect 14600 6259 14610 6285
rect 14582 6258 14610 6259
rect 14634 6285 14662 6286
rect 14634 6259 14636 6285
rect 14636 6259 14662 6285
rect 14634 6258 14662 6259
rect 14686 6285 14714 6286
rect 14738 6285 14766 6286
rect 14686 6259 14698 6285
rect 14698 6259 14714 6285
rect 14738 6259 14760 6285
rect 14760 6259 14766 6285
rect 14686 6258 14714 6259
rect 14738 6258 14766 6259
rect 14790 6258 14818 6286
rect 14842 6285 14870 6286
rect 14894 6285 14922 6286
rect 14842 6259 14848 6285
rect 14848 6259 14870 6285
rect 14894 6259 14910 6285
rect 14910 6259 14922 6285
rect 14842 6258 14870 6259
rect 14894 6258 14922 6259
rect 14946 6285 14974 6286
rect 14946 6259 14972 6285
rect 14972 6259 14974 6285
rect 14946 6258 14974 6259
rect 14998 6285 15026 6286
rect 14998 6259 15008 6285
rect 15008 6259 15026 6285
rect 14998 6258 15026 6259
rect 14582 5501 14610 5502
rect 14582 5475 14600 5501
rect 14600 5475 14610 5501
rect 14582 5474 14610 5475
rect 14634 5501 14662 5502
rect 14634 5475 14636 5501
rect 14636 5475 14662 5501
rect 14634 5474 14662 5475
rect 14686 5501 14714 5502
rect 14738 5501 14766 5502
rect 14686 5475 14698 5501
rect 14698 5475 14714 5501
rect 14738 5475 14760 5501
rect 14760 5475 14766 5501
rect 14686 5474 14714 5475
rect 14738 5474 14766 5475
rect 14790 5474 14818 5502
rect 14842 5501 14870 5502
rect 14894 5501 14922 5502
rect 14842 5475 14848 5501
rect 14848 5475 14870 5501
rect 14894 5475 14910 5501
rect 14910 5475 14922 5501
rect 14842 5474 14870 5475
rect 14894 5474 14922 5475
rect 14946 5501 14974 5502
rect 14946 5475 14972 5501
rect 14972 5475 14974 5501
rect 14946 5474 14974 5475
rect 14998 5501 15026 5502
rect 14998 5475 15008 5501
rect 15008 5475 15026 5501
rect 14998 5474 15026 5475
rect 13286 5305 13314 5306
rect 13286 5279 13287 5305
rect 13287 5279 13313 5305
rect 13313 5279 13314 5305
rect 13286 5278 13314 5279
rect 13510 5305 13538 5306
rect 13510 5279 13511 5305
rect 13511 5279 13537 5305
rect 13537 5279 13538 5305
rect 13510 5278 13538 5279
rect 14582 4717 14610 4718
rect 14582 4691 14600 4717
rect 14600 4691 14610 4717
rect 14582 4690 14610 4691
rect 14634 4717 14662 4718
rect 14634 4691 14636 4717
rect 14636 4691 14662 4717
rect 14634 4690 14662 4691
rect 14686 4717 14714 4718
rect 14738 4717 14766 4718
rect 14686 4691 14698 4717
rect 14698 4691 14714 4717
rect 14738 4691 14760 4717
rect 14760 4691 14766 4717
rect 14686 4690 14714 4691
rect 14738 4690 14766 4691
rect 14790 4690 14818 4718
rect 14842 4717 14870 4718
rect 14894 4717 14922 4718
rect 14842 4691 14848 4717
rect 14848 4691 14870 4717
rect 14894 4691 14910 4717
rect 14910 4691 14922 4717
rect 14842 4690 14870 4691
rect 14894 4690 14922 4691
rect 14946 4717 14974 4718
rect 14946 4691 14972 4717
rect 14972 4691 14974 4717
rect 14946 4690 14974 4691
rect 14998 4717 15026 4718
rect 14998 4691 15008 4717
rect 15008 4691 15026 4717
rect 14998 4690 15026 4691
rect 12950 4129 12978 4130
rect 12950 4103 12951 4129
rect 12951 4103 12977 4129
rect 12977 4103 12978 4129
rect 12950 4102 12978 4103
rect 13230 4129 13258 4130
rect 13230 4103 13231 4129
rect 13231 4103 13257 4129
rect 13257 4103 13258 4129
rect 13230 4102 13258 4103
rect 13230 3710 13258 3738
rect 13790 3737 13818 3738
rect 13790 3711 13791 3737
rect 13791 3711 13817 3737
rect 13817 3711 13818 3737
rect 13790 3710 13818 3711
rect 14070 3710 14098 3738
rect 14070 3374 14098 3402
rect 13174 2926 13202 2954
rect 16534 13537 16562 13538
rect 16534 13511 16535 13537
rect 16535 13511 16561 13537
rect 16561 13511 16562 13537
rect 16534 13510 16562 13511
rect 16534 11718 16562 11746
rect 16814 10401 16842 10402
rect 16814 10375 16815 10401
rect 16815 10375 16841 10401
rect 16841 10375 16842 10401
rect 16814 10374 16842 10375
rect 17082 18437 17110 18438
rect 17082 18411 17100 18437
rect 17100 18411 17110 18437
rect 17082 18410 17110 18411
rect 17134 18437 17162 18438
rect 17134 18411 17136 18437
rect 17136 18411 17162 18437
rect 17134 18410 17162 18411
rect 17186 18437 17214 18438
rect 17238 18437 17266 18438
rect 17186 18411 17198 18437
rect 17198 18411 17214 18437
rect 17238 18411 17260 18437
rect 17260 18411 17266 18437
rect 17186 18410 17214 18411
rect 17238 18410 17266 18411
rect 17290 18410 17318 18438
rect 17342 18437 17370 18438
rect 17394 18437 17422 18438
rect 17342 18411 17348 18437
rect 17348 18411 17370 18437
rect 17394 18411 17410 18437
rect 17410 18411 17422 18437
rect 17342 18410 17370 18411
rect 17394 18410 17422 18411
rect 17446 18437 17474 18438
rect 17446 18411 17472 18437
rect 17472 18411 17474 18437
rect 17446 18410 17474 18411
rect 17498 18437 17526 18438
rect 17498 18411 17508 18437
rect 17508 18411 17526 18437
rect 17498 18410 17526 18411
rect 19582 18045 19610 18046
rect 19582 18019 19600 18045
rect 19600 18019 19610 18045
rect 19582 18018 19610 18019
rect 19634 18045 19662 18046
rect 19634 18019 19636 18045
rect 19636 18019 19662 18045
rect 19634 18018 19662 18019
rect 19686 18045 19714 18046
rect 19738 18045 19766 18046
rect 19686 18019 19698 18045
rect 19698 18019 19714 18045
rect 19738 18019 19760 18045
rect 19760 18019 19766 18045
rect 19686 18018 19714 18019
rect 19738 18018 19766 18019
rect 19790 18018 19818 18046
rect 19842 18045 19870 18046
rect 19894 18045 19922 18046
rect 19842 18019 19848 18045
rect 19848 18019 19870 18045
rect 19894 18019 19910 18045
rect 19910 18019 19922 18045
rect 19842 18018 19870 18019
rect 19894 18018 19922 18019
rect 19946 18045 19974 18046
rect 19946 18019 19972 18045
rect 19972 18019 19974 18045
rect 19946 18018 19974 18019
rect 19998 18045 20026 18046
rect 19998 18019 20008 18045
rect 20008 18019 20026 18045
rect 19998 18018 20026 18019
rect 17082 17653 17110 17654
rect 17082 17627 17100 17653
rect 17100 17627 17110 17653
rect 17082 17626 17110 17627
rect 17134 17653 17162 17654
rect 17134 17627 17136 17653
rect 17136 17627 17162 17653
rect 17134 17626 17162 17627
rect 17186 17653 17214 17654
rect 17238 17653 17266 17654
rect 17186 17627 17198 17653
rect 17198 17627 17214 17653
rect 17238 17627 17260 17653
rect 17260 17627 17266 17653
rect 17186 17626 17214 17627
rect 17238 17626 17266 17627
rect 17290 17626 17318 17654
rect 17342 17653 17370 17654
rect 17394 17653 17422 17654
rect 17342 17627 17348 17653
rect 17348 17627 17370 17653
rect 17394 17627 17410 17653
rect 17410 17627 17422 17653
rect 17342 17626 17370 17627
rect 17394 17626 17422 17627
rect 17446 17653 17474 17654
rect 17446 17627 17472 17653
rect 17472 17627 17474 17653
rect 17446 17626 17474 17627
rect 17498 17653 17526 17654
rect 17498 17627 17508 17653
rect 17508 17627 17526 17653
rect 17498 17626 17526 17627
rect 19582 17261 19610 17262
rect 19582 17235 19600 17261
rect 19600 17235 19610 17261
rect 19582 17234 19610 17235
rect 19634 17261 19662 17262
rect 19634 17235 19636 17261
rect 19636 17235 19662 17261
rect 19634 17234 19662 17235
rect 19686 17261 19714 17262
rect 19738 17261 19766 17262
rect 19686 17235 19698 17261
rect 19698 17235 19714 17261
rect 19738 17235 19760 17261
rect 19760 17235 19766 17261
rect 19686 17234 19714 17235
rect 19738 17234 19766 17235
rect 19790 17234 19818 17262
rect 19842 17261 19870 17262
rect 19894 17261 19922 17262
rect 19842 17235 19848 17261
rect 19848 17235 19870 17261
rect 19894 17235 19910 17261
rect 19910 17235 19922 17261
rect 19842 17234 19870 17235
rect 19894 17234 19922 17235
rect 19946 17261 19974 17262
rect 19946 17235 19972 17261
rect 19972 17235 19974 17261
rect 19946 17234 19974 17235
rect 19998 17261 20026 17262
rect 19998 17235 20008 17261
rect 20008 17235 20026 17261
rect 19998 17234 20026 17235
rect 17082 16869 17110 16870
rect 17082 16843 17100 16869
rect 17100 16843 17110 16869
rect 17082 16842 17110 16843
rect 17134 16869 17162 16870
rect 17134 16843 17136 16869
rect 17136 16843 17162 16869
rect 17134 16842 17162 16843
rect 17186 16869 17214 16870
rect 17238 16869 17266 16870
rect 17186 16843 17198 16869
rect 17198 16843 17214 16869
rect 17238 16843 17260 16869
rect 17260 16843 17266 16869
rect 17186 16842 17214 16843
rect 17238 16842 17266 16843
rect 17290 16842 17318 16870
rect 17342 16869 17370 16870
rect 17394 16869 17422 16870
rect 17342 16843 17348 16869
rect 17348 16843 17370 16869
rect 17394 16843 17410 16869
rect 17410 16843 17422 16869
rect 17342 16842 17370 16843
rect 17394 16842 17422 16843
rect 17446 16869 17474 16870
rect 17446 16843 17472 16869
rect 17472 16843 17474 16869
rect 17446 16842 17474 16843
rect 17498 16869 17526 16870
rect 17498 16843 17508 16869
rect 17508 16843 17526 16869
rect 17498 16842 17526 16843
rect 19582 16477 19610 16478
rect 19582 16451 19600 16477
rect 19600 16451 19610 16477
rect 19582 16450 19610 16451
rect 19634 16477 19662 16478
rect 19634 16451 19636 16477
rect 19636 16451 19662 16477
rect 19634 16450 19662 16451
rect 19686 16477 19714 16478
rect 19738 16477 19766 16478
rect 19686 16451 19698 16477
rect 19698 16451 19714 16477
rect 19738 16451 19760 16477
rect 19760 16451 19766 16477
rect 19686 16450 19714 16451
rect 19738 16450 19766 16451
rect 19790 16450 19818 16478
rect 19842 16477 19870 16478
rect 19894 16477 19922 16478
rect 19842 16451 19848 16477
rect 19848 16451 19870 16477
rect 19894 16451 19910 16477
rect 19910 16451 19922 16477
rect 19842 16450 19870 16451
rect 19894 16450 19922 16451
rect 19946 16477 19974 16478
rect 19946 16451 19972 16477
rect 19972 16451 19974 16477
rect 19946 16450 19974 16451
rect 19998 16477 20026 16478
rect 19998 16451 20008 16477
rect 20008 16451 20026 16477
rect 19998 16450 20026 16451
rect 17082 16085 17110 16086
rect 17082 16059 17100 16085
rect 17100 16059 17110 16085
rect 17082 16058 17110 16059
rect 17134 16085 17162 16086
rect 17134 16059 17136 16085
rect 17136 16059 17162 16085
rect 17134 16058 17162 16059
rect 17186 16085 17214 16086
rect 17238 16085 17266 16086
rect 17186 16059 17198 16085
rect 17198 16059 17214 16085
rect 17238 16059 17260 16085
rect 17260 16059 17266 16085
rect 17186 16058 17214 16059
rect 17238 16058 17266 16059
rect 17290 16058 17318 16086
rect 17342 16085 17370 16086
rect 17394 16085 17422 16086
rect 17342 16059 17348 16085
rect 17348 16059 17370 16085
rect 17394 16059 17410 16085
rect 17410 16059 17422 16085
rect 17342 16058 17370 16059
rect 17394 16058 17422 16059
rect 17446 16085 17474 16086
rect 17446 16059 17472 16085
rect 17472 16059 17474 16085
rect 17446 16058 17474 16059
rect 17498 16085 17526 16086
rect 17498 16059 17508 16085
rect 17508 16059 17526 16085
rect 17498 16058 17526 16059
rect 16926 15918 16954 15946
rect 20286 15862 20314 15890
rect 19582 15693 19610 15694
rect 19582 15667 19600 15693
rect 19600 15667 19610 15693
rect 19582 15666 19610 15667
rect 19634 15693 19662 15694
rect 19634 15667 19636 15693
rect 19636 15667 19662 15693
rect 19634 15666 19662 15667
rect 19686 15693 19714 15694
rect 19738 15693 19766 15694
rect 19686 15667 19698 15693
rect 19698 15667 19714 15693
rect 19738 15667 19760 15693
rect 19760 15667 19766 15693
rect 19686 15666 19714 15667
rect 19738 15666 19766 15667
rect 19790 15666 19818 15694
rect 19842 15693 19870 15694
rect 19894 15693 19922 15694
rect 19842 15667 19848 15693
rect 19848 15667 19870 15693
rect 19894 15667 19910 15693
rect 19910 15667 19922 15693
rect 19842 15666 19870 15667
rect 19894 15666 19922 15667
rect 19946 15693 19974 15694
rect 19946 15667 19972 15693
rect 19972 15667 19974 15693
rect 19946 15666 19974 15667
rect 19998 15693 20026 15694
rect 19998 15667 20008 15693
rect 20008 15667 20026 15693
rect 19998 15666 20026 15667
rect 17082 15301 17110 15302
rect 17082 15275 17100 15301
rect 17100 15275 17110 15301
rect 17082 15274 17110 15275
rect 17134 15301 17162 15302
rect 17134 15275 17136 15301
rect 17136 15275 17162 15301
rect 17134 15274 17162 15275
rect 17186 15301 17214 15302
rect 17238 15301 17266 15302
rect 17186 15275 17198 15301
rect 17198 15275 17214 15301
rect 17238 15275 17260 15301
rect 17260 15275 17266 15301
rect 17186 15274 17214 15275
rect 17238 15274 17266 15275
rect 17290 15274 17318 15302
rect 17342 15301 17370 15302
rect 17394 15301 17422 15302
rect 17342 15275 17348 15301
rect 17348 15275 17370 15301
rect 17394 15275 17410 15301
rect 17410 15275 17422 15301
rect 17342 15274 17370 15275
rect 17394 15274 17422 15275
rect 17446 15301 17474 15302
rect 17446 15275 17472 15301
rect 17472 15275 17474 15301
rect 17446 15274 17474 15275
rect 17498 15301 17526 15302
rect 17498 15275 17508 15301
rect 17508 15275 17526 15301
rect 17498 15274 17526 15275
rect 17094 14713 17122 14714
rect 17094 14687 17095 14713
rect 17095 14687 17121 14713
rect 17121 14687 17122 14713
rect 17094 14686 17122 14687
rect 17082 14517 17110 14518
rect 17082 14491 17100 14517
rect 17100 14491 17110 14517
rect 17082 14490 17110 14491
rect 17134 14517 17162 14518
rect 17134 14491 17136 14517
rect 17136 14491 17162 14517
rect 17134 14490 17162 14491
rect 17186 14517 17214 14518
rect 17238 14517 17266 14518
rect 17186 14491 17198 14517
rect 17198 14491 17214 14517
rect 17238 14491 17260 14517
rect 17260 14491 17266 14517
rect 17186 14490 17214 14491
rect 17238 14490 17266 14491
rect 17290 14490 17318 14518
rect 17342 14517 17370 14518
rect 17394 14517 17422 14518
rect 17342 14491 17348 14517
rect 17348 14491 17370 14517
rect 17394 14491 17410 14517
rect 17410 14491 17422 14517
rect 17342 14490 17370 14491
rect 17394 14490 17422 14491
rect 17446 14517 17474 14518
rect 17446 14491 17472 14517
rect 17472 14491 17474 14517
rect 17446 14490 17474 14491
rect 17498 14517 17526 14518
rect 17498 14491 17508 14517
rect 17508 14491 17526 14517
rect 17498 14490 17526 14491
rect 17430 14265 17458 14266
rect 17430 14239 17431 14265
rect 17431 14239 17457 14265
rect 17457 14239 17458 14265
rect 17430 14238 17458 14239
rect 18270 14630 18298 14658
rect 18438 14686 18466 14714
rect 17766 14238 17794 14266
rect 17082 13733 17110 13734
rect 17082 13707 17100 13733
rect 17100 13707 17110 13733
rect 17082 13706 17110 13707
rect 17134 13733 17162 13734
rect 17134 13707 17136 13733
rect 17136 13707 17162 13733
rect 17134 13706 17162 13707
rect 17186 13733 17214 13734
rect 17238 13733 17266 13734
rect 17186 13707 17198 13733
rect 17198 13707 17214 13733
rect 17238 13707 17260 13733
rect 17260 13707 17266 13733
rect 17186 13706 17214 13707
rect 17238 13706 17266 13707
rect 17290 13706 17318 13734
rect 17342 13733 17370 13734
rect 17394 13733 17422 13734
rect 17342 13707 17348 13733
rect 17348 13707 17370 13733
rect 17394 13707 17410 13733
rect 17410 13707 17422 13733
rect 17342 13706 17370 13707
rect 17394 13706 17422 13707
rect 17446 13733 17474 13734
rect 17446 13707 17472 13733
rect 17472 13707 17474 13733
rect 17446 13706 17474 13707
rect 17498 13733 17526 13734
rect 17498 13707 17508 13733
rect 17508 13707 17526 13733
rect 17498 13706 17526 13707
rect 16982 13510 17010 13538
rect 17430 13481 17458 13482
rect 17430 13455 17431 13481
rect 17431 13455 17457 13481
rect 17457 13455 17458 13481
rect 17430 13454 17458 13455
rect 16982 13118 17010 13146
rect 17094 13145 17122 13146
rect 17094 13119 17095 13145
rect 17095 13119 17121 13145
rect 17121 13119 17122 13145
rect 17094 13118 17122 13119
rect 18718 14238 18746 14266
rect 18774 14630 18802 14658
rect 18774 14321 18802 14322
rect 18774 14295 18775 14321
rect 18775 14295 18801 14321
rect 18801 14295 18802 14321
rect 18774 14294 18802 14295
rect 19582 14909 19610 14910
rect 19582 14883 19600 14909
rect 19600 14883 19610 14909
rect 19582 14882 19610 14883
rect 19634 14909 19662 14910
rect 19634 14883 19636 14909
rect 19636 14883 19662 14909
rect 19634 14882 19662 14883
rect 19686 14909 19714 14910
rect 19738 14909 19766 14910
rect 19686 14883 19698 14909
rect 19698 14883 19714 14909
rect 19738 14883 19760 14909
rect 19760 14883 19766 14909
rect 19686 14882 19714 14883
rect 19738 14882 19766 14883
rect 19790 14882 19818 14910
rect 19842 14909 19870 14910
rect 19894 14909 19922 14910
rect 19842 14883 19848 14909
rect 19848 14883 19870 14909
rect 19894 14883 19910 14909
rect 19910 14883 19922 14909
rect 19842 14882 19870 14883
rect 19894 14882 19922 14883
rect 19946 14909 19974 14910
rect 19946 14883 19972 14909
rect 19972 14883 19974 14909
rect 19946 14882 19974 14883
rect 19998 14909 20026 14910
rect 19998 14883 20008 14909
rect 20008 14883 20026 14909
rect 19998 14882 20026 14883
rect 18942 14238 18970 14266
rect 20230 14321 20258 14322
rect 20230 14295 20231 14321
rect 20231 14295 20257 14321
rect 20257 14295 20258 14321
rect 20230 14294 20258 14295
rect 19582 14125 19610 14126
rect 19582 14099 19600 14125
rect 19600 14099 19610 14125
rect 19582 14098 19610 14099
rect 19634 14125 19662 14126
rect 19634 14099 19636 14125
rect 19636 14099 19662 14125
rect 19634 14098 19662 14099
rect 19686 14125 19714 14126
rect 19738 14125 19766 14126
rect 19686 14099 19698 14125
rect 19698 14099 19714 14125
rect 19738 14099 19760 14125
rect 19760 14099 19766 14125
rect 19686 14098 19714 14099
rect 19738 14098 19766 14099
rect 19790 14098 19818 14126
rect 19842 14125 19870 14126
rect 19894 14125 19922 14126
rect 19842 14099 19848 14125
rect 19848 14099 19870 14125
rect 19894 14099 19910 14125
rect 19910 14099 19922 14125
rect 19842 14098 19870 14099
rect 19894 14098 19922 14099
rect 19946 14125 19974 14126
rect 19946 14099 19972 14125
rect 19972 14099 19974 14125
rect 19946 14098 19974 14099
rect 19998 14125 20026 14126
rect 19998 14099 20008 14125
rect 20008 14099 20026 14125
rect 19998 14098 20026 14099
rect 18550 13510 18578 13538
rect 19054 13537 19082 13538
rect 19054 13511 19055 13537
rect 19055 13511 19081 13537
rect 19081 13511 19082 13537
rect 19054 13510 19082 13511
rect 19582 13341 19610 13342
rect 19582 13315 19600 13341
rect 19600 13315 19610 13341
rect 19582 13314 19610 13315
rect 19634 13341 19662 13342
rect 19634 13315 19636 13341
rect 19636 13315 19662 13341
rect 19634 13314 19662 13315
rect 19686 13341 19714 13342
rect 19738 13341 19766 13342
rect 19686 13315 19698 13341
rect 19698 13315 19714 13341
rect 19738 13315 19760 13341
rect 19760 13315 19766 13341
rect 19686 13314 19714 13315
rect 19738 13314 19766 13315
rect 19790 13314 19818 13342
rect 19842 13341 19870 13342
rect 19894 13341 19922 13342
rect 19842 13315 19848 13341
rect 19848 13315 19870 13341
rect 19894 13315 19910 13341
rect 19910 13315 19922 13341
rect 19842 13314 19870 13315
rect 19894 13314 19922 13315
rect 19946 13341 19974 13342
rect 19946 13315 19972 13341
rect 19972 13315 19974 13341
rect 19946 13314 19974 13315
rect 19998 13341 20026 13342
rect 19998 13315 20008 13341
rect 20008 13315 20026 13341
rect 19998 13314 20026 13315
rect 18550 13145 18578 13146
rect 18550 13119 18551 13145
rect 18551 13119 18577 13145
rect 18577 13119 18578 13145
rect 18550 13118 18578 13119
rect 17082 12949 17110 12950
rect 17082 12923 17100 12949
rect 17100 12923 17110 12949
rect 17082 12922 17110 12923
rect 17134 12949 17162 12950
rect 17134 12923 17136 12949
rect 17136 12923 17162 12949
rect 17134 12922 17162 12923
rect 17186 12949 17214 12950
rect 17238 12949 17266 12950
rect 17186 12923 17198 12949
rect 17198 12923 17214 12949
rect 17238 12923 17260 12949
rect 17260 12923 17266 12949
rect 17186 12922 17214 12923
rect 17238 12922 17266 12923
rect 17290 12922 17318 12950
rect 17342 12949 17370 12950
rect 17394 12949 17422 12950
rect 17342 12923 17348 12949
rect 17348 12923 17370 12949
rect 17394 12923 17410 12949
rect 17410 12923 17422 12949
rect 17342 12922 17370 12923
rect 17394 12922 17422 12923
rect 17446 12949 17474 12950
rect 17446 12923 17472 12949
rect 17472 12923 17474 12949
rect 17446 12922 17474 12923
rect 17498 12949 17526 12950
rect 17498 12923 17508 12949
rect 17508 12923 17526 12949
rect 17498 12922 17526 12923
rect 17082 12165 17110 12166
rect 17082 12139 17100 12165
rect 17100 12139 17110 12165
rect 17082 12138 17110 12139
rect 17134 12165 17162 12166
rect 17134 12139 17136 12165
rect 17136 12139 17162 12165
rect 17134 12138 17162 12139
rect 17186 12165 17214 12166
rect 17238 12165 17266 12166
rect 17186 12139 17198 12165
rect 17198 12139 17214 12165
rect 17238 12139 17260 12165
rect 17260 12139 17266 12165
rect 17186 12138 17214 12139
rect 17238 12138 17266 12139
rect 17290 12138 17318 12166
rect 17342 12165 17370 12166
rect 17394 12165 17422 12166
rect 17342 12139 17348 12165
rect 17348 12139 17370 12165
rect 17394 12139 17410 12165
rect 17410 12139 17422 12165
rect 17342 12138 17370 12139
rect 17394 12138 17422 12139
rect 17446 12165 17474 12166
rect 17446 12139 17472 12165
rect 17472 12139 17474 12165
rect 17446 12138 17474 12139
rect 17498 12165 17526 12166
rect 17498 12139 17508 12165
rect 17508 12139 17526 12165
rect 17498 12138 17526 12139
rect 17430 11969 17458 11970
rect 17430 11943 17431 11969
rect 17431 11943 17457 11969
rect 17457 11943 17458 11969
rect 17430 11942 17458 11943
rect 18550 12614 18578 12642
rect 17598 11942 17626 11970
rect 19054 12614 19082 12642
rect 17990 11942 18018 11970
rect 17082 11381 17110 11382
rect 17082 11355 17100 11381
rect 17100 11355 17110 11381
rect 17082 11354 17110 11355
rect 17134 11381 17162 11382
rect 17134 11355 17136 11381
rect 17136 11355 17162 11381
rect 17134 11354 17162 11355
rect 17186 11381 17214 11382
rect 17238 11381 17266 11382
rect 17186 11355 17198 11381
rect 17198 11355 17214 11381
rect 17238 11355 17260 11381
rect 17260 11355 17266 11381
rect 17186 11354 17214 11355
rect 17238 11354 17266 11355
rect 17290 11354 17318 11382
rect 17342 11381 17370 11382
rect 17394 11381 17422 11382
rect 17342 11355 17348 11381
rect 17348 11355 17370 11381
rect 17394 11355 17410 11381
rect 17410 11355 17422 11381
rect 17342 11354 17370 11355
rect 17394 11354 17422 11355
rect 17446 11381 17474 11382
rect 17446 11355 17472 11381
rect 17472 11355 17474 11381
rect 17446 11354 17474 11355
rect 17498 11381 17526 11382
rect 17498 11355 17508 11381
rect 17508 11355 17526 11381
rect 17498 11354 17526 11355
rect 16926 10766 16954 10794
rect 17262 10793 17290 10794
rect 17262 10767 17263 10793
rect 17263 10767 17289 10793
rect 17289 10767 17290 10793
rect 17262 10766 17290 10767
rect 17486 10793 17514 10794
rect 17486 10767 17487 10793
rect 17487 10767 17513 10793
rect 17513 10767 17514 10793
rect 17486 10766 17514 10767
rect 17082 10597 17110 10598
rect 17082 10571 17100 10597
rect 17100 10571 17110 10597
rect 17082 10570 17110 10571
rect 17134 10597 17162 10598
rect 17134 10571 17136 10597
rect 17136 10571 17162 10597
rect 17134 10570 17162 10571
rect 17186 10597 17214 10598
rect 17238 10597 17266 10598
rect 17186 10571 17198 10597
rect 17198 10571 17214 10597
rect 17238 10571 17260 10597
rect 17260 10571 17266 10597
rect 17186 10570 17214 10571
rect 17238 10570 17266 10571
rect 17290 10570 17318 10598
rect 17342 10597 17370 10598
rect 17394 10597 17422 10598
rect 17342 10571 17348 10597
rect 17348 10571 17370 10597
rect 17394 10571 17410 10597
rect 17410 10571 17422 10597
rect 17342 10570 17370 10571
rect 17394 10570 17422 10571
rect 17446 10597 17474 10598
rect 17446 10571 17472 10597
rect 17472 10571 17474 10597
rect 17446 10570 17474 10571
rect 17498 10597 17526 10598
rect 17498 10571 17508 10597
rect 17508 10571 17526 10597
rect 17498 10570 17526 10571
rect 16926 10401 16954 10402
rect 16926 10375 16927 10401
rect 16927 10375 16953 10401
rect 16953 10375 16954 10401
rect 16926 10374 16954 10375
rect 16758 10038 16786 10066
rect 16814 9617 16842 9618
rect 16814 9591 16815 9617
rect 16815 9591 16841 9617
rect 16841 9591 16842 9617
rect 16814 9590 16842 9591
rect 16814 8441 16842 8442
rect 16814 8415 16815 8441
rect 16815 8415 16841 8441
rect 16841 8415 16842 8441
rect 16814 8414 16842 8415
rect 16366 4606 16394 4634
rect 16422 5166 16450 5194
rect 16758 5166 16786 5194
rect 16870 5558 16898 5586
rect 14582 3933 14610 3934
rect 14582 3907 14600 3933
rect 14600 3907 14610 3933
rect 14582 3906 14610 3907
rect 14634 3933 14662 3934
rect 14634 3907 14636 3933
rect 14636 3907 14662 3933
rect 14634 3906 14662 3907
rect 14686 3933 14714 3934
rect 14738 3933 14766 3934
rect 14686 3907 14698 3933
rect 14698 3907 14714 3933
rect 14738 3907 14760 3933
rect 14760 3907 14766 3933
rect 14686 3906 14714 3907
rect 14738 3906 14766 3907
rect 14790 3906 14818 3934
rect 14842 3933 14870 3934
rect 14894 3933 14922 3934
rect 14842 3907 14848 3933
rect 14848 3907 14870 3933
rect 14894 3907 14910 3933
rect 14910 3907 14922 3933
rect 14842 3906 14870 3907
rect 14894 3906 14922 3907
rect 14946 3933 14974 3934
rect 14946 3907 14972 3933
rect 14972 3907 14974 3933
rect 14946 3906 14974 3907
rect 14998 3933 15026 3934
rect 14998 3907 15008 3933
rect 15008 3907 15026 3933
rect 14998 3906 15026 3907
rect 14406 3289 14434 3290
rect 14406 3263 14407 3289
rect 14407 3263 14433 3289
rect 14433 3263 14434 3289
rect 14406 3262 14434 3263
rect 15078 3262 15106 3290
rect 14582 3149 14610 3150
rect 14582 3123 14600 3149
rect 14600 3123 14610 3149
rect 14582 3122 14610 3123
rect 14634 3149 14662 3150
rect 14634 3123 14636 3149
rect 14636 3123 14662 3149
rect 14634 3122 14662 3123
rect 14686 3149 14714 3150
rect 14738 3149 14766 3150
rect 14686 3123 14698 3149
rect 14698 3123 14714 3149
rect 14738 3123 14760 3149
rect 14760 3123 14766 3149
rect 14686 3122 14714 3123
rect 14738 3122 14766 3123
rect 14790 3122 14818 3150
rect 14842 3149 14870 3150
rect 14894 3149 14922 3150
rect 14842 3123 14848 3149
rect 14848 3123 14870 3149
rect 14894 3123 14910 3149
rect 14910 3123 14922 3149
rect 14842 3122 14870 3123
rect 14894 3122 14922 3123
rect 14946 3149 14974 3150
rect 14946 3123 14972 3149
rect 14972 3123 14974 3149
rect 14946 3122 14974 3123
rect 14998 3149 15026 3150
rect 14998 3123 15008 3149
rect 15008 3123 15026 3149
rect 14998 3122 15026 3123
rect 14406 2982 14434 3010
rect 13062 2198 13090 2226
rect 13790 2198 13818 2226
rect 13790 2086 13818 2114
rect 14238 2169 14266 2170
rect 14238 2143 14239 2169
rect 14239 2143 14265 2169
rect 14265 2143 14266 2169
rect 14238 2142 14266 2143
rect 13510 1694 13538 1722
rect 13734 1694 13762 1722
rect 14238 1694 14266 1722
rect 14966 2953 14994 2954
rect 14966 2927 14967 2953
rect 14967 2927 14993 2953
rect 14993 2927 14994 2953
rect 14966 2926 14994 2927
rect 15078 2926 15106 2954
rect 15246 3737 15274 3738
rect 15246 3711 15247 3737
rect 15247 3711 15273 3737
rect 15273 3711 15274 3737
rect 15246 3710 15274 3711
rect 15526 3710 15554 3738
rect 15246 3374 15274 3402
rect 15750 3374 15778 3402
rect 14582 2365 14610 2366
rect 14582 2339 14600 2365
rect 14600 2339 14610 2365
rect 14582 2338 14610 2339
rect 14634 2365 14662 2366
rect 14634 2339 14636 2365
rect 14636 2339 14662 2365
rect 14634 2338 14662 2339
rect 14686 2365 14714 2366
rect 14738 2365 14766 2366
rect 14686 2339 14698 2365
rect 14698 2339 14714 2365
rect 14738 2339 14760 2365
rect 14760 2339 14766 2365
rect 14686 2338 14714 2339
rect 14738 2338 14766 2339
rect 14790 2338 14818 2366
rect 14842 2365 14870 2366
rect 14894 2365 14922 2366
rect 14842 2339 14848 2365
rect 14848 2339 14870 2365
rect 14894 2339 14910 2365
rect 14910 2339 14922 2365
rect 14842 2338 14870 2339
rect 14894 2338 14922 2339
rect 14946 2365 14974 2366
rect 14946 2339 14972 2365
rect 14972 2339 14974 2365
rect 14946 2338 14974 2339
rect 14998 2365 15026 2366
rect 14998 2339 15008 2365
rect 15008 2339 15026 2365
rect 14998 2338 15026 2339
rect 14462 2169 14490 2170
rect 14462 2143 14463 2169
rect 14463 2143 14489 2169
rect 14489 2143 14490 2169
rect 14462 2142 14490 2143
rect 15694 2953 15722 2954
rect 15694 2927 15695 2953
rect 15695 2927 15721 2953
rect 15721 2927 15722 2953
rect 15694 2926 15722 2927
rect 15526 2870 15554 2898
rect 14582 1581 14610 1582
rect 14582 1555 14600 1581
rect 14600 1555 14610 1581
rect 14582 1554 14610 1555
rect 14634 1581 14662 1582
rect 14634 1555 14636 1581
rect 14636 1555 14662 1581
rect 14634 1554 14662 1555
rect 14686 1581 14714 1582
rect 14738 1581 14766 1582
rect 14686 1555 14698 1581
rect 14698 1555 14714 1581
rect 14738 1555 14760 1581
rect 14760 1555 14766 1581
rect 14686 1554 14714 1555
rect 14738 1554 14766 1555
rect 14790 1554 14818 1582
rect 14842 1581 14870 1582
rect 14894 1581 14922 1582
rect 14842 1555 14848 1581
rect 14848 1555 14870 1581
rect 14894 1555 14910 1581
rect 14910 1555 14922 1581
rect 14842 1554 14870 1555
rect 14894 1554 14922 1555
rect 14946 1581 14974 1582
rect 14946 1555 14972 1581
rect 14972 1555 14974 1581
rect 14946 1554 14974 1555
rect 14998 1581 15026 1582
rect 14998 1555 15008 1581
rect 15008 1555 15026 1581
rect 14998 1554 15026 1555
rect 15582 1777 15610 1778
rect 15582 1751 15583 1777
rect 15583 1751 15609 1777
rect 15609 1751 15610 1777
rect 15582 1750 15610 1751
rect 16422 2953 16450 2954
rect 16422 2927 16423 2953
rect 16423 2927 16449 2953
rect 16449 2927 16450 2953
rect 16422 2926 16450 2927
rect 16758 2926 16786 2954
rect 16758 2561 16786 2562
rect 16758 2535 16759 2561
rect 16759 2535 16785 2561
rect 16785 2535 16786 2561
rect 16758 2534 16786 2535
rect 18830 11214 18858 11242
rect 19054 11158 19082 11186
rect 19222 11214 19250 11242
rect 19582 12557 19610 12558
rect 19582 12531 19600 12557
rect 19600 12531 19610 12557
rect 19582 12530 19610 12531
rect 19634 12557 19662 12558
rect 19634 12531 19636 12557
rect 19636 12531 19662 12557
rect 19634 12530 19662 12531
rect 19686 12557 19714 12558
rect 19738 12557 19766 12558
rect 19686 12531 19698 12557
rect 19698 12531 19714 12557
rect 19738 12531 19760 12557
rect 19760 12531 19766 12557
rect 19686 12530 19714 12531
rect 19738 12530 19766 12531
rect 19790 12530 19818 12558
rect 19842 12557 19870 12558
rect 19894 12557 19922 12558
rect 19842 12531 19848 12557
rect 19848 12531 19870 12557
rect 19894 12531 19910 12557
rect 19910 12531 19922 12557
rect 19842 12530 19870 12531
rect 19894 12530 19922 12531
rect 19946 12557 19974 12558
rect 19946 12531 19972 12557
rect 19972 12531 19974 12557
rect 19946 12530 19974 12531
rect 19998 12557 20026 12558
rect 19998 12531 20008 12557
rect 20008 12531 20026 12557
rect 19998 12530 20026 12531
rect 19334 11214 19362 11242
rect 19502 11886 19530 11914
rect 18830 10766 18858 10794
rect 17082 9813 17110 9814
rect 17082 9787 17100 9813
rect 17100 9787 17110 9813
rect 17082 9786 17110 9787
rect 17134 9813 17162 9814
rect 17134 9787 17136 9813
rect 17136 9787 17162 9813
rect 17134 9786 17162 9787
rect 17186 9813 17214 9814
rect 17238 9813 17266 9814
rect 17186 9787 17198 9813
rect 17198 9787 17214 9813
rect 17238 9787 17260 9813
rect 17260 9787 17266 9813
rect 17186 9786 17214 9787
rect 17238 9786 17266 9787
rect 17290 9786 17318 9814
rect 17342 9813 17370 9814
rect 17394 9813 17422 9814
rect 17342 9787 17348 9813
rect 17348 9787 17370 9813
rect 17394 9787 17410 9813
rect 17410 9787 17422 9813
rect 17342 9786 17370 9787
rect 17394 9786 17422 9787
rect 17446 9813 17474 9814
rect 17446 9787 17472 9813
rect 17472 9787 17474 9813
rect 17446 9786 17474 9787
rect 17498 9813 17526 9814
rect 17498 9787 17508 9813
rect 17508 9787 17526 9813
rect 17498 9786 17526 9787
rect 17990 9281 18018 9282
rect 17990 9255 17991 9281
rect 17991 9255 18017 9281
rect 18017 9255 18018 9281
rect 17990 9254 18018 9255
rect 17082 9029 17110 9030
rect 17082 9003 17100 9029
rect 17100 9003 17110 9029
rect 17082 9002 17110 9003
rect 17134 9029 17162 9030
rect 17134 9003 17136 9029
rect 17136 9003 17162 9029
rect 17134 9002 17162 9003
rect 17186 9029 17214 9030
rect 17238 9029 17266 9030
rect 17186 9003 17198 9029
rect 17198 9003 17214 9029
rect 17238 9003 17260 9029
rect 17260 9003 17266 9029
rect 17186 9002 17214 9003
rect 17238 9002 17266 9003
rect 17290 9002 17318 9030
rect 17342 9029 17370 9030
rect 17394 9029 17422 9030
rect 17342 9003 17348 9029
rect 17348 9003 17370 9029
rect 17394 9003 17410 9029
rect 17410 9003 17422 9029
rect 17342 9002 17370 9003
rect 17394 9002 17422 9003
rect 17446 9029 17474 9030
rect 17446 9003 17472 9029
rect 17472 9003 17474 9029
rect 17446 9002 17474 9003
rect 17498 9029 17526 9030
rect 17498 9003 17508 9029
rect 17508 9003 17526 9029
rect 17498 9002 17526 9003
rect 18214 10318 18242 10346
rect 17082 8245 17110 8246
rect 17082 8219 17100 8245
rect 17100 8219 17110 8245
rect 17082 8218 17110 8219
rect 17134 8245 17162 8246
rect 17134 8219 17136 8245
rect 17136 8219 17162 8245
rect 17134 8218 17162 8219
rect 17186 8245 17214 8246
rect 17238 8245 17266 8246
rect 17186 8219 17198 8245
rect 17198 8219 17214 8245
rect 17238 8219 17260 8245
rect 17260 8219 17266 8245
rect 17186 8218 17214 8219
rect 17238 8218 17266 8219
rect 17290 8218 17318 8246
rect 17342 8245 17370 8246
rect 17394 8245 17422 8246
rect 17342 8219 17348 8245
rect 17348 8219 17370 8245
rect 17394 8219 17410 8245
rect 17410 8219 17422 8245
rect 17342 8218 17370 8219
rect 17394 8218 17422 8219
rect 17446 8245 17474 8246
rect 17446 8219 17472 8245
rect 17472 8219 17474 8245
rect 17446 8218 17474 8219
rect 17498 8245 17526 8246
rect 17498 8219 17508 8245
rect 17508 8219 17526 8245
rect 17498 8218 17526 8219
rect 17082 7461 17110 7462
rect 17082 7435 17100 7461
rect 17100 7435 17110 7461
rect 17082 7434 17110 7435
rect 17134 7461 17162 7462
rect 17134 7435 17136 7461
rect 17136 7435 17162 7461
rect 17134 7434 17162 7435
rect 17186 7461 17214 7462
rect 17238 7461 17266 7462
rect 17186 7435 17198 7461
rect 17198 7435 17214 7461
rect 17238 7435 17260 7461
rect 17260 7435 17266 7461
rect 17186 7434 17214 7435
rect 17238 7434 17266 7435
rect 17290 7434 17318 7462
rect 17342 7461 17370 7462
rect 17394 7461 17422 7462
rect 17342 7435 17348 7461
rect 17348 7435 17370 7461
rect 17394 7435 17410 7461
rect 17410 7435 17422 7461
rect 17342 7434 17370 7435
rect 17394 7434 17422 7435
rect 17446 7461 17474 7462
rect 17446 7435 17472 7461
rect 17472 7435 17474 7461
rect 17446 7434 17474 7435
rect 17498 7461 17526 7462
rect 17498 7435 17508 7461
rect 17508 7435 17526 7461
rect 17498 7434 17526 7435
rect 17082 6677 17110 6678
rect 17082 6651 17100 6677
rect 17100 6651 17110 6677
rect 17082 6650 17110 6651
rect 17134 6677 17162 6678
rect 17134 6651 17136 6677
rect 17136 6651 17162 6677
rect 17134 6650 17162 6651
rect 17186 6677 17214 6678
rect 17238 6677 17266 6678
rect 17186 6651 17198 6677
rect 17198 6651 17214 6677
rect 17238 6651 17260 6677
rect 17260 6651 17266 6677
rect 17186 6650 17214 6651
rect 17238 6650 17266 6651
rect 17290 6650 17318 6678
rect 17342 6677 17370 6678
rect 17394 6677 17422 6678
rect 17342 6651 17348 6677
rect 17348 6651 17370 6677
rect 17394 6651 17410 6677
rect 17410 6651 17422 6677
rect 17342 6650 17370 6651
rect 17394 6650 17422 6651
rect 17446 6677 17474 6678
rect 17446 6651 17472 6677
rect 17472 6651 17474 6677
rect 17446 6650 17474 6651
rect 17498 6677 17526 6678
rect 17498 6651 17508 6677
rect 17508 6651 17526 6677
rect 17498 6650 17526 6651
rect 17486 6481 17514 6482
rect 17486 6455 17487 6481
rect 17487 6455 17513 6481
rect 17513 6455 17514 6481
rect 17486 6454 17514 6455
rect 17082 5893 17110 5894
rect 17082 5867 17100 5893
rect 17100 5867 17110 5893
rect 17082 5866 17110 5867
rect 17134 5893 17162 5894
rect 17134 5867 17136 5893
rect 17136 5867 17162 5893
rect 17134 5866 17162 5867
rect 17186 5893 17214 5894
rect 17238 5893 17266 5894
rect 17186 5867 17198 5893
rect 17198 5867 17214 5893
rect 17238 5867 17260 5893
rect 17260 5867 17266 5893
rect 17186 5866 17214 5867
rect 17238 5866 17266 5867
rect 17290 5866 17318 5894
rect 17342 5893 17370 5894
rect 17394 5893 17422 5894
rect 17342 5867 17348 5893
rect 17348 5867 17370 5893
rect 17394 5867 17410 5893
rect 17410 5867 17422 5893
rect 17342 5866 17370 5867
rect 17394 5866 17422 5867
rect 17446 5893 17474 5894
rect 17446 5867 17472 5893
rect 17472 5867 17474 5893
rect 17446 5866 17474 5867
rect 17498 5893 17526 5894
rect 17498 5867 17508 5893
rect 17508 5867 17526 5893
rect 17498 5866 17526 5867
rect 17082 5109 17110 5110
rect 17082 5083 17100 5109
rect 17100 5083 17110 5109
rect 17082 5082 17110 5083
rect 17134 5109 17162 5110
rect 17134 5083 17136 5109
rect 17136 5083 17162 5109
rect 17134 5082 17162 5083
rect 17186 5109 17214 5110
rect 17238 5109 17266 5110
rect 17186 5083 17198 5109
rect 17198 5083 17214 5109
rect 17238 5083 17260 5109
rect 17260 5083 17266 5109
rect 17186 5082 17214 5083
rect 17238 5082 17266 5083
rect 17290 5082 17318 5110
rect 17342 5109 17370 5110
rect 17394 5109 17422 5110
rect 17342 5083 17348 5109
rect 17348 5083 17370 5109
rect 17394 5083 17410 5109
rect 17410 5083 17422 5109
rect 17342 5082 17370 5083
rect 17394 5082 17422 5083
rect 17446 5109 17474 5110
rect 17446 5083 17472 5109
rect 17472 5083 17474 5109
rect 17446 5082 17474 5083
rect 17498 5109 17526 5110
rect 17498 5083 17508 5109
rect 17508 5083 17526 5109
rect 17498 5082 17526 5083
rect 16982 4438 17010 4466
rect 17082 4325 17110 4326
rect 17082 4299 17100 4325
rect 17100 4299 17110 4325
rect 17082 4298 17110 4299
rect 17134 4325 17162 4326
rect 17134 4299 17136 4325
rect 17136 4299 17162 4325
rect 17134 4298 17162 4299
rect 17186 4325 17214 4326
rect 17238 4325 17266 4326
rect 17186 4299 17198 4325
rect 17198 4299 17214 4325
rect 17238 4299 17260 4325
rect 17260 4299 17266 4325
rect 17186 4298 17214 4299
rect 17238 4298 17266 4299
rect 17290 4298 17318 4326
rect 17342 4325 17370 4326
rect 17394 4325 17422 4326
rect 17342 4299 17348 4325
rect 17348 4299 17370 4325
rect 17394 4299 17410 4325
rect 17410 4299 17422 4325
rect 17342 4298 17370 4299
rect 17394 4298 17422 4299
rect 17446 4325 17474 4326
rect 17446 4299 17472 4325
rect 17472 4299 17474 4325
rect 17446 4298 17474 4299
rect 17498 4325 17526 4326
rect 17498 4299 17508 4325
rect 17508 4299 17526 4325
rect 17498 4298 17526 4299
rect 17082 3541 17110 3542
rect 17082 3515 17100 3541
rect 17100 3515 17110 3541
rect 17082 3514 17110 3515
rect 17134 3541 17162 3542
rect 17134 3515 17136 3541
rect 17136 3515 17162 3541
rect 17134 3514 17162 3515
rect 17186 3541 17214 3542
rect 17238 3541 17266 3542
rect 17186 3515 17198 3541
rect 17198 3515 17214 3541
rect 17238 3515 17260 3541
rect 17260 3515 17266 3541
rect 17186 3514 17214 3515
rect 17238 3514 17266 3515
rect 17290 3514 17318 3542
rect 17342 3541 17370 3542
rect 17394 3541 17422 3542
rect 17342 3515 17348 3541
rect 17348 3515 17370 3541
rect 17394 3515 17410 3541
rect 17410 3515 17422 3541
rect 17342 3514 17370 3515
rect 17394 3514 17422 3515
rect 17446 3541 17474 3542
rect 17446 3515 17472 3541
rect 17472 3515 17474 3541
rect 17446 3514 17474 3515
rect 17498 3541 17526 3542
rect 17498 3515 17508 3541
rect 17508 3515 17526 3541
rect 17498 3514 17526 3515
rect 17598 3374 17626 3402
rect 18270 8441 18298 8442
rect 18270 8415 18271 8441
rect 18271 8415 18297 8441
rect 18297 8415 18298 8441
rect 18270 8414 18298 8415
rect 20846 14294 20874 14322
rect 20790 13929 20818 13930
rect 20790 13903 20791 13929
rect 20791 13903 20817 13929
rect 20817 13903 20818 13929
rect 20790 13902 20818 13903
rect 20510 13510 20538 13538
rect 21406 13510 21434 13538
rect 21238 13454 21266 13482
rect 19950 11913 19978 11914
rect 19950 11887 19951 11913
rect 19951 11887 19977 11913
rect 19977 11887 19978 11913
rect 19950 11886 19978 11887
rect 19582 11773 19610 11774
rect 19582 11747 19600 11773
rect 19600 11747 19610 11773
rect 19582 11746 19610 11747
rect 19634 11773 19662 11774
rect 19634 11747 19636 11773
rect 19636 11747 19662 11773
rect 19634 11746 19662 11747
rect 19686 11773 19714 11774
rect 19738 11773 19766 11774
rect 19686 11747 19698 11773
rect 19698 11747 19714 11773
rect 19738 11747 19760 11773
rect 19760 11747 19766 11773
rect 19686 11746 19714 11747
rect 19738 11746 19766 11747
rect 19790 11746 19818 11774
rect 19842 11773 19870 11774
rect 19894 11773 19922 11774
rect 19842 11747 19848 11773
rect 19848 11747 19870 11773
rect 19894 11747 19910 11773
rect 19910 11747 19922 11773
rect 19842 11746 19870 11747
rect 19894 11746 19922 11747
rect 19946 11773 19974 11774
rect 19946 11747 19972 11773
rect 19972 11747 19974 11773
rect 19946 11746 19974 11747
rect 19998 11773 20026 11774
rect 19998 11747 20008 11773
rect 20008 11747 20026 11773
rect 19998 11746 20026 11747
rect 19950 11214 19978 11242
rect 20230 11185 20258 11186
rect 20230 11159 20231 11185
rect 20231 11159 20257 11185
rect 20257 11159 20258 11185
rect 20230 11158 20258 11159
rect 20790 11158 20818 11186
rect 19950 11046 19978 11074
rect 19582 10989 19610 10990
rect 19582 10963 19600 10989
rect 19600 10963 19610 10989
rect 19582 10962 19610 10963
rect 19634 10989 19662 10990
rect 19634 10963 19636 10989
rect 19636 10963 19662 10989
rect 19634 10962 19662 10963
rect 19686 10989 19714 10990
rect 19738 10989 19766 10990
rect 19686 10963 19698 10989
rect 19698 10963 19714 10989
rect 19738 10963 19760 10989
rect 19760 10963 19766 10989
rect 19686 10962 19714 10963
rect 19738 10962 19766 10963
rect 19790 10962 19818 10990
rect 19842 10989 19870 10990
rect 19894 10989 19922 10990
rect 19842 10963 19848 10989
rect 19848 10963 19870 10989
rect 19894 10963 19910 10989
rect 19910 10963 19922 10989
rect 19842 10962 19870 10963
rect 19894 10962 19922 10963
rect 19946 10989 19974 10990
rect 19946 10963 19972 10989
rect 19972 10963 19974 10989
rect 19946 10962 19974 10963
rect 19998 10989 20026 10990
rect 19998 10963 20008 10989
rect 20008 10963 20026 10989
rect 19998 10962 20026 10963
rect 20958 12334 20986 12362
rect 19582 10205 19610 10206
rect 19582 10179 19600 10205
rect 19600 10179 19610 10205
rect 19582 10178 19610 10179
rect 19634 10205 19662 10206
rect 19634 10179 19636 10205
rect 19636 10179 19662 10205
rect 19634 10178 19662 10179
rect 19686 10205 19714 10206
rect 19738 10205 19766 10206
rect 19686 10179 19698 10205
rect 19698 10179 19714 10205
rect 19738 10179 19760 10205
rect 19760 10179 19766 10205
rect 19686 10178 19714 10179
rect 19738 10178 19766 10179
rect 19790 10178 19818 10206
rect 19842 10205 19870 10206
rect 19894 10205 19922 10206
rect 19842 10179 19848 10205
rect 19848 10179 19870 10205
rect 19894 10179 19910 10205
rect 19910 10179 19922 10205
rect 19842 10178 19870 10179
rect 19894 10178 19922 10179
rect 19946 10205 19974 10206
rect 19946 10179 19972 10205
rect 19972 10179 19974 10205
rect 19946 10178 19974 10179
rect 19998 10205 20026 10206
rect 19998 10179 20008 10205
rect 20008 10179 20026 10205
rect 19998 10178 20026 10179
rect 19582 9421 19610 9422
rect 19582 9395 19600 9421
rect 19600 9395 19610 9421
rect 19582 9394 19610 9395
rect 19634 9421 19662 9422
rect 19634 9395 19636 9421
rect 19636 9395 19662 9421
rect 19634 9394 19662 9395
rect 19686 9421 19714 9422
rect 19738 9421 19766 9422
rect 19686 9395 19698 9421
rect 19698 9395 19714 9421
rect 19738 9395 19760 9421
rect 19760 9395 19766 9421
rect 19686 9394 19714 9395
rect 19738 9394 19766 9395
rect 19790 9394 19818 9422
rect 19842 9421 19870 9422
rect 19894 9421 19922 9422
rect 19842 9395 19848 9421
rect 19848 9395 19870 9421
rect 19894 9395 19910 9421
rect 19910 9395 19922 9421
rect 19842 9394 19870 9395
rect 19894 9394 19922 9395
rect 19946 9421 19974 9422
rect 19946 9395 19972 9421
rect 19972 9395 19974 9421
rect 19946 9394 19974 9395
rect 19998 9421 20026 9422
rect 19998 9395 20008 9421
rect 20008 9395 20026 9421
rect 19998 9394 20026 9395
rect 19278 9254 19306 9282
rect 18774 8414 18802 8442
rect 19582 8637 19610 8638
rect 19582 8611 19600 8637
rect 19600 8611 19610 8637
rect 19582 8610 19610 8611
rect 19634 8637 19662 8638
rect 19634 8611 19636 8637
rect 19636 8611 19662 8637
rect 19634 8610 19662 8611
rect 19686 8637 19714 8638
rect 19738 8637 19766 8638
rect 19686 8611 19698 8637
rect 19698 8611 19714 8637
rect 19738 8611 19760 8637
rect 19760 8611 19766 8637
rect 19686 8610 19714 8611
rect 19738 8610 19766 8611
rect 19790 8610 19818 8638
rect 19842 8637 19870 8638
rect 19894 8637 19922 8638
rect 19842 8611 19848 8637
rect 19848 8611 19870 8637
rect 19894 8611 19910 8637
rect 19910 8611 19922 8637
rect 19842 8610 19870 8611
rect 19894 8610 19922 8611
rect 19946 8637 19974 8638
rect 19946 8611 19972 8637
rect 19972 8611 19974 8637
rect 19946 8610 19974 8611
rect 19998 8637 20026 8638
rect 19998 8611 20008 8637
rect 20008 8611 20026 8637
rect 19998 8610 20026 8611
rect 20230 8470 20258 8498
rect 19446 8441 19474 8442
rect 19446 8415 19447 8441
rect 19447 8415 19473 8441
rect 19473 8415 19474 8441
rect 19446 8414 19474 8415
rect 19950 8414 19978 8442
rect 20902 10766 20930 10794
rect 21742 13510 21770 13538
rect 21462 13454 21490 13482
rect 21798 12222 21826 12250
rect 21294 11046 21322 11074
rect 21350 11886 21378 11914
rect 22082 18437 22110 18438
rect 22082 18411 22100 18437
rect 22100 18411 22110 18437
rect 22082 18410 22110 18411
rect 22134 18437 22162 18438
rect 22134 18411 22136 18437
rect 22136 18411 22162 18437
rect 22134 18410 22162 18411
rect 22186 18437 22214 18438
rect 22238 18437 22266 18438
rect 22186 18411 22198 18437
rect 22198 18411 22214 18437
rect 22238 18411 22260 18437
rect 22260 18411 22266 18437
rect 22186 18410 22214 18411
rect 22238 18410 22266 18411
rect 22290 18410 22318 18438
rect 22342 18437 22370 18438
rect 22394 18437 22422 18438
rect 22342 18411 22348 18437
rect 22348 18411 22370 18437
rect 22394 18411 22410 18437
rect 22410 18411 22422 18437
rect 22342 18410 22370 18411
rect 22394 18410 22422 18411
rect 22446 18437 22474 18438
rect 22446 18411 22472 18437
rect 22472 18411 22474 18437
rect 22446 18410 22474 18411
rect 22498 18437 22526 18438
rect 22498 18411 22508 18437
rect 22508 18411 22526 18437
rect 22498 18410 22526 18411
rect 24582 18045 24610 18046
rect 24582 18019 24600 18045
rect 24600 18019 24610 18045
rect 24582 18018 24610 18019
rect 24634 18045 24662 18046
rect 24634 18019 24636 18045
rect 24636 18019 24662 18045
rect 24634 18018 24662 18019
rect 24686 18045 24714 18046
rect 24738 18045 24766 18046
rect 24686 18019 24698 18045
rect 24698 18019 24714 18045
rect 24738 18019 24760 18045
rect 24760 18019 24766 18045
rect 24686 18018 24714 18019
rect 24738 18018 24766 18019
rect 24790 18018 24818 18046
rect 24842 18045 24870 18046
rect 24894 18045 24922 18046
rect 24842 18019 24848 18045
rect 24848 18019 24870 18045
rect 24894 18019 24910 18045
rect 24910 18019 24922 18045
rect 24842 18018 24870 18019
rect 24894 18018 24922 18019
rect 24946 18045 24974 18046
rect 24946 18019 24972 18045
rect 24972 18019 24974 18045
rect 24946 18018 24974 18019
rect 24998 18045 25026 18046
rect 24998 18019 25008 18045
rect 25008 18019 25026 18045
rect 24998 18018 25026 18019
rect 22082 17653 22110 17654
rect 22082 17627 22100 17653
rect 22100 17627 22110 17653
rect 22082 17626 22110 17627
rect 22134 17653 22162 17654
rect 22134 17627 22136 17653
rect 22136 17627 22162 17653
rect 22134 17626 22162 17627
rect 22186 17653 22214 17654
rect 22238 17653 22266 17654
rect 22186 17627 22198 17653
rect 22198 17627 22214 17653
rect 22238 17627 22260 17653
rect 22260 17627 22266 17653
rect 22186 17626 22214 17627
rect 22238 17626 22266 17627
rect 22290 17626 22318 17654
rect 22342 17653 22370 17654
rect 22394 17653 22422 17654
rect 22342 17627 22348 17653
rect 22348 17627 22370 17653
rect 22394 17627 22410 17653
rect 22410 17627 22422 17653
rect 22342 17626 22370 17627
rect 22394 17626 22422 17627
rect 22446 17653 22474 17654
rect 22446 17627 22472 17653
rect 22472 17627 22474 17653
rect 22446 17626 22474 17627
rect 22498 17653 22526 17654
rect 22498 17627 22508 17653
rect 22508 17627 22526 17653
rect 22498 17626 22526 17627
rect 23926 17318 23954 17346
rect 22082 16869 22110 16870
rect 22082 16843 22100 16869
rect 22100 16843 22110 16869
rect 22082 16842 22110 16843
rect 22134 16869 22162 16870
rect 22134 16843 22136 16869
rect 22136 16843 22162 16869
rect 22134 16842 22162 16843
rect 22186 16869 22214 16870
rect 22238 16869 22266 16870
rect 22186 16843 22198 16869
rect 22198 16843 22214 16869
rect 22238 16843 22260 16869
rect 22260 16843 22266 16869
rect 22186 16842 22214 16843
rect 22238 16842 22266 16843
rect 22290 16842 22318 16870
rect 22342 16869 22370 16870
rect 22394 16869 22422 16870
rect 22342 16843 22348 16869
rect 22348 16843 22370 16869
rect 22394 16843 22410 16869
rect 22410 16843 22422 16869
rect 22342 16842 22370 16843
rect 22394 16842 22422 16843
rect 22446 16869 22474 16870
rect 22446 16843 22472 16869
rect 22472 16843 22474 16869
rect 22446 16842 22474 16843
rect 22498 16869 22526 16870
rect 22498 16843 22508 16869
rect 22508 16843 22526 16869
rect 22498 16842 22526 16843
rect 22082 16085 22110 16086
rect 22082 16059 22100 16085
rect 22100 16059 22110 16085
rect 22082 16058 22110 16059
rect 22134 16085 22162 16086
rect 22134 16059 22136 16085
rect 22136 16059 22162 16085
rect 22134 16058 22162 16059
rect 22186 16085 22214 16086
rect 22238 16085 22266 16086
rect 22186 16059 22198 16085
rect 22198 16059 22214 16085
rect 22238 16059 22260 16085
rect 22260 16059 22266 16085
rect 22186 16058 22214 16059
rect 22238 16058 22266 16059
rect 22290 16058 22318 16086
rect 22342 16085 22370 16086
rect 22394 16085 22422 16086
rect 22342 16059 22348 16085
rect 22348 16059 22370 16085
rect 22394 16059 22410 16085
rect 22410 16059 22422 16085
rect 22342 16058 22370 16059
rect 22394 16058 22422 16059
rect 22446 16085 22474 16086
rect 22446 16059 22472 16085
rect 22472 16059 22474 16085
rect 22446 16058 22474 16059
rect 22498 16085 22526 16086
rect 22498 16059 22508 16085
rect 22508 16059 22526 16085
rect 22498 16058 22526 16059
rect 22082 15301 22110 15302
rect 22082 15275 22100 15301
rect 22100 15275 22110 15301
rect 22082 15274 22110 15275
rect 22134 15301 22162 15302
rect 22134 15275 22136 15301
rect 22136 15275 22162 15301
rect 22134 15274 22162 15275
rect 22186 15301 22214 15302
rect 22238 15301 22266 15302
rect 22186 15275 22198 15301
rect 22198 15275 22214 15301
rect 22238 15275 22260 15301
rect 22260 15275 22266 15301
rect 22186 15274 22214 15275
rect 22238 15274 22266 15275
rect 22290 15274 22318 15302
rect 22342 15301 22370 15302
rect 22394 15301 22422 15302
rect 22342 15275 22348 15301
rect 22348 15275 22370 15301
rect 22394 15275 22410 15301
rect 22410 15275 22422 15301
rect 22342 15274 22370 15275
rect 22394 15274 22422 15275
rect 22446 15301 22474 15302
rect 22446 15275 22472 15301
rect 22472 15275 22474 15301
rect 22446 15274 22474 15275
rect 22498 15301 22526 15302
rect 22498 15275 22508 15301
rect 22508 15275 22526 15301
rect 22498 15274 22526 15275
rect 22082 14517 22110 14518
rect 22082 14491 22100 14517
rect 22100 14491 22110 14517
rect 22082 14490 22110 14491
rect 22134 14517 22162 14518
rect 22134 14491 22136 14517
rect 22136 14491 22162 14517
rect 22134 14490 22162 14491
rect 22186 14517 22214 14518
rect 22238 14517 22266 14518
rect 22186 14491 22198 14517
rect 22198 14491 22214 14517
rect 22238 14491 22260 14517
rect 22260 14491 22266 14517
rect 22186 14490 22214 14491
rect 22238 14490 22266 14491
rect 22290 14490 22318 14518
rect 22342 14517 22370 14518
rect 22394 14517 22422 14518
rect 22342 14491 22348 14517
rect 22348 14491 22370 14517
rect 22394 14491 22410 14517
rect 22410 14491 22422 14517
rect 22342 14490 22370 14491
rect 22394 14490 22422 14491
rect 22446 14517 22474 14518
rect 22446 14491 22472 14517
rect 22472 14491 22474 14517
rect 22446 14490 22474 14491
rect 22498 14517 22526 14518
rect 22498 14491 22508 14517
rect 22508 14491 22526 14517
rect 22498 14490 22526 14491
rect 22582 13846 22610 13874
rect 22082 13733 22110 13734
rect 22082 13707 22100 13733
rect 22100 13707 22110 13733
rect 22082 13706 22110 13707
rect 22134 13733 22162 13734
rect 22134 13707 22136 13733
rect 22136 13707 22162 13733
rect 22134 13706 22162 13707
rect 22186 13733 22214 13734
rect 22238 13733 22266 13734
rect 22186 13707 22198 13733
rect 22198 13707 22214 13733
rect 22238 13707 22260 13733
rect 22260 13707 22266 13733
rect 22186 13706 22214 13707
rect 22238 13706 22266 13707
rect 22290 13706 22318 13734
rect 22342 13733 22370 13734
rect 22394 13733 22422 13734
rect 22342 13707 22348 13733
rect 22348 13707 22370 13733
rect 22394 13707 22410 13733
rect 22410 13707 22422 13733
rect 22342 13706 22370 13707
rect 22394 13706 22422 13707
rect 22446 13733 22474 13734
rect 22446 13707 22472 13733
rect 22472 13707 22474 13733
rect 22446 13706 22474 13707
rect 22498 13733 22526 13734
rect 22498 13707 22508 13733
rect 22508 13707 22526 13733
rect 22498 13706 22526 13707
rect 22526 13454 22554 13482
rect 23870 14265 23898 14266
rect 23870 14239 23871 14265
rect 23871 14239 23897 14265
rect 23897 14239 23898 14265
rect 23870 14238 23898 14239
rect 23030 13454 23058 13482
rect 23422 13510 23450 13538
rect 22082 12949 22110 12950
rect 22082 12923 22100 12949
rect 22100 12923 22110 12949
rect 22082 12922 22110 12923
rect 22134 12949 22162 12950
rect 22134 12923 22136 12949
rect 22136 12923 22162 12949
rect 22134 12922 22162 12923
rect 22186 12949 22214 12950
rect 22238 12949 22266 12950
rect 22186 12923 22198 12949
rect 22198 12923 22214 12949
rect 22238 12923 22260 12949
rect 22260 12923 22266 12949
rect 22186 12922 22214 12923
rect 22238 12922 22266 12923
rect 22290 12922 22318 12950
rect 22342 12949 22370 12950
rect 22394 12949 22422 12950
rect 22342 12923 22348 12949
rect 22348 12923 22370 12949
rect 22394 12923 22410 12949
rect 22410 12923 22422 12949
rect 22342 12922 22370 12923
rect 22394 12922 22422 12923
rect 22446 12949 22474 12950
rect 22446 12923 22472 12949
rect 22472 12923 22474 12949
rect 22446 12922 22474 12923
rect 22498 12949 22526 12950
rect 22498 12923 22508 12949
rect 22508 12923 22526 12949
rect 22498 12922 22526 12923
rect 23870 13537 23898 13538
rect 23870 13511 23871 13537
rect 23871 13511 23897 13537
rect 23897 13511 23898 13537
rect 23870 13510 23898 13511
rect 23870 12697 23898 12698
rect 23870 12671 23871 12697
rect 23871 12671 23897 12697
rect 23897 12671 23898 12697
rect 23870 12670 23898 12671
rect 22526 12361 22554 12362
rect 22526 12335 22527 12361
rect 22527 12335 22553 12361
rect 22553 12335 22554 12361
rect 22526 12334 22554 12335
rect 22082 12165 22110 12166
rect 22082 12139 22100 12165
rect 22100 12139 22110 12165
rect 22082 12138 22110 12139
rect 22134 12165 22162 12166
rect 22134 12139 22136 12165
rect 22136 12139 22162 12165
rect 22134 12138 22162 12139
rect 22186 12165 22214 12166
rect 22238 12165 22266 12166
rect 22186 12139 22198 12165
rect 22198 12139 22214 12165
rect 22238 12139 22260 12165
rect 22260 12139 22266 12165
rect 22186 12138 22214 12139
rect 22238 12138 22266 12139
rect 22290 12138 22318 12166
rect 22342 12165 22370 12166
rect 22394 12165 22422 12166
rect 22342 12139 22348 12165
rect 22348 12139 22370 12165
rect 22394 12139 22410 12165
rect 22410 12139 22422 12165
rect 22342 12138 22370 12139
rect 22394 12138 22422 12139
rect 22446 12165 22474 12166
rect 22446 12139 22472 12165
rect 22472 12139 22474 12165
rect 22446 12138 22474 12139
rect 22498 12165 22526 12166
rect 22498 12139 22508 12165
rect 22508 12139 22526 12165
rect 22498 12138 22526 12139
rect 23422 12222 23450 12250
rect 22582 11942 22610 11970
rect 23030 11969 23058 11970
rect 23030 11943 23031 11969
rect 23031 11943 23057 11969
rect 23057 11943 23058 11969
rect 23030 11942 23058 11943
rect 22082 11381 22110 11382
rect 22082 11355 22100 11381
rect 22100 11355 22110 11381
rect 22082 11354 22110 11355
rect 22134 11381 22162 11382
rect 22134 11355 22136 11381
rect 22136 11355 22162 11381
rect 22134 11354 22162 11355
rect 22186 11381 22214 11382
rect 22238 11381 22266 11382
rect 22186 11355 22198 11381
rect 22198 11355 22214 11381
rect 22238 11355 22260 11381
rect 22260 11355 22266 11381
rect 22186 11354 22214 11355
rect 22238 11354 22266 11355
rect 22290 11354 22318 11382
rect 22342 11381 22370 11382
rect 22394 11381 22422 11382
rect 22342 11355 22348 11381
rect 22348 11355 22370 11381
rect 22394 11355 22410 11381
rect 22410 11355 22422 11381
rect 22342 11354 22370 11355
rect 22394 11354 22422 11355
rect 22446 11381 22474 11382
rect 22446 11355 22472 11381
rect 22472 11355 22474 11381
rect 22446 11354 22474 11355
rect 22498 11381 22526 11382
rect 22498 11355 22508 11381
rect 22508 11355 22526 11381
rect 22498 11354 22526 11355
rect 21854 11158 21882 11186
rect 20846 9982 20874 10010
rect 20790 8470 20818 8498
rect 21406 8414 21434 8442
rect 21406 8302 21434 8330
rect 21798 8302 21826 8330
rect 19582 7853 19610 7854
rect 19582 7827 19600 7853
rect 19600 7827 19610 7853
rect 19582 7826 19610 7827
rect 19634 7853 19662 7854
rect 19634 7827 19636 7853
rect 19636 7827 19662 7853
rect 19634 7826 19662 7827
rect 19686 7853 19714 7854
rect 19738 7853 19766 7854
rect 19686 7827 19698 7853
rect 19698 7827 19714 7853
rect 19738 7827 19760 7853
rect 19760 7827 19766 7853
rect 19686 7826 19714 7827
rect 19738 7826 19766 7827
rect 19790 7826 19818 7854
rect 19842 7853 19870 7854
rect 19894 7853 19922 7854
rect 19842 7827 19848 7853
rect 19848 7827 19870 7853
rect 19894 7827 19910 7853
rect 19910 7827 19922 7853
rect 19842 7826 19870 7827
rect 19894 7826 19922 7827
rect 19946 7853 19974 7854
rect 19946 7827 19972 7853
rect 19972 7827 19974 7853
rect 19946 7826 19974 7827
rect 19998 7853 20026 7854
rect 19998 7827 20008 7853
rect 20008 7827 20026 7853
rect 19998 7826 20026 7827
rect 22526 10793 22554 10794
rect 22526 10767 22527 10793
rect 22527 10767 22553 10793
rect 22553 10767 22554 10793
rect 22526 10766 22554 10767
rect 23030 10766 23058 10794
rect 22082 10597 22110 10598
rect 22082 10571 22100 10597
rect 22100 10571 22110 10597
rect 22082 10570 22110 10571
rect 22134 10597 22162 10598
rect 22134 10571 22136 10597
rect 22136 10571 22162 10597
rect 22134 10570 22162 10571
rect 22186 10597 22214 10598
rect 22238 10597 22266 10598
rect 22186 10571 22198 10597
rect 22198 10571 22214 10597
rect 22238 10571 22260 10597
rect 22260 10571 22266 10597
rect 22186 10570 22214 10571
rect 22238 10570 22266 10571
rect 22290 10570 22318 10598
rect 22342 10597 22370 10598
rect 22394 10597 22422 10598
rect 22342 10571 22348 10597
rect 22348 10571 22370 10597
rect 22394 10571 22410 10597
rect 22410 10571 22422 10597
rect 22342 10570 22370 10571
rect 22394 10570 22422 10571
rect 22446 10597 22474 10598
rect 22446 10571 22472 10597
rect 22472 10571 22474 10597
rect 22446 10570 22474 10571
rect 22498 10597 22526 10598
rect 22498 10571 22508 10597
rect 22508 10571 22526 10597
rect 22498 10570 22526 10571
rect 23030 10262 23058 10290
rect 22246 10009 22274 10010
rect 22246 9983 22247 10009
rect 22247 9983 22273 10009
rect 22273 9983 22274 10009
rect 22246 9982 22274 9983
rect 22582 9982 22610 10010
rect 22082 9813 22110 9814
rect 22082 9787 22100 9813
rect 22100 9787 22110 9813
rect 22082 9786 22110 9787
rect 22134 9813 22162 9814
rect 22134 9787 22136 9813
rect 22136 9787 22162 9813
rect 22134 9786 22162 9787
rect 22186 9813 22214 9814
rect 22238 9813 22266 9814
rect 22186 9787 22198 9813
rect 22198 9787 22214 9813
rect 22238 9787 22260 9813
rect 22260 9787 22266 9813
rect 22186 9786 22214 9787
rect 22238 9786 22266 9787
rect 22290 9786 22318 9814
rect 22342 9813 22370 9814
rect 22394 9813 22422 9814
rect 22342 9787 22348 9813
rect 22348 9787 22370 9813
rect 22394 9787 22410 9813
rect 22410 9787 22422 9813
rect 22342 9786 22370 9787
rect 22394 9786 22422 9787
rect 22446 9813 22474 9814
rect 22446 9787 22472 9813
rect 22472 9787 22474 9813
rect 22446 9786 22474 9787
rect 22498 9813 22526 9814
rect 22498 9787 22508 9813
rect 22508 9787 22526 9813
rect 22498 9786 22526 9787
rect 23422 10009 23450 10010
rect 23422 9983 23423 10009
rect 23423 9983 23449 10009
rect 23449 9983 23450 10009
rect 23422 9982 23450 9983
rect 23870 9982 23898 10010
rect 22082 9029 22110 9030
rect 22082 9003 22100 9029
rect 22100 9003 22110 9029
rect 22082 9002 22110 9003
rect 22134 9029 22162 9030
rect 22134 9003 22136 9029
rect 22136 9003 22162 9029
rect 22134 9002 22162 9003
rect 22186 9029 22214 9030
rect 22238 9029 22266 9030
rect 22186 9003 22198 9029
rect 22198 9003 22214 9029
rect 22238 9003 22260 9029
rect 22260 9003 22266 9029
rect 22186 9002 22214 9003
rect 22238 9002 22266 9003
rect 22290 9002 22318 9030
rect 22342 9029 22370 9030
rect 22394 9029 22422 9030
rect 22342 9003 22348 9029
rect 22348 9003 22370 9029
rect 22394 9003 22410 9029
rect 22410 9003 22422 9029
rect 22342 9002 22370 9003
rect 22394 9002 22422 9003
rect 22446 9029 22474 9030
rect 22446 9003 22472 9029
rect 22472 9003 22474 9029
rect 22446 9002 22474 9003
rect 22498 9029 22526 9030
rect 22498 9003 22508 9029
rect 22508 9003 22526 9029
rect 22498 9002 22526 9003
rect 23870 9561 23898 9562
rect 23870 9535 23871 9561
rect 23871 9535 23897 9561
rect 23897 9535 23898 9561
rect 23870 9534 23898 9535
rect 22082 8245 22110 8246
rect 22082 8219 22100 8245
rect 22100 8219 22110 8245
rect 22082 8218 22110 8219
rect 22134 8245 22162 8246
rect 22134 8219 22136 8245
rect 22136 8219 22162 8245
rect 22134 8218 22162 8219
rect 22186 8245 22214 8246
rect 22238 8245 22266 8246
rect 22186 8219 22198 8245
rect 22198 8219 22214 8245
rect 22238 8219 22260 8245
rect 22260 8219 22266 8245
rect 22186 8218 22214 8219
rect 22238 8218 22266 8219
rect 22290 8218 22318 8246
rect 22342 8245 22370 8246
rect 22394 8245 22422 8246
rect 22342 8219 22348 8245
rect 22348 8219 22370 8245
rect 22394 8219 22410 8245
rect 22410 8219 22422 8245
rect 22342 8218 22370 8219
rect 22394 8218 22422 8219
rect 22446 8245 22474 8246
rect 22446 8219 22472 8245
rect 22472 8219 22474 8245
rect 22446 8218 22474 8219
rect 22498 8245 22526 8246
rect 22498 8219 22508 8245
rect 22508 8219 22526 8245
rect 22498 8218 22526 8219
rect 23422 8862 23450 8890
rect 23870 8862 23898 8890
rect 20006 7657 20034 7658
rect 20006 7631 20007 7657
rect 20007 7631 20033 7657
rect 20033 7631 20034 7657
rect 20006 7630 20034 7631
rect 20510 7265 20538 7266
rect 20510 7239 20511 7265
rect 20511 7239 20537 7265
rect 20537 7239 20538 7265
rect 20510 7238 20538 7239
rect 21406 7630 21434 7658
rect 20958 7238 20986 7266
rect 19582 7069 19610 7070
rect 19582 7043 19600 7069
rect 19600 7043 19610 7069
rect 19582 7042 19610 7043
rect 19634 7069 19662 7070
rect 19634 7043 19636 7069
rect 19636 7043 19662 7069
rect 19634 7042 19662 7043
rect 19686 7069 19714 7070
rect 19738 7069 19766 7070
rect 19686 7043 19698 7069
rect 19698 7043 19714 7069
rect 19738 7043 19760 7069
rect 19760 7043 19766 7069
rect 19686 7042 19714 7043
rect 19738 7042 19766 7043
rect 19790 7042 19818 7070
rect 19842 7069 19870 7070
rect 19894 7069 19922 7070
rect 19842 7043 19848 7069
rect 19848 7043 19870 7069
rect 19894 7043 19910 7069
rect 19910 7043 19922 7069
rect 19842 7042 19870 7043
rect 19894 7042 19922 7043
rect 19946 7069 19974 7070
rect 19946 7043 19972 7069
rect 19972 7043 19974 7069
rect 19946 7042 19974 7043
rect 19998 7069 20026 7070
rect 19998 7043 20008 7069
rect 20008 7043 20026 7069
rect 19998 7042 20026 7043
rect 20958 6873 20986 6874
rect 20958 6847 20959 6873
rect 20959 6847 20985 6873
rect 20985 6847 20986 6873
rect 20958 6846 20986 6847
rect 21350 7209 21378 7210
rect 21350 7183 21351 7209
rect 21351 7183 21377 7209
rect 21377 7183 21378 7209
rect 21350 7182 21378 7183
rect 19582 6285 19610 6286
rect 19582 6259 19600 6285
rect 19600 6259 19610 6285
rect 19582 6258 19610 6259
rect 19634 6285 19662 6286
rect 19634 6259 19636 6285
rect 19636 6259 19662 6285
rect 19634 6258 19662 6259
rect 19686 6285 19714 6286
rect 19738 6285 19766 6286
rect 19686 6259 19698 6285
rect 19698 6259 19714 6285
rect 19738 6259 19760 6285
rect 19760 6259 19766 6285
rect 19686 6258 19714 6259
rect 19738 6258 19766 6259
rect 19790 6258 19818 6286
rect 19842 6285 19870 6286
rect 19894 6285 19922 6286
rect 19842 6259 19848 6285
rect 19848 6259 19870 6285
rect 19894 6259 19910 6285
rect 19910 6259 19922 6285
rect 19842 6258 19870 6259
rect 19894 6258 19922 6259
rect 19946 6285 19974 6286
rect 19946 6259 19972 6285
rect 19972 6259 19974 6285
rect 19946 6258 19974 6259
rect 19998 6285 20026 6286
rect 19998 6259 20008 6285
rect 20008 6259 20026 6285
rect 19998 6258 20026 6259
rect 19110 6089 19138 6090
rect 19110 6063 19111 6089
rect 19111 6063 19137 6089
rect 19137 6063 19138 6089
rect 19110 6062 19138 6063
rect 18438 5166 18466 5194
rect 18438 5054 18466 5082
rect 19582 5501 19610 5502
rect 19582 5475 19600 5501
rect 19600 5475 19610 5501
rect 19582 5474 19610 5475
rect 19634 5501 19662 5502
rect 19634 5475 19636 5501
rect 19636 5475 19662 5501
rect 19634 5474 19662 5475
rect 19686 5501 19714 5502
rect 19738 5501 19766 5502
rect 19686 5475 19698 5501
rect 19698 5475 19714 5501
rect 19738 5475 19760 5501
rect 19760 5475 19766 5501
rect 19686 5474 19714 5475
rect 19738 5474 19766 5475
rect 19790 5474 19818 5502
rect 19842 5501 19870 5502
rect 19894 5501 19922 5502
rect 19842 5475 19848 5501
rect 19848 5475 19870 5501
rect 19894 5475 19910 5501
rect 19910 5475 19922 5501
rect 19842 5474 19870 5475
rect 19894 5474 19922 5475
rect 19946 5501 19974 5502
rect 19946 5475 19972 5501
rect 19972 5475 19974 5501
rect 19946 5474 19974 5475
rect 19998 5501 20026 5502
rect 19998 5475 20008 5501
rect 20008 5475 20026 5501
rect 19998 5474 20026 5475
rect 20006 5305 20034 5306
rect 20006 5279 20007 5305
rect 20007 5279 20033 5305
rect 20033 5279 20034 5305
rect 20006 5278 20034 5279
rect 20118 5278 20146 5306
rect 19950 5054 19978 5082
rect 18214 2982 18242 3010
rect 19582 4717 19610 4718
rect 19582 4691 19600 4717
rect 19600 4691 19610 4717
rect 19582 4690 19610 4691
rect 19634 4717 19662 4718
rect 19634 4691 19636 4717
rect 19636 4691 19662 4717
rect 19634 4690 19662 4691
rect 19686 4717 19714 4718
rect 19738 4717 19766 4718
rect 19686 4691 19698 4717
rect 19698 4691 19714 4717
rect 19738 4691 19760 4717
rect 19760 4691 19766 4717
rect 19686 4690 19714 4691
rect 19738 4690 19766 4691
rect 19790 4690 19818 4718
rect 19842 4717 19870 4718
rect 19894 4717 19922 4718
rect 19842 4691 19848 4717
rect 19848 4691 19870 4717
rect 19894 4691 19910 4717
rect 19910 4691 19922 4717
rect 19842 4690 19870 4691
rect 19894 4690 19922 4691
rect 19946 4717 19974 4718
rect 19946 4691 19972 4717
rect 19972 4691 19974 4717
rect 19946 4690 19974 4691
rect 19998 4717 20026 4718
rect 19998 4691 20008 4717
rect 20008 4691 20026 4717
rect 19998 4690 20026 4691
rect 19582 3933 19610 3934
rect 19582 3907 19600 3933
rect 19600 3907 19610 3933
rect 19582 3906 19610 3907
rect 19634 3933 19662 3934
rect 19634 3907 19636 3933
rect 19636 3907 19662 3933
rect 19634 3906 19662 3907
rect 19686 3933 19714 3934
rect 19738 3933 19766 3934
rect 19686 3907 19698 3933
rect 19698 3907 19714 3933
rect 19738 3907 19760 3933
rect 19760 3907 19766 3933
rect 19686 3906 19714 3907
rect 19738 3906 19766 3907
rect 19790 3906 19818 3934
rect 19842 3933 19870 3934
rect 19894 3933 19922 3934
rect 19842 3907 19848 3933
rect 19848 3907 19870 3933
rect 19894 3907 19910 3933
rect 19910 3907 19922 3933
rect 19842 3906 19870 3907
rect 19894 3906 19922 3907
rect 19946 3933 19974 3934
rect 19946 3907 19972 3933
rect 19972 3907 19974 3933
rect 19946 3906 19974 3907
rect 19998 3933 20026 3934
rect 19998 3907 20008 3933
rect 20008 3907 20026 3933
rect 19998 3906 20026 3907
rect 20510 6062 20538 6090
rect 21798 7657 21826 7658
rect 21798 7631 21799 7657
rect 21799 7631 21825 7657
rect 21825 7631 21826 7657
rect 21798 7630 21826 7631
rect 22082 7461 22110 7462
rect 22082 7435 22100 7461
rect 22100 7435 22110 7461
rect 22082 7434 22110 7435
rect 22134 7461 22162 7462
rect 22134 7435 22136 7461
rect 22136 7435 22162 7461
rect 22134 7434 22162 7435
rect 22186 7461 22214 7462
rect 22238 7461 22266 7462
rect 22186 7435 22198 7461
rect 22198 7435 22214 7461
rect 22238 7435 22260 7461
rect 22260 7435 22266 7461
rect 22186 7434 22214 7435
rect 22238 7434 22266 7435
rect 22290 7434 22318 7462
rect 22342 7461 22370 7462
rect 22394 7461 22422 7462
rect 22342 7435 22348 7461
rect 22348 7435 22370 7461
rect 22394 7435 22410 7461
rect 22410 7435 22422 7461
rect 22342 7434 22370 7435
rect 22394 7434 22422 7435
rect 22446 7461 22474 7462
rect 22446 7435 22472 7461
rect 22472 7435 22474 7461
rect 22446 7434 22474 7435
rect 22498 7461 22526 7462
rect 22498 7435 22508 7461
rect 22508 7435 22526 7461
rect 22498 7434 22526 7435
rect 23422 8302 23450 8330
rect 22750 7265 22778 7266
rect 22750 7239 22751 7265
rect 22751 7239 22777 7265
rect 22777 7239 22778 7265
rect 22750 7238 22778 7239
rect 21742 7182 21770 7210
rect 23534 7574 23562 7602
rect 23870 7574 23898 7602
rect 22526 6873 22554 6874
rect 22526 6847 22527 6873
rect 22527 6847 22553 6873
rect 22553 6847 22554 6873
rect 22526 6846 22554 6847
rect 22082 6677 22110 6678
rect 22082 6651 22100 6677
rect 22100 6651 22110 6677
rect 22082 6650 22110 6651
rect 22134 6677 22162 6678
rect 22134 6651 22136 6677
rect 22136 6651 22162 6677
rect 22134 6650 22162 6651
rect 22186 6677 22214 6678
rect 22238 6677 22266 6678
rect 22186 6651 22198 6677
rect 22198 6651 22214 6677
rect 22238 6651 22260 6677
rect 22260 6651 22266 6677
rect 22186 6650 22214 6651
rect 22238 6650 22266 6651
rect 22290 6650 22318 6678
rect 22342 6677 22370 6678
rect 22394 6677 22422 6678
rect 22342 6651 22348 6677
rect 22348 6651 22370 6677
rect 22394 6651 22410 6677
rect 22410 6651 22422 6677
rect 22342 6650 22370 6651
rect 22394 6650 22422 6651
rect 22446 6677 22474 6678
rect 22446 6651 22472 6677
rect 22472 6651 22474 6677
rect 22446 6650 22474 6651
rect 22498 6677 22526 6678
rect 22498 6651 22508 6677
rect 22508 6651 22526 6677
rect 22498 6650 22526 6651
rect 22082 5893 22110 5894
rect 22082 5867 22100 5893
rect 22100 5867 22110 5893
rect 22082 5866 22110 5867
rect 22134 5893 22162 5894
rect 22134 5867 22136 5893
rect 22136 5867 22162 5893
rect 22134 5866 22162 5867
rect 22186 5893 22214 5894
rect 22238 5893 22266 5894
rect 22186 5867 22198 5893
rect 22198 5867 22214 5893
rect 22238 5867 22260 5893
rect 22260 5867 22266 5893
rect 22186 5866 22214 5867
rect 22238 5866 22266 5867
rect 22290 5866 22318 5894
rect 22342 5893 22370 5894
rect 22394 5893 22422 5894
rect 22342 5867 22348 5893
rect 22348 5867 22370 5893
rect 22394 5867 22410 5893
rect 22410 5867 22422 5893
rect 22342 5866 22370 5867
rect 22394 5866 22422 5867
rect 22446 5893 22474 5894
rect 22446 5867 22472 5893
rect 22472 5867 22474 5893
rect 22446 5866 22474 5867
rect 22498 5893 22526 5894
rect 22498 5867 22508 5893
rect 22508 5867 22526 5893
rect 22498 5866 22526 5867
rect 21798 5782 21826 5810
rect 21854 5782 21882 5810
rect 21462 5305 21490 5306
rect 21462 5279 21463 5305
rect 21463 5279 21489 5305
rect 21489 5279 21490 5305
rect 21462 5278 21490 5279
rect 21350 4550 21378 4578
rect 20510 4129 20538 4130
rect 20510 4103 20511 4129
rect 20511 4103 20537 4129
rect 20537 4103 20538 4129
rect 20510 4102 20538 4103
rect 19110 3374 19138 3402
rect 20510 3374 20538 3402
rect 17082 2757 17110 2758
rect 17082 2731 17100 2757
rect 17100 2731 17110 2757
rect 17082 2730 17110 2731
rect 17134 2757 17162 2758
rect 17134 2731 17136 2757
rect 17136 2731 17162 2757
rect 17134 2730 17162 2731
rect 17186 2757 17214 2758
rect 17238 2757 17266 2758
rect 17186 2731 17198 2757
rect 17198 2731 17214 2757
rect 17238 2731 17260 2757
rect 17260 2731 17266 2757
rect 17186 2730 17214 2731
rect 17238 2730 17266 2731
rect 17290 2730 17318 2758
rect 17342 2757 17370 2758
rect 17394 2757 17422 2758
rect 17342 2731 17348 2757
rect 17348 2731 17370 2757
rect 17394 2731 17410 2757
rect 17410 2731 17422 2757
rect 17342 2730 17370 2731
rect 17394 2730 17422 2731
rect 17446 2757 17474 2758
rect 17446 2731 17472 2757
rect 17472 2731 17474 2757
rect 17446 2730 17474 2731
rect 17498 2757 17526 2758
rect 17498 2731 17508 2757
rect 17508 2731 17526 2757
rect 17498 2730 17526 2731
rect 16870 2590 16898 2618
rect 16254 2142 16282 2170
rect 15694 1777 15722 1778
rect 15694 1751 15695 1777
rect 15695 1751 15721 1777
rect 15721 1751 15722 1777
rect 15694 1750 15722 1751
rect 19582 3149 19610 3150
rect 19582 3123 19600 3149
rect 19600 3123 19610 3149
rect 19582 3122 19610 3123
rect 19634 3149 19662 3150
rect 19634 3123 19636 3149
rect 19636 3123 19662 3149
rect 19634 3122 19662 3123
rect 19686 3149 19714 3150
rect 19738 3149 19766 3150
rect 19686 3123 19698 3149
rect 19698 3123 19714 3149
rect 19738 3123 19760 3149
rect 19760 3123 19766 3149
rect 19686 3122 19714 3123
rect 19738 3122 19766 3123
rect 19790 3122 19818 3150
rect 19842 3149 19870 3150
rect 19894 3149 19922 3150
rect 19842 3123 19848 3149
rect 19848 3123 19870 3149
rect 19894 3123 19910 3149
rect 19910 3123 19922 3149
rect 19842 3122 19870 3123
rect 19894 3122 19922 3123
rect 19946 3149 19974 3150
rect 19946 3123 19972 3149
rect 19972 3123 19974 3149
rect 19946 3122 19974 3123
rect 19998 3149 20026 3150
rect 19998 3123 20008 3149
rect 20008 3123 20026 3149
rect 19998 3122 20026 3123
rect 20006 2953 20034 2954
rect 20006 2927 20007 2953
rect 20007 2927 20033 2953
rect 20033 2927 20034 2953
rect 20006 2926 20034 2927
rect 18270 2561 18298 2562
rect 18270 2535 18271 2561
rect 18271 2535 18297 2561
rect 18297 2535 18298 2561
rect 18270 2534 18298 2535
rect 17082 1973 17110 1974
rect 17082 1947 17100 1973
rect 17100 1947 17110 1973
rect 17082 1946 17110 1947
rect 17134 1973 17162 1974
rect 17134 1947 17136 1973
rect 17136 1947 17162 1973
rect 17134 1946 17162 1947
rect 17186 1973 17214 1974
rect 17238 1973 17266 1974
rect 17186 1947 17198 1973
rect 17198 1947 17214 1973
rect 17238 1947 17260 1973
rect 17260 1947 17266 1973
rect 17186 1946 17214 1947
rect 17238 1946 17266 1947
rect 17290 1946 17318 1974
rect 17342 1973 17370 1974
rect 17394 1973 17422 1974
rect 17342 1947 17348 1973
rect 17348 1947 17370 1973
rect 17394 1947 17410 1973
rect 17410 1947 17422 1973
rect 17342 1946 17370 1947
rect 17394 1946 17422 1947
rect 17446 1973 17474 1974
rect 17446 1947 17472 1973
rect 17472 1947 17474 1973
rect 17446 1946 17474 1947
rect 17498 1973 17526 1974
rect 17498 1947 17508 1973
rect 17508 1947 17526 1973
rect 17498 1946 17526 1947
rect 18102 2254 18130 2282
rect 19502 2534 19530 2562
rect 20118 2926 20146 2954
rect 19950 2561 19978 2562
rect 19950 2535 19951 2561
rect 19951 2535 19977 2561
rect 19977 2535 19978 2561
rect 19950 2534 19978 2535
rect 20958 4102 20986 4130
rect 20958 3737 20986 3738
rect 20958 3711 20959 3737
rect 20959 3711 20985 3737
rect 20985 3711 20986 3737
rect 20958 3710 20986 3711
rect 21798 4577 21826 4578
rect 21798 4551 21799 4577
rect 21799 4551 21825 4577
rect 21825 4551 21826 4577
rect 21798 4550 21826 4551
rect 22526 5390 22554 5418
rect 23030 5390 23058 5418
rect 22082 5109 22110 5110
rect 22082 5083 22100 5109
rect 22100 5083 22110 5109
rect 22082 5082 22110 5083
rect 22134 5109 22162 5110
rect 22134 5083 22136 5109
rect 22136 5083 22162 5109
rect 22134 5082 22162 5083
rect 22186 5109 22214 5110
rect 22238 5109 22266 5110
rect 22186 5083 22198 5109
rect 22198 5083 22214 5109
rect 22238 5083 22260 5109
rect 22260 5083 22266 5109
rect 22186 5082 22214 5083
rect 22238 5082 22266 5083
rect 22290 5082 22318 5110
rect 22342 5109 22370 5110
rect 22394 5109 22422 5110
rect 22342 5083 22348 5109
rect 22348 5083 22370 5109
rect 22394 5083 22410 5109
rect 22410 5083 22422 5109
rect 22342 5082 22370 5083
rect 22394 5082 22422 5083
rect 22446 5109 22474 5110
rect 22446 5083 22472 5109
rect 22472 5083 22474 5109
rect 22446 5082 22474 5083
rect 22498 5109 22526 5110
rect 22498 5083 22508 5109
rect 22508 5083 22526 5109
rect 22498 5082 22526 5083
rect 21854 4494 21882 4522
rect 22082 4325 22110 4326
rect 22082 4299 22100 4325
rect 22100 4299 22110 4325
rect 22082 4298 22110 4299
rect 22134 4325 22162 4326
rect 22134 4299 22136 4325
rect 22136 4299 22162 4325
rect 22134 4298 22162 4299
rect 22186 4325 22214 4326
rect 22238 4325 22266 4326
rect 22186 4299 22198 4325
rect 22198 4299 22214 4325
rect 22238 4299 22260 4325
rect 22260 4299 22266 4325
rect 22186 4298 22214 4299
rect 22238 4298 22266 4299
rect 22290 4298 22318 4326
rect 22342 4325 22370 4326
rect 22394 4325 22422 4326
rect 22342 4299 22348 4325
rect 22348 4299 22370 4325
rect 22394 4299 22410 4325
rect 22410 4299 22422 4325
rect 22342 4298 22370 4299
rect 22394 4298 22422 4299
rect 22446 4325 22474 4326
rect 22446 4299 22472 4325
rect 22472 4299 22474 4325
rect 22446 4298 22474 4299
rect 22498 4325 22526 4326
rect 22498 4299 22508 4325
rect 22508 4299 22526 4325
rect 22498 4298 22526 4299
rect 22694 4521 22722 4522
rect 22694 4495 22695 4521
rect 22695 4495 22721 4521
rect 22721 4495 22722 4521
rect 22694 4494 22722 4495
rect 22526 3737 22554 3738
rect 22526 3711 22527 3737
rect 22527 3711 22553 3737
rect 22553 3711 22554 3737
rect 22526 3710 22554 3711
rect 23198 6481 23226 6482
rect 23198 6455 23199 6481
rect 23199 6455 23225 6481
rect 23225 6455 23226 6481
rect 23198 6454 23226 6455
rect 23534 6481 23562 6482
rect 23534 6455 23535 6481
rect 23535 6455 23561 6481
rect 23561 6455 23562 6481
rect 23534 6454 23562 6455
rect 23422 5782 23450 5810
rect 23422 5305 23450 5306
rect 23422 5279 23423 5305
rect 23423 5279 23449 5305
rect 23449 5279 23450 5305
rect 23422 5278 23450 5279
rect 23870 5782 23898 5810
rect 23198 4886 23226 4914
rect 22082 3541 22110 3542
rect 22082 3515 22100 3541
rect 22100 3515 22110 3541
rect 22082 3514 22110 3515
rect 22134 3541 22162 3542
rect 22134 3515 22136 3541
rect 22136 3515 22162 3541
rect 22134 3514 22162 3515
rect 22186 3541 22214 3542
rect 22238 3541 22266 3542
rect 22186 3515 22198 3541
rect 22198 3515 22214 3541
rect 22238 3515 22260 3541
rect 22260 3515 22266 3541
rect 22186 3514 22214 3515
rect 22238 3514 22266 3515
rect 22290 3514 22318 3542
rect 22342 3541 22370 3542
rect 22394 3541 22422 3542
rect 22342 3515 22348 3541
rect 22348 3515 22370 3541
rect 22394 3515 22410 3541
rect 22410 3515 22422 3541
rect 22342 3514 22370 3515
rect 22394 3514 22422 3515
rect 22446 3541 22474 3542
rect 22446 3515 22472 3541
rect 22472 3515 22474 3541
rect 22446 3514 22474 3515
rect 22498 3541 22526 3542
rect 22498 3515 22508 3541
rect 22508 3515 22526 3541
rect 22498 3514 22526 3515
rect 22918 4521 22946 4522
rect 22918 4495 22919 4521
rect 22919 4495 22945 4521
rect 22945 4495 22946 4521
rect 22918 4494 22946 4495
rect 23198 4494 23226 4522
rect 23030 3710 23058 3738
rect 21350 2953 21378 2954
rect 21350 2927 21351 2953
rect 21351 2927 21377 2953
rect 21377 2927 21378 2953
rect 21350 2926 21378 2927
rect 22082 2757 22110 2758
rect 22082 2731 22100 2757
rect 22100 2731 22110 2757
rect 22082 2730 22110 2731
rect 22134 2757 22162 2758
rect 22134 2731 22136 2757
rect 22136 2731 22162 2757
rect 22134 2730 22162 2731
rect 22186 2757 22214 2758
rect 22238 2757 22266 2758
rect 22186 2731 22198 2757
rect 22198 2731 22214 2757
rect 22238 2731 22260 2757
rect 22260 2731 22266 2757
rect 22186 2730 22214 2731
rect 22238 2730 22266 2731
rect 22290 2730 22318 2758
rect 22342 2757 22370 2758
rect 22394 2757 22422 2758
rect 22342 2731 22348 2757
rect 22348 2731 22370 2757
rect 22394 2731 22410 2757
rect 22410 2731 22422 2757
rect 22342 2730 22370 2731
rect 22394 2730 22422 2731
rect 22446 2757 22474 2758
rect 22446 2731 22472 2757
rect 22472 2731 22474 2757
rect 22446 2730 22474 2731
rect 22498 2757 22526 2758
rect 22498 2731 22508 2757
rect 22508 2731 22526 2757
rect 22498 2730 22526 2731
rect 21798 2534 21826 2562
rect 19582 2365 19610 2366
rect 19582 2339 19600 2365
rect 19600 2339 19610 2365
rect 19582 2338 19610 2339
rect 19634 2365 19662 2366
rect 19634 2339 19636 2365
rect 19636 2339 19662 2365
rect 19634 2338 19662 2339
rect 19686 2365 19714 2366
rect 19738 2365 19766 2366
rect 19686 2339 19698 2365
rect 19698 2339 19714 2365
rect 19738 2339 19760 2365
rect 19760 2339 19766 2365
rect 19686 2338 19714 2339
rect 19738 2338 19766 2339
rect 19790 2338 19818 2366
rect 19842 2365 19870 2366
rect 19894 2365 19922 2366
rect 19842 2339 19848 2365
rect 19848 2339 19870 2365
rect 19894 2339 19910 2365
rect 19910 2339 19922 2365
rect 19842 2338 19870 2339
rect 19894 2338 19922 2339
rect 19946 2365 19974 2366
rect 19946 2339 19972 2365
rect 19972 2339 19974 2365
rect 19946 2338 19974 2339
rect 19998 2365 20026 2366
rect 19998 2339 20008 2365
rect 20008 2339 20026 2365
rect 19998 2338 20026 2339
rect 19334 2030 19362 2058
rect 19334 1694 19362 1722
rect 18102 1638 18130 1666
rect 20510 2086 20538 2114
rect 20790 2086 20818 2114
rect 21630 2086 21658 2114
rect 20566 1806 20594 1834
rect 19582 1581 19610 1582
rect 19582 1555 19600 1581
rect 19600 1555 19610 1581
rect 19582 1554 19610 1555
rect 19634 1581 19662 1582
rect 19634 1555 19636 1581
rect 19636 1555 19662 1581
rect 19634 1554 19662 1555
rect 19686 1581 19714 1582
rect 19738 1581 19766 1582
rect 19686 1555 19698 1581
rect 19698 1555 19714 1581
rect 19738 1555 19760 1581
rect 19760 1555 19766 1581
rect 19686 1554 19714 1555
rect 19738 1554 19766 1555
rect 19790 1554 19818 1582
rect 19842 1581 19870 1582
rect 19894 1581 19922 1582
rect 19842 1555 19848 1581
rect 19848 1555 19870 1581
rect 19894 1555 19910 1581
rect 19910 1555 19922 1581
rect 19842 1554 19870 1555
rect 19894 1554 19922 1555
rect 19946 1581 19974 1582
rect 19946 1555 19972 1581
rect 19972 1555 19974 1581
rect 19946 1554 19974 1555
rect 19998 1581 20026 1582
rect 19998 1555 20008 1581
rect 20008 1555 20026 1581
rect 19998 1554 20026 1555
rect 22246 2086 22274 2114
rect 22582 2086 22610 2114
rect 22082 1973 22110 1974
rect 22082 1947 22100 1973
rect 22100 1947 22110 1973
rect 22082 1946 22110 1947
rect 22134 1973 22162 1974
rect 22134 1947 22136 1973
rect 22136 1947 22162 1973
rect 22134 1946 22162 1947
rect 22186 1973 22214 1974
rect 22238 1973 22266 1974
rect 22186 1947 22198 1973
rect 22198 1947 22214 1973
rect 22238 1947 22260 1973
rect 22260 1947 22266 1973
rect 22186 1946 22214 1947
rect 22238 1946 22266 1947
rect 22290 1946 22318 1974
rect 22342 1973 22370 1974
rect 22394 1973 22422 1974
rect 22342 1947 22348 1973
rect 22348 1947 22370 1973
rect 22394 1947 22410 1973
rect 22410 1947 22422 1973
rect 22342 1946 22370 1947
rect 22394 1946 22422 1947
rect 22446 1973 22474 1974
rect 22446 1947 22472 1973
rect 22472 1947 22474 1973
rect 22446 1946 22474 1947
rect 22498 1973 22526 1974
rect 22498 1947 22508 1973
rect 22508 1947 22526 1973
rect 22498 1946 22526 1947
rect 22470 1806 22498 1834
rect 23870 3430 23898 3458
rect 23422 2534 23450 2562
rect 24582 17261 24610 17262
rect 24582 17235 24600 17261
rect 24600 17235 24610 17261
rect 24582 17234 24610 17235
rect 24634 17261 24662 17262
rect 24634 17235 24636 17261
rect 24636 17235 24662 17261
rect 24634 17234 24662 17235
rect 24686 17261 24714 17262
rect 24738 17261 24766 17262
rect 24686 17235 24698 17261
rect 24698 17235 24714 17261
rect 24738 17235 24760 17261
rect 24760 17235 24766 17261
rect 24686 17234 24714 17235
rect 24738 17234 24766 17235
rect 24790 17234 24818 17262
rect 24842 17261 24870 17262
rect 24894 17261 24922 17262
rect 24842 17235 24848 17261
rect 24848 17235 24870 17261
rect 24894 17235 24910 17261
rect 24910 17235 24922 17261
rect 24842 17234 24870 17235
rect 24894 17234 24922 17235
rect 24946 17261 24974 17262
rect 24946 17235 24972 17261
rect 24972 17235 24974 17261
rect 24946 17234 24974 17235
rect 24998 17261 25026 17262
rect 24998 17235 25008 17261
rect 25008 17235 25026 17261
rect 24998 17234 25026 17235
rect 24582 16477 24610 16478
rect 24582 16451 24600 16477
rect 24600 16451 24610 16477
rect 24582 16450 24610 16451
rect 24634 16477 24662 16478
rect 24634 16451 24636 16477
rect 24636 16451 24662 16477
rect 24634 16450 24662 16451
rect 24686 16477 24714 16478
rect 24738 16477 24766 16478
rect 24686 16451 24698 16477
rect 24698 16451 24714 16477
rect 24738 16451 24760 16477
rect 24760 16451 24766 16477
rect 24686 16450 24714 16451
rect 24738 16450 24766 16451
rect 24790 16450 24818 16478
rect 24842 16477 24870 16478
rect 24894 16477 24922 16478
rect 24842 16451 24848 16477
rect 24848 16451 24870 16477
rect 24894 16451 24910 16477
rect 24910 16451 24922 16477
rect 24842 16450 24870 16451
rect 24894 16450 24922 16451
rect 24946 16477 24974 16478
rect 24946 16451 24972 16477
rect 24972 16451 24974 16477
rect 24946 16450 24974 16451
rect 24998 16477 25026 16478
rect 24998 16451 25008 16477
rect 25008 16451 25026 16477
rect 24998 16450 25026 16451
rect 24582 15693 24610 15694
rect 24582 15667 24600 15693
rect 24600 15667 24610 15693
rect 24582 15666 24610 15667
rect 24634 15693 24662 15694
rect 24634 15667 24636 15693
rect 24636 15667 24662 15693
rect 24634 15666 24662 15667
rect 24686 15693 24714 15694
rect 24738 15693 24766 15694
rect 24686 15667 24698 15693
rect 24698 15667 24714 15693
rect 24738 15667 24760 15693
rect 24760 15667 24766 15693
rect 24686 15666 24714 15667
rect 24738 15666 24766 15667
rect 24790 15666 24818 15694
rect 24842 15693 24870 15694
rect 24894 15693 24922 15694
rect 24842 15667 24848 15693
rect 24848 15667 24870 15693
rect 24894 15667 24910 15693
rect 24910 15667 24922 15693
rect 24842 15666 24870 15667
rect 24894 15666 24922 15667
rect 24946 15693 24974 15694
rect 24946 15667 24972 15693
rect 24972 15667 24974 15693
rect 24946 15666 24974 15667
rect 24998 15693 25026 15694
rect 24998 15667 25008 15693
rect 25008 15667 25026 15693
rect 24998 15666 25026 15667
rect 24486 15134 24514 15162
rect 24430 13454 24458 13482
rect 27082 18437 27110 18438
rect 27082 18411 27100 18437
rect 27100 18411 27110 18437
rect 27082 18410 27110 18411
rect 27134 18437 27162 18438
rect 27134 18411 27136 18437
rect 27136 18411 27162 18437
rect 27134 18410 27162 18411
rect 27186 18437 27214 18438
rect 27238 18437 27266 18438
rect 27186 18411 27198 18437
rect 27198 18411 27214 18437
rect 27238 18411 27260 18437
rect 27260 18411 27266 18437
rect 27186 18410 27214 18411
rect 27238 18410 27266 18411
rect 27290 18410 27318 18438
rect 27342 18437 27370 18438
rect 27394 18437 27422 18438
rect 27342 18411 27348 18437
rect 27348 18411 27370 18437
rect 27394 18411 27410 18437
rect 27410 18411 27422 18437
rect 27342 18410 27370 18411
rect 27394 18410 27422 18411
rect 27446 18437 27474 18438
rect 27446 18411 27472 18437
rect 27472 18411 27474 18437
rect 27446 18410 27474 18411
rect 27498 18437 27526 18438
rect 27498 18411 27508 18437
rect 27508 18411 27526 18437
rect 27498 18410 27526 18411
rect 29582 18045 29610 18046
rect 29582 18019 29600 18045
rect 29600 18019 29610 18045
rect 29582 18018 29610 18019
rect 29634 18045 29662 18046
rect 29634 18019 29636 18045
rect 29636 18019 29662 18045
rect 29634 18018 29662 18019
rect 29686 18045 29714 18046
rect 29738 18045 29766 18046
rect 29686 18019 29698 18045
rect 29698 18019 29714 18045
rect 29738 18019 29760 18045
rect 29760 18019 29766 18045
rect 29686 18018 29714 18019
rect 29738 18018 29766 18019
rect 29790 18018 29818 18046
rect 29842 18045 29870 18046
rect 29894 18045 29922 18046
rect 29842 18019 29848 18045
rect 29848 18019 29870 18045
rect 29894 18019 29910 18045
rect 29910 18019 29922 18045
rect 29842 18018 29870 18019
rect 29894 18018 29922 18019
rect 29946 18045 29974 18046
rect 29946 18019 29972 18045
rect 29972 18019 29974 18045
rect 29946 18018 29974 18019
rect 29998 18045 30026 18046
rect 29998 18019 30008 18045
rect 30008 18019 30026 18045
rect 29998 18018 30026 18019
rect 27082 17653 27110 17654
rect 27082 17627 27100 17653
rect 27100 17627 27110 17653
rect 27082 17626 27110 17627
rect 27134 17653 27162 17654
rect 27134 17627 27136 17653
rect 27136 17627 27162 17653
rect 27134 17626 27162 17627
rect 27186 17653 27214 17654
rect 27238 17653 27266 17654
rect 27186 17627 27198 17653
rect 27198 17627 27214 17653
rect 27238 17627 27260 17653
rect 27260 17627 27266 17653
rect 27186 17626 27214 17627
rect 27238 17626 27266 17627
rect 27290 17626 27318 17654
rect 27342 17653 27370 17654
rect 27394 17653 27422 17654
rect 27342 17627 27348 17653
rect 27348 17627 27370 17653
rect 27394 17627 27410 17653
rect 27410 17627 27422 17653
rect 27342 17626 27370 17627
rect 27394 17626 27422 17627
rect 27446 17653 27474 17654
rect 27446 17627 27472 17653
rect 27472 17627 27474 17653
rect 27446 17626 27474 17627
rect 27498 17653 27526 17654
rect 27498 17627 27508 17653
rect 27508 17627 27526 17653
rect 27498 17626 27526 17627
rect 29582 17261 29610 17262
rect 29582 17235 29600 17261
rect 29600 17235 29610 17261
rect 29582 17234 29610 17235
rect 29634 17261 29662 17262
rect 29634 17235 29636 17261
rect 29636 17235 29662 17261
rect 29634 17234 29662 17235
rect 29686 17261 29714 17262
rect 29738 17261 29766 17262
rect 29686 17235 29698 17261
rect 29698 17235 29714 17261
rect 29738 17235 29760 17261
rect 29760 17235 29766 17261
rect 29686 17234 29714 17235
rect 29738 17234 29766 17235
rect 29790 17234 29818 17262
rect 29842 17261 29870 17262
rect 29894 17261 29922 17262
rect 29842 17235 29848 17261
rect 29848 17235 29870 17261
rect 29894 17235 29910 17261
rect 29910 17235 29922 17261
rect 29842 17234 29870 17235
rect 29894 17234 29922 17235
rect 29946 17261 29974 17262
rect 29946 17235 29972 17261
rect 29972 17235 29974 17261
rect 29946 17234 29974 17235
rect 29998 17261 30026 17262
rect 29998 17235 30008 17261
rect 30008 17235 30026 17261
rect 29998 17234 30026 17235
rect 27082 16869 27110 16870
rect 27082 16843 27100 16869
rect 27100 16843 27110 16869
rect 27082 16842 27110 16843
rect 27134 16869 27162 16870
rect 27134 16843 27136 16869
rect 27136 16843 27162 16869
rect 27134 16842 27162 16843
rect 27186 16869 27214 16870
rect 27238 16869 27266 16870
rect 27186 16843 27198 16869
rect 27198 16843 27214 16869
rect 27238 16843 27260 16869
rect 27260 16843 27266 16869
rect 27186 16842 27214 16843
rect 27238 16842 27266 16843
rect 27290 16842 27318 16870
rect 27342 16869 27370 16870
rect 27394 16869 27422 16870
rect 27342 16843 27348 16869
rect 27348 16843 27370 16869
rect 27394 16843 27410 16869
rect 27410 16843 27422 16869
rect 27342 16842 27370 16843
rect 27394 16842 27422 16843
rect 27446 16869 27474 16870
rect 27446 16843 27472 16869
rect 27472 16843 27474 16869
rect 27446 16842 27474 16843
rect 27498 16869 27526 16870
rect 27498 16843 27508 16869
rect 27508 16843 27526 16869
rect 27498 16842 27526 16843
rect 29582 16477 29610 16478
rect 29582 16451 29600 16477
rect 29600 16451 29610 16477
rect 29582 16450 29610 16451
rect 29634 16477 29662 16478
rect 29634 16451 29636 16477
rect 29636 16451 29662 16477
rect 29634 16450 29662 16451
rect 29686 16477 29714 16478
rect 29738 16477 29766 16478
rect 29686 16451 29698 16477
rect 29698 16451 29714 16477
rect 29738 16451 29760 16477
rect 29760 16451 29766 16477
rect 29686 16450 29714 16451
rect 29738 16450 29766 16451
rect 29790 16450 29818 16478
rect 29842 16477 29870 16478
rect 29894 16477 29922 16478
rect 29842 16451 29848 16477
rect 29848 16451 29870 16477
rect 29894 16451 29910 16477
rect 29910 16451 29922 16477
rect 29842 16450 29870 16451
rect 29894 16450 29922 16451
rect 29946 16477 29974 16478
rect 29946 16451 29972 16477
rect 29972 16451 29974 16477
rect 29946 16450 29974 16451
rect 29998 16477 30026 16478
rect 29998 16451 30008 16477
rect 30008 16451 30026 16477
rect 29998 16450 30026 16451
rect 27082 16085 27110 16086
rect 27082 16059 27100 16085
rect 27100 16059 27110 16085
rect 27082 16058 27110 16059
rect 27134 16085 27162 16086
rect 27134 16059 27136 16085
rect 27136 16059 27162 16085
rect 27134 16058 27162 16059
rect 27186 16085 27214 16086
rect 27238 16085 27266 16086
rect 27186 16059 27198 16085
rect 27198 16059 27214 16085
rect 27238 16059 27260 16085
rect 27260 16059 27266 16085
rect 27186 16058 27214 16059
rect 27238 16058 27266 16059
rect 27290 16058 27318 16086
rect 27342 16085 27370 16086
rect 27394 16085 27422 16086
rect 27342 16059 27348 16085
rect 27348 16059 27370 16085
rect 27394 16059 27410 16085
rect 27410 16059 27422 16085
rect 27342 16058 27370 16059
rect 27394 16058 27422 16059
rect 27446 16085 27474 16086
rect 27446 16059 27472 16085
rect 27472 16059 27474 16085
rect 27446 16058 27474 16059
rect 27498 16085 27526 16086
rect 27498 16059 27508 16085
rect 27508 16059 27526 16085
rect 27498 16058 27526 16059
rect 29582 15693 29610 15694
rect 29582 15667 29600 15693
rect 29600 15667 29610 15693
rect 29582 15666 29610 15667
rect 29634 15693 29662 15694
rect 29634 15667 29636 15693
rect 29636 15667 29662 15693
rect 29634 15666 29662 15667
rect 29686 15693 29714 15694
rect 29738 15693 29766 15694
rect 29686 15667 29698 15693
rect 29698 15667 29714 15693
rect 29738 15667 29760 15693
rect 29760 15667 29766 15693
rect 29686 15666 29714 15667
rect 29738 15666 29766 15667
rect 29790 15666 29818 15694
rect 29842 15693 29870 15694
rect 29894 15693 29922 15694
rect 29842 15667 29848 15693
rect 29848 15667 29870 15693
rect 29894 15667 29910 15693
rect 29910 15667 29922 15693
rect 29842 15666 29870 15667
rect 29894 15666 29922 15667
rect 29946 15693 29974 15694
rect 29946 15667 29972 15693
rect 29972 15667 29974 15693
rect 29946 15666 29974 15667
rect 29998 15693 30026 15694
rect 29998 15667 30008 15693
rect 30008 15667 30026 15693
rect 29998 15666 30026 15667
rect 27082 15301 27110 15302
rect 27082 15275 27100 15301
rect 27100 15275 27110 15301
rect 27082 15274 27110 15275
rect 27134 15301 27162 15302
rect 27134 15275 27136 15301
rect 27136 15275 27162 15301
rect 27134 15274 27162 15275
rect 27186 15301 27214 15302
rect 27238 15301 27266 15302
rect 27186 15275 27198 15301
rect 27198 15275 27214 15301
rect 27238 15275 27260 15301
rect 27260 15275 27266 15301
rect 27186 15274 27214 15275
rect 27238 15274 27266 15275
rect 27290 15274 27318 15302
rect 27342 15301 27370 15302
rect 27394 15301 27422 15302
rect 27342 15275 27348 15301
rect 27348 15275 27370 15301
rect 27394 15275 27410 15301
rect 27410 15275 27422 15301
rect 27342 15274 27370 15275
rect 27394 15274 27422 15275
rect 27446 15301 27474 15302
rect 27446 15275 27472 15301
rect 27472 15275 27474 15301
rect 27446 15274 27474 15275
rect 27498 15301 27526 15302
rect 27498 15275 27508 15301
rect 27508 15275 27526 15301
rect 27498 15274 27526 15275
rect 26894 15134 26922 15162
rect 24582 14909 24610 14910
rect 24582 14883 24600 14909
rect 24600 14883 24610 14909
rect 24582 14882 24610 14883
rect 24634 14909 24662 14910
rect 24634 14883 24636 14909
rect 24636 14883 24662 14909
rect 24634 14882 24662 14883
rect 24686 14909 24714 14910
rect 24738 14909 24766 14910
rect 24686 14883 24698 14909
rect 24698 14883 24714 14909
rect 24738 14883 24760 14909
rect 24760 14883 24766 14909
rect 24686 14882 24714 14883
rect 24738 14882 24766 14883
rect 24790 14882 24818 14910
rect 24842 14909 24870 14910
rect 24894 14909 24922 14910
rect 24842 14883 24848 14909
rect 24848 14883 24870 14909
rect 24894 14883 24910 14909
rect 24910 14883 24922 14909
rect 24842 14882 24870 14883
rect 24894 14882 24922 14883
rect 24946 14909 24974 14910
rect 24946 14883 24972 14909
rect 24972 14883 24974 14909
rect 24946 14882 24974 14883
rect 24998 14909 25026 14910
rect 24998 14883 25008 14909
rect 25008 14883 25026 14909
rect 24998 14882 25026 14883
rect 29582 14909 29610 14910
rect 29582 14883 29600 14909
rect 29600 14883 29610 14909
rect 29582 14882 29610 14883
rect 29634 14909 29662 14910
rect 29634 14883 29636 14909
rect 29636 14883 29662 14909
rect 29634 14882 29662 14883
rect 29686 14909 29714 14910
rect 29738 14909 29766 14910
rect 29686 14883 29698 14909
rect 29698 14883 29714 14909
rect 29738 14883 29760 14909
rect 29760 14883 29766 14909
rect 29686 14882 29714 14883
rect 29738 14882 29766 14883
rect 29790 14882 29818 14910
rect 29842 14909 29870 14910
rect 29894 14909 29922 14910
rect 29842 14883 29848 14909
rect 29848 14883 29870 14909
rect 29894 14883 29910 14909
rect 29910 14883 29922 14909
rect 29842 14882 29870 14883
rect 29894 14882 29922 14883
rect 29946 14909 29974 14910
rect 29946 14883 29972 14909
rect 29972 14883 29974 14909
rect 29946 14882 29974 14883
rect 29998 14909 30026 14910
rect 29998 14883 30008 14909
rect 30008 14883 30026 14909
rect 29998 14882 30026 14883
rect 27082 14517 27110 14518
rect 27082 14491 27100 14517
rect 27100 14491 27110 14517
rect 27082 14490 27110 14491
rect 27134 14517 27162 14518
rect 27134 14491 27136 14517
rect 27136 14491 27162 14517
rect 27134 14490 27162 14491
rect 27186 14517 27214 14518
rect 27238 14517 27266 14518
rect 27186 14491 27198 14517
rect 27198 14491 27214 14517
rect 27238 14491 27260 14517
rect 27260 14491 27266 14517
rect 27186 14490 27214 14491
rect 27238 14490 27266 14491
rect 27290 14490 27318 14518
rect 27342 14517 27370 14518
rect 27394 14517 27422 14518
rect 27342 14491 27348 14517
rect 27348 14491 27370 14517
rect 27394 14491 27410 14517
rect 27410 14491 27422 14517
rect 27342 14490 27370 14491
rect 27394 14490 27422 14491
rect 27446 14517 27474 14518
rect 27446 14491 27472 14517
rect 27472 14491 27474 14517
rect 27446 14490 27474 14491
rect 27498 14517 27526 14518
rect 27498 14491 27508 14517
rect 27508 14491 27526 14517
rect 27498 14490 27526 14491
rect 25158 14238 25186 14266
rect 24582 14125 24610 14126
rect 24582 14099 24600 14125
rect 24600 14099 24610 14125
rect 24582 14098 24610 14099
rect 24634 14125 24662 14126
rect 24634 14099 24636 14125
rect 24636 14099 24662 14125
rect 24634 14098 24662 14099
rect 24686 14125 24714 14126
rect 24738 14125 24766 14126
rect 24686 14099 24698 14125
rect 24698 14099 24714 14125
rect 24738 14099 24760 14125
rect 24760 14099 24766 14125
rect 24686 14098 24714 14099
rect 24738 14098 24766 14099
rect 24790 14098 24818 14126
rect 24842 14125 24870 14126
rect 24894 14125 24922 14126
rect 24842 14099 24848 14125
rect 24848 14099 24870 14125
rect 24894 14099 24910 14125
rect 24910 14099 24922 14125
rect 24842 14098 24870 14099
rect 24894 14098 24922 14099
rect 24946 14125 24974 14126
rect 24946 14099 24972 14125
rect 24972 14099 24974 14125
rect 24946 14098 24974 14099
rect 24998 14125 25026 14126
rect 24998 14099 25008 14125
rect 25008 14099 25026 14125
rect 24998 14098 25026 14099
rect 29582 14125 29610 14126
rect 29582 14099 29600 14125
rect 29600 14099 29610 14125
rect 29582 14098 29610 14099
rect 29634 14125 29662 14126
rect 29634 14099 29636 14125
rect 29636 14099 29662 14125
rect 29634 14098 29662 14099
rect 29686 14125 29714 14126
rect 29738 14125 29766 14126
rect 29686 14099 29698 14125
rect 29698 14099 29714 14125
rect 29738 14099 29760 14125
rect 29760 14099 29766 14125
rect 29686 14098 29714 14099
rect 29738 14098 29766 14099
rect 29790 14098 29818 14126
rect 29842 14125 29870 14126
rect 29894 14125 29922 14126
rect 29842 14099 29848 14125
rect 29848 14099 29870 14125
rect 29894 14099 29910 14125
rect 29910 14099 29922 14125
rect 29842 14098 29870 14099
rect 29894 14098 29922 14099
rect 29946 14125 29974 14126
rect 29946 14099 29972 14125
rect 29972 14099 29974 14125
rect 29946 14098 29974 14099
rect 29998 14125 30026 14126
rect 29998 14099 30008 14125
rect 30008 14099 30026 14125
rect 29998 14098 30026 14099
rect 24486 13398 24514 13426
rect 24582 13341 24610 13342
rect 24374 12334 24402 12362
rect 24430 13286 24458 13314
rect 24582 13315 24600 13341
rect 24600 13315 24610 13341
rect 24582 13314 24610 13315
rect 24634 13341 24662 13342
rect 24634 13315 24636 13341
rect 24636 13315 24662 13341
rect 24634 13314 24662 13315
rect 24686 13341 24714 13342
rect 24738 13341 24766 13342
rect 24686 13315 24698 13341
rect 24698 13315 24714 13341
rect 24738 13315 24760 13341
rect 24760 13315 24766 13341
rect 24686 13314 24714 13315
rect 24738 13314 24766 13315
rect 24790 13314 24818 13342
rect 24842 13341 24870 13342
rect 24894 13341 24922 13342
rect 24842 13315 24848 13341
rect 24848 13315 24870 13341
rect 24894 13315 24910 13341
rect 24910 13315 24922 13341
rect 24842 13314 24870 13315
rect 24894 13314 24922 13315
rect 24946 13341 24974 13342
rect 24946 13315 24972 13341
rect 24972 13315 24974 13341
rect 24946 13314 24974 13315
rect 24998 13341 25026 13342
rect 24998 13315 25008 13341
rect 25008 13315 25026 13341
rect 24998 13314 25026 13315
rect 24582 12557 24610 12558
rect 24582 12531 24600 12557
rect 24600 12531 24610 12557
rect 24582 12530 24610 12531
rect 24634 12557 24662 12558
rect 24634 12531 24636 12557
rect 24636 12531 24662 12557
rect 24634 12530 24662 12531
rect 24686 12557 24714 12558
rect 24738 12557 24766 12558
rect 24686 12531 24698 12557
rect 24698 12531 24714 12557
rect 24738 12531 24760 12557
rect 24760 12531 24766 12557
rect 24686 12530 24714 12531
rect 24738 12530 24766 12531
rect 24790 12530 24818 12558
rect 24842 12557 24870 12558
rect 24894 12557 24922 12558
rect 24842 12531 24848 12557
rect 24848 12531 24870 12557
rect 24894 12531 24910 12557
rect 24910 12531 24922 12557
rect 24842 12530 24870 12531
rect 24894 12530 24922 12531
rect 24946 12557 24974 12558
rect 24946 12531 24972 12557
rect 24972 12531 24974 12557
rect 24946 12530 24974 12531
rect 24998 12557 25026 12558
rect 24998 12531 25008 12557
rect 25008 12531 25026 12557
rect 24998 12530 25026 12531
rect 24486 12334 24514 12362
rect 24766 12361 24794 12362
rect 24766 12335 24767 12361
rect 24767 12335 24793 12361
rect 24793 12335 24794 12361
rect 24766 12334 24794 12335
rect 27082 13733 27110 13734
rect 27082 13707 27100 13733
rect 27100 13707 27110 13733
rect 27082 13706 27110 13707
rect 27134 13733 27162 13734
rect 27134 13707 27136 13733
rect 27136 13707 27162 13733
rect 27134 13706 27162 13707
rect 27186 13733 27214 13734
rect 27238 13733 27266 13734
rect 27186 13707 27198 13733
rect 27198 13707 27214 13733
rect 27238 13707 27260 13733
rect 27260 13707 27266 13733
rect 27186 13706 27214 13707
rect 27238 13706 27266 13707
rect 27290 13706 27318 13734
rect 27342 13733 27370 13734
rect 27394 13733 27422 13734
rect 27342 13707 27348 13733
rect 27348 13707 27370 13733
rect 27394 13707 27410 13733
rect 27410 13707 27422 13733
rect 27342 13706 27370 13707
rect 27394 13706 27422 13707
rect 27446 13733 27474 13734
rect 27446 13707 27472 13733
rect 27472 13707 27474 13733
rect 27446 13706 27474 13707
rect 27498 13733 27526 13734
rect 27498 13707 27508 13733
rect 27508 13707 27526 13733
rect 27498 13706 27526 13707
rect 25102 12334 25130 12362
rect 25158 12697 25186 12698
rect 25158 12671 25159 12697
rect 25159 12671 25185 12697
rect 25185 12671 25186 12697
rect 25158 12670 25186 12671
rect 25102 11942 25130 11970
rect 24582 11773 24610 11774
rect 24582 11747 24600 11773
rect 24600 11747 24610 11773
rect 24582 11746 24610 11747
rect 24634 11773 24662 11774
rect 24634 11747 24636 11773
rect 24636 11747 24662 11773
rect 24634 11746 24662 11747
rect 24686 11773 24714 11774
rect 24738 11773 24766 11774
rect 24686 11747 24698 11773
rect 24698 11747 24714 11773
rect 24738 11747 24760 11773
rect 24760 11747 24766 11773
rect 24686 11746 24714 11747
rect 24738 11746 24766 11747
rect 24790 11746 24818 11774
rect 24842 11773 24870 11774
rect 24894 11773 24922 11774
rect 24842 11747 24848 11773
rect 24848 11747 24870 11773
rect 24894 11747 24910 11773
rect 24910 11747 24922 11773
rect 24842 11746 24870 11747
rect 24894 11746 24922 11747
rect 24946 11773 24974 11774
rect 24946 11747 24972 11773
rect 24972 11747 24974 11773
rect 24946 11746 24974 11747
rect 24998 11773 25026 11774
rect 24998 11747 25008 11773
rect 25008 11747 25026 11773
rect 24998 11746 25026 11747
rect 24582 10989 24610 10990
rect 24582 10963 24600 10989
rect 24600 10963 24610 10989
rect 24582 10962 24610 10963
rect 24634 10989 24662 10990
rect 24634 10963 24636 10989
rect 24636 10963 24662 10989
rect 24634 10962 24662 10963
rect 24686 10989 24714 10990
rect 24738 10989 24766 10990
rect 24686 10963 24698 10989
rect 24698 10963 24714 10989
rect 24738 10963 24760 10989
rect 24760 10963 24766 10989
rect 24686 10962 24714 10963
rect 24738 10962 24766 10963
rect 24790 10962 24818 10990
rect 24842 10989 24870 10990
rect 24894 10989 24922 10990
rect 24842 10963 24848 10989
rect 24848 10963 24870 10989
rect 24894 10963 24910 10989
rect 24910 10963 24922 10989
rect 24842 10962 24870 10963
rect 24894 10962 24922 10963
rect 24946 10989 24974 10990
rect 24946 10963 24972 10989
rect 24972 10963 24974 10989
rect 24946 10962 24974 10963
rect 24998 10989 25026 10990
rect 24998 10963 25008 10989
rect 25008 10963 25026 10989
rect 24998 10962 25026 10963
rect 29582 13341 29610 13342
rect 29582 13315 29600 13341
rect 29600 13315 29610 13341
rect 29582 13314 29610 13315
rect 29634 13341 29662 13342
rect 29634 13315 29636 13341
rect 29636 13315 29662 13341
rect 29634 13314 29662 13315
rect 29686 13341 29714 13342
rect 29738 13341 29766 13342
rect 29686 13315 29698 13341
rect 29698 13315 29714 13341
rect 29738 13315 29760 13341
rect 29760 13315 29766 13341
rect 29686 13314 29714 13315
rect 29738 13314 29766 13315
rect 29790 13314 29818 13342
rect 29842 13341 29870 13342
rect 29894 13341 29922 13342
rect 29842 13315 29848 13341
rect 29848 13315 29870 13341
rect 29894 13315 29910 13341
rect 29910 13315 29922 13341
rect 29842 13314 29870 13315
rect 29894 13314 29922 13315
rect 29946 13341 29974 13342
rect 29946 13315 29972 13341
rect 29972 13315 29974 13341
rect 29946 13314 29974 13315
rect 29998 13341 30026 13342
rect 29998 13315 30008 13341
rect 30008 13315 30026 13341
rect 29998 13314 30026 13315
rect 25214 12222 25242 12250
rect 27082 12949 27110 12950
rect 27082 12923 27100 12949
rect 27100 12923 27110 12949
rect 27082 12922 27110 12923
rect 27134 12949 27162 12950
rect 27134 12923 27136 12949
rect 27136 12923 27162 12949
rect 27134 12922 27162 12923
rect 27186 12949 27214 12950
rect 27238 12949 27266 12950
rect 27186 12923 27198 12949
rect 27198 12923 27214 12949
rect 27238 12923 27260 12949
rect 27260 12923 27266 12949
rect 27186 12922 27214 12923
rect 27238 12922 27266 12923
rect 27290 12922 27318 12950
rect 27342 12949 27370 12950
rect 27394 12949 27422 12950
rect 27342 12923 27348 12949
rect 27348 12923 27370 12949
rect 27394 12923 27410 12949
rect 27410 12923 27422 12949
rect 27342 12922 27370 12923
rect 27394 12922 27422 12923
rect 27446 12949 27474 12950
rect 27446 12923 27472 12949
rect 27472 12923 27474 12949
rect 27446 12922 27474 12923
rect 27498 12949 27526 12950
rect 27498 12923 27508 12949
rect 27508 12923 27526 12949
rect 27498 12922 27526 12923
rect 25942 12417 25970 12418
rect 25942 12391 25943 12417
rect 25943 12391 25969 12417
rect 25969 12391 25970 12417
rect 25942 12390 25970 12391
rect 26502 12361 26530 12362
rect 26502 12335 26503 12361
rect 26503 12335 26529 12361
rect 26529 12335 26530 12361
rect 26502 12334 26530 12335
rect 25942 12222 25970 12250
rect 27398 12361 27426 12362
rect 27398 12335 27399 12361
rect 27399 12335 27425 12361
rect 27425 12335 27426 12361
rect 27398 12334 27426 12335
rect 27678 12334 27706 12362
rect 27082 12165 27110 12166
rect 27082 12139 27100 12165
rect 27100 12139 27110 12165
rect 27082 12138 27110 12139
rect 27134 12165 27162 12166
rect 27134 12139 27136 12165
rect 27136 12139 27162 12165
rect 27134 12138 27162 12139
rect 27186 12165 27214 12166
rect 27238 12165 27266 12166
rect 27186 12139 27198 12165
rect 27198 12139 27214 12165
rect 27238 12139 27260 12165
rect 27260 12139 27266 12165
rect 27186 12138 27214 12139
rect 27238 12138 27266 12139
rect 27290 12138 27318 12166
rect 27342 12165 27370 12166
rect 27394 12165 27422 12166
rect 27342 12139 27348 12165
rect 27348 12139 27370 12165
rect 27394 12139 27410 12165
rect 27410 12139 27422 12165
rect 27342 12138 27370 12139
rect 27394 12138 27422 12139
rect 27446 12165 27474 12166
rect 27446 12139 27472 12165
rect 27472 12139 27474 12165
rect 27446 12138 27474 12139
rect 27498 12165 27526 12166
rect 27498 12139 27508 12165
rect 27508 12139 27526 12165
rect 27498 12138 27526 12139
rect 27678 11969 27706 11970
rect 27678 11943 27679 11969
rect 27679 11943 27705 11969
rect 27705 11943 27706 11969
rect 27678 11942 27706 11943
rect 25158 11550 25186 11578
rect 25214 11577 25242 11578
rect 25214 11551 25215 11577
rect 25215 11551 25241 11577
rect 25241 11551 25242 11577
rect 25214 11550 25242 11551
rect 25158 11185 25186 11186
rect 25158 11159 25159 11185
rect 25159 11159 25185 11185
rect 25185 11159 25186 11185
rect 25158 11158 25186 11159
rect 24374 10318 24402 10346
rect 24430 10262 24458 10290
rect 24582 10205 24610 10206
rect 24582 10179 24600 10205
rect 24600 10179 24610 10205
rect 24582 10178 24610 10179
rect 24634 10205 24662 10206
rect 24634 10179 24636 10205
rect 24636 10179 24662 10205
rect 24634 10178 24662 10179
rect 24686 10205 24714 10206
rect 24738 10205 24766 10206
rect 24686 10179 24698 10205
rect 24698 10179 24714 10205
rect 24738 10179 24760 10205
rect 24760 10179 24766 10205
rect 24686 10178 24714 10179
rect 24738 10178 24766 10179
rect 24790 10178 24818 10206
rect 24842 10205 24870 10206
rect 24894 10205 24922 10206
rect 24842 10179 24848 10205
rect 24848 10179 24870 10205
rect 24894 10179 24910 10205
rect 24910 10179 24922 10205
rect 24842 10178 24870 10179
rect 24894 10178 24922 10179
rect 24946 10205 24974 10206
rect 24946 10179 24972 10205
rect 24972 10179 24974 10205
rect 24946 10178 24974 10179
rect 24998 10205 25026 10206
rect 24998 10179 25008 10205
rect 25008 10179 25026 10205
rect 24998 10178 25026 10179
rect 24582 9421 24610 9422
rect 24582 9395 24600 9421
rect 24600 9395 24610 9421
rect 24582 9394 24610 9395
rect 24634 9421 24662 9422
rect 24634 9395 24636 9421
rect 24636 9395 24662 9421
rect 24634 9394 24662 9395
rect 24686 9421 24714 9422
rect 24738 9421 24766 9422
rect 24686 9395 24698 9421
rect 24698 9395 24714 9421
rect 24738 9395 24760 9421
rect 24760 9395 24766 9421
rect 24686 9394 24714 9395
rect 24738 9394 24766 9395
rect 24790 9394 24818 9422
rect 24842 9421 24870 9422
rect 24894 9421 24922 9422
rect 24842 9395 24848 9421
rect 24848 9395 24870 9421
rect 24894 9395 24910 9421
rect 24910 9395 24922 9421
rect 24842 9394 24870 9395
rect 24894 9394 24922 9395
rect 24946 9421 24974 9422
rect 24946 9395 24972 9421
rect 24972 9395 24974 9421
rect 24946 9394 24974 9395
rect 24998 9421 25026 9422
rect 24998 9395 25008 9421
rect 25008 9395 25026 9421
rect 24998 9394 25026 9395
rect 24430 8358 24458 8386
rect 24582 8637 24610 8638
rect 24582 8611 24600 8637
rect 24600 8611 24610 8637
rect 24582 8610 24610 8611
rect 24634 8637 24662 8638
rect 24634 8611 24636 8637
rect 24636 8611 24662 8637
rect 24634 8610 24662 8611
rect 24686 8637 24714 8638
rect 24738 8637 24766 8638
rect 24686 8611 24698 8637
rect 24698 8611 24714 8637
rect 24738 8611 24760 8637
rect 24760 8611 24766 8637
rect 24686 8610 24714 8611
rect 24738 8610 24766 8611
rect 24790 8610 24818 8638
rect 24842 8637 24870 8638
rect 24894 8637 24922 8638
rect 24842 8611 24848 8637
rect 24848 8611 24870 8637
rect 24894 8611 24910 8637
rect 24910 8611 24922 8637
rect 24842 8610 24870 8611
rect 24894 8610 24922 8611
rect 24946 8637 24974 8638
rect 24946 8611 24972 8637
rect 24972 8611 24974 8637
rect 24946 8610 24974 8611
rect 24998 8637 25026 8638
rect 24998 8611 25008 8637
rect 25008 8611 25026 8637
rect 24998 8610 25026 8611
rect 24582 7853 24610 7854
rect 24582 7827 24600 7853
rect 24600 7827 24610 7853
rect 24582 7826 24610 7827
rect 24634 7853 24662 7854
rect 24634 7827 24636 7853
rect 24636 7827 24662 7853
rect 24634 7826 24662 7827
rect 24686 7853 24714 7854
rect 24738 7853 24766 7854
rect 24686 7827 24698 7853
rect 24698 7827 24714 7853
rect 24738 7827 24760 7853
rect 24760 7827 24766 7853
rect 24686 7826 24714 7827
rect 24738 7826 24766 7827
rect 24790 7826 24818 7854
rect 24842 7853 24870 7854
rect 24894 7853 24922 7854
rect 24842 7827 24848 7853
rect 24848 7827 24870 7853
rect 24894 7827 24910 7853
rect 24910 7827 24922 7853
rect 24842 7826 24870 7827
rect 24894 7826 24922 7827
rect 24946 7853 24974 7854
rect 24946 7827 24972 7853
rect 24972 7827 24974 7853
rect 24946 7826 24974 7827
rect 24998 7853 25026 7854
rect 24998 7827 25008 7853
rect 25008 7827 25026 7853
rect 24998 7826 25026 7827
rect 24654 7574 24682 7602
rect 24374 7518 24402 7546
rect 24374 7265 24402 7266
rect 24374 7239 24375 7265
rect 24375 7239 24401 7265
rect 24401 7239 24402 7265
rect 24374 7238 24402 7239
rect 25438 11577 25466 11578
rect 25438 11551 25439 11577
rect 25439 11551 25465 11577
rect 25465 11551 25466 11577
rect 25438 11550 25466 11551
rect 28574 11886 28602 11914
rect 29358 11913 29386 11914
rect 29358 11887 29359 11913
rect 29359 11887 29385 11913
rect 29385 11887 29386 11913
rect 29358 11886 29386 11887
rect 28350 11577 28378 11578
rect 28350 11551 28351 11577
rect 28351 11551 28377 11577
rect 28377 11551 28378 11577
rect 28350 11550 28378 11551
rect 27082 11381 27110 11382
rect 27082 11355 27100 11381
rect 27100 11355 27110 11381
rect 27082 11354 27110 11355
rect 27134 11381 27162 11382
rect 27134 11355 27136 11381
rect 27136 11355 27162 11381
rect 27134 11354 27162 11355
rect 27186 11381 27214 11382
rect 27238 11381 27266 11382
rect 27186 11355 27198 11381
rect 27198 11355 27214 11381
rect 27238 11355 27260 11381
rect 27260 11355 27266 11381
rect 27186 11354 27214 11355
rect 27238 11354 27266 11355
rect 27290 11354 27318 11382
rect 27342 11381 27370 11382
rect 27394 11381 27422 11382
rect 27342 11355 27348 11381
rect 27348 11355 27370 11381
rect 27394 11355 27410 11381
rect 27410 11355 27422 11381
rect 27342 11354 27370 11355
rect 27394 11354 27422 11355
rect 27446 11381 27474 11382
rect 27446 11355 27472 11381
rect 27472 11355 27474 11381
rect 27446 11354 27474 11355
rect 27498 11381 27526 11382
rect 27498 11355 27508 11381
rect 27508 11355 27526 11381
rect 27498 11354 27526 11355
rect 25214 8862 25242 8890
rect 27082 10597 27110 10598
rect 27082 10571 27100 10597
rect 27100 10571 27110 10597
rect 27082 10570 27110 10571
rect 27134 10597 27162 10598
rect 27134 10571 27136 10597
rect 27136 10571 27162 10597
rect 27134 10570 27162 10571
rect 27186 10597 27214 10598
rect 27238 10597 27266 10598
rect 27186 10571 27198 10597
rect 27198 10571 27214 10597
rect 27238 10571 27260 10597
rect 27260 10571 27266 10597
rect 27186 10570 27214 10571
rect 27238 10570 27266 10571
rect 27290 10570 27318 10598
rect 27342 10597 27370 10598
rect 27394 10597 27422 10598
rect 27342 10571 27348 10597
rect 27348 10571 27370 10597
rect 27394 10571 27410 10597
rect 27410 10571 27422 10597
rect 27342 10570 27370 10571
rect 27394 10570 27422 10571
rect 27446 10597 27474 10598
rect 27446 10571 27472 10597
rect 27472 10571 27474 10597
rect 27446 10570 27474 10571
rect 27498 10597 27526 10598
rect 27498 10571 27508 10597
rect 27508 10571 27526 10597
rect 27498 10570 27526 10571
rect 25942 10065 25970 10066
rect 25942 10039 25943 10065
rect 25943 10039 25969 10065
rect 25969 10039 25970 10065
rect 25942 10038 25970 10039
rect 26838 10009 26866 10010
rect 26838 9983 26839 10009
rect 26839 9983 26865 10009
rect 26865 9983 26866 10009
rect 26838 9982 26866 9983
rect 28070 10878 28098 10906
rect 27566 9982 27594 10010
rect 27678 10401 27706 10402
rect 27678 10375 27679 10401
rect 27679 10375 27705 10401
rect 27705 10375 27706 10401
rect 27678 10374 27706 10375
rect 27082 9813 27110 9814
rect 27082 9787 27100 9813
rect 27100 9787 27110 9813
rect 27082 9786 27110 9787
rect 27134 9813 27162 9814
rect 27134 9787 27136 9813
rect 27136 9787 27162 9813
rect 27134 9786 27162 9787
rect 27186 9813 27214 9814
rect 27238 9813 27266 9814
rect 27186 9787 27198 9813
rect 27198 9787 27214 9813
rect 27238 9787 27260 9813
rect 27260 9787 27266 9813
rect 27186 9786 27214 9787
rect 27238 9786 27266 9787
rect 27290 9786 27318 9814
rect 27342 9813 27370 9814
rect 27394 9813 27422 9814
rect 27342 9787 27348 9813
rect 27348 9787 27370 9813
rect 27394 9787 27410 9813
rect 27410 9787 27422 9813
rect 27342 9786 27370 9787
rect 27394 9786 27422 9787
rect 27446 9813 27474 9814
rect 27446 9787 27472 9813
rect 27472 9787 27474 9813
rect 27446 9786 27474 9787
rect 27498 9813 27526 9814
rect 27498 9787 27508 9813
rect 27508 9787 27526 9813
rect 27498 9786 27526 9787
rect 25382 9561 25410 9562
rect 25382 9535 25383 9561
rect 25383 9535 25409 9561
rect 25409 9535 25410 9561
rect 25382 9534 25410 9535
rect 25158 8358 25186 8386
rect 25382 8302 25410 8330
rect 28350 10878 28378 10906
rect 29582 12557 29610 12558
rect 29582 12531 29600 12557
rect 29600 12531 29610 12557
rect 29582 12530 29610 12531
rect 29634 12557 29662 12558
rect 29634 12531 29636 12557
rect 29636 12531 29662 12557
rect 29634 12530 29662 12531
rect 29686 12557 29714 12558
rect 29738 12557 29766 12558
rect 29686 12531 29698 12557
rect 29698 12531 29714 12557
rect 29738 12531 29760 12557
rect 29760 12531 29766 12557
rect 29686 12530 29714 12531
rect 29738 12530 29766 12531
rect 29790 12530 29818 12558
rect 29842 12557 29870 12558
rect 29894 12557 29922 12558
rect 29842 12531 29848 12557
rect 29848 12531 29870 12557
rect 29894 12531 29910 12557
rect 29910 12531 29922 12557
rect 29842 12530 29870 12531
rect 29894 12530 29922 12531
rect 29946 12557 29974 12558
rect 29946 12531 29972 12557
rect 29972 12531 29974 12557
rect 29946 12530 29974 12531
rect 29998 12557 30026 12558
rect 29998 12531 30008 12557
rect 30008 12531 30026 12557
rect 29998 12530 30026 12531
rect 30198 12334 30226 12362
rect 30366 12361 30394 12362
rect 30366 12335 30367 12361
rect 30367 12335 30393 12361
rect 30393 12335 30394 12361
rect 30366 12334 30394 12335
rect 30702 12361 30730 12362
rect 30702 12335 30703 12361
rect 30703 12335 30729 12361
rect 30729 12335 30730 12361
rect 30702 12334 30730 12335
rect 29918 11886 29946 11914
rect 29582 11773 29610 11774
rect 29582 11747 29600 11773
rect 29600 11747 29610 11773
rect 29582 11746 29610 11747
rect 29634 11773 29662 11774
rect 29634 11747 29636 11773
rect 29636 11747 29662 11773
rect 29634 11746 29662 11747
rect 29686 11773 29714 11774
rect 29738 11773 29766 11774
rect 29686 11747 29698 11773
rect 29698 11747 29714 11773
rect 29738 11747 29760 11773
rect 29760 11747 29766 11773
rect 29686 11746 29714 11747
rect 29738 11746 29766 11747
rect 29790 11746 29818 11774
rect 29842 11773 29870 11774
rect 29894 11773 29922 11774
rect 29842 11747 29848 11773
rect 29848 11747 29870 11773
rect 29894 11747 29910 11773
rect 29910 11747 29922 11773
rect 29842 11746 29870 11747
rect 29894 11746 29922 11747
rect 29946 11773 29974 11774
rect 29946 11747 29972 11773
rect 29972 11747 29974 11773
rect 29946 11746 29974 11747
rect 29998 11773 30026 11774
rect 29998 11747 30008 11773
rect 30008 11747 30026 11773
rect 29998 11746 30026 11747
rect 29414 11577 29442 11578
rect 29414 11551 29415 11577
rect 29415 11551 29441 11577
rect 29441 11551 29442 11577
rect 29414 11550 29442 11551
rect 28070 10401 28098 10402
rect 28070 10375 28071 10401
rect 28071 10375 28097 10401
rect 28097 10375 28098 10401
rect 28070 10374 28098 10375
rect 27678 10038 27706 10066
rect 27902 10038 27930 10066
rect 28406 10038 28434 10066
rect 25942 8302 25970 8330
rect 25158 7630 25186 7658
rect 26222 8358 26250 8386
rect 26222 8022 26250 8050
rect 26726 8049 26754 8050
rect 26726 8023 26727 8049
rect 26727 8023 26753 8049
rect 26753 8023 26754 8049
rect 26726 8022 26754 8023
rect 25942 7574 25970 7602
rect 24766 7518 24794 7546
rect 24582 7069 24610 7070
rect 24582 7043 24600 7069
rect 24600 7043 24610 7069
rect 24582 7042 24610 7043
rect 24634 7069 24662 7070
rect 24634 7043 24636 7069
rect 24636 7043 24662 7069
rect 24634 7042 24662 7043
rect 24686 7069 24714 7070
rect 24738 7069 24766 7070
rect 24686 7043 24698 7069
rect 24698 7043 24714 7069
rect 24738 7043 24760 7069
rect 24760 7043 24766 7069
rect 24686 7042 24714 7043
rect 24738 7042 24766 7043
rect 24790 7042 24818 7070
rect 24842 7069 24870 7070
rect 24894 7069 24922 7070
rect 24842 7043 24848 7069
rect 24848 7043 24870 7069
rect 24894 7043 24910 7069
rect 24910 7043 24922 7069
rect 24842 7042 24870 7043
rect 24894 7042 24922 7043
rect 24946 7069 24974 7070
rect 24946 7043 24972 7069
rect 24972 7043 24974 7069
rect 24946 7042 24974 7043
rect 24998 7069 25026 7070
rect 24998 7043 25008 7069
rect 25008 7043 25026 7069
rect 24998 7042 25026 7043
rect 23926 2590 23954 2618
rect 24262 3374 24290 3402
rect 24582 6285 24610 6286
rect 24582 6259 24600 6285
rect 24600 6259 24610 6285
rect 24582 6258 24610 6259
rect 24634 6285 24662 6286
rect 24634 6259 24636 6285
rect 24636 6259 24662 6285
rect 24634 6258 24662 6259
rect 24686 6285 24714 6286
rect 24738 6285 24766 6286
rect 24686 6259 24698 6285
rect 24698 6259 24714 6285
rect 24738 6259 24760 6285
rect 24760 6259 24766 6285
rect 24686 6258 24714 6259
rect 24738 6258 24766 6259
rect 24790 6258 24818 6286
rect 24842 6285 24870 6286
rect 24894 6285 24922 6286
rect 24842 6259 24848 6285
rect 24848 6259 24870 6285
rect 24894 6259 24910 6285
rect 24910 6259 24922 6285
rect 24842 6258 24870 6259
rect 24894 6258 24922 6259
rect 24946 6285 24974 6286
rect 24946 6259 24972 6285
rect 24972 6259 24974 6285
rect 24946 6258 24974 6259
rect 24998 6285 25026 6286
rect 24998 6259 25008 6285
rect 25008 6259 25026 6285
rect 24998 6258 25026 6259
rect 24486 5614 24514 5642
rect 25158 5782 25186 5810
rect 25046 5614 25074 5642
rect 24582 5501 24610 5502
rect 24582 5475 24600 5501
rect 24600 5475 24610 5501
rect 24582 5474 24610 5475
rect 24634 5501 24662 5502
rect 24634 5475 24636 5501
rect 24636 5475 24662 5501
rect 24634 5474 24662 5475
rect 24686 5501 24714 5502
rect 24738 5501 24766 5502
rect 24686 5475 24698 5501
rect 24698 5475 24714 5501
rect 24738 5475 24760 5501
rect 24760 5475 24766 5501
rect 24686 5474 24714 5475
rect 24738 5474 24766 5475
rect 24790 5474 24818 5502
rect 24842 5501 24870 5502
rect 24894 5501 24922 5502
rect 24842 5475 24848 5501
rect 24848 5475 24870 5501
rect 24894 5475 24910 5501
rect 24910 5475 24922 5501
rect 24842 5474 24870 5475
rect 24894 5474 24922 5475
rect 24946 5501 24974 5502
rect 24946 5475 24972 5501
rect 24972 5475 24974 5501
rect 24946 5474 24974 5475
rect 24998 5501 25026 5502
rect 24998 5475 25008 5501
rect 25008 5475 25026 5501
rect 24998 5474 25026 5475
rect 24430 5390 24458 5418
rect 25046 5390 25074 5418
rect 24654 4913 24682 4914
rect 24654 4887 24655 4913
rect 24655 4887 24681 4913
rect 24681 4887 24682 4913
rect 24654 4886 24682 4887
rect 24878 4913 24906 4914
rect 24878 4887 24879 4913
rect 24879 4887 24905 4913
rect 24905 4887 24906 4913
rect 24878 4886 24906 4887
rect 24582 4717 24610 4718
rect 24582 4691 24600 4717
rect 24600 4691 24610 4717
rect 24582 4690 24610 4691
rect 24634 4717 24662 4718
rect 24634 4691 24636 4717
rect 24636 4691 24662 4717
rect 24634 4690 24662 4691
rect 24686 4717 24714 4718
rect 24738 4717 24766 4718
rect 24686 4691 24698 4717
rect 24698 4691 24714 4717
rect 24738 4691 24760 4717
rect 24760 4691 24766 4717
rect 24686 4690 24714 4691
rect 24738 4690 24766 4691
rect 24790 4690 24818 4718
rect 24842 4717 24870 4718
rect 24894 4717 24922 4718
rect 24842 4691 24848 4717
rect 24848 4691 24870 4717
rect 24894 4691 24910 4717
rect 24910 4691 24922 4717
rect 24842 4690 24870 4691
rect 24894 4690 24922 4691
rect 24946 4717 24974 4718
rect 24946 4691 24972 4717
rect 24972 4691 24974 4717
rect 24946 4690 24974 4691
rect 24998 4717 25026 4718
rect 24998 4691 25008 4717
rect 25008 4691 25026 4717
rect 24998 4690 25026 4691
rect 24374 2422 24402 2450
rect 24374 2254 24402 2282
rect 24486 4129 24514 4130
rect 24486 4103 24487 4129
rect 24487 4103 24513 4129
rect 24513 4103 24514 4129
rect 24486 4102 24514 4103
rect 25158 4886 25186 4914
rect 25438 4521 25466 4522
rect 25438 4495 25439 4521
rect 25439 4495 25465 4521
rect 25465 4495 25466 4521
rect 25438 4494 25466 4495
rect 25102 4102 25130 4130
rect 24582 3933 24610 3934
rect 24582 3907 24600 3933
rect 24600 3907 24610 3933
rect 24582 3906 24610 3907
rect 24634 3933 24662 3934
rect 24634 3907 24636 3933
rect 24636 3907 24662 3933
rect 24634 3906 24662 3907
rect 24686 3933 24714 3934
rect 24738 3933 24766 3934
rect 24686 3907 24698 3933
rect 24698 3907 24714 3933
rect 24738 3907 24760 3933
rect 24760 3907 24766 3933
rect 24686 3906 24714 3907
rect 24738 3906 24766 3907
rect 24790 3906 24818 3934
rect 24842 3933 24870 3934
rect 24894 3933 24922 3934
rect 24842 3907 24848 3933
rect 24848 3907 24870 3933
rect 24894 3907 24910 3933
rect 24910 3907 24922 3933
rect 24842 3906 24870 3907
rect 24894 3906 24922 3907
rect 24946 3933 24974 3934
rect 24946 3907 24972 3933
rect 24972 3907 24974 3933
rect 24946 3906 24974 3907
rect 24998 3933 25026 3934
rect 24998 3907 25008 3933
rect 25008 3907 25026 3933
rect 24998 3906 25026 3907
rect 26502 5614 26530 5642
rect 26894 5558 26922 5586
rect 26894 4998 26922 5026
rect 26502 4718 26530 4746
rect 26894 4718 26922 4746
rect 26894 4521 26922 4522
rect 26894 4495 26895 4521
rect 26895 4495 26921 4521
rect 26921 4495 26922 4521
rect 26894 4494 26922 4495
rect 26894 4214 26922 4242
rect 26502 4102 26530 4130
rect 26838 4129 26866 4130
rect 26838 4103 26839 4129
rect 26839 4103 26865 4129
rect 26865 4103 26866 4129
rect 26838 4102 26866 4103
rect 26166 3822 26194 3850
rect 25382 3430 25410 3458
rect 24582 3149 24610 3150
rect 24582 3123 24600 3149
rect 24600 3123 24610 3149
rect 24582 3122 24610 3123
rect 24634 3149 24662 3150
rect 24634 3123 24636 3149
rect 24636 3123 24662 3149
rect 24634 3122 24662 3123
rect 24686 3149 24714 3150
rect 24738 3149 24766 3150
rect 24686 3123 24698 3149
rect 24698 3123 24714 3149
rect 24738 3123 24760 3149
rect 24760 3123 24766 3149
rect 24686 3122 24714 3123
rect 24738 3122 24766 3123
rect 24790 3122 24818 3150
rect 24842 3149 24870 3150
rect 24894 3149 24922 3150
rect 24842 3123 24848 3149
rect 24848 3123 24870 3149
rect 24894 3123 24910 3149
rect 24910 3123 24922 3149
rect 24842 3122 24870 3123
rect 24894 3122 24922 3123
rect 24946 3149 24974 3150
rect 24946 3123 24972 3149
rect 24972 3123 24974 3149
rect 24946 3122 24974 3123
rect 24998 3149 25026 3150
rect 24998 3123 25008 3149
rect 25008 3123 25026 3149
rect 24998 3122 25026 3123
rect 24430 2478 24458 2506
rect 24766 2478 24794 2506
rect 24582 2365 24610 2366
rect 24582 2339 24600 2365
rect 24600 2339 24610 2365
rect 24582 2338 24610 2339
rect 24634 2365 24662 2366
rect 24634 2339 24636 2365
rect 24636 2339 24662 2365
rect 24634 2338 24662 2339
rect 24686 2365 24714 2366
rect 24738 2365 24766 2366
rect 24686 2339 24698 2365
rect 24698 2339 24714 2365
rect 24738 2339 24760 2365
rect 24760 2339 24766 2365
rect 24686 2338 24714 2339
rect 24738 2338 24766 2339
rect 24790 2338 24818 2366
rect 24842 2365 24870 2366
rect 24894 2365 24922 2366
rect 24842 2339 24848 2365
rect 24848 2339 24870 2365
rect 24894 2339 24910 2365
rect 24910 2339 24922 2365
rect 24842 2338 24870 2339
rect 24894 2338 24922 2339
rect 24946 2365 24974 2366
rect 24946 2339 24972 2365
rect 24972 2339 24974 2365
rect 24946 2338 24974 2339
rect 24998 2365 25026 2366
rect 24998 2339 25008 2365
rect 25008 2339 25026 2365
rect 24998 2338 25026 2339
rect 24430 1806 24458 1834
rect 24766 2169 24794 2170
rect 24766 2143 24767 2169
rect 24767 2143 24793 2169
rect 24793 2143 24794 2169
rect 24766 2142 24794 2143
rect 26166 3374 26194 3402
rect 25942 2646 25970 2674
rect 24766 1806 24794 1834
rect 25998 3318 26026 3346
rect 26894 3878 26922 3906
rect 26222 2534 26250 2562
rect 26726 2561 26754 2562
rect 26726 2535 26727 2561
rect 26727 2535 26753 2561
rect 26753 2535 26754 2561
rect 26726 2534 26754 2535
rect 26222 2169 26250 2170
rect 26222 2143 26223 2169
rect 26223 2143 26249 2169
rect 26249 2143 26250 2169
rect 26222 2142 26250 2143
rect 26390 2478 26418 2506
rect 26390 1694 26418 1722
rect 26726 2254 26754 2282
rect 24582 1581 24610 1582
rect 24582 1555 24600 1581
rect 24600 1555 24610 1581
rect 24582 1554 24610 1555
rect 24634 1581 24662 1582
rect 24634 1555 24636 1581
rect 24636 1555 24662 1581
rect 24634 1554 24662 1555
rect 24686 1581 24714 1582
rect 24738 1581 24766 1582
rect 24686 1555 24698 1581
rect 24698 1555 24714 1581
rect 24738 1555 24760 1581
rect 24760 1555 24766 1581
rect 24686 1554 24714 1555
rect 24738 1554 24766 1555
rect 24790 1554 24818 1582
rect 24842 1581 24870 1582
rect 24894 1581 24922 1582
rect 24842 1555 24848 1581
rect 24848 1555 24870 1581
rect 24894 1555 24910 1581
rect 24910 1555 24922 1581
rect 24842 1554 24870 1555
rect 24894 1554 24922 1555
rect 24946 1581 24974 1582
rect 24946 1555 24972 1581
rect 24972 1555 24974 1581
rect 24946 1554 24974 1555
rect 24998 1581 25026 1582
rect 24998 1555 25008 1581
rect 25008 1555 25026 1581
rect 24998 1554 25026 1555
rect 27082 9029 27110 9030
rect 27082 9003 27100 9029
rect 27100 9003 27110 9029
rect 27082 9002 27110 9003
rect 27134 9029 27162 9030
rect 27134 9003 27136 9029
rect 27136 9003 27162 9029
rect 27134 9002 27162 9003
rect 27186 9029 27214 9030
rect 27238 9029 27266 9030
rect 27186 9003 27198 9029
rect 27198 9003 27214 9029
rect 27238 9003 27260 9029
rect 27260 9003 27266 9029
rect 27186 9002 27214 9003
rect 27238 9002 27266 9003
rect 27290 9002 27318 9030
rect 27342 9029 27370 9030
rect 27394 9029 27422 9030
rect 27342 9003 27348 9029
rect 27348 9003 27370 9029
rect 27394 9003 27410 9029
rect 27410 9003 27422 9029
rect 27342 9002 27370 9003
rect 27394 9002 27422 9003
rect 27446 9029 27474 9030
rect 27446 9003 27472 9029
rect 27472 9003 27474 9029
rect 27446 9002 27474 9003
rect 27498 9029 27526 9030
rect 27498 9003 27508 9029
rect 27508 9003 27526 9029
rect 27498 9002 27526 9003
rect 27566 8862 27594 8890
rect 27398 8358 27426 8386
rect 27082 8245 27110 8246
rect 27082 8219 27100 8245
rect 27100 8219 27110 8245
rect 27082 8218 27110 8219
rect 27134 8245 27162 8246
rect 27134 8219 27136 8245
rect 27136 8219 27162 8245
rect 27134 8218 27162 8219
rect 27186 8245 27214 8246
rect 27238 8245 27266 8246
rect 27186 8219 27198 8245
rect 27198 8219 27214 8245
rect 27238 8219 27260 8245
rect 27260 8219 27266 8245
rect 27186 8218 27214 8219
rect 27238 8218 27266 8219
rect 27290 8218 27318 8246
rect 27342 8245 27370 8246
rect 27394 8245 27422 8246
rect 27342 8219 27348 8245
rect 27348 8219 27370 8245
rect 27394 8219 27410 8245
rect 27410 8219 27422 8245
rect 27342 8218 27370 8219
rect 27394 8218 27422 8219
rect 27446 8245 27474 8246
rect 27446 8219 27472 8245
rect 27472 8219 27474 8245
rect 27446 8218 27474 8219
rect 27498 8245 27526 8246
rect 27498 8219 27508 8245
rect 27508 8219 27526 8245
rect 27498 8218 27526 8219
rect 27082 7461 27110 7462
rect 27082 7435 27100 7461
rect 27100 7435 27110 7461
rect 27082 7434 27110 7435
rect 27134 7461 27162 7462
rect 27134 7435 27136 7461
rect 27136 7435 27162 7461
rect 27134 7434 27162 7435
rect 27186 7461 27214 7462
rect 27238 7461 27266 7462
rect 27186 7435 27198 7461
rect 27198 7435 27214 7461
rect 27238 7435 27260 7461
rect 27260 7435 27266 7461
rect 27186 7434 27214 7435
rect 27238 7434 27266 7435
rect 27290 7434 27318 7462
rect 27342 7461 27370 7462
rect 27394 7461 27422 7462
rect 27342 7435 27348 7461
rect 27348 7435 27370 7461
rect 27394 7435 27410 7461
rect 27410 7435 27422 7461
rect 27342 7434 27370 7435
rect 27394 7434 27422 7435
rect 27446 7461 27474 7462
rect 27446 7435 27472 7461
rect 27472 7435 27474 7461
rect 27446 7434 27474 7435
rect 27498 7461 27526 7462
rect 27498 7435 27508 7461
rect 27508 7435 27526 7461
rect 27498 7434 27526 7435
rect 27678 8358 27706 8386
rect 27958 9982 27986 10010
rect 28350 10009 28378 10010
rect 28350 9983 28351 10009
rect 28351 9983 28377 10009
rect 28377 9983 28378 10009
rect 28350 9982 28378 9983
rect 29582 10989 29610 10990
rect 29582 10963 29600 10989
rect 29600 10963 29610 10989
rect 29582 10962 29610 10963
rect 29634 10989 29662 10990
rect 29634 10963 29636 10989
rect 29636 10963 29662 10989
rect 29634 10962 29662 10963
rect 29686 10989 29714 10990
rect 29738 10989 29766 10990
rect 29686 10963 29698 10989
rect 29698 10963 29714 10989
rect 29738 10963 29760 10989
rect 29760 10963 29766 10989
rect 29686 10962 29714 10963
rect 29738 10962 29766 10963
rect 29790 10962 29818 10990
rect 29842 10989 29870 10990
rect 29894 10989 29922 10990
rect 29842 10963 29848 10989
rect 29848 10963 29870 10989
rect 29894 10963 29910 10989
rect 29910 10963 29922 10989
rect 29842 10962 29870 10963
rect 29894 10962 29922 10963
rect 29946 10989 29974 10990
rect 29946 10963 29972 10989
rect 29972 10963 29974 10989
rect 29946 10962 29974 10963
rect 29998 10989 30026 10990
rect 29998 10963 30008 10989
rect 30008 10963 30026 10989
rect 29998 10962 30026 10963
rect 29582 10205 29610 10206
rect 29582 10179 29600 10205
rect 29600 10179 29610 10205
rect 29582 10178 29610 10179
rect 29634 10205 29662 10206
rect 29634 10179 29636 10205
rect 29636 10179 29662 10205
rect 29634 10178 29662 10179
rect 29686 10205 29714 10206
rect 29738 10205 29766 10206
rect 29686 10179 29698 10205
rect 29698 10179 29714 10205
rect 29738 10179 29760 10205
rect 29760 10179 29766 10205
rect 29686 10178 29714 10179
rect 29738 10178 29766 10179
rect 29790 10178 29818 10206
rect 29842 10205 29870 10206
rect 29894 10205 29922 10206
rect 29842 10179 29848 10205
rect 29848 10179 29870 10205
rect 29894 10179 29910 10205
rect 29910 10179 29922 10205
rect 29842 10178 29870 10179
rect 29894 10178 29922 10179
rect 29946 10205 29974 10206
rect 29946 10179 29972 10205
rect 29972 10179 29974 10205
rect 29946 10178 29974 10179
rect 29998 10205 30026 10206
rect 29998 10179 30008 10205
rect 30008 10179 30026 10205
rect 29998 10178 30026 10179
rect 29470 10038 29498 10066
rect 29806 10038 29834 10066
rect 28798 9982 28826 10010
rect 27958 9142 27986 9170
rect 27566 6873 27594 6874
rect 27566 6847 27567 6873
rect 27567 6847 27593 6873
rect 27593 6847 27594 6873
rect 27566 6846 27594 6847
rect 27082 6677 27110 6678
rect 27082 6651 27100 6677
rect 27100 6651 27110 6677
rect 27082 6650 27110 6651
rect 27134 6677 27162 6678
rect 27134 6651 27136 6677
rect 27136 6651 27162 6677
rect 27134 6650 27162 6651
rect 27186 6677 27214 6678
rect 27238 6677 27266 6678
rect 27186 6651 27198 6677
rect 27198 6651 27214 6677
rect 27238 6651 27260 6677
rect 27260 6651 27266 6677
rect 27186 6650 27214 6651
rect 27238 6650 27266 6651
rect 27290 6650 27318 6678
rect 27342 6677 27370 6678
rect 27394 6677 27422 6678
rect 27342 6651 27348 6677
rect 27348 6651 27370 6677
rect 27394 6651 27410 6677
rect 27410 6651 27422 6677
rect 27342 6650 27370 6651
rect 27394 6650 27422 6651
rect 27446 6677 27474 6678
rect 27446 6651 27472 6677
rect 27472 6651 27474 6677
rect 27446 6650 27474 6651
rect 27498 6677 27526 6678
rect 27498 6651 27508 6677
rect 27508 6651 27526 6677
rect 27498 6650 27526 6651
rect 27678 6846 27706 6874
rect 27790 6873 27818 6874
rect 27790 6847 27791 6873
rect 27791 6847 27817 6873
rect 27817 6847 27818 6873
rect 27790 6846 27818 6847
rect 27082 5893 27110 5894
rect 27082 5867 27100 5893
rect 27100 5867 27110 5893
rect 27082 5866 27110 5867
rect 27134 5893 27162 5894
rect 27134 5867 27136 5893
rect 27136 5867 27162 5893
rect 27134 5866 27162 5867
rect 27186 5893 27214 5894
rect 27238 5893 27266 5894
rect 27186 5867 27198 5893
rect 27198 5867 27214 5893
rect 27238 5867 27260 5893
rect 27260 5867 27266 5893
rect 27186 5866 27214 5867
rect 27238 5866 27266 5867
rect 27290 5866 27318 5894
rect 27342 5893 27370 5894
rect 27394 5893 27422 5894
rect 27342 5867 27348 5893
rect 27348 5867 27370 5893
rect 27394 5867 27410 5893
rect 27410 5867 27422 5893
rect 27342 5866 27370 5867
rect 27394 5866 27422 5867
rect 27446 5893 27474 5894
rect 27446 5867 27472 5893
rect 27472 5867 27474 5893
rect 27446 5866 27474 5867
rect 27498 5893 27526 5894
rect 27498 5867 27508 5893
rect 27508 5867 27526 5893
rect 27498 5866 27526 5867
rect 27006 5558 27034 5586
rect 27082 5109 27110 5110
rect 27082 5083 27100 5109
rect 27100 5083 27110 5109
rect 27082 5082 27110 5083
rect 27134 5109 27162 5110
rect 27134 5083 27136 5109
rect 27136 5083 27162 5109
rect 27134 5082 27162 5083
rect 27186 5109 27214 5110
rect 27238 5109 27266 5110
rect 27186 5083 27198 5109
rect 27198 5083 27214 5109
rect 27238 5083 27260 5109
rect 27260 5083 27266 5109
rect 27186 5082 27214 5083
rect 27238 5082 27266 5083
rect 27290 5082 27318 5110
rect 27342 5109 27370 5110
rect 27394 5109 27422 5110
rect 27342 5083 27348 5109
rect 27348 5083 27370 5109
rect 27394 5083 27410 5109
rect 27410 5083 27422 5109
rect 27342 5082 27370 5083
rect 27394 5082 27422 5083
rect 27446 5109 27474 5110
rect 27446 5083 27472 5109
rect 27472 5083 27474 5109
rect 27446 5082 27474 5083
rect 27498 5109 27526 5110
rect 27498 5083 27508 5109
rect 27508 5083 27526 5109
rect 27498 5082 27526 5083
rect 27006 4886 27034 4914
rect 27174 4998 27202 5026
rect 27174 4494 27202 4522
rect 27082 4325 27110 4326
rect 27082 4299 27100 4325
rect 27100 4299 27110 4325
rect 27082 4298 27110 4299
rect 27134 4325 27162 4326
rect 27134 4299 27136 4325
rect 27136 4299 27162 4325
rect 27134 4298 27162 4299
rect 27186 4325 27214 4326
rect 27238 4325 27266 4326
rect 27186 4299 27198 4325
rect 27198 4299 27214 4325
rect 27238 4299 27260 4325
rect 27260 4299 27266 4325
rect 27186 4298 27214 4299
rect 27238 4298 27266 4299
rect 27290 4298 27318 4326
rect 27342 4325 27370 4326
rect 27394 4325 27422 4326
rect 27342 4299 27348 4325
rect 27348 4299 27370 4325
rect 27394 4299 27410 4325
rect 27410 4299 27422 4325
rect 27342 4298 27370 4299
rect 27394 4298 27422 4299
rect 27446 4325 27474 4326
rect 27446 4299 27472 4325
rect 27472 4299 27474 4325
rect 27446 4298 27474 4299
rect 27498 4325 27526 4326
rect 27498 4299 27508 4325
rect 27508 4299 27526 4325
rect 27498 4298 27526 4299
rect 27510 4214 27538 4242
rect 27174 3878 27202 3906
rect 27082 3541 27110 3542
rect 27082 3515 27100 3541
rect 27100 3515 27110 3541
rect 27082 3514 27110 3515
rect 27134 3541 27162 3542
rect 27134 3515 27136 3541
rect 27136 3515 27162 3541
rect 27134 3514 27162 3515
rect 27186 3541 27214 3542
rect 27238 3541 27266 3542
rect 27186 3515 27198 3541
rect 27198 3515 27214 3541
rect 27238 3515 27260 3541
rect 27260 3515 27266 3541
rect 27186 3514 27214 3515
rect 27238 3514 27266 3515
rect 27290 3514 27318 3542
rect 27342 3541 27370 3542
rect 27394 3541 27422 3542
rect 27342 3515 27348 3541
rect 27348 3515 27370 3541
rect 27394 3515 27410 3541
rect 27410 3515 27422 3541
rect 27342 3514 27370 3515
rect 27394 3514 27422 3515
rect 27446 3541 27474 3542
rect 27446 3515 27472 3541
rect 27472 3515 27474 3541
rect 27446 3514 27474 3515
rect 27498 3541 27526 3542
rect 27498 3515 27508 3541
rect 27508 3515 27526 3541
rect 27498 3514 27526 3515
rect 27082 2757 27110 2758
rect 27082 2731 27100 2757
rect 27100 2731 27110 2757
rect 27082 2730 27110 2731
rect 27134 2757 27162 2758
rect 27134 2731 27136 2757
rect 27136 2731 27162 2757
rect 27134 2730 27162 2731
rect 27186 2757 27214 2758
rect 27238 2757 27266 2758
rect 27186 2731 27198 2757
rect 27198 2731 27214 2757
rect 27238 2731 27260 2757
rect 27260 2731 27266 2757
rect 27186 2730 27214 2731
rect 27238 2730 27266 2731
rect 27290 2730 27318 2758
rect 27342 2757 27370 2758
rect 27394 2757 27422 2758
rect 27342 2731 27348 2757
rect 27348 2731 27370 2757
rect 27394 2731 27410 2757
rect 27410 2731 27422 2757
rect 27342 2730 27370 2731
rect 27394 2730 27422 2731
rect 27446 2757 27474 2758
rect 27446 2731 27472 2757
rect 27472 2731 27474 2757
rect 27446 2730 27474 2731
rect 27498 2757 27526 2758
rect 27498 2731 27508 2757
rect 27508 2731 27526 2757
rect 27498 2730 27526 2731
rect 26950 2254 26978 2282
rect 27622 2646 27650 2674
rect 27398 2225 27426 2226
rect 27398 2199 27399 2225
rect 27399 2199 27425 2225
rect 27425 2199 27426 2225
rect 27398 2198 27426 2199
rect 27082 1973 27110 1974
rect 27082 1947 27100 1973
rect 27100 1947 27110 1973
rect 27082 1946 27110 1947
rect 27134 1973 27162 1974
rect 27134 1947 27136 1973
rect 27136 1947 27162 1973
rect 27134 1946 27162 1947
rect 27186 1973 27214 1974
rect 27238 1973 27266 1974
rect 27186 1947 27198 1973
rect 27198 1947 27214 1973
rect 27238 1947 27260 1973
rect 27260 1947 27266 1973
rect 27186 1946 27214 1947
rect 27238 1946 27266 1947
rect 27290 1946 27318 1974
rect 27342 1973 27370 1974
rect 27394 1973 27422 1974
rect 27342 1947 27348 1973
rect 27348 1947 27370 1973
rect 27394 1947 27410 1973
rect 27410 1947 27422 1973
rect 27342 1946 27370 1947
rect 27394 1946 27422 1947
rect 27446 1973 27474 1974
rect 27446 1947 27472 1973
rect 27472 1947 27474 1973
rect 27446 1946 27474 1947
rect 27498 1973 27526 1974
rect 27498 1947 27508 1973
rect 27508 1947 27526 1973
rect 27498 1946 27526 1947
rect 27678 4214 27706 4242
rect 27678 2198 27706 2226
rect 28350 6734 28378 6762
rect 28238 4998 28266 5026
rect 28182 4718 28210 4746
rect 28070 4577 28098 4578
rect 28070 4551 28071 4577
rect 28071 4551 28097 4577
rect 28097 4551 28098 4577
rect 28070 4550 28098 4551
rect 28070 4438 28098 4466
rect 28462 4913 28490 4914
rect 28462 4887 28463 4913
rect 28463 4887 28489 4913
rect 28489 4887 28490 4913
rect 28462 4886 28490 4887
rect 28238 4577 28266 4578
rect 28238 4551 28239 4577
rect 28239 4551 28265 4577
rect 28265 4551 28266 4577
rect 28238 4550 28266 4551
rect 28294 4830 28322 4858
rect 28238 4158 28266 4186
rect 28462 4494 28490 4522
rect 28742 4521 28770 4522
rect 28742 4495 28743 4521
rect 28743 4495 28769 4521
rect 28769 4495 28770 4521
rect 28742 4494 28770 4495
rect 28686 4214 28714 4242
rect 28462 4129 28490 4130
rect 28462 4103 28463 4129
rect 28463 4103 28489 4129
rect 28489 4103 28490 4129
rect 28462 4102 28490 4103
rect 28350 3009 28378 3010
rect 28350 2983 28351 3009
rect 28351 2983 28377 3009
rect 28377 2983 28378 3009
rect 28350 2982 28378 2983
rect 28070 2590 28098 2618
rect 28518 2982 28546 3010
rect 28462 2561 28490 2562
rect 28462 2535 28463 2561
rect 28463 2535 28489 2561
rect 28489 2535 28490 2561
rect 28462 2534 28490 2535
rect 28742 2534 28770 2562
rect 28350 2086 28378 2114
rect 28518 1777 28546 1778
rect 28518 1751 28519 1777
rect 28519 1751 28545 1777
rect 28545 1751 28546 1777
rect 28518 1750 28546 1751
rect 30030 10038 30058 10066
rect 30086 9870 30114 9898
rect 29582 9421 29610 9422
rect 29582 9395 29600 9421
rect 29600 9395 29610 9421
rect 29582 9394 29610 9395
rect 29634 9421 29662 9422
rect 29634 9395 29636 9421
rect 29636 9395 29662 9421
rect 29634 9394 29662 9395
rect 29686 9421 29714 9422
rect 29738 9421 29766 9422
rect 29686 9395 29698 9421
rect 29698 9395 29714 9421
rect 29738 9395 29760 9421
rect 29760 9395 29766 9421
rect 29686 9394 29714 9395
rect 29738 9394 29766 9395
rect 29790 9394 29818 9422
rect 29842 9421 29870 9422
rect 29894 9421 29922 9422
rect 29842 9395 29848 9421
rect 29848 9395 29870 9421
rect 29894 9395 29910 9421
rect 29910 9395 29922 9421
rect 29842 9394 29870 9395
rect 29894 9394 29922 9395
rect 29946 9421 29974 9422
rect 29946 9395 29972 9421
rect 29972 9395 29974 9421
rect 29946 9394 29974 9395
rect 29998 9421 30026 9422
rect 29998 9395 30008 9421
rect 30008 9395 30026 9421
rect 29998 9394 30026 9395
rect 29414 9198 29442 9226
rect 29526 9225 29554 9226
rect 29526 9199 29527 9225
rect 29527 9199 29553 9225
rect 29553 9199 29554 9225
rect 29526 9198 29554 9199
rect 28854 8833 28882 8834
rect 28854 8807 28855 8833
rect 28855 8807 28881 8833
rect 28881 8807 28882 8833
rect 28854 8806 28882 8807
rect 29414 8833 29442 8834
rect 29414 8807 29415 8833
rect 29415 8807 29441 8833
rect 29441 8807 29442 8833
rect 29414 8806 29442 8807
rect 29582 8637 29610 8638
rect 29582 8611 29600 8637
rect 29600 8611 29610 8637
rect 29582 8610 29610 8611
rect 29634 8637 29662 8638
rect 29634 8611 29636 8637
rect 29636 8611 29662 8637
rect 29634 8610 29662 8611
rect 29686 8637 29714 8638
rect 29738 8637 29766 8638
rect 29686 8611 29698 8637
rect 29698 8611 29714 8637
rect 29738 8611 29760 8637
rect 29760 8611 29766 8637
rect 29686 8610 29714 8611
rect 29738 8610 29766 8611
rect 29790 8610 29818 8638
rect 29842 8637 29870 8638
rect 29894 8637 29922 8638
rect 29842 8611 29848 8637
rect 29848 8611 29870 8637
rect 29894 8611 29910 8637
rect 29910 8611 29922 8637
rect 29842 8610 29870 8611
rect 29894 8610 29922 8611
rect 29946 8637 29974 8638
rect 29946 8611 29972 8637
rect 29972 8611 29974 8637
rect 29946 8610 29974 8611
rect 29998 8637 30026 8638
rect 29998 8611 30008 8637
rect 30008 8611 30026 8637
rect 29998 8610 30026 8611
rect 30198 8833 30226 8834
rect 30198 8807 30199 8833
rect 30199 8807 30225 8833
rect 30225 8807 30226 8833
rect 30198 8806 30226 8807
rect 29582 7853 29610 7854
rect 29582 7827 29600 7853
rect 29600 7827 29610 7853
rect 29582 7826 29610 7827
rect 29634 7853 29662 7854
rect 29634 7827 29636 7853
rect 29636 7827 29662 7853
rect 29634 7826 29662 7827
rect 29686 7853 29714 7854
rect 29738 7853 29766 7854
rect 29686 7827 29698 7853
rect 29698 7827 29714 7853
rect 29738 7827 29760 7853
rect 29760 7827 29766 7853
rect 29686 7826 29714 7827
rect 29738 7826 29766 7827
rect 29790 7826 29818 7854
rect 29842 7853 29870 7854
rect 29894 7853 29922 7854
rect 29842 7827 29848 7853
rect 29848 7827 29870 7853
rect 29894 7827 29910 7853
rect 29910 7827 29922 7853
rect 29842 7826 29870 7827
rect 29894 7826 29922 7827
rect 29946 7853 29974 7854
rect 29946 7827 29972 7853
rect 29972 7827 29974 7853
rect 29946 7826 29974 7827
rect 29998 7853 30026 7854
rect 29998 7827 30008 7853
rect 30008 7827 30026 7853
rect 29998 7826 30026 7827
rect 28854 6734 28882 6762
rect 29582 7069 29610 7070
rect 29582 7043 29600 7069
rect 29600 7043 29610 7069
rect 29582 7042 29610 7043
rect 29634 7069 29662 7070
rect 29634 7043 29636 7069
rect 29636 7043 29662 7069
rect 29634 7042 29662 7043
rect 29686 7069 29714 7070
rect 29738 7069 29766 7070
rect 29686 7043 29698 7069
rect 29698 7043 29714 7069
rect 29738 7043 29760 7069
rect 29760 7043 29766 7069
rect 29686 7042 29714 7043
rect 29738 7042 29766 7043
rect 29790 7042 29818 7070
rect 29842 7069 29870 7070
rect 29894 7069 29922 7070
rect 29842 7043 29848 7069
rect 29848 7043 29870 7069
rect 29894 7043 29910 7069
rect 29910 7043 29922 7069
rect 29842 7042 29870 7043
rect 29894 7042 29922 7043
rect 29946 7069 29974 7070
rect 29946 7043 29972 7069
rect 29972 7043 29974 7069
rect 29946 7042 29974 7043
rect 29998 7069 30026 7070
rect 29998 7043 30008 7069
rect 30008 7043 30026 7069
rect 29998 7042 30026 7043
rect 29358 6734 29386 6762
rect 29582 6285 29610 6286
rect 29582 6259 29600 6285
rect 29600 6259 29610 6285
rect 29582 6258 29610 6259
rect 29634 6285 29662 6286
rect 29634 6259 29636 6285
rect 29636 6259 29662 6285
rect 29634 6258 29662 6259
rect 29686 6285 29714 6286
rect 29738 6285 29766 6286
rect 29686 6259 29698 6285
rect 29698 6259 29714 6285
rect 29738 6259 29760 6285
rect 29760 6259 29766 6285
rect 29686 6258 29714 6259
rect 29738 6258 29766 6259
rect 29790 6258 29818 6286
rect 29842 6285 29870 6286
rect 29894 6285 29922 6286
rect 29842 6259 29848 6285
rect 29848 6259 29870 6285
rect 29894 6259 29910 6285
rect 29910 6259 29922 6285
rect 29842 6258 29870 6259
rect 29894 6258 29922 6259
rect 29946 6285 29974 6286
rect 29946 6259 29972 6285
rect 29972 6259 29974 6285
rect 29946 6258 29974 6259
rect 29998 6285 30026 6286
rect 29998 6259 30008 6285
rect 30008 6259 30026 6285
rect 29998 6258 30026 6259
rect 30198 5838 30226 5866
rect 29582 5501 29610 5502
rect 29582 5475 29600 5501
rect 29600 5475 29610 5501
rect 29582 5474 29610 5475
rect 29634 5501 29662 5502
rect 29634 5475 29636 5501
rect 29636 5475 29662 5501
rect 29634 5474 29662 5475
rect 29686 5501 29714 5502
rect 29738 5501 29766 5502
rect 29686 5475 29698 5501
rect 29698 5475 29714 5501
rect 29738 5475 29760 5501
rect 29760 5475 29766 5501
rect 29686 5474 29714 5475
rect 29738 5474 29766 5475
rect 29790 5474 29818 5502
rect 29842 5501 29870 5502
rect 29894 5501 29922 5502
rect 29842 5475 29848 5501
rect 29848 5475 29870 5501
rect 29894 5475 29910 5501
rect 29910 5475 29922 5501
rect 29842 5474 29870 5475
rect 29894 5474 29922 5475
rect 29946 5501 29974 5502
rect 29946 5475 29972 5501
rect 29972 5475 29974 5501
rect 29946 5474 29974 5475
rect 29998 5501 30026 5502
rect 29998 5475 30008 5501
rect 30008 5475 30026 5501
rect 29998 5474 30026 5475
rect 29358 5305 29386 5306
rect 29358 5279 29359 5305
rect 29359 5279 29385 5305
rect 29385 5279 29386 5305
rect 29358 5278 29386 5279
rect 30254 10038 30282 10066
rect 30142 4998 30170 5026
rect 30030 4857 30058 4858
rect 30030 4831 30031 4857
rect 30031 4831 30057 4857
rect 30057 4831 30058 4857
rect 30030 4830 30058 4831
rect 29582 4717 29610 4718
rect 29582 4691 29600 4717
rect 29600 4691 29610 4717
rect 29582 4690 29610 4691
rect 29634 4717 29662 4718
rect 29634 4691 29636 4717
rect 29636 4691 29662 4717
rect 29634 4690 29662 4691
rect 29686 4717 29714 4718
rect 29738 4717 29766 4718
rect 29686 4691 29698 4717
rect 29698 4691 29714 4717
rect 29738 4691 29760 4717
rect 29760 4691 29766 4717
rect 29686 4690 29714 4691
rect 29738 4690 29766 4691
rect 29790 4690 29818 4718
rect 29842 4717 29870 4718
rect 29894 4717 29922 4718
rect 29842 4691 29848 4717
rect 29848 4691 29870 4717
rect 29894 4691 29910 4717
rect 29910 4691 29922 4717
rect 29842 4690 29870 4691
rect 29894 4690 29922 4691
rect 29946 4717 29974 4718
rect 29946 4691 29972 4717
rect 29972 4691 29974 4717
rect 29946 4690 29974 4691
rect 29998 4717 30026 4718
rect 29998 4691 30008 4717
rect 30008 4691 30026 4717
rect 29998 4690 30026 4691
rect 28910 4214 28938 4242
rect 29414 4214 29442 4242
rect 28966 2422 28994 2450
rect 28966 1750 28994 1778
rect 29358 2926 29386 2954
rect 29358 2646 29386 2674
rect 29582 3933 29610 3934
rect 29582 3907 29600 3933
rect 29600 3907 29610 3933
rect 29582 3906 29610 3907
rect 29634 3933 29662 3934
rect 29634 3907 29636 3933
rect 29636 3907 29662 3933
rect 29634 3906 29662 3907
rect 29686 3933 29714 3934
rect 29738 3933 29766 3934
rect 29686 3907 29698 3933
rect 29698 3907 29714 3933
rect 29738 3907 29760 3933
rect 29760 3907 29766 3933
rect 29686 3906 29714 3907
rect 29738 3906 29766 3907
rect 29790 3906 29818 3934
rect 29842 3933 29870 3934
rect 29894 3933 29922 3934
rect 29842 3907 29848 3933
rect 29848 3907 29870 3933
rect 29894 3907 29910 3933
rect 29910 3907 29922 3933
rect 29842 3906 29870 3907
rect 29894 3906 29922 3907
rect 29946 3933 29974 3934
rect 29946 3907 29972 3933
rect 29972 3907 29974 3933
rect 29946 3906 29974 3907
rect 29998 3933 30026 3934
rect 29998 3907 30008 3933
rect 30008 3907 30026 3933
rect 29998 3906 30026 3907
rect 30030 3289 30058 3290
rect 30030 3263 30031 3289
rect 30031 3263 30057 3289
rect 30057 3263 30058 3289
rect 30030 3262 30058 3263
rect 29582 3149 29610 3150
rect 29582 3123 29600 3149
rect 29600 3123 29610 3149
rect 29582 3122 29610 3123
rect 29634 3149 29662 3150
rect 29634 3123 29636 3149
rect 29636 3123 29662 3149
rect 29634 3122 29662 3123
rect 29686 3149 29714 3150
rect 29738 3149 29766 3150
rect 29686 3123 29698 3149
rect 29698 3123 29714 3149
rect 29738 3123 29760 3149
rect 29760 3123 29766 3149
rect 29686 3122 29714 3123
rect 29738 3122 29766 3123
rect 29790 3122 29818 3150
rect 29842 3149 29870 3150
rect 29894 3149 29922 3150
rect 29842 3123 29848 3149
rect 29848 3123 29870 3149
rect 29894 3123 29910 3149
rect 29910 3123 29922 3149
rect 29842 3122 29870 3123
rect 29894 3122 29922 3123
rect 29946 3149 29974 3150
rect 29946 3123 29972 3149
rect 29972 3123 29974 3149
rect 29946 3122 29974 3123
rect 29998 3149 30026 3150
rect 29998 3123 30008 3149
rect 30008 3123 30026 3149
rect 29998 3122 30026 3123
rect 29470 2926 29498 2954
rect 29918 2953 29946 2954
rect 29918 2927 29919 2953
rect 29919 2927 29945 2953
rect 29945 2927 29946 2953
rect 29918 2926 29946 2927
rect 30086 2982 30114 3010
rect 30142 4073 30170 4074
rect 30142 4047 30143 4073
rect 30143 4047 30169 4073
rect 30169 4047 30170 4073
rect 30142 4046 30170 4047
rect 30142 2590 30170 2618
rect 29582 2365 29610 2366
rect 29582 2339 29600 2365
rect 29600 2339 29610 2365
rect 29582 2338 29610 2339
rect 29634 2365 29662 2366
rect 29634 2339 29636 2365
rect 29636 2339 29662 2365
rect 29634 2338 29662 2339
rect 29686 2365 29714 2366
rect 29738 2365 29766 2366
rect 29686 2339 29698 2365
rect 29698 2339 29714 2365
rect 29738 2339 29760 2365
rect 29760 2339 29766 2365
rect 29686 2338 29714 2339
rect 29738 2338 29766 2339
rect 29790 2338 29818 2366
rect 29842 2365 29870 2366
rect 29894 2365 29922 2366
rect 29842 2339 29848 2365
rect 29848 2339 29870 2365
rect 29894 2339 29910 2365
rect 29910 2339 29922 2365
rect 29842 2338 29870 2339
rect 29894 2338 29922 2339
rect 29946 2365 29974 2366
rect 29946 2339 29972 2365
rect 29972 2339 29974 2365
rect 29946 2338 29974 2339
rect 29998 2365 30026 2366
rect 29998 2339 30008 2365
rect 30008 2339 30026 2365
rect 29998 2338 30026 2339
rect 29414 2142 29442 2170
rect 29918 2169 29946 2170
rect 29918 2143 29919 2169
rect 29919 2143 29945 2169
rect 29945 2143 29946 2169
rect 29918 2142 29946 2143
rect 29582 1581 29610 1582
rect 29582 1555 29600 1581
rect 29600 1555 29610 1581
rect 29582 1554 29610 1555
rect 29634 1581 29662 1582
rect 29634 1555 29636 1581
rect 29636 1555 29662 1581
rect 29634 1554 29662 1555
rect 29686 1581 29714 1582
rect 29738 1581 29766 1582
rect 29686 1555 29698 1581
rect 29698 1555 29714 1581
rect 29738 1555 29760 1581
rect 29760 1555 29766 1581
rect 29686 1554 29714 1555
rect 29738 1554 29766 1555
rect 29790 1554 29818 1582
rect 29842 1581 29870 1582
rect 29894 1581 29922 1582
rect 29842 1555 29848 1581
rect 29848 1555 29870 1581
rect 29894 1555 29910 1581
rect 29910 1555 29922 1581
rect 29842 1554 29870 1555
rect 29894 1554 29922 1555
rect 29946 1581 29974 1582
rect 29946 1555 29972 1581
rect 29972 1555 29974 1581
rect 29946 1554 29974 1555
rect 29998 1581 30026 1582
rect 29998 1555 30008 1581
rect 30008 1555 30026 1581
rect 29998 1554 30026 1555
rect 30310 9982 30338 10010
rect 31486 11633 31514 11634
rect 31486 11607 31487 11633
rect 31487 11607 31513 11633
rect 31513 11607 31514 11633
rect 31486 11606 31514 11607
rect 32082 18437 32110 18438
rect 32082 18411 32100 18437
rect 32100 18411 32110 18437
rect 32082 18410 32110 18411
rect 32134 18437 32162 18438
rect 32134 18411 32136 18437
rect 32136 18411 32162 18437
rect 32134 18410 32162 18411
rect 32186 18437 32214 18438
rect 32238 18437 32266 18438
rect 32186 18411 32198 18437
rect 32198 18411 32214 18437
rect 32238 18411 32260 18437
rect 32260 18411 32266 18437
rect 32186 18410 32214 18411
rect 32238 18410 32266 18411
rect 32290 18410 32318 18438
rect 32342 18437 32370 18438
rect 32394 18437 32422 18438
rect 32342 18411 32348 18437
rect 32348 18411 32370 18437
rect 32394 18411 32410 18437
rect 32410 18411 32422 18437
rect 32342 18410 32370 18411
rect 32394 18410 32422 18411
rect 32446 18437 32474 18438
rect 32446 18411 32472 18437
rect 32472 18411 32474 18437
rect 32446 18410 32474 18411
rect 32498 18437 32526 18438
rect 32498 18411 32508 18437
rect 32508 18411 32526 18437
rect 32498 18410 32526 18411
rect 34582 18045 34610 18046
rect 34582 18019 34600 18045
rect 34600 18019 34610 18045
rect 34582 18018 34610 18019
rect 34634 18045 34662 18046
rect 34634 18019 34636 18045
rect 34636 18019 34662 18045
rect 34634 18018 34662 18019
rect 34686 18045 34714 18046
rect 34738 18045 34766 18046
rect 34686 18019 34698 18045
rect 34698 18019 34714 18045
rect 34738 18019 34760 18045
rect 34760 18019 34766 18045
rect 34686 18018 34714 18019
rect 34738 18018 34766 18019
rect 34790 18018 34818 18046
rect 34842 18045 34870 18046
rect 34894 18045 34922 18046
rect 34842 18019 34848 18045
rect 34848 18019 34870 18045
rect 34894 18019 34910 18045
rect 34910 18019 34922 18045
rect 34842 18018 34870 18019
rect 34894 18018 34922 18019
rect 34946 18045 34974 18046
rect 34946 18019 34972 18045
rect 34972 18019 34974 18045
rect 34946 18018 34974 18019
rect 34998 18045 35026 18046
rect 34998 18019 35008 18045
rect 35008 18019 35026 18045
rect 34998 18018 35026 18019
rect 32082 17653 32110 17654
rect 32082 17627 32100 17653
rect 32100 17627 32110 17653
rect 32082 17626 32110 17627
rect 32134 17653 32162 17654
rect 32134 17627 32136 17653
rect 32136 17627 32162 17653
rect 32134 17626 32162 17627
rect 32186 17653 32214 17654
rect 32238 17653 32266 17654
rect 32186 17627 32198 17653
rect 32198 17627 32214 17653
rect 32238 17627 32260 17653
rect 32260 17627 32266 17653
rect 32186 17626 32214 17627
rect 32238 17626 32266 17627
rect 32290 17626 32318 17654
rect 32342 17653 32370 17654
rect 32394 17653 32422 17654
rect 32342 17627 32348 17653
rect 32348 17627 32370 17653
rect 32394 17627 32410 17653
rect 32410 17627 32422 17653
rect 32342 17626 32370 17627
rect 32394 17626 32422 17627
rect 32446 17653 32474 17654
rect 32446 17627 32472 17653
rect 32472 17627 32474 17653
rect 32446 17626 32474 17627
rect 32498 17653 32526 17654
rect 32498 17627 32508 17653
rect 32508 17627 32526 17653
rect 32498 17626 32526 17627
rect 34582 17261 34610 17262
rect 34582 17235 34600 17261
rect 34600 17235 34610 17261
rect 34582 17234 34610 17235
rect 34634 17261 34662 17262
rect 34634 17235 34636 17261
rect 34636 17235 34662 17261
rect 34634 17234 34662 17235
rect 34686 17261 34714 17262
rect 34738 17261 34766 17262
rect 34686 17235 34698 17261
rect 34698 17235 34714 17261
rect 34738 17235 34760 17261
rect 34760 17235 34766 17261
rect 34686 17234 34714 17235
rect 34738 17234 34766 17235
rect 34790 17234 34818 17262
rect 34842 17261 34870 17262
rect 34894 17261 34922 17262
rect 34842 17235 34848 17261
rect 34848 17235 34870 17261
rect 34894 17235 34910 17261
rect 34910 17235 34922 17261
rect 34842 17234 34870 17235
rect 34894 17234 34922 17235
rect 34946 17261 34974 17262
rect 34946 17235 34972 17261
rect 34972 17235 34974 17261
rect 34946 17234 34974 17235
rect 34998 17261 35026 17262
rect 34998 17235 35008 17261
rect 35008 17235 35026 17261
rect 34998 17234 35026 17235
rect 32082 16869 32110 16870
rect 32082 16843 32100 16869
rect 32100 16843 32110 16869
rect 32082 16842 32110 16843
rect 32134 16869 32162 16870
rect 32134 16843 32136 16869
rect 32136 16843 32162 16869
rect 32134 16842 32162 16843
rect 32186 16869 32214 16870
rect 32238 16869 32266 16870
rect 32186 16843 32198 16869
rect 32198 16843 32214 16869
rect 32238 16843 32260 16869
rect 32260 16843 32266 16869
rect 32186 16842 32214 16843
rect 32238 16842 32266 16843
rect 32290 16842 32318 16870
rect 32342 16869 32370 16870
rect 32394 16869 32422 16870
rect 32342 16843 32348 16869
rect 32348 16843 32370 16869
rect 32394 16843 32410 16869
rect 32410 16843 32422 16869
rect 32342 16842 32370 16843
rect 32394 16842 32422 16843
rect 32446 16869 32474 16870
rect 32446 16843 32472 16869
rect 32472 16843 32474 16869
rect 32446 16842 32474 16843
rect 32498 16869 32526 16870
rect 32498 16843 32508 16869
rect 32508 16843 32526 16869
rect 32498 16842 32526 16843
rect 34582 16477 34610 16478
rect 34582 16451 34600 16477
rect 34600 16451 34610 16477
rect 34582 16450 34610 16451
rect 34634 16477 34662 16478
rect 34634 16451 34636 16477
rect 34636 16451 34662 16477
rect 34634 16450 34662 16451
rect 34686 16477 34714 16478
rect 34738 16477 34766 16478
rect 34686 16451 34698 16477
rect 34698 16451 34714 16477
rect 34738 16451 34760 16477
rect 34760 16451 34766 16477
rect 34686 16450 34714 16451
rect 34738 16450 34766 16451
rect 34790 16450 34818 16478
rect 34842 16477 34870 16478
rect 34894 16477 34922 16478
rect 34842 16451 34848 16477
rect 34848 16451 34870 16477
rect 34894 16451 34910 16477
rect 34910 16451 34922 16477
rect 34842 16450 34870 16451
rect 34894 16450 34922 16451
rect 34946 16477 34974 16478
rect 34946 16451 34972 16477
rect 34972 16451 34974 16477
rect 34946 16450 34974 16451
rect 34998 16477 35026 16478
rect 34998 16451 35008 16477
rect 35008 16451 35026 16477
rect 34998 16450 35026 16451
rect 32082 16085 32110 16086
rect 32082 16059 32100 16085
rect 32100 16059 32110 16085
rect 32082 16058 32110 16059
rect 32134 16085 32162 16086
rect 32134 16059 32136 16085
rect 32136 16059 32162 16085
rect 32134 16058 32162 16059
rect 32186 16085 32214 16086
rect 32238 16085 32266 16086
rect 32186 16059 32198 16085
rect 32198 16059 32214 16085
rect 32238 16059 32260 16085
rect 32260 16059 32266 16085
rect 32186 16058 32214 16059
rect 32238 16058 32266 16059
rect 32290 16058 32318 16086
rect 32342 16085 32370 16086
rect 32394 16085 32422 16086
rect 32342 16059 32348 16085
rect 32348 16059 32370 16085
rect 32394 16059 32410 16085
rect 32410 16059 32422 16085
rect 32342 16058 32370 16059
rect 32394 16058 32422 16059
rect 32446 16085 32474 16086
rect 32446 16059 32472 16085
rect 32472 16059 32474 16085
rect 32446 16058 32474 16059
rect 32498 16085 32526 16086
rect 32498 16059 32508 16085
rect 32508 16059 32526 16085
rect 32498 16058 32526 16059
rect 34582 15693 34610 15694
rect 34582 15667 34600 15693
rect 34600 15667 34610 15693
rect 34582 15666 34610 15667
rect 34634 15693 34662 15694
rect 34634 15667 34636 15693
rect 34636 15667 34662 15693
rect 34634 15666 34662 15667
rect 34686 15693 34714 15694
rect 34738 15693 34766 15694
rect 34686 15667 34698 15693
rect 34698 15667 34714 15693
rect 34738 15667 34760 15693
rect 34760 15667 34766 15693
rect 34686 15666 34714 15667
rect 34738 15666 34766 15667
rect 34790 15666 34818 15694
rect 34842 15693 34870 15694
rect 34894 15693 34922 15694
rect 34842 15667 34848 15693
rect 34848 15667 34870 15693
rect 34894 15667 34910 15693
rect 34910 15667 34922 15693
rect 34842 15666 34870 15667
rect 34894 15666 34922 15667
rect 34946 15693 34974 15694
rect 34946 15667 34972 15693
rect 34972 15667 34974 15693
rect 34946 15666 34974 15667
rect 34998 15693 35026 15694
rect 34998 15667 35008 15693
rect 35008 15667 35026 15693
rect 34998 15666 35026 15667
rect 32082 15301 32110 15302
rect 32082 15275 32100 15301
rect 32100 15275 32110 15301
rect 32082 15274 32110 15275
rect 32134 15301 32162 15302
rect 32134 15275 32136 15301
rect 32136 15275 32162 15301
rect 32134 15274 32162 15275
rect 32186 15301 32214 15302
rect 32238 15301 32266 15302
rect 32186 15275 32198 15301
rect 32198 15275 32214 15301
rect 32238 15275 32260 15301
rect 32260 15275 32266 15301
rect 32186 15274 32214 15275
rect 32238 15274 32266 15275
rect 32290 15274 32318 15302
rect 32342 15301 32370 15302
rect 32394 15301 32422 15302
rect 32342 15275 32348 15301
rect 32348 15275 32370 15301
rect 32394 15275 32410 15301
rect 32410 15275 32422 15301
rect 32342 15274 32370 15275
rect 32394 15274 32422 15275
rect 32446 15301 32474 15302
rect 32446 15275 32472 15301
rect 32472 15275 32474 15301
rect 32446 15274 32474 15275
rect 32498 15301 32526 15302
rect 32498 15275 32508 15301
rect 32508 15275 32526 15301
rect 32498 15274 32526 15275
rect 34582 14909 34610 14910
rect 34582 14883 34600 14909
rect 34600 14883 34610 14909
rect 34582 14882 34610 14883
rect 34634 14909 34662 14910
rect 34634 14883 34636 14909
rect 34636 14883 34662 14909
rect 34634 14882 34662 14883
rect 34686 14909 34714 14910
rect 34738 14909 34766 14910
rect 34686 14883 34698 14909
rect 34698 14883 34714 14909
rect 34738 14883 34760 14909
rect 34760 14883 34766 14909
rect 34686 14882 34714 14883
rect 34738 14882 34766 14883
rect 34790 14882 34818 14910
rect 34842 14909 34870 14910
rect 34894 14909 34922 14910
rect 34842 14883 34848 14909
rect 34848 14883 34870 14909
rect 34894 14883 34910 14909
rect 34910 14883 34922 14909
rect 34842 14882 34870 14883
rect 34894 14882 34922 14883
rect 34946 14909 34974 14910
rect 34946 14883 34972 14909
rect 34972 14883 34974 14909
rect 34946 14882 34974 14883
rect 34998 14909 35026 14910
rect 34998 14883 35008 14909
rect 35008 14883 35026 14909
rect 34998 14882 35026 14883
rect 32082 14517 32110 14518
rect 32082 14491 32100 14517
rect 32100 14491 32110 14517
rect 32082 14490 32110 14491
rect 32134 14517 32162 14518
rect 32134 14491 32136 14517
rect 32136 14491 32162 14517
rect 32134 14490 32162 14491
rect 32186 14517 32214 14518
rect 32238 14517 32266 14518
rect 32186 14491 32198 14517
rect 32198 14491 32214 14517
rect 32238 14491 32260 14517
rect 32260 14491 32266 14517
rect 32186 14490 32214 14491
rect 32238 14490 32266 14491
rect 32290 14490 32318 14518
rect 32342 14517 32370 14518
rect 32394 14517 32422 14518
rect 32342 14491 32348 14517
rect 32348 14491 32370 14517
rect 32394 14491 32410 14517
rect 32410 14491 32422 14517
rect 32342 14490 32370 14491
rect 32394 14490 32422 14491
rect 32446 14517 32474 14518
rect 32446 14491 32472 14517
rect 32472 14491 32474 14517
rect 32446 14490 32474 14491
rect 32498 14517 32526 14518
rect 32498 14491 32508 14517
rect 32508 14491 32526 14517
rect 32498 14490 32526 14491
rect 34582 14125 34610 14126
rect 34582 14099 34600 14125
rect 34600 14099 34610 14125
rect 34582 14098 34610 14099
rect 34634 14125 34662 14126
rect 34634 14099 34636 14125
rect 34636 14099 34662 14125
rect 34634 14098 34662 14099
rect 34686 14125 34714 14126
rect 34738 14125 34766 14126
rect 34686 14099 34698 14125
rect 34698 14099 34714 14125
rect 34738 14099 34760 14125
rect 34760 14099 34766 14125
rect 34686 14098 34714 14099
rect 34738 14098 34766 14099
rect 34790 14098 34818 14126
rect 34842 14125 34870 14126
rect 34894 14125 34922 14126
rect 34842 14099 34848 14125
rect 34848 14099 34870 14125
rect 34894 14099 34910 14125
rect 34910 14099 34922 14125
rect 34842 14098 34870 14099
rect 34894 14098 34922 14099
rect 34946 14125 34974 14126
rect 34946 14099 34972 14125
rect 34972 14099 34974 14125
rect 34946 14098 34974 14099
rect 34998 14125 35026 14126
rect 34998 14099 35008 14125
rect 35008 14099 35026 14125
rect 34998 14098 35026 14099
rect 32082 13733 32110 13734
rect 32082 13707 32100 13733
rect 32100 13707 32110 13733
rect 32082 13706 32110 13707
rect 32134 13733 32162 13734
rect 32134 13707 32136 13733
rect 32136 13707 32162 13733
rect 32134 13706 32162 13707
rect 32186 13733 32214 13734
rect 32238 13733 32266 13734
rect 32186 13707 32198 13733
rect 32198 13707 32214 13733
rect 32238 13707 32260 13733
rect 32260 13707 32266 13733
rect 32186 13706 32214 13707
rect 32238 13706 32266 13707
rect 32290 13706 32318 13734
rect 32342 13733 32370 13734
rect 32394 13733 32422 13734
rect 32342 13707 32348 13733
rect 32348 13707 32370 13733
rect 32394 13707 32410 13733
rect 32410 13707 32422 13733
rect 32342 13706 32370 13707
rect 32394 13706 32422 13707
rect 32446 13733 32474 13734
rect 32446 13707 32472 13733
rect 32472 13707 32474 13733
rect 32446 13706 32474 13707
rect 32498 13733 32526 13734
rect 32498 13707 32508 13733
rect 32508 13707 32526 13733
rect 32498 13706 32526 13707
rect 34582 13341 34610 13342
rect 34582 13315 34600 13341
rect 34600 13315 34610 13341
rect 34582 13314 34610 13315
rect 34634 13341 34662 13342
rect 34634 13315 34636 13341
rect 34636 13315 34662 13341
rect 34634 13314 34662 13315
rect 34686 13341 34714 13342
rect 34738 13341 34766 13342
rect 34686 13315 34698 13341
rect 34698 13315 34714 13341
rect 34738 13315 34760 13341
rect 34760 13315 34766 13341
rect 34686 13314 34714 13315
rect 34738 13314 34766 13315
rect 34790 13314 34818 13342
rect 34842 13341 34870 13342
rect 34894 13341 34922 13342
rect 34842 13315 34848 13341
rect 34848 13315 34870 13341
rect 34894 13315 34910 13341
rect 34910 13315 34922 13341
rect 34842 13314 34870 13315
rect 34894 13314 34922 13315
rect 34946 13341 34974 13342
rect 34946 13315 34972 13341
rect 34972 13315 34974 13341
rect 34946 13314 34974 13315
rect 34998 13341 35026 13342
rect 34998 13315 35008 13341
rect 35008 13315 35026 13341
rect 34998 13314 35026 13315
rect 32082 12949 32110 12950
rect 32082 12923 32100 12949
rect 32100 12923 32110 12949
rect 32082 12922 32110 12923
rect 32134 12949 32162 12950
rect 32134 12923 32136 12949
rect 32136 12923 32162 12949
rect 32134 12922 32162 12923
rect 32186 12949 32214 12950
rect 32238 12949 32266 12950
rect 32186 12923 32198 12949
rect 32198 12923 32214 12949
rect 32238 12923 32260 12949
rect 32260 12923 32266 12949
rect 32186 12922 32214 12923
rect 32238 12922 32266 12923
rect 32290 12922 32318 12950
rect 32342 12949 32370 12950
rect 32394 12949 32422 12950
rect 32342 12923 32348 12949
rect 32348 12923 32370 12949
rect 32394 12923 32410 12949
rect 32410 12923 32422 12949
rect 32342 12922 32370 12923
rect 32394 12922 32422 12923
rect 32446 12949 32474 12950
rect 32446 12923 32472 12949
rect 32472 12923 32474 12949
rect 32446 12922 32474 12923
rect 32498 12949 32526 12950
rect 32498 12923 32508 12949
rect 32508 12923 32526 12949
rect 32498 12922 32526 12923
rect 34582 12557 34610 12558
rect 34582 12531 34600 12557
rect 34600 12531 34610 12557
rect 34582 12530 34610 12531
rect 34634 12557 34662 12558
rect 34634 12531 34636 12557
rect 34636 12531 34662 12557
rect 34634 12530 34662 12531
rect 34686 12557 34714 12558
rect 34738 12557 34766 12558
rect 34686 12531 34698 12557
rect 34698 12531 34714 12557
rect 34738 12531 34760 12557
rect 34760 12531 34766 12557
rect 34686 12530 34714 12531
rect 34738 12530 34766 12531
rect 34790 12530 34818 12558
rect 34842 12557 34870 12558
rect 34894 12557 34922 12558
rect 34842 12531 34848 12557
rect 34848 12531 34870 12557
rect 34894 12531 34910 12557
rect 34910 12531 34922 12557
rect 34842 12530 34870 12531
rect 34894 12530 34922 12531
rect 34946 12557 34974 12558
rect 34946 12531 34972 12557
rect 34972 12531 34974 12557
rect 34946 12530 34974 12531
rect 34998 12557 35026 12558
rect 34998 12531 35008 12557
rect 35008 12531 35026 12557
rect 34998 12530 35026 12531
rect 32082 12165 32110 12166
rect 32082 12139 32100 12165
rect 32100 12139 32110 12165
rect 32082 12138 32110 12139
rect 32134 12165 32162 12166
rect 32134 12139 32136 12165
rect 32136 12139 32162 12165
rect 32134 12138 32162 12139
rect 32186 12165 32214 12166
rect 32238 12165 32266 12166
rect 32186 12139 32198 12165
rect 32198 12139 32214 12165
rect 32238 12139 32260 12165
rect 32260 12139 32266 12165
rect 32186 12138 32214 12139
rect 32238 12138 32266 12139
rect 32290 12138 32318 12166
rect 32342 12165 32370 12166
rect 32394 12165 32422 12166
rect 32342 12139 32348 12165
rect 32348 12139 32370 12165
rect 32394 12139 32410 12165
rect 32410 12139 32422 12165
rect 32342 12138 32370 12139
rect 32394 12138 32422 12139
rect 32446 12165 32474 12166
rect 32446 12139 32472 12165
rect 32472 12139 32474 12165
rect 32446 12138 32474 12139
rect 32498 12165 32526 12166
rect 32498 12139 32508 12165
rect 32508 12139 32526 12165
rect 32498 12138 32526 12139
rect 31934 11606 31962 11634
rect 32830 11969 32858 11970
rect 32830 11943 32831 11969
rect 32831 11943 32857 11969
rect 32857 11943 32858 11969
rect 32830 11942 32858 11943
rect 33110 11942 33138 11970
rect 32438 11550 32466 11578
rect 32774 11577 32802 11578
rect 32774 11551 32775 11577
rect 32775 11551 32801 11577
rect 32801 11551 32802 11577
rect 32774 11550 32802 11551
rect 32082 11381 32110 11382
rect 32082 11355 32100 11381
rect 32100 11355 32110 11381
rect 32082 11354 32110 11355
rect 32134 11381 32162 11382
rect 32134 11355 32136 11381
rect 32136 11355 32162 11381
rect 32134 11354 32162 11355
rect 32186 11381 32214 11382
rect 32238 11381 32266 11382
rect 32186 11355 32198 11381
rect 32198 11355 32214 11381
rect 32238 11355 32260 11381
rect 32260 11355 32266 11381
rect 32186 11354 32214 11355
rect 32238 11354 32266 11355
rect 32290 11354 32318 11382
rect 32342 11381 32370 11382
rect 32394 11381 32422 11382
rect 32342 11355 32348 11381
rect 32348 11355 32370 11381
rect 32394 11355 32410 11381
rect 32410 11355 32422 11381
rect 32342 11354 32370 11355
rect 32394 11354 32422 11355
rect 32446 11381 32474 11382
rect 32446 11355 32472 11381
rect 32472 11355 32474 11381
rect 32446 11354 32474 11355
rect 32498 11381 32526 11382
rect 32498 11355 32508 11381
rect 32508 11355 32526 11381
rect 32498 11354 32526 11355
rect 30758 10038 30786 10066
rect 30702 9982 30730 10010
rect 30814 10009 30842 10010
rect 30814 9983 30815 10009
rect 30815 9983 30841 10009
rect 30841 9983 30842 10009
rect 30814 9982 30842 9983
rect 30814 9702 30842 9730
rect 32438 11185 32466 11186
rect 32438 11159 32439 11185
rect 32439 11159 32465 11185
rect 32465 11159 32466 11185
rect 32438 11158 32466 11159
rect 34582 11773 34610 11774
rect 34582 11747 34600 11773
rect 34600 11747 34610 11773
rect 34582 11746 34610 11747
rect 34634 11773 34662 11774
rect 34634 11747 34636 11773
rect 34636 11747 34662 11773
rect 34634 11746 34662 11747
rect 34686 11773 34714 11774
rect 34738 11773 34766 11774
rect 34686 11747 34698 11773
rect 34698 11747 34714 11773
rect 34738 11747 34760 11773
rect 34760 11747 34766 11773
rect 34686 11746 34714 11747
rect 34738 11746 34766 11747
rect 34790 11746 34818 11774
rect 34842 11773 34870 11774
rect 34894 11773 34922 11774
rect 34842 11747 34848 11773
rect 34848 11747 34870 11773
rect 34894 11747 34910 11773
rect 34910 11747 34922 11773
rect 34842 11746 34870 11747
rect 34894 11746 34922 11747
rect 34946 11773 34974 11774
rect 34946 11747 34972 11773
rect 34972 11747 34974 11773
rect 34946 11746 34974 11747
rect 34998 11773 35026 11774
rect 34998 11747 35008 11773
rect 35008 11747 35026 11773
rect 34998 11746 35026 11747
rect 33166 11577 33194 11578
rect 33166 11551 33167 11577
rect 33167 11551 33193 11577
rect 33193 11551 33194 11577
rect 33166 11550 33194 11551
rect 33614 11577 33642 11578
rect 33614 11551 33615 11577
rect 33615 11551 33641 11577
rect 33641 11551 33642 11577
rect 33614 11550 33642 11551
rect 34510 11550 34538 11578
rect 34510 11214 34538 11242
rect 32774 11158 32802 11186
rect 32082 10597 32110 10598
rect 32082 10571 32100 10597
rect 32100 10571 32110 10597
rect 32082 10570 32110 10571
rect 32134 10597 32162 10598
rect 32134 10571 32136 10597
rect 32136 10571 32162 10597
rect 32134 10570 32162 10571
rect 32186 10597 32214 10598
rect 32238 10597 32266 10598
rect 32186 10571 32198 10597
rect 32198 10571 32214 10597
rect 32238 10571 32260 10597
rect 32260 10571 32266 10597
rect 32186 10570 32214 10571
rect 32238 10570 32266 10571
rect 32290 10570 32318 10598
rect 32342 10597 32370 10598
rect 32394 10597 32422 10598
rect 32342 10571 32348 10597
rect 32348 10571 32370 10597
rect 32394 10571 32410 10597
rect 32410 10571 32422 10597
rect 32342 10570 32370 10571
rect 32394 10570 32422 10571
rect 32446 10597 32474 10598
rect 32446 10571 32472 10597
rect 32472 10571 32474 10597
rect 32446 10570 32474 10571
rect 32498 10597 32526 10598
rect 32498 10571 32508 10597
rect 32508 10571 32526 10597
rect 32498 10570 32526 10571
rect 32158 10038 32186 10066
rect 31094 9870 31122 9898
rect 30982 9225 31010 9226
rect 30982 9199 30983 9225
rect 30983 9199 31009 9225
rect 31009 9199 31010 9225
rect 30982 9198 31010 9199
rect 31374 9617 31402 9618
rect 31374 9591 31375 9617
rect 31375 9591 31401 9617
rect 31401 9591 31402 9617
rect 31374 9590 31402 9591
rect 31038 8441 31066 8442
rect 31038 8415 31039 8441
rect 31039 8415 31065 8441
rect 31065 8415 31066 8441
rect 31038 8414 31066 8415
rect 31150 8833 31178 8834
rect 31150 8807 31151 8833
rect 31151 8807 31177 8833
rect 31177 8807 31178 8833
rect 31150 8806 31178 8807
rect 32830 10038 32858 10066
rect 32886 9982 32914 10010
rect 32774 9870 32802 9898
rect 32082 9813 32110 9814
rect 32082 9787 32100 9813
rect 32100 9787 32110 9813
rect 32082 9786 32110 9787
rect 32134 9813 32162 9814
rect 32134 9787 32136 9813
rect 32136 9787 32162 9813
rect 32134 9786 32162 9787
rect 32186 9813 32214 9814
rect 32238 9813 32266 9814
rect 32186 9787 32198 9813
rect 32198 9787 32214 9813
rect 32238 9787 32260 9813
rect 32260 9787 32266 9813
rect 32186 9786 32214 9787
rect 32238 9786 32266 9787
rect 32290 9786 32318 9814
rect 32342 9813 32370 9814
rect 32394 9813 32422 9814
rect 32342 9787 32348 9813
rect 32348 9787 32370 9813
rect 32394 9787 32410 9813
rect 32410 9787 32422 9813
rect 32342 9786 32370 9787
rect 32394 9786 32422 9787
rect 32446 9813 32474 9814
rect 32446 9787 32472 9813
rect 32472 9787 32474 9813
rect 32446 9786 32474 9787
rect 32498 9813 32526 9814
rect 32498 9787 32508 9813
rect 32508 9787 32526 9813
rect 32498 9786 32526 9787
rect 31374 8833 31402 8834
rect 31374 8807 31375 8833
rect 31375 8807 31401 8833
rect 31401 8807 31402 8833
rect 31374 8806 31402 8807
rect 31990 9702 32018 9730
rect 32158 9702 32186 9730
rect 32082 9029 32110 9030
rect 32082 9003 32100 9029
rect 32100 9003 32110 9029
rect 32082 9002 32110 9003
rect 32134 9029 32162 9030
rect 32134 9003 32136 9029
rect 32136 9003 32162 9029
rect 32134 9002 32162 9003
rect 32186 9029 32214 9030
rect 32238 9029 32266 9030
rect 32186 9003 32198 9029
rect 32198 9003 32214 9029
rect 32238 9003 32260 9029
rect 32260 9003 32266 9029
rect 32186 9002 32214 9003
rect 32238 9002 32266 9003
rect 32290 9002 32318 9030
rect 32342 9029 32370 9030
rect 32394 9029 32422 9030
rect 32342 9003 32348 9029
rect 32348 9003 32370 9029
rect 32394 9003 32410 9029
rect 32410 9003 32422 9029
rect 32342 9002 32370 9003
rect 32394 9002 32422 9003
rect 32446 9029 32474 9030
rect 32446 9003 32472 9029
rect 32472 9003 32474 9029
rect 32446 9002 32474 9003
rect 32498 9029 32526 9030
rect 32498 9003 32508 9029
rect 32508 9003 32526 9029
rect 32498 9002 32526 9003
rect 31430 8470 31458 8498
rect 31934 8414 31962 8442
rect 32158 8414 32186 8442
rect 32718 8441 32746 8442
rect 32718 8415 32719 8441
rect 32719 8415 32745 8441
rect 32745 8415 32746 8441
rect 32718 8414 32746 8415
rect 32082 8245 32110 8246
rect 32082 8219 32100 8245
rect 32100 8219 32110 8245
rect 32082 8218 32110 8219
rect 32134 8245 32162 8246
rect 32134 8219 32136 8245
rect 32136 8219 32162 8245
rect 32134 8218 32162 8219
rect 32186 8245 32214 8246
rect 32238 8245 32266 8246
rect 32186 8219 32198 8245
rect 32198 8219 32214 8245
rect 32238 8219 32260 8245
rect 32260 8219 32266 8245
rect 32186 8218 32214 8219
rect 32238 8218 32266 8219
rect 32290 8218 32318 8246
rect 32342 8245 32370 8246
rect 32394 8245 32422 8246
rect 32342 8219 32348 8245
rect 32348 8219 32370 8245
rect 32394 8219 32410 8245
rect 32410 8219 32422 8245
rect 32342 8218 32370 8219
rect 32394 8218 32422 8219
rect 32446 8245 32474 8246
rect 32446 8219 32472 8245
rect 32472 8219 32474 8245
rect 32446 8218 32474 8219
rect 32498 8245 32526 8246
rect 32498 8219 32508 8245
rect 32508 8219 32526 8245
rect 32498 8218 32526 8219
rect 31934 8022 31962 8050
rect 32438 8049 32466 8050
rect 32438 8023 32439 8049
rect 32439 8023 32465 8049
rect 32465 8023 32466 8049
rect 32438 8022 32466 8023
rect 32830 9617 32858 9618
rect 32830 9591 32831 9617
rect 32831 9591 32857 9617
rect 32857 9591 32858 9617
rect 32830 9590 32858 9591
rect 32830 9142 32858 9170
rect 32942 10038 32970 10066
rect 32942 9422 32970 9450
rect 35126 11214 35154 11242
rect 34958 11185 34986 11186
rect 34958 11159 34959 11185
rect 34959 11159 34985 11185
rect 34985 11159 34986 11185
rect 34958 11158 34986 11159
rect 35350 11214 35378 11242
rect 34582 10989 34610 10990
rect 34582 10963 34600 10989
rect 34600 10963 34610 10989
rect 34582 10962 34610 10963
rect 34634 10989 34662 10990
rect 34634 10963 34636 10989
rect 34636 10963 34662 10989
rect 34634 10962 34662 10963
rect 34686 10989 34714 10990
rect 34738 10989 34766 10990
rect 34686 10963 34698 10989
rect 34698 10963 34714 10989
rect 34738 10963 34760 10989
rect 34760 10963 34766 10989
rect 34686 10962 34714 10963
rect 34738 10962 34766 10963
rect 34790 10962 34818 10990
rect 34842 10989 34870 10990
rect 34894 10989 34922 10990
rect 34842 10963 34848 10989
rect 34848 10963 34870 10989
rect 34894 10963 34910 10989
rect 34910 10963 34922 10989
rect 34842 10962 34870 10963
rect 34894 10962 34922 10963
rect 34946 10989 34974 10990
rect 34946 10963 34972 10989
rect 34972 10963 34974 10989
rect 34946 10962 34974 10963
rect 34998 10989 35026 10990
rect 34998 10963 35008 10989
rect 35008 10963 35026 10989
rect 34998 10962 35026 10963
rect 34454 10374 34482 10402
rect 34958 10401 34986 10402
rect 34958 10375 34959 10401
rect 34959 10375 34985 10401
rect 34985 10375 34986 10401
rect 34958 10374 34986 10375
rect 36134 11185 36162 11186
rect 36134 11159 36135 11185
rect 36135 11159 36161 11185
rect 36161 11159 36162 11185
rect 36134 11158 36162 11159
rect 36694 10710 36722 10738
rect 36246 10374 36274 10402
rect 35350 10318 35378 10346
rect 34582 10205 34610 10206
rect 34582 10179 34600 10205
rect 34600 10179 34610 10205
rect 34582 10178 34610 10179
rect 34634 10205 34662 10206
rect 34634 10179 34636 10205
rect 34636 10179 34662 10205
rect 34634 10178 34662 10179
rect 34686 10205 34714 10206
rect 34738 10205 34766 10206
rect 34686 10179 34698 10205
rect 34698 10179 34714 10205
rect 34738 10179 34760 10205
rect 34760 10179 34766 10205
rect 34686 10178 34714 10179
rect 34738 10178 34766 10179
rect 34790 10178 34818 10206
rect 34842 10205 34870 10206
rect 34894 10205 34922 10206
rect 34842 10179 34848 10205
rect 34848 10179 34870 10205
rect 34894 10179 34910 10205
rect 34910 10179 34922 10205
rect 34842 10178 34870 10179
rect 34894 10178 34922 10179
rect 34946 10205 34974 10206
rect 34946 10179 34972 10205
rect 34972 10179 34974 10205
rect 34946 10178 34974 10179
rect 34998 10205 35026 10206
rect 34998 10179 35008 10205
rect 35008 10179 35026 10205
rect 34998 10178 35026 10179
rect 34454 10094 34482 10122
rect 32886 8862 32914 8890
rect 32774 7966 32802 7994
rect 32830 8750 32858 8778
rect 33110 9590 33138 9618
rect 33110 8777 33138 8778
rect 33110 8751 33111 8777
rect 33111 8751 33137 8777
rect 33137 8751 33138 8777
rect 33110 8750 33138 8751
rect 32830 8470 32858 8498
rect 32438 7574 32466 7602
rect 32606 7574 32634 7602
rect 32082 7461 32110 7462
rect 32082 7435 32100 7461
rect 32100 7435 32110 7461
rect 32082 7434 32110 7435
rect 32134 7461 32162 7462
rect 32134 7435 32136 7461
rect 32136 7435 32162 7461
rect 32134 7434 32162 7435
rect 32186 7461 32214 7462
rect 32238 7461 32266 7462
rect 32186 7435 32198 7461
rect 32198 7435 32214 7461
rect 32238 7435 32260 7461
rect 32260 7435 32266 7461
rect 32186 7434 32214 7435
rect 32238 7434 32266 7435
rect 32290 7434 32318 7462
rect 32342 7461 32370 7462
rect 32394 7461 32422 7462
rect 32342 7435 32348 7461
rect 32348 7435 32370 7461
rect 32394 7435 32410 7461
rect 32410 7435 32422 7461
rect 32342 7434 32370 7435
rect 32394 7434 32422 7435
rect 32446 7461 32474 7462
rect 32446 7435 32472 7461
rect 32472 7435 32474 7461
rect 32446 7434 32474 7435
rect 32498 7461 32526 7462
rect 32498 7435 32508 7461
rect 32508 7435 32526 7461
rect 32498 7434 32526 7435
rect 33166 8358 33194 8386
rect 34622 10009 34650 10010
rect 34622 9983 34623 10009
rect 34623 9983 34649 10009
rect 34649 9983 34650 10009
rect 34622 9982 34650 9983
rect 34846 10009 34874 10010
rect 34846 9983 34847 10009
rect 34847 9983 34873 10009
rect 34873 9983 34874 10009
rect 34846 9982 34874 9983
rect 35126 9982 35154 10010
rect 34454 9870 34482 9898
rect 34454 9478 34482 9506
rect 35350 9617 35378 9618
rect 35350 9591 35351 9617
rect 35351 9591 35377 9617
rect 35377 9591 35378 9617
rect 35350 9590 35378 9591
rect 36414 9926 36442 9954
rect 36694 9926 36722 9954
rect 34958 9478 34986 9506
rect 36414 9478 36442 9506
rect 34174 9422 34202 9450
rect 34582 9421 34610 9422
rect 34582 9395 34600 9421
rect 34600 9395 34610 9421
rect 34582 9394 34610 9395
rect 34634 9421 34662 9422
rect 34634 9395 34636 9421
rect 34636 9395 34662 9421
rect 34634 9394 34662 9395
rect 34686 9421 34714 9422
rect 34738 9421 34766 9422
rect 34686 9395 34698 9421
rect 34698 9395 34714 9421
rect 34738 9395 34760 9421
rect 34760 9395 34766 9421
rect 34686 9394 34714 9395
rect 34738 9394 34766 9395
rect 34790 9394 34818 9422
rect 34842 9421 34870 9422
rect 34894 9421 34922 9422
rect 34842 9395 34848 9421
rect 34848 9395 34870 9421
rect 34894 9395 34910 9421
rect 34910 9395 34922 9421
rect 34842 9394 34870 9395
rect 34894 9394 34922 9395
rect 34946 9421 34974 9422
rect 34946 9395 34972 9421
rect 34972 9395 34974 9421
rect 34946 9394 34974 9395
rect 34998 9421 35026 9422
rect 34998 9395 35008 9421
rect 35008 9395 35026 9421
rect 34998 9394 35026 9395
rect 34174 9254 34202 9282
rect 34678 9254 34706 9282
rect 34398 8414 34426 8442
rect 33614 8358 33642 8386
rect 32830 7238 32858 7266
rect 32998 7574 33026 7602
rect 32998 6734 33026 6762
rect 33390 7657 33418 7658
rect 33390 7631 33391 7657
rect 33391 7631 33417 7657
rect 33417 7631 33418 7657
rect 33390 7630 33418 7631
rect 32082 6677 32110 6678
rect 32082 6651 32100 6677
rect 32100 6651 32110 6677
rect 32082 6650 32110 6651
rect 32134 6677 32162 6678
rect 32134 6651 32136 6677
rect 32136 6651 32162 6677
rect 32134 6650 32162 6651
rect 32186 6677 32214 6678
rect 32238 6677 32266 6678
rect 32186 6651 32198 6677
rect 32198 6651 32214 6677
rect 32238 6651 32260 6677
rect 32260 6651 32266 6677
rect 32186 6650 32214 6651
rect 32238 6650 32266 6651
rect 32290 6650 32318 6678
rect 32342 6677 32370 6678
rect 32394 6677 32422 6678
rect 32342 6651 32348 6677
rect 32348 6651 32370 6677
rect 32394 6651 32410 6677
rect 32410 6651 32422 6677
rect 32342 6650 32370 6651
rect 32394 6650 32422 6651
rect 32446 6677 32474 6678
rect 32446 6651 32472 6677
rect 32472 6651 32474 6677
rect 32446 6650 32474 6651
rect 32498 6677 32526 6678
rect 32498 6651 32508 6677
rect 32508 6651 32526 6677
rect 32498 6650 32526 6651
rect 33334 7265 33362 7266
rect 33334 7239 33335 7265
rect 33335 7239 33361 7265
rect 33361 7239 33362 7265
rect 33334 7238 33362 7239
rect 33334 6734 33362 6762
rect 31822 5838 31850 5866
rect 32082 5893 32110 5894
rect 32082 5867 32100 5893
rect 32100 5867 32110 5893
rect 32082 5866 32110 5867
rect 32134 5893 32162 5894
rect 32134 5867 32136 5893
rect 32136 5867 32162 5893
rect 32134 5866 32162 5867
rect 32186 5893 32214 5894
rect 32238 5893 32266 5894
rect 32186 5867 32198 5893
rect 32198 5867 32214 5893
rect 32238 5867 32260 5893
rect 32260 5867 32266 5893
rect 32186 5866 32214 5867
rect 32238 5866 32266 5867
rect 32290 5866 32318 5894
rect 32342 5893 32370 5894
rect 32394 5893 32422 5894
rect 32342 5867 32348 5893
rect 32348 5867 32370 5893
rect 32394 5867 32410 5893
rect 32410 5867 32422 5893
rect 32342 5866 32370 5867
rect 32394 5866 32422 5867
rect 32446 5893 32474 5894
rect 32446 5867 32472 5893
rect 32472 5867 32474 5893
rect 32446 5866 32474 5867
rect 32498 5893 32526 5894
rect 32498 5867 32508 5893
rect 32508 5867 32526 5893
rect 32498 5866 32526 5867
rect 32438 5697 32466 5698
rect 32438 5671 32439 5697
rect 32439 5671 32465 5697
rect 32465 5671 32466 5697
rect 32438 5670 32466 5671
rect 32718 5670 32746 5698
rect 30926 5305 30954 5306
rect 30926 5279 30927 5305
rect 30927 5279 30953 5305
rect 30953 5279 30954 5305
rect 30926 5278 30954 5279
rect 30366 4998 30394 5026
rect 30310 4073 30338 4074
rect 30310 4047 30311 4073
rect 30311 4047 30337 4073
rect 30337 4047 30338 4073
rect 30310 4046 30338 4047
rect 32718 5305 32746 5306
rect 32718 5279 32719 5305
rect 32719 5279 32745 5305
rect 32745 5279 32746 5305
rect 32718 5278 32746 5279
rect 32082 5109 32110 5110
rect 32082 5083 32100 5109
rect 32100 5083 32110 5109
rect 32082 5082 32110 5083
rect 32134 5109 32162 5110
rect 32134 5083 32136 5109
rect 32136 5083 32162 5109
rect 32134 5082 32162 5083
rect 32186 5109 32214 5110
rect 32238 5109 32266 5110
rect 32186 5083 32198 5109
rect 32198 5083 32214 5109
rect 32238 5083 32260 5109
rect 32260 5083 32266 5109
rect 32186 5082 32214 5083
rect 32238 5082 32266 5083
rect 32290 5082 32318 5110
rect 32342 5109 32370 5110
rect 32394 5109 32422 5110
rect 32342 5083 32348 5109
rect 32348 5083 32370 5109
rect 32394 5083 32410 5109
rect 32410 5083 32422 5109
rect 32342 5082 32370 5083
rect 32394 5082 32422 5083
rect 32446 5109 32474 5110
rect 32446 5083 32472 5109
rect 32472 5083 32474 5109
rect 32446 5082 32474 5083
rect 32498 5109 32526 5110
rect 32498 5083 32508 5109
rect 32508 5083 32526 5109
rect 32498 5082 32526 5083
rect 30982 4214 31010 4242
rect 30478 3374 30506 3402
rect 30814 3822 30842 3850
rect 30702 3345 30730 3346
rect 30702 3319 30703 3345
rect 30703 3319 30729 3345
rect 30729 3319 30730 3345
rect 30702 3318 30730 3319
rect 30310 2982 30338 3010
rect 30310 2590 30338 2618
rect 30702 2534 30730 2562
rect 31934 4830 31962 4858
rect 31934 4494 31962 4522
rect 32046 4521 32074 4522
rect 32046 4495 32047 4521
rect 32047 4495 32073 4521
rect 32073 4495 32074 4521
rect 32046 4494 32074 4495
rect 32158 4438 32186 4466
rect 32326 4438 32354 4466
rect 33390 5222 33418 5250
rect 33670 5894 33698 5922
rect 33726 6481 33754 6482
rect 33726 6455 33727 6481
rect 33727 6455 33753 6481
rect 33753 6455 33754 6481
rect 33726 6454 33754 6455
rect 33670 5054 33698 5082
rect 32082 4325 32110 4326
rect 32082 4299 32100 4325
rect 32100 4299 32110 4325
rect 32082 4298 32110 4299
rect 32134 4325 32162 4326
rect 32134 4299 32136 4325
rect 32136 4299 32162 4325
rect 32134 4298 32162 4299
rect 32186 4325 32214 4326
rect 32238 4325 32266 4326
rect 32186 4299 32198 4325
rect 32198 4299 32214 4325
rect 32238 4299 32260 4325
rect 32260 4299 32266 4325
rect 32186 4298 32214 4299
rect 32238 4298 32266 4299
rect 32290 4298 32318 4326
rect 32342 4325 32370 4326
rect 32394 4325 32422 4326
rect 32342 4299 32348 4325
rect 32348 4299 32370 4325
rect 32394 4299 32410 4325
rect 32410 4299 32422 4325
rect 32342 4298 32370 4299
rect 32394 4298 32422 4299
rect 32446 4325 32474 4326
rect 32446 4299 32472 4325
rect 32472 4299 32474 4325
rect 32446 4298 32474 4299
rect 32498 4325 32526 4326
rect 32498 4299 32508 4325
rect 32508 4299 32526 4325
rect 32498 4298 32526 4299
rect 31990 4214 32018 4242
rect 32158 4214 32186 4242
rect 32718 4214 32746 4242
rect 30982 3374 31010 3402
rect 31598 3318 31626 3346
rect 31318 2926 31346 2954
rect 31262 2142 31290 2170
rect 31486 2142 31514 2170
rect 30310 1777 30338 1778
rect 30310 1751 30311 1777
rect 30311 1751 30337 1777
rect 30337 1751 30338 1777
rect 30310 1750 30338 1751
rect 31486 1721 31514 1722
rect 31486 1695 31487 1721
rect 31487 1695 31513 1721
rect 31513 1695 31514 1721
rect 31486 1694 31514 1695
rect 32158 3737 32186 3738
rect 32158 3711 32159 3737
rect 32159 3711 32185 3737
rect 32185 3711 32186 3737
rect 32158 3710 32186 3711
rect 32326 3737 32354 3738
rect 32326 3711 32327 3737
rect 32327 3711 32353 3737
rect 32353 3711 32354 3737
rect 32326 3710 32354 3711
rect 32082 3541 32110 3542
rect 32082 3515 32100 3541
rect 32100 3515 32110 3541
rect 32082 3514 32110 3515
rect 32134 3541 32162 3542
rect 32134 3515 32136 3541
rect 32136 3515 32162 3541
rect 32134 3514 32162 3515
rect 32186 3541 32214 3542
rect 32238 3541 32266 3542
rect 32186 3515 32198 3541
rect 32198 3515 32214 3541
rect 32238 3515 32260 3541
rect 32260 3515 32266 3541
rect 32186 3514 32214 3515
rect 32238 3514 32266 3515
rect 32290 3514 32318 3542
rect 32342 3541 32370 3542
rect 32394 3541 32422 3542
rect 32342 3515 32348 3541
rect 32348 3515 32370 3541
rect 32394 3515 32410 3541
rect 32410 3515 32422 3541
rect 32342 3514 32370 3515
rect 32394 3514 32422 3515
rect 32446 3541 32474 3542
rect 32446 3515 32472 3541
rect 32472 3515 32474 3541
rect 32446 3514 32474 3515
rect 32498 3541 32526 3542
rect 32498 3515 32508 3541
rect 32508 3515 32526 3541
rect 32498 3514 32526 3515
rect 32158 3009 32186 3010
rect 32158 2983 32159 3009
rect 32159 2983 32185 3009
rect 32185 2983 32186 3009
rect 32158 2982 32186 2983
rect 32326 3009 32354 3010
rect 32326 2983 32327 3009
rect 32327 2983 32353 3009
rect 32353 2983 32354 3009
rect 32326 2982 32354 2983
rect 32830 2926 32858 2954
rect 32886 2982 32914 3010
rect 32438 2870 32466 2898
rect 32082 2757 32110 2758
rect 32082 2731 32100 2757
rect 32100 2731 32110 2757
rect 32082 2730 32110 2731
rect 32134 2757 32162 2758
rect 32134 2731 32136 2757
rect 32136 2731 32162 2757
rect 32134 2730 32162 2731
rect 32186 2757 32214 2758
rect 32238 2757 32266 2758
rect 32186 2731 32198 2757
rect 32198 2731 32214 2757
rect 32238 2731 32260 2757
rect 32260 2731 32266 2757
rect 32186 2730 32214 2731
rect 32238 2730 32266 2731
rect 32290 2730 32318 2758
rect 32342 2757 32370 2758
rect 32394 2757 32422 2758
rect 32342 2731 32348 2757
rect 32348 2731 32370 2757
rect 32394 2731 32410 2757
rect 32410 2731 32422 2757
rect 32342 2730 32370 2731
rect 32394 2730 32422 2731
rect 32446 2757 32474 2758
rect 32446 2731 32472 2757
rect 32472 2731 32474 2757
rect 32446 2730 32474 2731
rect 32498 2757 32526 2758
rect 32498 2731 32508 2757
rect 32508 2731 32526 2757
rect 32498 2730 32526 2731
rect 32158 2561 32186 2562
rect 32158 2535 32159 2561
rect 32159 2535 32185 2561
rect 32185 2535 32186 2561
rect 32158 2534 32186 2535
rect 32606 2534 32634 2562
rect 32158 2225 32186 2226
rect 32158 2199 32159 2225
rect 32159 2199 32185 2225
rect 32185 2199 32186 2225
rect 32158 2198 32186 2199
rect 32326 2225 32354 2226
rect 32326 2199 32327 2225
rect 32327 2199 32353 2225
rect 32353 2199 32354 2225
rect 32326 2198 32354 2199
rect 32102 2169 32130 2170
rect 32102 2143 32103 2169
rect 32103 2143 32129 2169
rect 32129 2143 32130 2169
rect 32102 2142 32130 2143
rect 32082 1973 32110 1974
rect 32082 1947 32100 1973
rect 32100 1947 32110 1973
rect 32082 1946 32110 1947
rect 32134 1973 32162 1974
rect 32134 1947 32136 1973
rect 32136 1947 32162 1973
rect 32134 1946 32162 1947
rect 32186 1973 32214 1974
rect 32238 1973 32266 1974
rect 32186 1947 32198 1973
rect 32198 1947 32214 1973
rect 32238 1947 32260 1973
rect 32260 1947 32266 1973
rect 32186 1946 32214 1947
rect 32238 1946 32266 1947
rect 32290 1946 32318 1974
rect 32342 1973 32370 1974
rect 32394 1973 32422 1974
rect 32342 1947 32348 1973
rect 32348 1947 32370 1973
rect 32394 1947 32410 1973
rect 32410 1947 32422 1973
rect 32342 1946 32370 1947
rect 32394 1946 32422 1947
rect 32446 1973 32474 1974
rect 32446 1947 32472 1973
rect 32472 1947 32474 1973
rect 32446 1946 32474 1947
rect 32498 1973 32526 1974
rect 32498 1947 32508 1973
rect 32508 1947 32526 1973
rect 32498 1946 32526 1947
rect 31878 1750 31906 1778
rect 33166 2953 33194 2954
rect 33166 2927 33167 2953
rect 33167 2927 33193 2953
rect 33193 2927 33194 2953
rect 33166 2926 33194 2927
rect 32998 2870 33026 2898
rect 33390 2953 33418 2954
rect 33390 2927 33391 2953
rect 33391 2927 33417 2953
rect 33417 2927 33418 2953
rect 33390 2926 33418 2927
rect 33334 2505 33362 2506
rect 33334 2479 33335 2505
rect 33335 2479 33361 2505
rect 33361 2479 33362 2505
rect 33334 2478 33362 2479
rect 33894 6734 33922 6762
rect 33894 6481 33922 6482
rect 33894 6455 33895 6481
rect 33895 6455 33921 6481
rect 33921 6455 33922 6481
rect 33894 6454 33922 6455
rect 33782 4998 33810 5026
rect 33894 3737 33922 3738
rect 33894 3711 33895 3737
rect 33895 3711 33921 3737
rect 33921 3711 33922 3737
rect 33894 3710 33922 3711
rect 33726 2198 33754 2226
rect 33838 2478 33866 2506
rect 34582 8637 34610 8638
rect 34582 8611 34600 8637
rect 34600 8611 34610 8637
rect 34582 8610 34610 8611
rect 34634 8637 34662 8638
rect 34634 8611 34636 8637
rect 34636 8611 34662 8637
rect 34634 8610 34662 8611
rect 34686 8637 34714 8638
rect 34738 8637 34766 8638
rect 34686 8611 34698 8637
rect 34698 8611 34714 8637
rect 34738 8611 34760 8637
rect 34760 8611 34766 8637
rect 34686 8610 34714 8611
rect 34738 8610 34766 8611
rect 34790 8610 34818 8638
rect 34842 8637 34870 8638
rect 34894 8637 34922 8638
rect 34842 8611 34848 8637
rect 34848 8611 34870 8637
rect 34894 8611 34910 8637
rect 34910 8611 34922 8637
rect 34842 8610 34870 8611
rect 34894 8610 34922 8611
rect 34946 8637 34974 8638
rect 34946 8611 34972 8637
rect 34972 8611 34974 8637
rect 34946 8610 34974 8611
rect 34998 8637 35026 8638
rect 34998 8611 35008 8637
rect 35008 8611 35026 8637
rect 34998 8610 35026 8611
rect 34678 8049 34706 8050
rect 34678 8023 34679 8049
rect 34679 8023 34705 8049
rect 34705 8023 34706 8049
rect 34678 8022 34706 8023
rect 34582 7853 34610 7854
rect 34582 7827 34600 7853
rect 34600 7827 34610 7853
rect 34582 7826 34610 7827
rect 34634 7853 34662 7854
rect 34634 7827 34636 7853
rect 34636 7827 34662 7853
rect 34634 7826 34662 7827
rect 34686 7853 34714 7854
rect 34738 7853 34766 7854
rect 34686 7827 34698 7853
rect 34698 7827 34714 7853
rect 34738 7827 34760 7853
rect 34760 7827 34766 7853
rect 34686 7826 34714 7827
rect 34738 7826 34766 7827
rect 34790 7826 34818 7854
rect 34842 7853 34870 7854
rect 34894 7853 34922 7854
rect 34842 7827 34848 7853
rect 34848 7827 34870 7853
rect 34894 7827 34910 7853
rect 34910 7827 34922 7853
rect 34842 7826 34870 7827
rect 34894 7826 34922 7827
rect 34946 7853 34974 7854
rect 34946 7827 34972 7853
rect 34972 7827 34974 7853
rect 34946 7826 34974 7827
rect 34998 7853 35026 7854
rect 34998 7827 35008 7853
rect 35008 7827 35026 7853
rect 34998 7826 35026 7827
rect 36190 9142 36218 9170
rect 35854 8777 35882 8778
rect 35854 8751 35855 8777
rect 35855 8751 35881 8777
rect 35881 8751 35882 8777
rect 35854 8750 35882 8751
rect 35238 7657 35266 7658
rect 35238 7631 35239 7657
rect 35239 7631 35265 7657
rect 35265 7631 35266 7657
rect 35238 7630 35266 7631
rect 35798 7630 35826 7658
rect 34398 7238 34426 7266
rect 34958 7265 34986 7266
rect 34958 7239 34959 7265
rect 34959 7239 34985 7265
rect 34985 7239 34986 7265
rect 34958 7238 34986 7239
rect 34582 7069 34610 7070
rect 34582 7043 34600 7069
rect 34600 7043 34610 7069
rect 34582 7042 34610 7043
rect 34634 7069 34662 7070
rect 34634 7043 34636 7069
rect 34636 7043 34662 7069
rect 34634 7042 34662 7043
rect 34686 7069 34714 7070
rect 34738 7069 34766 7070
rect 34686 7043 34698 7069
rect 34698 7043 34714 7069
rect 34738 7043 34760 7069
rect 34760 7043 34766 7069
rect 34686 7042 34714 7043
rect 34738 7042 34766 7043
rect 34790 7042 34818 7070
rect 34842 7069 34870 7070
rect 34894 7069 34922 7070
rect 34842 7043 34848 7069
rect 34848 7043 34870 7069
rect 34894 7043 34910 7069
rect 34910 7043 34922 7069
rect 34842 7042 34870 7043
rect 34894 7042 34922 7043
rect 34946 7069 34974 7070
rect 34946 7043 34972 7069
rect 34972 7043 34974 7069
rect 34946 7042 34974 7043
rect 34998 7069 35026 7070
rect 34998 7043 35008 7069
rect 35008 7043 35026 7069
rect 34998 7042 35026 7043
rect 35350 7518 35378 7546
rect 35518 7518 35546 7546
rect 35182 6902 35210 6930
rect 35294 6873 35322 6874
rect 35294 6847 35295 6873
rect 35295 6847 35321 6873
rect 35321 6847 35322 6873
rect 35294 6846 35322 6847
rect 34398 6678 34426 6706
rect 35854 7518 35882 7546
rect 36134 8049 36162 8050
rect 36134 8023 36135 8049
rect 36135 8023 36161 8049
rect 36161 8023 36162 8049
rect 36134 8022 36162 8023
rect 36134 7630 36162 7658
rect 37082 18437 37110 18438
rect 37082 18411 37100 18437
rect 37100 18411 37110 18437
rect 37082 18410 37110 18411
rect 37134 18437 37162 18438
rect 37134 18411 37136 18437
rect 37136 18411 37162 18437
rect 37134 18410 37162 18411
rect 37186 18437 37214 18438
rect 37238 18437 37266 18438
rect 37186 18411 37198 18437
rect 37198 18411 37214 18437
rect 37238 18411 37260 18437
rect 37260 18411 37266 18437
rect 37186 18410 37214 18411
rect 37238 18410 37266 18411
rect 37290 18410 37318 18438
rect 37342 18437 37370 18438
rect 37394 18437 37422 18438
rect 37342 18411 37348 18437
rect 37348 18411 37370 18437
rect 37394 18411 37410 18437
rect 37410 18411 37422 18437
rect 37342 18410 37370 18411
rect 37394 18410 37422 18411
rect 37446 18437 37474 18438
rect 37446 18411 37472 18437
rect 37472 18411 37474 18437
rect 37446 18410 37474 18411
rect 37498 18437 37526 18438
rect 37498 18411 37508 18437
rect 37508 18411 37526 18437
rect 37498 18410 37526 18411
rect 37082 17653 37110 17654
rect 37082 17627 37100 17653
rect 37100 17627 37110 17653
rect 37082 17626 37110 17627
rect 37134 17653 37162 17654
rect 37134 17627 37136 17653
rect 37136 17627 37162 17653
rect 37134 17626 37162 17627
rect 37186 17653 37214 17654
rect 37238 17653 37266 17654
rect 37186 17627 37198 17653
rect 37198 17627 37214 17653
rect 37238 17627 37260 17653
rect 37260 17627 37266 17653
rect 37186 17626 37214 17627
rect 37238 17626 37266 17627
rect 37290 17626 37318 17654
rect 37342 17653 37370 17654
rect 37394 17653 37422 17654
rect 37342 17627 37348 17653
rect 37348 17627 37370 17653
rect 37394 17627 37410 17653
rect 37410 17627 37422 17653
rect 37342 17626 37370 17627
rect 37394 17626 37422 17627
rect 37446 17653 37474 17654
rect 37446 17627 37472 17653
rect 37472 17627 37474 17653
rect 37446 17626 37474 17627
rect 37498 17653 37526 17654
rect 37498 17627 37508 17653
rect 37508 17627 37526 17653
rect 37498 17626 37526 17627
rect 37082 16869 37110 16870
rect 37082 16843 37100 16869
rect 37100 16843 37110 16869
rect 37082 16842 37110 16843
rect 37134 16869 37162 16870
rect 37134 16843 37136 16869
rect 37136 16843 37162 16869
rect 37134 16842 37162 16843
rect 37186 16869 37214 16870
rect 37238 16869 37266 16870
rect 37186 16843 37198 16869
rect 37198 16843 37214 16869
rect 37238 16843 37260 16869
rect 37260 16843 37266 16869
rect 37186 16842 37214 16843
rect 37238 16842 37266 16843
rect 37290 16842 37318 16870
rect 37342 16869 37370 16870
rect 37394 16869 37422 16870
rect 37342 16843 37348 16869
rect 37348 16843 37370 16869
rect 37394 16843 37410 16869
rect 37410 16843 37422 16869
rect 37342 16842 37370 16843
rect 37394 16842 37422 16843
rect 37446 16869 37474 16870
rect 37446 16843 37472 16869
rect 37472 16843 37474 16869
rect 37446 16842 37474 16843
rect 37498 16869 37526 16870
rect 37498 16843 37508 16869
rect 37508 16843 37526 16869
rect 37498 16842 37526 16843
rect 37082 16085 37110 16086
rect 37082 16059 37100 16085
rect 37100 16059 37110 16085
rect 37082 16058 37110 16059
rect 37134 16085 37162 16086
rect 37134 16059 37136 16085
rect 37136 16059 37162 16085
rect 37134 16058 37162 16059
rect 37186 16085 37214 16086
rect 37238 16085 37266 16086
rect 37186 16059 37198 16085
rect 37198 16059 37214 16085
rect 37238 16059 37260 16085
rect 37260 16059 37266 16085
rect 37186 16058 37214 16059
rect 37238 16058 37266 16059
rect 37290 16058 37318 16086
rect 37342 16085 37370 16086
rect 37394 16085 37422 16086
rect 37342 16059 37348 16085
rect 37348 16059 37370 16085
rect 37394 16059 37410 16085
rect 37410 16059 37422 16085
rect 37342 16058 37370 16059
rect 37394 16058 37422 16059
rect 37446 16085 37474 16086
rect 37446 16059 37472 16085
rect 37472 16059 37474 16085
rect 37446 16058 37474 16059
rect 37498 16085 37526 16086
rect 37498 16059 37508 16085
rect 37508 16059 37526 16085
rect 37498 16058 37526 16059
rect 37082 15301 37110 15302
rect 37082 15275 37100 15301
rect 37100 15275 37110 15301
rect 37082 15274 37110 15275
rect 37134 15301 37162 15302
rect 37134 15275 37136 15301
rect 37136 15275 37162 15301
rect 37134 15274 37162 15275
rect 37186 15301 37214 15302
rect 37238 15301 37266 15302
rect 37186 15275 37198 15301
rect 37198 15275 37214 15301
rect 37238 15275 37260 15301
rect 37260 15275 37266 15301
rect 37186 15274 37214 15275
rect 37238 15274 37266 15275
rect 37290 15274 37318 15302
rect 37342 15301 37370 15302
rect 37394 15301 37422 15302
rect 37342 15275 37348 15301
rect 37348 15275 37370 15301
rect 37394 15275 37410 15301
rect 37410 15275 37422 15301
rect 37342 15274 37370 15275
rect 37394 15274 37422 15275
rect 37446 15301 37474 15302
rect 37446 15275 37472 15301
rect 37472 15275 37474 15301
rect 37446 15274 37474 15275
rect 37498 15301 37526 15302
rect 37498 15275 37508 15301
rect 37508 15275 37526 15301
rect 37498 15274 37526 15275
rect 37082 14517 37110 14518
rect 37082 14491 37100 14517
rect 37100 14491 37110 14517
rect 37082 14490 37110 14491
rect 37134 14517 37162 14518
rect 37134 14491 37136 14517
rect 37136 14491 37162 14517
rect 37134 14490 37162 14491
rect 37186 14517 37214 14518
rect 37238 14517 37266 14518
rect 37186 14491 37198 14517
rect 37198 14491 37214 14517
rect 37238 14491 37260 14517
rect 37260 14491 37266 14517
rect 37186 14490 37214 14491
rect 37238 14490 37266 14491
rect 37290 14490 37318 14518
rect 37342 14517 37370 14518
rect 37394 14517 37422 14518
rect 37342 14491 37348 14517
rect 37348 14491 37370 14517
rect 37394 14491 37410 14517
rect 37410 14491 37422 14517
rect 37342 14490 37370 14491
rect 37394 14490 37422 14491
rect 37446 14517 37474 14518
rect 37446 14491 37472 14517
rect 37472 14491 37474 14517
rect 37446 14490 37474 14491
rect 37498 14517 37526 14518
rect 37498 14491 37508 14517
rect 37508 14491 37526 14517
rect 37498 14490 37526 14491
rect 37082 13733 37110 13734
rect 37082 13707 37100 13733
rect 37100 13707 37110 13733
rect 37082 13706 37110 13707
rect 37134 13733 37162 13734
rect 37134 13707 37136 13733
rect 37136 13707 37162 13733
rect 37134 13706 37162 13707
rect 37186 13733 37214 13734
rect 37238 13733 37266 13734
rect 37186 13707 37198 13733
rect 37198 13707 37214 13733
rect 37238 13707 37260 13733
rect 37260 13707 37266 13733
rect 37186 13706 37214 13707
rect 37238 13706 37266 13707
rect 37290 13706 37318 13734
rect 37342 13733 37370 13734
rect 37394 13733 37422 13734
rect 37342 13707 37348 13733
rect 37348 13707 37370 13733
rect 37394 13707 37410 13733
rect 37410 13707 37422 13733
rect 37342 13706 37370 13707
rect 37394 13706 37422 13707
rect 37446 13733 37474 13734
rect 37446 13707 37472 13733
rect 37472 13707 37474 13733
rect 37446 13706 37474 13707
rect 37498 13733 37526 13734
rect 37498 13707 37508 13733
rect 37508 13707 37526 13733
rect 37498 13706 37526 13707
rect 37082 12949 37110 12950
rect 37082 12923 37100 12949
rect 37100 12923 37110 12949
rect 37082 12922 37110 12923
rect 37134 12949 37162 12950
rect 37134 12923 37136 12949
rect 37136 12923 37162 12949
rect 37134 12922 37162 12923
rect 37186 12949 37214 12950
rect 37238 12949 37266 12950
rect 37186 12923 37198 12949
rect 37198 12923 37214 12949
rect 37238 12923 37260 12949
rect 37260 12923 37266 12949
rect 37186 12922 37214 12923
rect 37238 12922 37266 12923
rect 37290 12922 37318 12950
rect 37342 12949 37370 12950
rect 37394 12949 37422 12950
rect 37342 12923 37348 12949
rect 37348 12923 37370 12949
rect 37394 12923 37410 12949
rect 37410 12923 37422 12949
rect 37342 12922 37370 12923
rect 37394 12922 37422 12923
rect 37446 12949 37474 12950
rect 37446 12923 37472 12949
rect 37472 12923 37474 12949
rect 37446 12922 37474 12923
rect 37498 12949 37526 12950
rect 37498 12923 37508 12949
rect 37508 12923 37526 12949
rect 37498 12922 37526 12923
rect 37082 12165 37110 12166
rect 37082 12139 37100 12165
rect 37100 12139 37110 12165
rect 37082 12138 37110 12139
rect 37134 12165 37162 12166
rect 37134 12139 37136 12165
rect 37136 12139 37162 12165
rect 37134 12138 37162 12139
rect 37186 12165 37214 12166
rect 37238 12165 37266 12166
rect 37186 12139 37198 12165
rect 37198 12139 37214 12165
rect 37238 12139 37260 12165
rect 37260 12139 37266 12165
rect 37186 12138 37214 12139
rect 37238 12138 37266 12139
rect 37290 12138 37318 12166
rect 37342 12165 37370 12166
rect 37394 12165 37422 12166
rect 37342 12139 37348 12165
rect 37348 12139 37370 12165
rect 37394 12139 37410 12165
rect 37410 12139 37422 12165
rect 37342 12138 37370 12139
rect 37394 12138 37422 12139
rect 37446 12165 37474 12166
rect 37446 12139 37472 12165
rect 37472 12139 37474 12165
rect 37446 12138 37474 12139
rect 37498 12165 37526 12166
rect 37498 12139 37508 12165
rect 37508 12139 37526 12165
rect 37498 12138 37526 12139
rect 37082 11381 37110 11382
rect 37082 11355 37100 11381
rect 37100 11355 37110 11381
rect 37082 11354 37110 11355
rect 37134 11381 37162 11382
rect 37134 11355 37136 11381
rect 37136 11355 37162 11381
rect 37134 11354 37162 11355
rect 37186 11381 37214 11382
rect 37238 11381 37266 11382
rect 37186 11355 37198 11381
rect 37198 11355 37214 11381
rect 37238 11355 37260 11381
rect 37260 11355 37266 11381
rect 37186 11354 37214 11355
rect 37238 11354 37266 11355
rect 37290 11354 37318 11382
rect 37342 11381 37370 11382
rect 37394 11381 37422 11382
rect 37342 11355 37348 11381
rect 37348 11355 37370 11381
rect 37394 11355 37410 11381
rect 37410 11355 37422 11381
rect 37342 11354 37370 11355
rect 37394 11354 37422 11355
rect 37446 11381 37474 11382
rect 37446 11355 37472 11381
rect 37472 11355 37474 11381
rect 37446 11354 37474 11355
rect 37498 11381 37526 11382
rect 37498 11355 37508 11381
rect 37508 11355 37526 11381
rect 37498 11354 37526 11355
rect 37082 10597 37110 10598
rect 37082 10571 37100 10597
rect 37100 10571 37110 10597
rect 37082 10570 37110 10571
rect 37134 10597 37162 10598
rect 37134 10571 37136 10597
rect 37136 10571 37162 10597
rect 37134 10570 37162 10571
rect 37186 10597 37214 10598
rect 37238 10597 37266 10598
rect 37186 10571 37198 10597
rect 37198 10571 37214 10597
rect 37238 10571 37260 10597
rect 37260 10571 37266 10597
rect 37186 10570 37214 10571
rect 37238 10570 37266 10571
rect 37290 10570 37318 10598
rect 37342 10597 37370 10598
rect 37394 10597 37422 10598
rect 37342 10571 37348 10597
rect 37348 10571 37370 10597
rect 37394 10571 37410 10597
rect 37410 10571 37422 10597
rect 37342 10570 37370 10571
rect 37394 10570 37422 10571
rect 37446 10597 37474 10598
rect 37446 10571 37472 10597
rect 37472 10571 37474 10597
rect 37446 10570 37474 10571
rect 37498 10597 37526 10598
rect 37498 10571 37508 10597
rect 37508 10571 37526 10597
rect 37498 10570 37526 10571
rect 37310 10345 37338 10346
rect 37310 10319 37311 10345
rect 37311 10319 37337 10345
rect 37337 10319 37338 10345
rect 37310 10318 37338 10319
rect 37590 10318 37618 10346
rect 37082 9813 37110 9814
rect 37082 9787 37100 9813
rect 37100 9787 37110 9813
rect 37082 9786 37110 9787
rect 37134 9813 37162 9814
rect 37134 9787 37136 9813
rect 37136 9787 37162 9813
rect 37134 9786 37162 9787
rect 37186 9813 37214 9814
rect 37238 9813 37266 9814
rect 37186 9787 37198 9813
rect 37198 9787 37214 9813
rect 37238 9787 37260 9813
rect 37260 9787 37266 9813
rect 37186 9786 37214 9787
rect 37238 9786 37266 9787
rect 37290 9786 37318 9814
rect 37342 9813 37370 9814
rect 37394 9813 37422 9814
rect 37342 9787 37348 9813
rect 37348 9787 37370 9813
rect 37394 9787 37410 9813
rect 37410 9787 37422 9813
rect 37342 9786 37370 9787
rect 37394 9786 37422 9787
rect 37446 9813 37474 9814
rect 37446 9787 37472 9813
rect 37472 9787 37474 9813
rect 37446 9786 37474 9787
rect 37498 9813 37526 9814
rect 37498 9787 37508 9813
rect 37508 9787 37526 9813
rect 37498 9786 37526 9787
rect 37310 9561 37338 9562
rect 37310 9535 37311 9561
rect 37311 9535 37337 9561
rect 37337 9535 37338 9561
rect 37310 9534 37338 9535
rect 37082 9029 37110 9030
rect 37082 9003 37100 9029
rect 37100 9003 37110 9029
rect 37082 9002 37110 9003
rect 37134 9029 37162 9030
rect 37134 9003 37136 9029
rect 37136 9003 37162 9029
rect 37134 9002 37162 9003
rect 37186 9029 37214 9030
rect 37238 9029 37266 9030
rect 37186 9003 37198 9029
rect 37198 9003 37214 9029
rect 37238 9003 37260 9029
rect 37260 9003 37266 9029
rect 37186 9002 37214 9003
rect 37238 9002 37266 9003
rect 37290 9002 37318 9030
rect 37342 9029 37370 9030
rect 37394 9029 37422 9030
rect 37342 9003 37348 9029
rect 37348 9003 37370 9029
rect 37394 9003 37410 9029
rect 37410 9003 37422 9029
rect 37342 9002 37370 9003
rect 37394 9002 37422 9003
rect 37446 9029 37474 9030
rect 37446 9003 37472 9029
rect 37472 9003 37474 9029
rect 37446 9002 37474 9003
rect 37498 9029 37526 9030
rect 37498 9003 37508 9029
rect 37508 9003 37526 9029
rect 37498 9002 37526 9003
rect 36974 8750 37002 8778
rect 37646 9534 37674 9562
rect 37082 8245 37110 8246
rect 37082 8219 37100 8245
rect 37100 8219 37110 8245
rect 37082 8218 37110 8219
rect 37134 8245 37162 8246
rect 37134 8219 37136 8245
rect 37136 8219 37162 8245
rect 37134 8218 37162 8219
rect 37186 8245 37214 8246
rect 37238 8245 37266 8246
rect 37186 8219 37198 8245
rect 37198 8219 37214 8245
rect 37238 8219 37260 8245
rect 37260 8219 37266 8245
rect 37186 8218 37214 8219
rect 37238 8218 37266 8219
rect 37290 8218 37318 8246
rect 37342 8245 37370 8246
rect 37394 8245 37422 8246
rect 37342 8219 37348 8245
rect 37348 8219 37370 8245
rect 37394 8219 37410 8245
rect 37410 8219 37422 8245
rect 37342 8218 37370 8219
rect 37394 8218 37422 8219
rect 37446 8245 37474 8246
rect 37446 8219 37472 8245
rect 37472 8219 37474 8245
rect 37446 8218 37474 8219
rect 37498 8245 37526 8246
rect 37498 8219 37508 8245
rect 37508 8219 37526 8245
rect 37498 8218 37526 8219
rect 36694 7657 36722 7658
rect 36694 7631 36695 7657
rect 36695 7631 36721 7657
rect 36721 7631 36722 7657
rect 36694 7630 36722 7631
rect 35854 7182 35882 7210
rect 35350 6734 35378 6762
rect 35630 6846 35658 6874
rect 34582 6285 34610 6286
rect 34582 6259 34600 6285
rect 34600 6259 34610 6285
rect 34582 6258 34610 6259
rect 34634 6285 34662 6286
rect 34634 6259 34636 6285
rect 34636 6259 34662 6285
rect 34634 6258 34662 6259
rect 34686 6285 34714 6286
rect 34738 6285 34766 6286
rect 34686 6259 34698 6285
rect 34698 6259 34714 6285
rect 34738 6259 34760 6285
rect 34760 6259 34766 6285
rect 34686 6258 34714 6259
rect 34738 6258 34766 6259
rect 34790 6258 34818 6286
rect 34842 6285 34870 6286
rect 34894 6285 34922 6286
rect 34842 6259 34848 6285
rect 34848 6259 34870 6285
rect 34894 6259 34910 6285
rect 34910 6259 34922 6285
rect 34842 6258 34870 6259
rect 34894 6258 34922 6259
rect 34946 6285 34974 6286
rect 34946 6259 34972 6285
rect 34972 6259 34974 6285
rect 34946 6258 34974 6259
rect 34998 6285 35026 6286
rect 34998 6259 35008 6285
rect 35008 6259 35026 6285
rect 34998 6258 35026 6259
rect 35574 5894 35602 5922
rect 34174 5305 34202 5306
rect 34174 5279 34175 5305
rect 34175 5279 34201 5305
rect 34201 5279 34202 5305
rect 34174 5278 34202 5279
rect 34582 5501 34610 5502
rect 34582 5475 34600 5501
rect 34600 5475 34610 5501
rect 34582 5474 34610 5475
rect 34634 5501 34662 5502
rect 34634 5475 34636 5501
rect 34636 5475 34662 5501
rect 34634 5474 34662 5475
rect 34686 5501 34714 5502
rect 34738 5501 34766 5502
rect 34686 5475 34698 5501
rect 34698 5475 34714 5501
rect 34738 5475 34760 5501
rect 34760 5475 34766 5501
rect 34686 5474 34714 5475
rect 34738 5474 34766 5475
rect 34790 5474 34818 5502
rect 34842 5501 34870 5502
rect 34894 5501 34922 5502
rect 34842 5475 34848 5501
rect 34848 5475 34870 5501
rect 34894 5475 34910 5501
rect 34910 5475 34922 5501
rect 34842 5474 34870 5475
rect 34894 5474 34922 5475
rect 34946 5501 34974 5502
rect 34946 5475 34972 5501
rect 34972 5475 34974 5501
rect 34946 5474 34974 5475
rect 34998 5501 35026 5502
rect 34998 5475 35008 5501
rect 35008 5475 35026 5501
rect 34998 5474 35026 5475
rect 34622 5222 34650 5250
rect 34846 5222 34874 5250
rect 34582 4717 34610 4718
rect 34582 4691 34600 4717
rect 34600 4691 34610 4717
rect 34582 4690 34610 4691
rect 34634 4717 34662 4718
rect 34634 4691 34636 4717
rect 34636 4691 34662 4717
rect 34634 4690 34662 4691
rect 34686 4717 34714 4718
rect 34738 4717 34766 4718
rect 34686 4691 34698 4717
rect 34698 4691 34714 4717
rect 34738 4691 34760 4717
rect 34760 4691 34766 4717
rect 34686 4690 34714 4691
rect 34738 4690 34766 4691
rect 34790 4690 34818 4718
rect 34842 4717 34870 4718
rect 34894 4717 34922 4718
rect 34842 4691 34848 4717
rect 34848 4691 34870 4717
rect 34894 4691 34910 4717
rect 34910 4691 34922 4717
rect 34842 4690 34870 4691
rect 34894 4690 34922 4691
rect 34946 4717 34974 4718
rect 34946 4691 34972 4717
rect 34972 4691 34974 4717
rect 34946 4690 34974 4691
rect 34998 4717 35026 4718
rect 34998 4691 35008 4717
rect 35008 4691 35026 4717
rect 34998 4690 35026 4691
rect 34174 3318 34202 3346
rect 34174 2982 34202 3010
rect 34454 3710 34482 3738
rect 33950 2422 33978 2450
rect 34230 2870 34258 2898
rect 33670 2142 33698 2170
rect 34118 2086 34146 2114
rect 33446 1777 33474 1778
rect 33446 1751 33447 1777
rect 33447 1751 33473 1777
rect 33473 1751 33474 1777
rect 33446 1750 33474 1751
rect 34582 3933 34610 3934
rect 34582 3907 34600 3933
rect 34600 3907 34610 3933
rect 34582 3906 34610 3907
rect 34634 3933 34662 3934
rect 34634 3907 34636 3933
rect 34636 3907 34662 3933
rect 34634 3906 34662 3907
rect 34686 3933 34714 3934
rect 34738 3933 34766 3934
rect 34686 3907 34698 3933
rect 34698 3907 34714 3933
rect 34738 3907 34760 3933
rect 34760 3907 34766 3933
rect 34686 3906 34714 3907
rect 34738 3906 34766 3907
rect 34790 3906 34818 3934
rect 34842 3933 34870 3934
rect 34894 3933 34922 3934
rect 34842 3907 34848 3933
rect 34848 3907 34870 3933
rect 34894 3907 34910 3933
rect 34910 3907 34922 3933
rect 34842 3906 34870 3907
rect 34894 3906 34922 3907
rect 34946 3933 34974 3934
rect 34946 3907 34972 3933
rect 34972 3907 34974 3933
rect 34946 3906 34974 3907
rect 34998 3933 35026 3934
rect 34998 3907 35008 3933
rect 35008 3907 35026 3933
rect 34998 3906 35026 3907
rect 37082 7461 37110 7462
rect 37082 7435 37100 7461
rect 37100 7435 37110 7461
rect 37082 7434 37110 7435
rect 37134 7461 37162 7462
rect 37134 7435 37136 7461
rect 37136 7435 37162 7461
rect 37134 7434 37162 7435
rect 37186 7461 37214 7462
rect 37238 7461 37266 7462
rect 37186 7435 37198 7461
rect 37198 7435 37214 7461
rect 37238 7435 37260 7461
rect 37260 7435 37266 7461
rect 37186 7434 37214 7435
rect 37238 7434 37266 7435
rect 37290 7434 37318 7462
rect 37342 7461 37370 7462
rect 37394 7461 37422 7462
rect 37342 7435 37348 7461
rect 37348 7435 37370 7461
rect 37394 7435 37410 7461
rect 37410 7435 37422 7461
rect 37342 7434 37370 7435
rect 37394 7434 37422 7435
rect 37446 7461 37474 7462
rect 37446 7435 37472 7461
rect 37472 7435 37474 7461
rect 37446 7434 37474 7435
rect 37498 7461 37526 7462
rect 37498 7435 37508 7461
rect 37508 7435 37526 7461
rect 37498 7434 37526 7435
rect 36750 7238 36778 7266
rect 35798 6454 35826 6482
rect 35686 5726 35714 5754
rect 35630 5054 35658 5082
rect 35742 4998 35770 5026
rect 35574 4886 35602 4914
rect 35350 3737 35378 3738
rect 35350 3711 35351 3737
rect 35351 3711 35377 3737
rect 35377 3711 35378 3737
rect 35350 3710 35378 3711
rect 34510 3318 34538 3346
rect 34678 3345 34706 3346
rect 34678 3319 34679 3345
rect 34679 3319 34705 3345
rect 34705 3319 34706 3345
rect 34678 3318 34706 3319
rect 34582 3149 34610 3150
rect 34582 3123 34600 3149
rect 34600 3123 34610 3149
rect 34582 3122 34610 3123
rect 34634 3149 34662 3150
rect 34634 3123 34636 3149
rect 34636 3123 34662 3149
rect 34634 3122 34662 3123
rect 34686 3149 34714 3150
rect 34738 3149 34766 3150
rect 34686 3123 34698 3149
rect 34698 3123 34714 3149
rect 34738 3123 34760 3149
rect 34760 3123 34766 3149
rect 34686 3122 34714 3123
rect 34738 3122 34766 3123
rect 34790 3122 34818 3150
rect 34842 3149 34870 3150
rect 34894 3149 34922 3150
rect 34842 3123 34848 3149
rect 34848 3123 34870 3149
rect 34894 3123 34910 3149
rect 34910 3123 34922 3149
rect 34842 3122 34870 3123
rect 34894 3122 34922 3123
rect 34946 3149 34974 3150
rect 34946 3123 34972 3149
rect 34972 3123 34974 3149
rect 34946 3122 34974 3123
rect 34998 3149 35026 3150
rect 34998 3123 35008 3149
rect 35008 3123 35026 3149
rect 34998 3122 35026 3123
rect 34678 2982 34706 3010
rect 35630 4158 35658 4186
rect 35630 3710 35658 3738
rect 35686 3262 35714 3290
rect 35854 4158 35882 4186
rect 36134 3345 36162 3346
rect 36134 3319 36135 3345
rect 36135 3319 36161 3345
rect 36161 3319 36162 3345
rect 36134 3318 36162 3319
rect 36694 3318 36722 3346
rect 37310 7209 37338 7210
rect 37310 7183 37311 7209
rect 37311 7183 37337 7209
rect 37337 7183 37338 7209
rect 37310 7182 37338 7183
rect 37646 7182 37674 7210
rect 37082 6677 37110 6678
rect 37082 6651 37100 6677
rect 37100 6651 37110 6677
rect 37082 6650 37110 6651
rect 37134 6677 37162 6678
rect 37134 6651 37136 6677
rect 37136 6651 37162 6677
rect 37134 6650 37162 6651
rect 37186 6677 37214 6678
rect 37238 6677 37266 6678
rect 37186 6651 37198 6677
rect 37198 6651 37214 6677
rect 37238 6651 37260 6677
rect 37260 6651 37266 6677
rect 37186 6650 37214 6651
rect 37238 6650 37266 6651
rect 37290 6650 37318 6678
rect 37342 6677 37370 6678
rect 37394 6677 37422 6678
rect 37342 6651 37348 6677
rect 37348 6651 37370 6677
rect 37394 6651 37410 6677
rect 37410 6651 37422 6677
rect 37342 6650 37370 6651
rect 37394 6650 37422 6651
rect 37446 6677 37474 6678
rect 37446 6651 37472 6677
rect 37472 6651 37474 6677
rect 37446 6650 37474 6651
rect 37498 6677 37526 6678
rect 37498 6651 37508 6677
rect 37508 6651 37526 6677
rect 37498 6650 37526 6651
rect 37366 6089 37394 6090
rect 37366 6063 37367 6089
rect 37367 6063 37393 6089
rect 37393 6063 37394 6089
rect 37366 6062 37394 6063
rect 37646 6062 37674 6090
rect 37082 5893 37110 5894
rect 37082 5867 37100 5893
rect 37100 5867 37110 5893
rect 37082 5866 37110 5867
rect 37134 5893 37162 5894
rect 37134 5867 37136 5893
rect 37136 5867 37162 5893
rect 37134 5866 37162 5867
rect 37186 5893 37214 5894
rect 37238 5893 37266 5894
rect 37186 5867 37198 5893
rect 37198 5867 37214 5893
rect 37238 5867 37260 5893
rect 37260 5867 37266 5893
rect 37186 5866 37214 5867
rect 37238 5866 37266 5867
rect 37290 5866 37318 5894
rect 37342 5893 37370 5894
rect 37394 5893 37422 5894
rect 37342 5867 37348 5893
rect 37348 5867 37370 5893
rect 37394 5867 37410 5893
rect 37410 5867 37422 5893
rect 37342 5866 37370 5867
rect 37394 5866 37422 5867
rect 37446 5893 37474 5894
rect 37446 5867 37472 5893
rect 37472 5867 37474 5893
rect 37446 5866 37474 5867
rect 37498 5893 37526 5894
rect 37498 5867 37508 5893
rect 37508 5867 37526 5893
rect 37498 5866 37526 5867
rect 37590 5641 37618 5642
rect 37590 5615 37591 5641
rect 37591 5615 37617 5641
rect 37617 5615 37618 5641
rect 37590 5614 37618 5615
rect 37082 5109 37110 5110
rect 37082 5083 37100 5109
rect 37100 5083 37110 5109
rect 37082 5082 37110 5083
rect 37134 5109 37162 5110
rect 37134 5083 37136 5109
rect 37136 5083 37162 5109
rect 37134 5082 37162 5083
rect 37186 5109 37214 5110
rect 37238 5109 37266 5110
rect 37186 5083 37198 5109
rect 37198 5083 37214 5109
rect 37238 5083 37260 5109
rect 37260 5083 37266 5109
rect 37186 5082 37214 5083
rect 37238 5082 37266 5083
rect 37290 5082 37318 5110
rect 37342 5109 37370 5110
rect 37394 5109 37422 5110
rect 37342 5083 37348 5109
rect 37348 5083 37370 5109
rect 37394 5083 37410 5109
rect 37410 5083 37422 5109
rect 37342 5082 37370 5083
rect 37394 5082 37422 5083
rect 37446 5109 37474 5110
rect 37446 5083 37472 5109
rect 37472 5083 37474 5109
rect 37446 5082 37474 5083
rect 37498 5109 37526 5110
rect 37498 5083 37508 5109
rect 37508 5083 37526 5109
rect 37498 5082 37526 5083
rect 37590 4857 37618 4858
rect 37590 4831 37591 4857
rect 37591 4831 37617 4857
rect 37617 4831 37618 4857
rect 37590 4830 37618 4831
rect 37082 4325 37110 4326
rect 37082 4299 37100 4325
rect 37100 4299 37110 4325
rect 37082 4298 37110 4299
rect 37134 4325 37162 4326
rect 37134 4299 37136 4325
rect 37136 4299 37162 4325
rect 37134 4298 37162 4299
rect 37186 4325 37214 4326
rect 37238 4325 37266 4326
rect 37186 4299 37198 4325
rect 37198 4299 37214 4325
rect 37238 4299 37260 4325
rect 37260 4299 37266 4325
rect 37186 4298 37214 4299
rect 37238 4298 37266 4299
rect 37290 4298 37318 4326
rect 37342 4325 37370 4326
rect 37394 4325 37422 4326
rect 37342 4299 37348 4325
rect 37348 4299 37370 4325
rect 37394 4299 37410 4325
rect 37410 4299 37422 4325
rect 37342 4298 37370 4299
rect 37394 4298 37422 4299
rect 37446 4325 37474 4326
rect 37446 4299 37472 4325
rect 37472 4299 37474 4325
rect 37446 4298 37474 4299
rect 37498 4325 37526 4326
rect 37498 4299 37508 4325
rect 37508 4299 37526 4325
rect 37498 4298 37526 4299
rect 37086 4129 37114 4130
rect 37086 4103 37087 4129
rect 37087 4103 37113 4129
rect 37113 4103 37114 4129
rect 37086 4102 37114 4103
rect 37590 3710 37618 3738
rect 37082 3541 37110 3542
rect 37082 3515 37100 3541
rect 37100 3515 37110 3541
rect 37082 3514 37110 3515
rect 37134 3541 37162 3542
rect 37134 3515 37136 3541
rect 37136 3515 37162 3541
rect 37134 3514 37162 3515
rect 37186 3541 37214 3542
rect 37238 3541 37266 3542
rect 37186 3515 37198 3541
rect 37198 3515 37214 3541
rect 37238 3515 37260 3541
rect 37260 3515 37266 3541
rect 37186 3514 37214 3515
rect 37238 3514 37266 3515
rect 37290 3514 37318 3542
rect 37342 3541 37370 3542
rect 37394 3541 37422 3542
rect 37342 3515 37348 3541
rect 37348 3515 37370 3541
rect 37394 3515 37410 3541
rect 37410 3515 37422 3541
rect 37342 3514 37370 3515
rect 37394 3514 37422 3515
rect 37446 3541 37474 3542
rect 37446 3515 37472 3541
rect 37472 3515 37474 3541
rect 37446 3514 37474 3515
rect 37498 3541 37526 3542
rect 37498 3515 37508 3541
rect 37508 3515 37526 3541
rect 37498 3514 37526 3515
rect 37142 3374 37170 3402
rect 37310 3038 37338 3066
rect 35910 2870 35938 2898
rect 35854 2505 35882 2506
rect 35854 2479 35855 2505
rect 35855 2479 35881 2505
rect 35881 2479 35882 2505
rect 35854 2478 35882 2479
rect 34582 2365 34610 2366
rect 34582 2339 34600 2365
rect 34600 2339 34610 2365
rect 34582 2338 34610 2339
rect 34634 2365 34662 2366
rect 34634 2339 34636 2365
rect 34636 2339 34662 2365
rect 34634 2338 34662 2339
rect 34686 2365 34714 2366
rect 34738 2365 34766 2366
rect 34686 2339 34698 2365
rect 34698 2339 34714 2365
rect 34738 2339 34760 2365
rect 34760 2339 34766 2365
rect 34686 2338 34714 2339
rect 34738 2338 34766 2339
rect 34790 2338 34818 2366
rect 34842 2365 34870 2366
rect 34894 2365 34922 2366
rect 34842 2339 34848 2365
rect 34848 2339 34870 2365
rect 34894 2339 34910 2365
rect 34910 2339 34922 2365
rect 34842 2338 34870 2339
rect 34894 2338 34922 2339
rect 34946 2365 34974 2366
rect 34946 2339 34972 2365
rect 34972 2339 34974 2365
rect 34946 2338 34974 2339
rect 34998 2365 35026 2366
rect 34998 2339 35008 2365
rect 35008 2339 35026 2365
rect 34998 2338 35026 2339
rect 37082 2757 37110 2758
rect 37082 2731 37100 2757
rect 37100 2731 37110 2757
rect 37082 2730 37110 2731
rect 37134 2757 37162 2758
rect 37134 2731 37136 2757
rect 37136 2731 37162 2757
rect 37134 2730 37162 2731
rect 37186 2757 37214 2758
rect 37238 2757 37266 2758
rect 37186 2731 37198 2757
rect 37198 2731 37214 2757
rect 37238 2731 37260 2757
rect 37260 2731 37266 2757
rect 37186 2730 37214 2731
rect 37238 2730 37266 2731
rect 37290 2730 37318 2758
rect 37342 2757 37370 2758
rect 37394 2757 37422 2758
rect 37342 2731 37348 2757
rect 37348 2731 37370 2757
rect 37394 2731 37410 2757
rect 37410 2731 37422 2757
rect 37342 2730 37370 2731
rect 37394 2730 37422 2731
rect 37446 2757 37474 2758
rect 37446 2731 37472 2757
rect 37472 2731 37474 2757
rect 37446 2730 37474 2731
rect 37498 2757 37526 2758
rect 37498 2731 37508 2757
rect 37508 2731 37526 2757
rect 37498 2730 37526 2731
rect 37646 3038 37674 3066
rect 36134 2254 36162 2282
rect 34454 1750 34482 1778
rect 35742 2225 35770 2226
rect 35742 2199 35743 2225
rect 35743 2199 35769 2225
rect 35769 2199 35770 2225
rect 35742 2198 35770 2199
rect 35910 2225 35938 2226
rect 35910 2199 35911 2225
rect 35911 2199 35937 2225
rect 35937 2199 35938 2225
rect 35910 2198 35938 2199
rect 35686 2169 35714 2170
rect 35686 2143 35687 2169
rect 35687 2143 35713 2169
rect 35713 2143 35714 2169
rect 35686 2142 35714 2143
rect 35182 1721 35210 1722
rect 35182 1695 35183 1721
rect 35183 1695 35209 1721
rect 35209 1695 35210 1721
rect 35182 1694 35210 1695
rect 35350 1750 35378 1778
rect 36582 2422 36610 2450
rect 34582 1581 34610 1582
rect 34582 1555 34600 1581
rect 34600 1555 34610 1581
rect 34582 1554 34610 1555
rect 34634 1581 34662 1582
rect 34634 1555 34636 1581
rect 34636 1555 34662 1581
rect 34634 1554 34662 1555
rect 34686 1581 34714 1582
rect 34738 1581 34766 1582
rect 34686 1555 34698 1581
rect 34698 1555 34714 1581
rect 34738 1555 34760 1581
rect 34760 1555 34766 1581
rect 34686 1554 34714 1555
rect 34738 1554 34766 1555
rect 34790 1554 34818 1582
rect 34842 1581 34870 1582
rect 34894 1581 34922 1582
rect 34842 1555 34848 1581
rect 34848 1555 34870 1581
rect 34894 1555 34910 1581
rect 34910 1555 34922 1581
rect 34842 1554 34870 1555
rect 34894 1554 34922 1555
rect 34946 1581 34974 1582
rect 34946 1555 34972 1581
rect 34972 1555 34974 1581
rect 34946 1554 34974 1555
rect 34998 1581 35026 1582
rect 34998 1555 35008 1581
rect 35008 1555 35026 1581
rect 34998 1554 35026 1555
rect 36694 2254 36722 2282
rect 37590 2366 37618 2394
rect 37646 2478 37674 2506
rect 37534 2142 37562 2170
rect 38990 5614 39018 5642
rect 37702 4998 37730 5026
rect 38206 4830 38234 4858
rect 38150 3737 38178 3738
rect 38150 3711 38151 3737
rect 38151 3711 38177 3737
rect 38177 3711 38178 3737
rect 38150 3710 38178 3711
rect 38206 2478 38234 2506
rect 37702 2198 37730 2226
rect 38150 2422 38178 2450
rect 38206 2366 38234 2394
rect 38598 4214 38626 4242
rect 38822 4214 38850 4242
rect 38654 3934 38682 3962
rect 38654 3737 38682 3738
rect 38654 3711 38655 3737
rect 38655 3711 38681 3737
rect 38681 3711 38682 3737
rect 38654 3710 38682 3711
rect 37814 2142 37842 2170
rect 37082 1973 37110 1974
rect 37082 1947 37100 1973
rect 37100 1947 37110 1973
rect 37082 1946 37110 1947
rect 37134 1973 37162 1974
rect 37134 1947 37136 1973
rect 37136 1947 37162 1973
rect 37134 1946 37162 1947
rect 37186 1973 37214 1974
rect 37238 1973 37266 1974
rect 37186 1947 37198 1973
rect 37198 1947 37214 1973
rect 37238 1947 37260 1973
rect 37260 1947 37266 1973
rect 37186 1946 37214 1947
rect 37238 1946 37266 1947
rect 37290 1946 37318 1974
rect 37342 1973 37370 1974
rect 37394 1973 37422 1974
rect 37342 1947 37348 1973
rect 37348 1947 37370 1973
rect 37394 1947 37410 1973
rect 37410 1947 37422 1973
rect 37342 1946 37370 1947
rect 37394 1946 37422 1947
rect 37446 1973 37474 1974
rect 37446 1947 37472 1973
rect 37472 1947 37474 1973
rect 37446 1946 37474 1947
rect 37498 1973 37526 1974
rect 37498 1947 37508 1973
rect 37508 1947 37526 1973
rect 37498 1946 37526 1947
rect 38150 2142 38178 2170
rect 38262 2198 38290 2226
rect 38318 2870 38346 2898
rect 38654 2870 38682 2898
rect 38934 3934 38962 3962
rect 38822 3737 38850 3738
rect 38822 3711 38823 3737
rect 38823 3711 38849 3737
rect 38849 3711 38850 3737
rect 38822 3710 38850 3711
rect 38822 2870 38850 2898
rect 38710 2225 38738 2226
rect 38710 2199 38711 2225
rect 38711 2199 38737 2225
rect 38737 2199 38738 2225
rect 38710 2198 38738 2199
rect 38878 2225 38906 2226
rect 38878 2199 38879 2225
rect 38879 2199 38905 2225
rect 38905 2199 38906 2225
rect 38878 2198 38906 2199
rect 38934 2169 38962 2170
rect 38934 2143 38935 2169
rect 38935 2143 38961 2169
rect 38961 2143 38962 2169
rect 38934 2142 38962 2143
rect 39046 2478 39074 2506
rect 38822 2086 38850 2114
rect 38934 1777 38962 1778
rect 38934 1751 38935 1777
rect 38935 1751 38961 1777
rect 38961 1751 38962 1777
rect 38934 1750 38962 1751
rect 39102 1750 39130 1778
<< metal3 >>
rect 2077 18410 2082 18438
rect 2110 18410 2134 18438
rect 2162 18410 2186 18438
rect 2214 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2394 18438
rect 2422 18410 2446 18438
rect 2474 18410 2498 18438
rect 2526 18410 2531 18438
rect 7077 18410 7082 18438
rect 7110 18410 7134 18438
rect 7162 18410 7186 18438
rect 7214 18410 7238 18438
rect 7266 18410 7290 18438
rect 7318 18410 7342 18438
rect 7370 18410 7394 18438
rect 7422 18410 7446 18438
rect 7474 18410 7498 18438
rect 7526 18410 7531 18438
rect 12077 18410 12082 18438
rect 12110 18410 12134 18438
rect 12162 18410 12186 18438
rect 12214 18410 12238 18438
rect 12266 18410 12290 18438
rect 12318 18410 12342 18438
rect 12370 18410 12394 18438
rect 12422 18410 12446 18438
rect 12474 18410 12498 18438
rect 12526 18410 12531 18438
rect 17077 18410 17082 18438
rect 17110 18410 17134 18438
rect 17162 18410 17186 18438
rect 17214 18410 17238 18438
rect 17266 18410 17290 18438
rect 17318 18410 17342 18438
rect 17370 18410 17394 18438
rect 17422 18410 17446 18438
rect 17474 18410 17498 18438
rect 17526 18410 17531 18438
rect 22077 18410 22082 18438
rect 22110 18410 22134 18438
rect 22162 18410 22186 18438
rect 22214 18410 22238 18438
rect 22266 18410 22290 18438
rect 22318 18410 22342 18438
rect 22370 18410 22394 18438
rect 22422 18410 22446 18438
rect 22474 18410 22498 18438
rect 22526 18410 22531 18438
rect 27077 18410 27082 18438
rect 27110 18410 27134 18438
rect 27162 18410 27186 18438
rect 27214 18410 27238 18438
rect 27266 18410 27290 18438
rect 27318 18410 27342 18438
rect 27370 18410 27394 18438
rect 27422 18410 27446 18438
rect 27474 18410 27498 18438
rect 27526 18410 27531 18438
rect 32077 18410 32082 18438
rect 32110 18410 32134 18438
rect 32162 18410 32186 18438
rect 32214 18410 32238 18438
rect 32266 18410 32290 18438
rect 32318 18410 32342 18438
rect 32370 18410 32394 18438
rect 32422 18410 32446 18438
rect 32474 18410 32498 18438
rect 32526 18410 32531 18438
rect 37077 18410 37082 18438
rect 37110 18410 37134 18438
rect 37162 18410 37186 18438
rect 37214 18410 37238 18438
rect 37266 18410 37290 18438
rect 37318 18410 37342 18438
rect 37370 18410 37394 18438
rect 37422 18410 37446 18438
rect 37474 18410 37498 18438
rect 37526 18410 37531 18438
rect 4577 18018 4582 18046
rect 4610 18018 4634 18046
rect 4662 18018 4686 18046
rect 4714 18018 4738 18046
rect 4766 18018 4790 18046
rect 4818 18018 4842 18046
rect 4870 18018 4894 18046
rect 4922 18018 4946 18046
rect 4974 18018 4998 18046
rect 5026 18018 5031 18046
rect 9577 18018 9582 18046
rect 9610 18018 9634 18046
rect 9662 18018 9686 18046
rect 9714 18018 9738 18046
rect 9766 18018 9790 18046
rect 9818 18018 9842 18046
rect 9870 18018 9894 18046
rect 9922 18018 9946 18046
rect 9974 18018 9998 18046
rect 10026 18018 10031 18046
rect 14577 18018 14582 18046
rect 14610 18018 14634 18046
rect 14662 18018 14686 18046
rect 14714 18018 14738 18046
rect 14766 18018 14790 18046
rect 14818 18018 14842 18046
rect 14870 18018 14894 18046
rect 14922 18018 14946 18046
rect 14974 18018 14998 18046
rect 15026 18018 15031 18046
rect 19577 18018 19582 18046
rect 19610 18018 19634 18046
rect 19662 18018 19686 18046
rect 19714 18018 19738 18046
rect 19766 18018 19790 18046
rect 19818 18018 19842 18046
rect 19870 18018 19894 18046
rect 19922 18018 19946 18046
rect 19974 18018 19998 18046
rect 20026 18018 20031 18046
rect 24577 18018 24582 18046
rect 24610 18018 24634 18046
rect 24662 18018 24686 18046
rect 24714 18018 24738 18046
rect 24766 18018 24790 18046
rect 24818 18018 24842 18046
rect 24870 18018 24894 18046
rect 24922 18018 24946 18046
rect 24974 18018 24998 18046
rect 25026 18018 25031 18046
rect 29577 18018 29582 18046
rect 29610 18018 29634 18046
rect 29662 18018 29686 18046
rect 29714 18018 29738 18046
rect 29766 18018 29790 18046
rect 29818 18018 29842 18046
rect 29870 18018 29894 18046
rect 29922 18018 29946 18046
rect 29974 18018 29998 18046
rect 30026 18018 30031 18046
rect 34577 18018 34582 18046
rect 34610 18018 34634 18046
rect 34662 18018 34686 18046
rect 34714 18018 34738 18046
rect 34766 18018 34790 18046
rect 34818 18018 34842 18046
rect 34870 18018 34894 18046
rect 34922 18018 34946 18046
rect 34974 18018 34998 18046
rect 35026 18018 35031 18046
rect 2077 17626 2082 17654
rect 2110 17626 2134 17654
rect 2162 17626 2186 17654
rect 2214 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2394 17654
rect 2422 17626 2446 17654
rect 2474 17626 2498 17654
rect 2526 17626 2531 17654
rect 7077 17626 7082 17654
rect 7110 17626 7134 17654
rect 7162 17626 7186 17654
rect 7214 17626 7238 17654
rect 7266 17626 7290 17654
rect 7318 17626 7342 17654
rect 7370 17626 7394 17654
rect 7422 17626 7446 17654
rect 7474 17626 7498 17654
rect 7526 17626 7531 17654
rect 12077 17626 12082 17654
rect 12110 17626 12134 17654
rect 12162 17626 12186 17654
rect 12214 17626 12238 17654
rect 12266 17626 12290 17654
rect 12318 17626 12342 17654
rect 12370 17626 12394 17654
rect 12422 17626 12446 17654
rect 12474 17626 12498 17654
rect 12526 17626 12531 17654
rect 17077 17626 17082 17654
rect 17110 17626 17134 17654
rect 17162 17626 17186 17654
rect 17214 17626 17238 17654
rect 17266 17626 17290 17654
rect 17318 17626 17342 17654
rect 17370 17626 17394 17654
rect 17422 17626 17446 17654
rect 17474 17626 17498 17654
rect 17526 17626 17531 17654
rect 22077 17626 22082 17654
rect 22110 17626 22134 17654
rect 22162 17626 22186 17654
rect 22214 17626 22238 17654
rect 22266 17626 22290 17654
rect 22318 17626 22342 17654
rect 22370 17626 22394 17654
rect 22422 17626 22446 17654
rect 22474 17626 22498 17654
rect 22526 17626 22531 17654
rect 27077 17626 27082 17654
rect 27110 17626 27134 17654
rect 27162 17626 27186 17654
rect 27214 17626 27238 17654
rect 27266 17626 27290 17654
rect 27318 17626 27342 17654
rect 27370 17626 27394 17654
rect 27422 17626 27446 17654
rect 27474 17626 27498 17654
rect 27526 17626 27531 17654
rect 32077 17626 32082 17654
rect 32110 17626 32134 17654
rect 32162 17626 32186 17654
rect 32214 17626 32238 17654
rect 32266 17626 32290 17654
rect 32318 17626 32342 17654
rect 32370 17626 32394 17654
rect 32422 17626 32446 17654
rect 32474 17626 32498 17654
rect 32526 17626 32531 17654
rect 37077 17626 37082 17654
rect 37110 17626 37134 17654
rect 37162 17626 37186 17654
rect 37214 17626 37238 17654
rect 37266 17626 37290 17654
rect 37318 17626 37342 17654
rect 37370 17626 37394 17654
rect 37422 17626 37446 17654
rect 37474 17626 37498 17654
rect 37526 17626 37531 17654
rect 12609 17318 12614 17346
rect 12642 17318 23926 17346
rect 23954 17318 23959 17346
rect 4577 17234 4582 17262
rect 4610 17234 4634 17262
rect 4662 17234 4686 17262
rect 4714 17234 4738 17262
rect 4766 17234 4790 17262
rect 4818 17234 4842 17262
rect 4870 17234 4894 17262
rect 4922 17234 4946 17262
rect 4974 17234 4998 17262
rect 5026 17234 5031 17262
rect 9577 17234 9582 17262
rect 9610 17234 9634 17262
rect 9662 17234 9686 17262
rect 9714 17234 9738 17262
rect 9766 17234 9790 17262
rect 9818 17234 9842 17262
rect 9870 17234 9894 17262
rect 9922 17234 9946 17262
rect 9974 17234 9998 17262
rect 10026 17234 10031 17262
rect 14577 17234 14582 17262
rect 14610 17234 14634 17262
rect 14662 17234 14686 17262
rect 14714 17234 14738 17262
rect 14766 17234 14790 17262
rect 14818 17234 14842 17262
rect 14870 17234 14894 17262
rect 14922 17234 14946 17262
rect 14974 17234 14998 17262
rect 15026 17234 15031 17262
rect 19577 17234 19582 17262
rect 19610 17234 19634 17262
rect 19662 17234 19686 17262
rect 19714 17234 19738 17262
rect 19766 17234 19790 17262
rect 19818 17234 19842 17262
rect 19870 17234 19894 17262
rect 19922 17234 19946 17262
rect 19974 17234 19998 17262
rect 20026 17234 20031 17262
rect 24577 17234 24582 17262
rect 24610 17234 24634 17262
rect 24662 17234 24686 17262
rect 24714 17234 24738 17262
rect 24766 17234 24790 17262
rect 24818 17234 24842 17262
rect 24870 17234 24894 17262
rect 24922 17234 24946 17262
rect 24974 17234 24998 17262
rect 25026 17234 25031 17262
rect 29577 17234 29582 17262
rect 29610 17234 29634 17262
rect 29662 17234 29686 17262
rect 29714 17234 29738 17262
rect 29766 17234 29790 17262
rect 29818 17234 29842 17262
rect 29870 17234 29894 17262
rect 29922 17234 29946 17262
rect 29974 17234 29998 17262
rect 30026 17234 30031 17262
rect 34577 17234 34582 17262
rect 34610 17234 34634 17262
rect 34662 17234 34686 17262
rect 34714 17234 34738 17262
rect 34766 17234 34790 17262
rect 34818 17234 34842 17262
rect 34870 17234 34894 17262
rect 34922 17234 34946 17262
rect 34974 17234 34998 17262
rect 35026 17234 35031 17262
rect 2077 16842 2082 16870
rect 2110 16842 2134 16870
rect 2162 16842 2186 16870
rect 2214 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2394 16870
rect 2422 16842 2446 16870
rect 2474 16842 2498 16870
rect 2526 16842 2531 16870
rect 7077 16842 7082 16870
rect 7110 16842 7134 16870
rect 7162 16842 7186 16870
rect 7214 16842 7238 16870
rect 7266 16842 7290 16870
rect 7318 16842 7342 16870
rect 7370 16842 7394 16870
rect 7422 16842 7446 16870
rect 7474 16842 7498 16870
rect 7526 16842 7531 16870
rect 12077 16842 12082 16870
rect 12110 16842 12134 16870
rect 12162 16842 12186 16870
rect 12214 16842 12238 16870
rect 12266 16842 12290 16870
rect 12318 16842 12342 16870
rect 12370 16842 12394 16870
rect 12422 16842 12446 16870
rect 12474 16842 12498 16870
rect 12526 16842 12531 16870
rect 17077 16842 17082 16870
rect 17110 16842 17134 16870
rect 17162 16842 17186 16870
rect 17214 16842 17238 16870
rect 17266 16842 17290 16870
rect 17318 16842 17342 16870
rect 17370 16842 17394 16870
rect 17422 16842 17446 16870
rect 17474 16842 17498 16870
rect 17526 16842 17531 16870
rect 22077 16842 22082 16870
rect 22110 16842 22134 16870
rect 22162 16842 22186 16870
rect 22214 16842 22238 16870
rect 22266 16842 22290 16870
rect 22318 16842 22342 16870
rect 22370 16842 22394 16870
rect 22422 16842 22446 16870
rect 22474 16842 22498 16870
rect 22526 16842 22531 16870
rect 27077 16842 27082 16870
rect 27110 16842 27134 16870
rect 27162 16842 27186 16870
rect 27214 16842 27238 16870
rect 27266 16842 27290 16870
rect 27318 16842 27342 16870
rect 27370 16842 27394 16870
rect 27422 16842 27446 16870
rect 27474 16842 27498 16870
rect 27526 16842 27531 16870
rect 32077 16842 32082 16870
rect 32110 16842 32134 16870
rect 32162 16842 32186 16870
rect 32214 16842 32238 16870
rect 32266 16842 32290 16870
rect 32318 16842 32342 16870
rect 32370 16842 32394 16870
rect 32422 16842 32446 16870
rect 32474 16842 32498 16870
rect 32526 16842 32531 16870
rect 37077 16842 37082 16870
rect 37110 16842 37134 16870
rect 37162 16842 37186 16870
rect 37214 16842 37238 16870
rect 37266 16842 37290 16870
rect 37318 16842 37342 16870
rect 37370 16842 37394 16870
rect 37422 16842 37446 16870
rect 37474 16842 37498 16870
rect 37526 16842 37531 16870
rect 11993 16590 11998 16618
rect 12026 16590 12334 16618
rect 12362 16590 13454 16618
rect 13482 16590 13790 16618
rect 13818 16590 13823 16618
rect 12614 16562 12642 16590
rect 12609 16534 12614 16562
rect 12642 16534 12647 16562
rect 4577 16450 4582 16478
rect 4610 16450 4634 16478
rect 4662 16450 4686 16478
rect 4714 16450 4738 16478
rect 4766 16450 4790 16478
rect 4818 16450 4842 16478
rect 4870 16450 4894 16478
rect 4922 16450 4946 16478
rect 4974 16450 4998 16478
rect 5026 16450 5031 16478
rect 9577 16450 9582 16478
rect 9610 16450 9634 16478
rect 9662 16450 9686 16478
rect 9714 16450 9738 16478
rect 9766 16450 9790 16478
rect 9818 16450 9842 16478
rect 9870 16450 9894 16478
rect 9922 16450 9946 16478
rect 9974 16450 9998 16478
rect 10026 16450 10031 16478
rect 14577 16450 14582 16478
rect 14610 16450 14634 16478
rect 14662 16450 14686 16478
rect 14714 16450 14738 16478
rect 14766 16450 14790 16478
rect 14818 16450 14842 16478
rect 14870 16450 14894 16478
rect 14922 16450 14946 16478
rect 14974 16450 14998 16478
rect 15026 16450 15031 16478
rect 19577 16450 19582 16478
rect 19610 16450 19634 16478
rect 19662 16450 19686 16478
rect 19714 16450 19738 16478
rect 19766 16450 19790 16478
rect 19818 16450 19842 16478
rect 19870 16450 19894 16478
rect 19922 16450 19946 16478
rect 19974 16450 19998 16478
rect 20026 16450 20031 16478
rect 24577 16450 24582 16478
rect 24610 16450 24634 16478
rect 24662 16450 24686 16478
rect 24714 16450 24738 16478
rect 24766 16450 24790 16478
rect 24818 16450 24842 16478
rect 24870 16450 24894 16478
rect 24922 16450 24946 16478
rect 24974 16450 24998 16478
rect 25026 16450 25031 16478
rect 29577 16450 29582 16478
rect 29610 16450 29634 16478
rect 29662 16450 29686 16478
rect 29714 16450 29738 16478
rect 29766 16450 29790 16478
rect 29818 16450 29842 16478
rect 29870 16450 29894 16478
rect 29922 16450 29946 16478
rect 29974 16450 29998 16478
rect 30026 16450 30031 16478
rect 34577 16450 34582 16478
rect 34610 16450 34634 16478
rect 34662 16450 34686 16478
rect 34714 16450 34738 16478
rect 34766 16450 34790 16478
rect 34818 16450 34842 16478
rect 34870 16450 34894 16478
rect 34922 16450 34946 16478
rect 34974 16450 34998 16478
rect 35026 16450 35031 16478
rect 10145 16310 10150 16338
rect 10178 16310 10822 16338
rect 10850 16310 11382 16338
rect 11410 16310 11415 16338
rect 5889 16254 5894 16282
rect 5922 16254 6118 16282
rect 6146 16254 7518 16282
rect 7546 16254 7551 16282
rect 9473 16254 9478 16282
rect 9506 16254 9982 16282
rect 10010 16254 10934 16282
rect 10962 16254 11158 16282
rect 11186 16254 11191 16282
rect 12945 16142 12950 16170
rect 12978 16142 13286 16170
rect 13314 16142 13319 16170
rect 2077 16058 2082 16086
rect 2110 16058 2134 16086
rect 2162 16058 2186 16086
rect 2214 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2394 16086
rect 2422 16058 2446 16086
rect 2474 16058 2498 16086
rect 2526 16058 2531 16086
rect 7077 16058 7082 16086
rect 7110 16058 7134 16086
rect 7162 16058 7186 16086
rect 7214 16058 7238 16086
rect 7266 16058 7290 16086
rect 7318 16058 7342 16086
rect 7370 16058 7394 16086
rect 7422 16058 7446 16086
rect 7474 16058 7498 16086
rect 7526 16058 7531 16086
rect 12077 16058 12082 16086
rect 12110 16058 12134 16086
rect 12162 16058 12186 16086
rect 12214 16058 12238 16086
rect 12266 16058 12290 16086
rect 12318 16058 12342 16086
rect 12370 16058 12394 16086
rect 12422 16058 12446 16086
rect 12474 16058 12498 16086
rect 12526 16058 12531 16086
rect 17077 16058 17082 16086
rect 17110 16058 17134 16086
rect 17162 16058 17186 16086
rect 17214 16058 17238 16086
rect 17266 16058 17290 16086
rect 17318 16058 17342 16086
rect 17370 16058 17394 16086
rect 17422 16058 17446 16086
rect 17474 16058 17498 16086
rect 17526 16058 17531 16086
rect 22077 16058 22082 16086
rect 22110 16058 22134 16086
rect 22162 16058 22186 16086
rect 22214 16058 22238 16086
rect 22266 16058 22290 16086
rect 22318 16058 22342 16086
rect 22370 16058 22394 16086
rect 22422 16058 22446 16086
rect 22474 16058 22498 16086
rect 22526 16058 22531 16086
rect 27077 16058 27082 16086
rect 27110 16058 27134 16086
rect 27162 16058 27186 16086
rect 27214 16058 27238 16086
rect 27266 16058 27290 16086
rect 27318 16058 27342 16086
rect 27370 16058 27394 16086
rect 27422 16058 27446 16086
rect 27474 16058 27498 16086
rect 27526 16058 27531 16086
rect 32077 16058 32082 16086
rect 32110 16058 32134 16086
rect 32162 16058 32186 16086
rect 32214 16058 32238 16086
rect 32266 16058 32290 16086
rect 32318 16058 32342 16086
rect 32370 16058 32394 16086
rect 32422 16058 32446 16086
rect 32474 16058 32498 16086
rect 32526 16058 32531 16086
rect 37077 16058 37082 16086
rect 37110 16058 37134 16086
rect 37162 16058 37186 16086
rect 37214 16058 37238 16086
rect 37266 16058 37290 16086
rect 37318 16058 37342 16086
rect 37370 16058 37394 16086
rect 37422 16058 37446 16086
rect 37474 16058 37498 16086
rect 37526 16058 37531 16086
rect 15409 15918 15414 15946
rect 15442 15918 16814 15946
rect 16842 15918 16926 15946
rect 16954 15918 16959 15946
rect 7793 15862 7798 15890
rect 7826 15862 9310 15890
rect 9338 15862 11102 15890
rect 11130 15862 15078 15890
rect 15106 15862 20286 15890
rect 20314 15862 20319 15890
rect 4577 15666 4582 15694
rect 4610 15666 4634 15694
rect 4662 15666 4686 15694
rect 4714 15666 4738 15694
rect 4766 15666 4790 15694
rect 4818 15666 4842 15694
rect 4870 15666 4894 15694
rect 4922 15666 4946 15694
rect 4974 15666 4998 15694
rect 5026 15666 5031 15694
rect 9577 15666 9582 15694
rect 9610 15666 9634 15694
rect 9662 15666 9686 15694
rect 9714 15666 9738 15694
rect 9766 15666 9790 15694
rect 9818 15666 9842 15694
rect 9870 15666 9894 15694
rect 9922 15666 9946 15694
rect 9974 15666 9998 15694
rect 10026 15666 10031 15694
rect 14577 15666 14582 15694
rect 14610 15666 14634 15694
rect 14662 15666 14686 15694
rect 14714 15666 14738 15694
rect 14766 15666 14790 15694
rect 14818 15666 14842 15694
rect 14870 15666 14894 15694
rect 14922 15666 14946 15694
rect 14974 15666 14998 15694
rect 15026 15666 15031 15694
rect 19577 15666 19582 15694
rect 19610 15666 19634 15694
rect 19662 15666 19686 15694
rect 19714 15666 19738 15694
rect 19766 15666 19790 15694
rect 19818 15666 19842 15694
rect 19870 15666 19894 15694
rect 19922 15666 19946 15694
rect 19974 15666 19998 15694
rect 20026 15666 20031 15694
rect 24577 15666 24582 15694
rect 24610 15666 24634 15694
rect 24662 15666 24686 15694
rect 24714 15666 24738 15694
rect 24766 15666 24790 15694
rect 24818 15666 24842 15694
rect 24870 15666 24894 15694
rect 24922 15666 24946 15694
rect 24974 15666 24998 15694
rect 25026 15666 25031 15694
rect 29577 15666 29582 15694
rect 29610 15666 29634 15694
rect 29662 15666 29686 15694
rect 29714 15666 29738 15694
rect 29766 15666 29790 15694
rect 29818 15666 29842 15694
rect 29870 15666 29894 15694
rect 29922 15666 29946 15694
rect 29974 15666 29998 15694
rect 30026 15666 30031 15694
rect 34577 15666 34582 15694
rect 34610 15666 34634 15694
rect 34662 15666 34686 15694
rect 34714 15666 34738 15694
rect 34766 15666 34790 15694
rect 34818 15666 34842 15694
rect 34870 15666 34894 15694
rect 34922 15666 34946 15694
rect 34974 15666 34998 15694
rect 35026 15666 35031 15694
rect 7009 15470 7014 15498
rect 7042 15470 7294 15498
rect 7322 15470 7798 15498
rect 7826 15470 7831 15498
rect 2077 15274 2082 15302
rect 2110 15274 2134 15302
rect 2162 15274 2186 15302
rect 2214 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2394 15302
rect 2422 15274 2446 15302
rect 2474 15274 2498 15302
rect 2526 15274 2531 15302
rect 7077 15274 7082 15302
rect 7110 15274 7134 15302
rect 7162 15274 7186 15302
rect 7214 15274 7238 15302
rect 7266 15274 7290 15302
rect 7318 15274 7342 15302
rect 7370 15274 7394 15302
rect 7422 15274 7446 15302
rect 7474 15274 7498 15302
rect 7526 15274 7531 15302
rect 12077 15274 12082 15302
rect 12110 15274 12134 15302
rect 12162 15274 12186 15302
rect 12214 15274 12238 15302
rect 12266 15274 12290 15302
rect 12318 15274 12342 15302
rect 12370 15274 12394 15302
rect 12422 15274 12446 15302
rect 12474 15274 12498 15302
rect 12526 15274 12531 15302
rect 17077 15274 17082 15302
rect 17110 15274 17134 15302
rect 17162 15274 17186 15302
rect 17214 15274 17238 15302
rect 17266 15274 17290 15302
rect 17318 15274 17342 15302
rect 17370 15274 17394 15302
rect 17422 15274 17446 15302
rect 17474 15274 17498 15302
rect 17526 15274 17531 15302
rect 22077 15274 22082 15302
rect 22110 15274 22134 15302
rect 22162 15274 22186 15302
rect 22214 15274 22238 15302
rect 22266 15274 22290 15302
rect 22318 15274 22342 15302
rect 22370 15274 22394 15302
rect 22422 15274 22446 15302
rect 22474 15274 22498 15302
rect 22526 15274 22531 15302
rect 27077 15274 27082 15302
rect 27110 15274 27134 15302
rect 27162 15274 27186 15302
rect 27214 15274 27238 15302
rect 27266 15274 27290 15302
rect 27318 15274 27342 15302
rect 27370 15274 27394 15302
rect 27422 15274 27446 15302
rect 27474 15274 27498 15302
rect 27526 15274 27531 15302
rect 32077 15274 32082 15302
rect 32110 15274 32134 15302
rect 32162 15274 32186 15302
rect 32214 15274 32238 15302
rect 32266 15274 32290 15302
rect 32318 15274 32342 15302
rect 32370 15274 32394 15302
rect 32422 15274 32446 15302
rect 32474 15274 32498 15302
rect 32526 15274 32531 15302
rect 37077 15274 37082 15302
rect 37110 15274 37134 15302
rect 37162 15274 37186 15302
rect 37214 15274 37238 15302
rect 37266 15274 37290 15302
rect 37318 15274 37342 15302
rect 37370 15274 37394 15302
rect 37422 15274 37446 15302
rect 37474 15274 37498 15302
rect 37526 15274 37531 15302
rect 10066 15134 10150 15162
rect 10178 15134 10183 15162
rect 24481 15134 24486 15162
rect 24514 15134 26894 15162
rect 26922 15134 26927 15162
rect 10066 15106 10094 15134
rect 8969 15078 8974 15106
rect 9002 15078 10094 15106
rect 13057 15078 13062 15106
rect 13090 15078 14294 15106
rect 14322 15078 14798 15106
rect 14826 15078 16534 15106
rect 16562 15078 16567 15106
rect 7569 15022 7574 15050
rect 7602 15022 16478 15050
rect 16506 15022 16511 15050
rect 4577 14882 4582 14910
rect 4610 14882 4634 14910
rect 4662 14882 4686 14910
rect 4714 14882 4738 14910
rect 4766 14882 4790 14910
rect 4818 14882 4842 14910
rect 4870 14882 4894 14910
rect 4922 14882 4946 14910
rect 4974 14882 4998 14910
rect 5026 14882 5031 14910
rect 9577 14882 9582 14910
rect 9610 14882 9634 14910
rect 9662 14882 9686 14910
rect 9714 14882 9738 14910
rect 9766 14882 9790 14910
rect 9818 14882 9842 14910
rect 9870 14882 9894 14910
rect 9922 14882 9946 14910
rect 9974 14882 9998 14910
rect 10026 14882 10031 14910
rect 14577 14882 14582 14910
rect 14610 14882 14634 14910
rect 14662 14882 14686 14910
rect 14714 14882 14738 14910
rect 14766 14882 14790 14910
rect 14818 14882 14842 14910
rect 14870 14882 14894 14910
rect 14922 14882 14946 14910
rect 14974 14882 14998 14910
rect 15026 14882 15031 14910
rect 19577 14882 19582 14910
rect 19610 14882 19634 14910
rect 19662 14882 19686 14910
rect 19714 14882 19738 14910
rect 19766 14882 19790 14910
rect 19818 14882 19842 14910
rect 19870 14882 19894 14910
rect 19922 14882 19946 14910
rect 19974 14882 19998 14910
rect 20026 14882 20031 14910
rect 24577 14882 24582 14910
rect 24610 14882 24634 14910
rect 24662 14882 24686 14910
rect 24714 14882 24738 14910
rect 24766 14882 24790 14910
rect 24818 14882 24842 14910
rect 24870 14882 24894 14910
rect 24922 14882 24946 14910
rect 24974 14882 24998 14910
rect 25026 14882 25031 14910
rect 29577 14882 29582 14910
rect 29610 14882 29634 14910
rect 29662 14882 29686 14910
rect 29714 14882 29738 14910
rect 29766 14882 29790 14910
rect 29818 14882 29842 14910
rect 29870 14882 29894 14910
rect 29922 14882 29946 14910
rect 29974 14882 29998 14910
rect 30026 14882 30031 14910
rect 34577 14882 34582 14910
rect 34610 14882 34634 14910
rect 34662 14882 34686 14910
rect 34714 14882 34738 14910
rect 34766 14882 34790 14910
rect 34818 14882 34842 14910
rect 34870 14882 34894 14910
rect 34922 14882 34946 14910
rect 34974 14882 34998 14910
rect 35026 14882 35031 14910
rect 6001 14742 6006 14770
rect 6034 14742 13062 14770
rect 13090 14742 13095 14770
rect 2417 14686 2422 14714
rect 2450 14686 2590 14714
rect 2618 14686 3038 14714
rect 3066 14686 3598 14714
rect 3626 14686 3631 14714
rect 5273 14686 5278 14714
rect 5306 14686 5838 14714
rect 5866 14686 5871 14714
rect 12441 14686 12446 14714
rect 12474 14686 12838 14714
rect 12866 14686 12871 14714
rect 16473 14686 16478 14714
rect 16506 14686 17094 14714
rect 17122 14686 18438 14714
rect 18466 14686 18471 14714
rect 3817 14630 3822 14658
rect 3850 14630 6846 14658
rect 6874 14630 18270 14658
rect 18298 14630 18774 14658
rect 18802 14630 18807 14658
rect 2077 14490 2082 14518
rect 2110 14490 2134 14518
rect 2162 14490 2186 14518
rect 2214 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2394 14518
rect 2422 14490 2446 14518
rect 2474 14490 2498 14518
rect 2526 14490 2531 14518
rect 7077 14490 7082 14518
rect 7110 14490 7134 14518
rect 7162 14490 7186 14518
rect 7214 14490 7238 14518
rect 7266 14490 7290 14518
rect 7318 14490 7342 14518
rect 7370 14490 7394 14518
rect 7422 14490 7446 14518
rect 7474 14490 7498 14518
rect 7526 14490 7531 14518
rect 12077 14490 12082 14518
rect 12110 14490 12134 14518
rect 12162 14490 12186 14518
rect 12214 14490 12238 14518
rect 12266 14490 12290 14518
rect 12318 14490 12342 14518
rect 12370 14490 12394 14518
rect 12422 14490 12446 14518
rect 12474 14490 12498 14518
rect 12526 14490 12531 14518
rect 17077 14490 17082 14518
rect 17110 14490 17134 14518
rect 17162 14490 17186 14518
rect 17214 14490 17238 14518
rect 17266 14490 17290 14518
rect 17318 14490 17342 14518
rect 17370 14490 17394 14518
rect 17422 14490 17446 14518
rect 17474 14490 17498 14518
rect 17526 14490 17531 14518
rect 22077 14490 22082 14518
rect 22110 14490 22134 14518
rect 22162 14490 22186 14518
rect 22214 14490 22238 14518
rect 22266 14490 22290 14518
rect 22318 14490 22342 14518
rect 22370 14490 22394 14518
rect 22422 14490 22446 14518
rect 22474 14490 22498 14518
rect 22526 14490 22531 14518
rect 27077 14490 27082 14518
rect 27110 14490 27134 14518
rect 27162 14490 27186 14518
rect 27214 14490 27238 14518
rect 27266 14490 27290 14518
rect 27318 14490 27342 14518
rect 27370 14490 27394 14518
rect 27422 14490 27446 14518
rect 27474 14490 27498 14518
rect 27526 14490 27531 14518
rect 32077 14490 32082 14518
rect 32110 14490 32134 14518
rect 32162 14490 32186 14518
rect 32214 14490 32238 14518
rect 32266 14490 32290 14518
rect 32318 14490 32342 14518
rect 32370 14490 32394 14518
rect 32422 14490 32446 14518
rect 32474 14490 32498 14518
rect 32526 14490 32531 14518
rect 37077 14490 37082 14518
rect 37110 14490 37134 14518
rect 37162 14490 37186 14518
rect 37214 14490 37238 14518
rect 37266 14490 37290 14518
rect 37318 14490 37342 14518
rect 37370 14490 37394 14518
rect 37422 14490 37446 14518
rect 37474 14490 37498 14518
rect 37526 14490 37531 14518
rect 2473 14350 2478 14378
rect 2506 14350 4494 14378
rect 4522 14350 4998 14378
rect 5026 14350 6398 14378
rect 6426 14350 6431 14378
rect 2417 14294 2422 14322
rect 2450 14294 2590 14322
rect 2618 14294 2623 14322
rect 3817 14294 3822 14322
rect 3850 14294 5278 14322
rect 5306 14294 5311 14322
rect 10873 14294 10878 14322
rect 10906 14294 12446 14322
rect 12474 14294 12894 14322
rect 12922 14294 14014 14322
rect 14042 14294 14047 14322
rect 18769 14294 18774 14322
rect 18802 14294 20230 14322
rect 20258 14294 20846 14322
rect 20874 14294 20879 14322
rect 17425 14238 17430 14266
rect 17458 14238 17766 14266
rect 17794 14238 18718 14266
rect 18746 14238 18942 14266
rect 18970 14238 18975 14266
rect 23865 14238 23870 14266
rect 23898 14238 25158 14266
rect 25186 14238 25191 14266
rect 4577 14098 4582 14126
rect 4610 14098 4634 14126
rect 4662 14098 4686 14126
rect 4714 14098 4738 14126
rect 4766 14098 4790 14126
rect 4818 14098 4842 14126
rect 4870 14098 4894 14126
rect 4922 14098 4946 14126
rect 4974 14098 4998 14126
rect 5026 14098 5031 14126
rect 9577 14098 9582 14126
rect 9610 14098 9634 14126
rect 9662 14098 9686 14126
rect 9714 14098 9738 14126
rect 9766 14098 9790 14126
rect 9818 14098 9842 14126
rect 9870 14098 9894 14126
rect 9922 14098 9946 14126
rect 9974 14098 9998 14126
rect 10026 14098 10031 14126
rect 14577 14098 14582 14126
rect 14610 14098 14634 14126
rect 14662 14098 14686 14126
rect 14714 14098 14738 14126
rect 14766 14098 14790 14126
rect 14818 14098 14842 14126
rect 14870 14098 14894 14126
rect 14922 14098 14946 14126
rect 14974 14098 14998 14126
rect 15026 14098 15031 14126
rect 19577 14098 19582 14126
rect 19610 14098 19634 14126
rect 19662 14098 19686 14126
rect 19714 14098 19738 14126
rect 19766 14098 19790 14126
rect 19818 14098 19842 14126
rect 19870 14098 19894 14126
rect 19922 14098 19946 14126
rect 19974 14098 19998 14126
rect 20026 14098 20031 14126
rect 24577 14098 24582 14126
rect 24610 14098 24634 14126
rect 24662 14098 24686 14126
rect 24714 14098 24738 14126
rect 24766 14098 24790 14126
rect 24818 14098 24842 14126
rect 24870 14098 24894 14126
rect 24922 14098 24946 14126
rect 24974 14098 24998 14126
rect 25026 14098 25031 14126
rect 29577 14098 29582 14126
rect 29610 14098 29634 14126
rect 29662 14098 29686 14126
rect 29714 14098 29738 14126
rect 29766 14098 29790 14126
rect 29818 14098 29842 14126
rect 29870 14098 29894 14126
rect 29922 14098 29946 14126
rect 29974 14098 29998 14126
rect 30026 14098 30031 14126
rect 34577 14098 34582 14126
rect 34610 14098 34634 14126
rect 34662 14098 34686 14126
rect 34714 14098 34738 14126
rect 34766 14098 34790 14126
rect 34818 14098 34842 14126
rect 34870 14098 34894 14126
rect 34922 14098 34946 14126
rect 34974 14098 34998 14126
rect 35026 14098 35031 14126
rect 6953 13958 6958 13986
rect 6986 13958 8470 13986
rect 8498 13958 8974 13986
rect 9002 13958 9007 13986
rect 5833 13902 5838 13930
rect 5866 13902 7014 13930
rect 7042 13902 7047 13930
rect 16361 13902 16366 13930
rect 16394 13902 20790 13930
rect 20818 13902 21854 13930
rect 21826 13874 21854 13902
rect 21826 13846 22582 13874
rect 22610 13846 22615 13874
rect 2077 13706 2082 13734
rect 2110 13706 2134 13734
rect 2162 13706 2186 13734
rect 2214 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2394 13734
rect 2422 13706 2446 13734
rect 2474 13706 2498 13734
rect 2526 13706 2531 13734
rect 7077 13706 7082 13734
rect 7110 13706 7134 13734
rect 7162 13706 7186 13734
rect 7214 13706 7238 13734
rect 7266 13706 7290 13734
rect 7318 13706 7342 13734
rect 7370 13706 7394 13734
rect 7422 13706 7446 13734
rect 7474 13706 7498 13734
rect 7526 13706 7531 13734
rect 12077 13706 12082 13734
rect 12110 13706 12134 13734
rect 12162 13706 12186 13734
rect 12214 13706 12238 13734
rect 12266 13706 12290 13734
rect 12318 13706 12342 13734
rect 12370 13706 12394 13734
rect 12422 13706 12446 13734
rect 12474 13706 12498 13734
rect 12526 13706 12531 13734
rect 17077 13706 17082 13734
rect 17110 13706 17134 13734
rect 17162 13706 17186 13734
rect 17214 13706 17238 13734
rect 17266 13706 17290 13734
rect 17318 13706 17342 13734
rect 17370 13706 17394 13734
rect 17422 13706 17446 13734
rect 17474 13706 17498 13734
rect 17526 13706 17531 13734
rect 22077 13706 22082 13734
rect 22110 13706 22134 13734
rect 22162 13706 22186 13734
rect 22214 13706 22238 13734
rect 22266 13706 22290 13734
rect 22318 13706 22342 13734
rect 22370 13706 22394 13734
rect 22422 13706 22446 13734
rect 22474 13706 22498 13734
rect 22526 13706 22531 13734
rect 27077 13706 27082 13734
rect 27110 13706 27134 13734
rect 27162 13706 27186 13734
rect 27214 13706 27238 13734
rect 27266 13706 27290 13734
rect 27318 13706 27342 13734
rect 27370 13706 27394 13734
rect 27422 13706 27446 13734
rect 27474 13706 27498 13734
rect 27526 13706 27531 13734
rect 32077 13706 32082 13734
rect 32110 13706 32134 13734
rect 32162 13706 32186 13734
rect 32214 13706 32238 13734
rect 32266 13706 32290 13734
rect 32318 13706 32342 13734
rect 32370 13706 32394 13734
rect 32422 13706 32446 13734
rect 32474 13706 32498 13734
rect 32526 13706 32531 13734
rect 37077 13706 37082 13734
rect 37110 13706 37134 13734
rect 37162 13706 37186 13734
rect 37214 13706 37238 13734
rect 37266 13706 37290 13734
rect 37318 13706 37342 13734
rect 37370 13706 37394 13734
rect 37422 13706 37446 13734
rect 37474 13706 37498 13734
rect 37526 13706 37531 13734
rect 4097 13510 4102 13538
rect 4130 13510 5278 13538
rect 5306 13510 5838 13538
rect 5866 13510 5871 13538
rect 6393 13510 6398 13538
rect 6426 13510 6902 13538
rect 6930 13510 6935 13538
rect 16529 13510 16534 13538
rect 16562 13510 16982 13538
rect 17010 13510 17015 13538
rect 18545 13510 18550 13538
rect 18578 13510 19054 13538
rect 19082 13510 20510 13538
rect 20538 13510 20543 13538
rect 21401 13510 21406 13538
rect 21434 13510 21742 13538
rect 21770 13510 23422 13538
rect 23450 13510 23870 13538
rect 23898 13510 23903 13538
rect 6449 13454 6454 13482
rect 6482 13454 6958 13482
rect 6986 13454 6991 13482
rect 15465 13454 15470 13482
rect 15498 13454 15862 13482
rect 15890 13454 17430 13482
rect 17458 13454 17463 13482
rect 21233 13454 21238 13482
rect 21266 13454 21462 13482
rect 21490 13454 21495 13482
rect 22521 13454 22526 13482
rect 22554 13454 23030 13482
rect 23058 13454 24430 13482
rect 24458 13454 24463 13482
rect 3369 13398 3374 13426
rect 3402 13398 3822 13426
rect 3850 13398 3855 13426
rect 11209 13398 11214 13426
rect 11242 13398 11550 13426
rect 11578 13398 11583 13426
rect 12665 13398 12670 13426
rect 12698 13398 13118 13426
rect 13146 13398 13151 13426
rect 24481 13398 24486 13426
rect 24514 13398 24519 13426
rect 4577 13314 4582 13342
rect 4610 13314 4634 13342
rect 4662 13314 4686 13342
rect 4714 13314 4738 13342
rect 4766 13314 4790 13342
rect 4818 13314 4842 13342
rect 4870 13314 4894 13342
rect 4922 13314 4946 13342
rect 4974 13314 4998 13342
rect 5026 13314 5031 13342
rect 9577 13314 9582 13342
rect 9610 13314 9634 13342
rect 9662 13314 9686 13342
rect 9714 13314 9738 13342
rect 9766 13314 9790 13342
rect 9818 13314 9842 13342
rect 9870 13314 9894 13342
rect 9922 13314 9946 13342
rect 9974 13314 9998 13342
rect 10026 13314 10031 13342
rect 14577 13314 14582 13342
rect 14610 13314 14634 13342
rect 14662 13314 14686 13342
rect 14714 13314 14738 13342
rect 14766 13314 14790 13342
rect 14818 13314 14842 13342
rect 14870 13314 14894 13342
rect 14922 13314 14946 13342
rect 14974 13314 14998 13342
rect 15026 13314 15031 13342
rect 19577 13314 19582 13342
rect 19610 13314 19634 13342
rect 19662 13314 19686 13342
rect 19714 13314 19738 13342
rect 19766 13314 19790 13342
rect 19818 13314 19842 13342
rect 19870 13314 19894 13342
rect 19922 13314 19946 13342
rect 19974 13314 19998 13342
rect 20026 13314 20031 13342
rect 24486 13314 24514 13398
rect 24577 13314 24582 13342
rect 24610 13314 24634 13342
rect 24662 13314 24686 13342
rect 24714 13314 24738 13342
rect 24766 13314 24790 13342
rect 24818 13314 24842 13342
rect 24870 13314 24894 13342
rect 24922 13314 24946 13342
rect 24974 13314 24998 13342
rect 25026 13314 25031 13342
rect 29577 13314 29582 13342
rect 29610 13314 29634 13342
rect 29662 13314 29686 13342
rect 29714 13314 29738 13342
rect 29766 13314 29790 13342
rect 29818 13314 29842 13342
rect 29870 13314 29894 13342
rect 29922 13314 29946 13342
rect 29974 13314 29998 13342
rect 30026 13314 30031 13342
rect 34577 13314 34582 13342
rect 34610 13314 34634 13342
rect 34662 13314 34686 13342
rect 34714 13314 34738 13342
rect 34766 13314 34790 13342
rect 34818 13314 34842 13342
rect 34870 13314 34894 13342
rect 34922 13314 34946 13342
rect 34974 13314 34998 13342
rect 35026 13314 35031 13342
rect 24425 13286 24430 13314
rect 24458 13286 24514 13314
rect 1969 13118 1974 13146
rect 2002 13118 2366 13146
rect 2394 13118 2399 13146
rect 2753 13118 2758 13146
rect 2786 13118 3318 13146
rect 3346 13118 3351 13146
rect 12945 13118 12950 13146
rect 12978 13118 13398 13146
rect 13426 13118 14014 13146
rect 14042 13118 15302 13146
rect 15330 13118 15335 13146
rect 16977 13118 16982 13146
rect 17010 13118 17094 13146
rect 17122 13118 18550 13146
rect 18578 13118 18583 13146
rect 2077 12922 2082 12950
rect 2110 12922 2134 12950
rect 2162 12922 2186 12950
rect 2214 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2394 12950
rect 2422 12922 2446 12950
rect 2474 12922 2498 12950
rect 2526 12922 2531 12950
rect 7077 12922 7082 12950
rect 7110 12922 7134 12950
rect 7162 12922 7186 12950
rect 7214 12922 7238 12950
rect 7266 12922 7290 12950
rect 7318 12922 7342 12950
rect 7370 12922 7394 12950
rect 7422 12922 7446 12950
rect 7474 12922 7498 12950
rect 7526 12922 7531 12950
rect 12077 12922 12082 12950
rect 12110 12922 12134 12950
rect 12162 12922 12186 12950
rect 12214 12922 12238 12950
rect 12266 12922 12290 12950
rect 12318 12922 12342 12950
rect 12370 12922 12394 12950
rect 12422 12922 12446 12950
rect 12474 12922 12498 12950
rect 12526 12922 12531 12950
rect 17077 12922 17082 12950
rect 17110 12922 17134 12950
rect 17162 12922 17186 12950
rect 17214 12922 17238 12950
rect 17266 12922 17290 12950
rect 17318 12922 17342 12950
rect 17370 12922 17394 12950
rect 17422 12922 17446 12950
rect 17474 12922 17498 12950
rect 17526 12922 17531 12950
rect 22077 12922 22082 12950
rect 22110 12922 22134 12950
rect 22162 12922 22186 12950
rect 22214 12922 22238 12950
rect 22266 12922 22290 12950
rect 22318 12922 22342 12950
rect 22370 12922 22394 12950
rect 22422 12922 22446 12950
rect 22474 12922 22498 12950
rect 22526 12922 22531 12950
rect 27077 12922 27082 12950
rect 27110 12922 27134 12950
rect 27162 12922 27186 12950
rect 27214 12922 27238 12950
rect 27266 12922 27290 12950
rect 27318 12922 27342 12950
rect 27370 12922 27394 12950
rect 27422 12922 27446 12950
rect 27474 12922 27498 12950
rect 27526 12922 27531 12950
rect 32077 12922 32082 12950
rect 32110 12922 32134 12950
rect 32162 12922 32186 12950
rect 32214 12922 32238 12950
rect 32266 12922 32290 12950
rect 32318 12922 32342 12950
rect 32370 12922 32394 12950
rect 32422 12922 32446 12950
rect 32474 12922 32498 12950
rect 32526 12922 32531 12950
rect 37077 12922 37082 12950
rect 37110 12922 37134 12950
rect 37162 12922 37186 12950
rect 37214 12922 37238 12950
rect 37266 12922 37290 12950
rect 37318 12922 37342 12950
rect 37370 12922 37394 12950
rect 37422 12922 37446 12950
rect 37474 12922 37498 12950
rect 37526 12922 37531 12950
rect 2193 12670 2198 12698
rect 2226 12670 2758 12698
rect 2786 12670 2791 12698
rect 23865 12670 23870 12698
rect 23898 12670 25158 12698
rect 25186 12670 25191 12698
rect 2641 12614 2646 12642
rect 2674 12614 4354 12642
rect 18545 12614 18550 12642
rect 18578 12614 19054 12642
rect 19082 12614 19087 12642
rect 4326 12586 4354 12614
rect 4321 12558 4326 12586
rect 4354 12558 4359 12586
rect 4577 12530 4582 12558
rect 4610 12530 4634 12558
rect 4662 12530 4686 12558
rect 4714 12530 4738 12558
rect 4766 12530 4790 12558
rect 4818 12530 4842 12558
rect 4870 12530 4894 12558
rect 4922 12530 4946 12558
rect 4974 12530 4998 12558
rect 5026 12530 5031 12558
rect 9577 12530 9582 12558
rect 9610 12530 9634 12558
rect 9662 12530 9686 12558
rect 9714 12530 9738 12558
rect 9766 12530 9790 12558
rect 9818 12530 9842 12558
rect 9870 12530 9894 12558
rect 9922 12530 9946 12558
rect 9974 12530 9998 12558
rect 10026 12530 10031 12558
rect 14577 12530 14582 12558
rect 14610 12530 14634 12558
rect 14662 12530 14686 12558
rect 14714 12530 14738 12558
rect 14766 12530 14790 12558
rect 14818 12530 14842 12558
rect 14870 12530 14894 12558
rect 14922 12530 14946 12558
rect 14974 12530 14998 12558
rect 15026 12530 15031 12558
rect 19577 12530 19582 12558
rect 19610 12530 19634 12558
rect 19662 12530 19686 12558
rect 19714 12530 19738 12558
rect 19766 12530 19790 12558
rect 19818 12530 19842 12558
rect 19870 12530 19894 12558
rect 19922 12530 19946 12558
rect 19974 12530 19998 12558
rect 20026 12530 20031 12558
rect 24577 12530 24582 12558
rect 24610 12530 24634 12558
rect 24662 12530 24686 12558
rect 24714 12530 24738 12558
rect 24766 12530 24790 12558
rect 24818 12530 24842 12558
rect 24870 12530 24894 12558
rect 24922 12530 24946 12558
rect 24974 12530 24998 12558
rect 25026 12530 25031 12558
rect 29577 12530 29582 12558
rect 29610 12530 29634 12558
rect 29662 12530 29686 12558
rect 29714 12530 29738 12558
rect 29766 12530 29790 12558
rect 29818 12530 29842 12558
rect 29870 12530 29894 12558
rect 29922 12530 29946 12558
rect 29974 12530 29998 12558
rect 30026 12530 30031 12558
rect 34577 12530 34582 12558
rect 34610 12530 34634 12558
rect 34662 12530 34686 12558
rect 34714 12530 34738 12558
rect 34766 12530 34790 12558
rect 34818 12530 34842 12558
rect 34870 12530 34894 12558
rect 34922 12530 34946 12558
rect 34974 12530 34998 12558
rect 35026 12530 35031 12558
rect 14233 12390 14238 12418
rect 14266 12390 14406 12418
rect 14434 12390 14439 12418
rect 25937 12390 25942 12418
rect 25970 12390 27426 12418
rect 27398 12362 27426 12390
rect 3033 12334 3038 12362
rect 3066 12334 3598 12362
rect 3626 12334 4102 12362
rect 4130 12334 4135 12362
rect 20953 12334 20958 12362
rect 20986 12334 22526 12362
rect 22554 12334 22559 12362
rect 24369 12334 24374 12362
rect 24402 12334 24486 12362
rect 24514 12334 24766 12362
rect 24794 12334 25102 12362
rect 25130 12334 26502 12362
rect 26530 12334 26535 12362
rect 27393 12334 27398 12362
rect 27426 12334 27678 12362
rect 27706 12334 27711 12362
rect 30193 12334 30198 12362
rect 30226 12334 30366 12362
rect 30394 12334 30702 12362
rect 30730 12334 30735 12362
rect 21793 12222 21798 12250
rect 21826 12222 23422 12250
rect 23450 12222 25214 12250
rect 25242 12222 25942 12250
rect 25970 12222 25975 12250
rect 2077 12138 2082 12166
rect 2110 12138 2134 12166
rect 2162 12138 2186 12166
rect 2214 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2394 12166
rect 2422 12138 2446 12166
rect 2474 12138 2498 12166
rect 2526 12138 2531 12166
rect 7077 12138 7082 12166
rect 7110 12138 7134 12166
rect 7162 12138 7186 12166
rect 7214 12138 7238 12166
rect 7266 12138 7290 12166
rect 7318 12138 7342 12166
rect 7370 12138 7394 12166
rect 7422 12138 7446 12166
rect 7474 12138 7498 12166
rect 7526 12138 7531 12166
rect 12077 12138 12082 12166
rect 12110 12138 12134 12166
rect 12162 12138 12186 12166
rect 12214 12138 12238 12166
rect 12266 12138 12290 12166
rect 12318 12138 12342 12166
rect 12370 12138 12394 12166
rect 12422 12138 12446 12166
rect 12474 12138 12498 12166
rect 12526 12138 12531 12166
rect 17077 12138 17082 12166
rect 17110 12138 17134 12166
rect 17162 12138 17186 12166
rect 17214 12138 17238 12166
rect 17266 12138 17290 12166
rect 17318 12138 17342 12166
rect 17370 12138 17394 12166
rect 17422 12138 17446 12166
rect 17474 12138 17498 12166
rect 17526 12138 17531 12166
rect 22077 12138 22082 12166
rect 22110 12138 22134 12166
rect 22162 12138 22186 12166
rect 22214 12138 22238 12166
rect 22266 12138 22290 12166
rect 22318 12138 22342 12166
rect 22370 12138 22394 12166
rect 22422 12138 22446 12166
rect 22474 12138 22498 12166
rect 22526 12138 22531 12166
rect 27077 12138 27082 12166
rect 27110 12138 27134 12166
rect 27162 12138 27186 12166
rect 27214 12138 27238 12166
rect 27266 12138 27290 12166
rect 27318 12138 27342 12166
rect 27370 12138 27394 12166
rect 27422 12138 27446 12166
rect 27474 12138 27498 12166
rect 27526 12138 27531 12166
rect 32077 12138 32082 12166
rect 32110 12138 32134 12166
rect 32162 12138 32186 12166
rect 32214 12138 32238 12166
rect 32266 12138 32290 12166
rect 32318 12138 32342 12166
rect 32370 12138 32394 12166
rect 32422 12138 32446 12166
rect 32474 12138 32498 12166
rect 32526 12138 32531 12166
rect 37077 12138 37082 12166
rect 37110 12138 37134 12166
rect 37162 12138 37186 12166
rect 37214 12138 37238 12166
rect 37266 12138 37290 12166
rect 37318 12138 37342 12166
rect 37370 12138 37394 12166
rect 37422 12138 37446 12166
rect 37474 12138 37498 12166
rect 37526 12138 37531 12166
rect 4097 11942 4102 11970
rect 4130 11942 5278 11970
rect 5306 11942 5311 11970
rect 8465 11942 8470 11970
rect 8498 11942 10430 11970
rect 10458 11942 10463 11970
rect 17425 11942 17430 11970
rect 17458 11942 17598 11970
rect 17626 11942 17990 11970
rect 18018 11942 18023 11970
rect 22577 11942 22582 11970
rect 22610 11942 23030 11970
rect 23058 11942 25102 11970
rect 25130 11942 25135 11970
rect 27673 11942 27678 11970
rect 27706 11942 32830 11970
rect 32858 11942 33110 11970
rect 33138 11942 33143 11970
rect 19497 11886 19502 11914
rect 19530 11886 19950 11914
rect 19978 11886 21350 11914
rect 21378 11886 21383 11914
rect 28569 11886 28574 11914
rect 28602 11886 29358 11914
rect 29386 11886 29918 11914
rect 29946 11886 29951 11914
rect 6393 11774 6398 11802
rect 6426 11774 7014 11802
rect 7042 11774 8358 11802
rect 8386 11774 8391 11802
rect 11993 11774 11998 11802
rect 12026 11774 13342 11802
rect 13370 11774 13375 11802
rect 4577 11746 4582 11774
rect 4610 11746 4634 11774
rect 4662 11746 4686 11774
rect 4714 11746 4738 11774
rect 4766 11746 4790 11774
rect 4818 11746 4842 11774
rect 4870 11746 4894 11774
rect 4922 11746 4946 11774
rect 4974 11746 4998 11774
rect 5026 11746 5031 11774
rect 9577 11746 9582 11774
rect 9610 11746 9634 11774
rect 9662 11746 9686 11774
rect 9714 11746 9738 11774
rect 9766 11746 9790 11774
rect 9818 11746 9842 11774
rect 9870 11746 9894 11774
rect 9922 11746 9946 11774
rect 9974 11746 9998 11774
rect 10026 11746 10031 11774
rect 14577 11746 14582 11774
rect 14610 11746 14634 11774
rect 14662 11746 14686 11774
rect 14714 11746 14738 11774
rect 14766 11746 14790 11774
rect 14818 11746 14842 11774
rect 14870 11746 14894 11774
rect 14922 11746 14946 11774
rect 14974 11746 14998 11774
rect 15026 11746 15031 11774
rect 19577 11746 19582 11774
rect 19610 11746 19634 11774
rect 19662 11746 19686 11774
rect 19714 11746 19738 11774
rect 19766 11746 19790 11774
rect 19818 11746 19842 11774
rect 19870 11746 19894 11774
rect 19922 11746 19946 11774
rect 19974 11746 19998 11774
rect 20026 11746 20031 11774
rect 24577 11746 24582 11774
rect 24610 11746 24634 11774
rect 24662 11746 24686 11774
rect 24714 11746 24738 11774
rect 24766 11746 24790 11774
rect 24818 11746 24842 11774
rect 24870 11746 24894 11774
rect 24922 11746 24946 11774
rect 24974 11746 24998 11774
rect 25026 11746 25031 11774
rect 29577 11746 29582 11774
rect 29610 11746 29634 11774
rect 29662 11746 29686 11774
rect 29714 11746 29738 11774
rect 29766 11746 29790 11774
rect 29818 11746 29842 11774
rect 29870 11746 29894 11774
rect 29922 11746 29946 11774
rect 29974 11746 29998 11774
rect 30026 11746 30031 11774
rect 34577 11746 34582 11774
rect 34610 11746 34634 11774
rect 34662 11746 34686 11774
rect 34714 11746 34738 11774
rect 34766 11746 34790 11774
rect 34818 11746 34842 11774
rect 34870 11746 34894 11774
rect 34922 11746 34946 11774
rect 34974 11746 34998 11774
rect 35026 11746 35031 11774
rect 15073 11718 15078 11746
rect 15106 11718 16534 11746
rect 16562 11718 16567 11746
rect 31481 11606 31486 11634
rect 31514 11606 31934 11634
rect 31962 11606 31967 11634
rect 25153 11550 25158 11578
rect 25186 11550 25214 11578
rect 25242 11550 25438 11578
rect 25466 11550 25471 11578
rect 28345 11550 28350 11578
rect 28378 11550 29414 11578
rect 29442 11550 29447 11578
rect 32433 11550 32438 11578
rect 32466 11550 32774 11578
rect 32802 11550 32807 11578
rect 33161 11550 33166 11578
rect 33194 11550 33614 11578
rect 33642 11550 34510 11578
rect 34538 11550 34543 11578
rect 2077 11354 2082 11382
rect 2110 11354 2134 11382
rect 2162 11354 2186 11382
rect 2214 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2394 11382
rect 2422 11354 2446 11382
rect 2474 11354 2498 11382
rect 2526 11354 2531 11382
rect 7077 11354 7082 11382
rect 7110 11354 7134 11382
rect 7162 11354 7186 11382
rect 7214 11354 7238 11382
rect 7266 11354 7290 11382
rect 7318 11354 7342 11382
rect 7370 11354 7394 11382
rect 7422 11354 7446 11382
rect 7474 11354 7498 11382
rect 7526 11354 7531 11382
rect 12077 11354 12082 11382
rect 12110 11354 12134 11382
rect 12162 11354 12186 11382
rect 12214 11354 12238 11382
rect 12266 11354 12290 11382
rect 12318 11354 12342 11382
rect 12370 11354 12394 11382
rect 12422 11354 12446 11382
rect 12474 11354 12498 11382
rect 12526 11354 12531 11382
rect 17077 11354 17082 11382
rect 17110 11354 17134 11382
rect 17162 11354 17186 11382
rect 17214 11354 17238 11382
rect 17266 11354 17290 11382
rect 17318 11354 17342 11382
rect 17370 11354 17394 11382
rect 17422 11354 17446 11382
rect 17474 11354 17498 11382
rect 17526 11354 17531 11382
rect 22077 11354 22082 11382
rect 22110 11354 22134 11382
rect 22162 11354 22186 11382
rect 22214 11354 22238 11382
rect 22266 11354 22290 11382
rect 22318 11354 22342 11382
rect 22370 11354 22394 11382
rect 22422 11354 22446 11382
rect 22474 11354 22498 11382
rect 22526 11354 22531 11382
rect 27077 11354 27082 11382
rect 27110 11354 27134 11382
rect 27162 11354 27186 11382
rect 27214 11354 27238 11382
rect 27266 11354 27290 11382
rect 27318 11354 27342 11382
rect 27370 11354 27394 11382
rect 27422 11354 27446 11382
rect 27474 11354 27498 11382
rect 27526 11354 27531 11382
rect 32077 11354 32082 11382
rect 32110 11354 32134 11382
rect 32162 11354 32186 11382
rect 32214 11354 32238 11382
rect 32266 11354 32290 11382
rect 32318 11354 32342 11382
rect 32370 11354 32394 11382
rect 32422 11354 32446 11382
rect 32474 11354 32498 11382
rect 32526 11354 32531 11382
rect 37077 11354 37082 11382
rect 37110 11354 37134 11382
rect 37162 11354 37186 11382
rect 37214 11354 37238 11382
rect 37266 11354 37290 11382
rect 37318 11354 37342 11382
rect 37370 11354 37394 11382
rect 37422 11354 37446 11382
rect 37474 11354 37498 11382
rect 37526 11354 37531 11382
rect 18825 11214 18830 11242
rect 18858 11214 19222 11242
rect 19250 11214 19334 11242
rect 19362 11214 19950 11242
rect 19978 11214 19983 11242
rect 34505 11214 34510 11242
rect 34538 11214 35126 11242
rect 35154 11214 35350 11242
rect 35378 11214 35383 11242
rect 19049 11158 19054 11186
rect 19082 11158 20230 11186
rect 20258 11158 20790 11186
rect 20818 11158 20823 11186
rect 21849 11158 21854 11186
rect 21882 11158 25158 11186
rect 25186 11158 25191 11186
rect 32433 11158 32438 11186
rect 32466 11158 32774 11186
rect 32802 11158 32807 11186
rect 34953 11158 34958 11186
rect 34986 11158 36134 11186
rect 36162 11158 36167 11186
rect 14289 11046 14294 11074
rect 14322 11046 14462 11074
rect 14490 11046 15862 11074
rect 15890 11046 15895 11074
rect 19945 11046 19950 11074
rect 19978 11046 21294 11074
rect 21322 11046 21327 11074
rect 4577 10962 4582 10990
rect 4610 10962 4634 10990
rect 4662 10962 4686 10990
rect 4714 10962 4738 10990
rect 4766 10962 4790 10990
rect 4818 10962 4842 10990
rect 4870 10962 4894 10990
rect 4922 10962 4946 10990
rect 4974 10962 4998 10990
rect 5026 10962 5031 10990
rect 9577 10962 9582 10990
rect 9610 10962 9634 10990
rect 9662 10962 9686 10990
rect 9714 10962 9738 10990
rect 9766 10962 9790 10990
rect 9818 10962 9842 10990
rect 9870 10962 9894 10990
rect 9922 10962 9946 10990
rect 9974 10962 9998 10990
rect 10026 10962 10031 10990
rect 14577 10962 14582 10990
rect 14610 10962 14634 10990
rect 14662 10962 14686 10990
rect 14714 10962 14738 10990
rect 14766 10962 14790 10990
rect 14818 10962 14842 10990
rect 14870 10962 14894 10990
rect 14922 10962 14946 10990
rect 14974 10962 14998 10990
rect 15026 10962 15031 10990
rect 19577 10962 19582 10990
rect 19610 10962 19634 10990
rect 19662 10962 19686 10990
rect 19714 10962 19738 10990
rect 19766 10962 19790 10990
rect 19818 10962 19842 10990
rect 19870 10962 19894 10990
rect 19922 10962 19946 10990
rect 19974 10962 19998 10990
rect 20026 10962 20031 10990
rect 24577 10962 24582 10990
rect 24610 10962 24634 10990
rect 24662 10962 24686 10990
rect 24714 10962 24738 10990
rect 24766 10962 24790 10990
rect 24818 10962 24842 10990
rect 24870 10962 24894 10990
rect 24922 10962 24946 10990
rect 24974 10962 24998 10990
rect 25026 10962 25031 10990
rect 29577 10962 29582 10990
rect 29610 10962 29634 10990
rect 29662 10962 29686 10990
rect 29714 10962 29738 10990
rect 29766 10962 29790 10990
rect 29818 10962 29842 10990
rect 29870 10962 29894 10990
rect 29922 10962 29946 10990
rect 29974 10962 29998 10990
rect 30026 10962 30031 10990
rect 34577 10962 34582 10990
rect 34610 10962 34634 10990
rect 34662 10962 34686 10990
rect 34714 10962 34738 10990
rect 34766 10962 34790 10990
rect 34818 10962 34842 10990
rect 34870 10962 34894 10990
rect 34922 10962 34946 10990
rect 34974 10962 34998 10990
rect 35026 10962 35031 10990
rect 5833 10934 5838 10962
rect 5866 10934 7294 10962
rect 7322 10934 7574 10962
rect 7602 10934 9254 10962
rect 9282 10934 9287 10962
rect 2473 10878 2478 10906
rect 2506 10878 2590 10906
rect 2618 10878 3038 10906
rect 3066 10878 3071 10906
rect 28065 10878 28070 10906
rect 28098 10878 28350 10906
rect 28378 10878 28383 10906
rect 1857 10766 1862 10794
rect 1890 10766 2086 10794
rect 2114 10766 2119 10794
rect 5273 10766 5278 10794
rect 5306 10766 5838 10794
rect 5866 10766 5871 10794
rect 16921 10766 16926 10794
rect 16954 10766 17262 10794
rect 17290 10766 17486 10794
rect 17514 10766 18830 10794
rect 18858 10766 18863 10794
rect 20897 10766 20902 10794
rect 20930 10766 22526 10794
rect 22554 10766 23030 10794
rect 23058 10766 23063 10794
rect 5441 10710 5446 10738
rect 5474 10710 36694 10738
rect 36722 10710 36727 10738
rect 2077 10570 2082 10598
rect 2110 10570 2134 10598
rect 2162 10570 2186 10598
rect 2214 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2394 10598
rect 2422 10570 2446 10598
rect 2474 10570 2498 10598
rect 2526 10570 2531 10598
rect 7077 10570 7082 10598
rect 7110 10570 7134 10598
rect 7162 10570 7186 10598
rect 7214 10570 7238 10598
rect 7266 10570 7290 10598
rect 7318 10570 7342 10598
rect 7370 10570 7394 10598
rect 7422 10570 7446 10598
rect 7474 10570 7498 10598
rect 7526 10570 7531 10598
rect 12077 10570 12082 10598
rect 12110 10570 12134 10598
rect 12162 10570 12186 10598
rect 12214 10570 12238 10598
rect 12266 10570 12290 10598
rect 12318 10570 12342 10598
rect 12370 10570 12394 10598
rect 12422 10570 12446 10598
rect 12474 10570 12498 10598
rect 12526 10570 12531 10598
rect 17077 10570 17082 10598
rect 17110 10570 17134 10598
rect 17162 10570 17186 10598
rect 17214 10570 17238 10598
rect 17266 10570 17290 10598
rect 17318 10570 17342 10598
rect 17370 10570 17394 10598
rect 17422 10570 17446 10598
rect 17474 10570 17498 10598
rect 17526 10570 17531 10598
rect 22077 10570 22082 10598
rect 22110 10570 22134 10598
rect 22162 10570 22186 10598
rect 22214 10570 22238 10598
rect 22266 10570 22290 10598
rect 22318 10570 22342 10598
rect 22370 10570 22394 10598
rect 22422 10570 22446 10598
rect 22474 10570 22498 10598
rect 22526 10570 22531 10598
rect 27077 10570 27082 10598
rect 27110 10570 27134 10598
rect 27162 10570 27186 10598
rect 27214 10570 27238 10598
rect 27266 10570 27290 10598
rect 27318 10570 27342 10598
rect 27370 10570 27394 10598
rect 27422 10570 27446 10598
rect 27474 10570 27498 10598
rect 27526 10570 27531 10598
rect 32077 10570 32082 10598
rect 32110 10570 32134 10598
rect 32162 10570 32186 10598
rect 32214 10570 32238 10598
rect 32266 10570 32290 10598
rect 32318 10570 32342 10598
rect 32370 10570 32394 10598
rect 32422 10570 32446 10598
rect 32474 10570 32498 10598
rect 32526 10570 32531 10598
rect 37077 10570 37082 10598
rect 37110 10570 37134 10598
rect 37162 10570 37186 10598
rect 37214 10570 37238 10598
rect 37266 10570 37290 10598
rect 37318 10570 37342 10598
rect 37370 10570 37394 10598
rect 37422 10570 37446 10598
rect 37474 10570 37498 10598
rect 37526 10570 37531 10598
rect 3817 10374 3822 10402
rect 3850 10374 5278 10402
rect 5306 10374 5311 10402
rect 16809 10374 16814 10402
rect 16842 10374 16926 10402
rect 16954 10374 16959 10402
rect 27673 10374 27678 10402
rect 27706 10374 28070 10402
rect 28098 10374 28103 10402
rect 34449 10374 34454 10402
rect 34482 10374 34958 10402
rect 34986 10374 36246 10402
rect 36274 10374 36279 10402
rect 18209 10318 18214 10346
rect 18242 10318 24374 10346
rect 24402 10318 24407 10346
rect 35345 10318 35350 10346
rect 35378 10318 37310 10346
rect 37338 10318 37590 10346
rect 37618 10318 37623 10346
rect 23025 10262 23030 10290
rect 23058 10262 24430 10290
rect 24458 10262 24463 10290
rect 4577 10178 4582 10206
rect 4610 10178 4634 10206
rect 4662 10178 4686 10206
rect 4714 10178 4738 10206
rect 4766 10178 4790 10206
rect 4818 10178 4842 10206
rect 4870 10178 4894 10206
rect 4922 10178 4946 10206
rect 4974 10178 4998 10206
rect 5026 10178 5031 10206
rect 9577 10178 9582 10206
rect 9610 10178 9634 10206
rect 9662 10178 9686 10206
rect 9714 10178 9738 10206
rect 9766 10178 9790 10206
rect 9818 10178 9842 10206
rect 9870 10178 9894 10206
rect 9922 10178 9946 10206
rect 9974 10178 9998 10206
rect 10026 10178 10031 10206
rect 14577 10178 14582 10206
rect 14610 10178 14634 10206
rect 14662 10178 14686 10206
rect 14714 10178 14738 10206
rect 14766 10178 14790 10206
rect 14818 10178 14842 10206
rect 14870 10178 14894 10206
rect 14922 10178 14946 10206
rect 14974 10178 14998 10206
rect 15026 10178 15031 10206
rect 19577 10178 19582 10206
rect 19610 10178 19634 10206
rect 19662 10178 19686 10206
rect 19714 10178 19738 10206
rect 19766 10178 19790 10206
rect 19818 10178 19842 10206
rect 19870 10178 19894 10206
rect 19922 10178 19946 10206
rect 19974 10178 19998 10206
rect 20026 10178 20031 10206
rect 24577 10178 24582 10206
rect 24610 10178 24634 10206
rect 24662 10178 24686 10206
rect 24714 10178 24738 10206
rect 24766 10178 24790 10206
rect 24818 10178 24842 10206
rect 24870 10178 24894 10206
rect 24922 10178 24946 10206
rect 24974 10178 24998 10206
rect 25026 10178 25031 10206
rect 29577 10178 29582 10206
rect 29610 10178 29634 10206
rect 29662 10178 29686 10206
rect 29714 10178 29738 10206
rect 29766 10178 29790 10206
rect 29818 10178 29842 10206
rect 29870 10178 29894 10206
rect 29922 10178 29946 10206
rect 29974 10178 29998 10206
rect 30026 10178 30031 10206
rect 34577 10178 34582 10206
rect 34610 10178 34634 10206
rect 34662 10178 34686 10206
rect 34714 10178 34738 10206
rect 34766 10178 34790 10206
rect 34818 10178 34842 10206
rect 34870 10178 34894 10206
rect 34922 10178 34946 10206
rect 34974 10178 34998 10206
rect 35026 10178 35031 10206
rect 8801 10094 8806 10122
rect 8834 10094 34454 10122
rect 34482 10094 34487 10122
rect 11993 10038 11998 10066
rect 12026 10038 12502 10066
rect 12530 10038 12950 10066
rect 12978 10038 12983 10066
rect 15745 10038 15750 10066
rect 15778 10038 16758 10066
rect 16786 10038 16791 10066
rect 25937 10038 25942 10066
rect 25970 10038 27678 10066
rect 27706 10038 27902 10066
rect 27930 10038 28406 10066
rect 28434 10038 28439 10066
rect 29465 10038 29470 10066
rect 29498 10038 29806 10066
rect 29834 10038 30030 10066
rect 30058 10038 30063 10066
rect 30249 10038 30254 10066
rect 30282 10038 30758 10066
rect 30786 10038 32158 10066
rect 32186 10038 32830 10066
rect 32858 10038 32942 10066
rect 32970 10038 32975 10066
rect 7009 9982 7014 10010
rect 7042 9982 8750 10010
rect 8778 9982 8783 10010
rect 13337 9982 13342 10010
rect 13370 9982 13622 10010
rect 13650 9982 13655 10010
rect 20841 9982 20846 10010
rect 20874 9982 22246 10010
rect 22274 9982 22582 10010
rect 22610 9982 22615 10010
rect 23417 9982 23422 10010
rect 23450 9982 23870 10010
rect 23898 9982 23903 10010
rect 26833 9982 26838 10010
rect 26866 9982 27566 10010
rect 27594 9982 27958 10010
rect 27986 9982 27991 10010
rect 28345 9982 28350 10010
rect 28378 9982 28798 10010
rect 28826 9982 30310 10010
rect 30338 9982 30702 10010
rect 30730 9982 30814 10010
rect 30842 9982 30847 10010
rect 32881 9982 32886 10010
rect 32914 9982 34622 10010
rect 34650 9982 34846 10010
rect 34874 9982 35126 10010
rect 35154 9982 35159 10010
rect 4041 9926 4046 9954
rect 4074 9926 36414 9954
rect 36442 9926 36694 9954
rect 36722 9926 36727 9954
rect 30081 9870 30086 9898
rect 30114 9870 31094 9898
rect 31122 9870 31127 9898
rect 32769 9870 32774 9898
rect 32802 9870 34454 9898
rect 34482 9870 34487 9898
rect 2077 9786 2082 9814
rect 2110 9786 2134 9814
rect 2162 9786 2186 9814
rect 2214 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2394 9814
rect 2422 9786 2446 9814
rect 2474 9786 2498 9814
rect 2526 9786 2531 9814
rect 7077 9786 7082 9814
rect 7110 9786 7134 9814
rect 7162 9786 7186 9814
rect 7214 9786 7238 9814
rect 7266 9786 7290 9814
rect 7318 9786 7342 9814
rect 7370 9786 7394 9814
rect 7422 9786 7446 9814
rect 7474 9786 7498 9814
rect 7526 9786 7531 9814
rect 12077 9786 12082 9814
rect 12110 9786 12134 9814
rect 12162 9786 12186 9814
rect 12214 9786 12238 9814
rect 12266 9786 12290 9814
rect 12318 9786 12342 9814
rect 12370 9786 12394 9814
rect 12422 9786 12446 9814
rect 12474 9786 12498 9814
rect 12526 9786 12531 9814
rect 17077 9786 17082 9814
rect 17110 9786 17134 9814
rect 17162 9786 17186 9814
rect 17214 9786 17238 9814
rect 17266 9786 17290 9814
rect 17318 9786 17342 9814
rect 17370 9786 17394 9814
rect 17422 9786 17446 9814
rect 17474 9786 17498 9814
rect 17526 9786 17531 9814
rect 22077 9786 22082 9814
rect 22110 9786 22134 9814
rect 22162 9786 22186 9814
rect 22214 9786 22238 9814
rect 22266 9786 22290 9814
rect 22318 9786 22342 9814
rect 22370 9786 22394 9814
rect 22422 9786 22446 9814
rect 22474 9786 22498 9814
rect 22526 9786 22531 9814
rect 27077 9786 27082 9814
rect 27110 9786 27134 9814
rect 27162 9786 27186 9814
rect 27214 9786 27238 9814
rect 27266 9786 27290 9814
rect 27318 9786 27342 9814
rect 27370 9786 27394 9814
rect 27422 9786 27446 9814
rect 27474 9786 27498 9814
rect 27526 9786 27531 9814
rect 32077 9786 32082 9814
rect 32110 9786 32134 9814
rect 32162 9786 32186 9814
rect 32214 9786 32238 9814
rect 32266 9786 32290 9814
rect 32318 9786 32342 9814
rect 32370 9786 32394 9814
rect 32422 9786 32446 9814
rect 32474 9786 32498 9814
rect 32526 9786 32531 9814
rect 37077 9786 37082 9814
rect 37110 9786 37134 9814
rect 37162 9786 37186 9814
rect 37214 9786 37238 9814
rect 37266 9786 37290 9814
rect 37318 9786 37342 9814
rect 37370 9786 37394 9814
rect 37422 9786 37446 9814
rect 37474 9786 37498 9814
rect 37526 9786 37531 9814
rect 30809 9702 30814 9730
rect 30842 9702 31990 9730
rect 32018 9702 32158 9730
rect 32186 9702 32191 9730
rect 3817 9590 3822 9618
rect 3850 9590 5950 9618
rect 5978 9590 6230 9618
rect 6258 9590 6263 9618
rect 14457 9590 14462 9618
rect 14490 9590 14798 9618
rect 14826 9590 15078 9618
rect 15106 9590 15111 9618
rect 15745 9590 15750 9618
rect 15778 9590 15862 9618
rect 15890 9590 16814 9618
rect 16842 9590 16847 9618
rect 31369 9590 31374 9618
rect 31402 9590 32830 9618
rect 32858 9590 33110 9618
rect 33138 9590 33143 9618
rect 35345 9590 35350 9618
rect 35378 9590 36974 9618
rect 36946 9562 36974 9590
rect 23865 9534 23870 9562
rect 23898 9534 25382 9562
rect 25410 9534 25415 9562
rect 36946 9534 37310 9562
rect 37338 9534 37646 9562
rect 37674 9534 37679 9562
rect 34449 9478 34454 9506
rect 34482 9478 34958 9506
rect 34986 9478 36414 9506
rect 36442 9478 36447 9506
rect 32937 9422 32942 9450
rect 32970 9422 34174 9450
rect 34202 9422 34207 9450
rect 4577 9394 4582 9422
rect 4610 9394 4634 9422
rect 4662 9394 4686 9422
rect 4714 9394 4738 9422
rect 4766 9394 4790 9422
rect 4818 9394 4842 9422
rect 4870 9394 4894 9422
rect 4922 9394 4946 9422
rect 4974 9394 4998 9422
rect 5026 9394 5031 9422
rect 9577 9394 9582 9422
rect 9610 9394 9634 9422
rect 9662 9394 9686 9422
rect 9714 9394 9738 9422
rect 9766 9394 9790 9422
rect 9818 9394 9842 9422
rect 9870 9394 9894 9422
rect 9922 9394 9946 9422
rect 9974 9394 9998 9422
rect 10026 9394 10031 9422
rect 14577 9394 14582 9422
rect 14610 9394 14634 9422
rect 14662 9394 14686 9422
rect 14714 9394 14738 9422
rect 14766 9394 14790 9422
rect 14818 9394 14842 9422
rect 14870 9394 14894 9422
rect 14922 9394 14946 9422
rect 14974 9394 14998 9422
rect 15026 9394 15031 9422
rect 19577 9394 19582 9422
rect 19610 9394 19634 9422
rect 19662 9394 19686 9422
rect 19714 9394 19738 9422
rect 19766 9394 19790 9422
rect 19818 9394 19842 9422
rect 19870 9394 19894 9422
rect 19922 9394 19946 9422
rect 19974 9394 19998 9422
rect 20026 9394 20031 9422
rect 24577 9394 24582 9422
rect 24610 9394 24634 9422
rect 24662 9394 24686 9422
rect 24714 9394 24738 9422
rect 24766 9394 24790 9422
rect 24818 9394 24842 9422
rect 24870 9394 24894 9422
rect 24922 9394 24946 9422
rect 24974 9394 24998 9422
rect 25026 9394 25031 9422
rect 29577 9394 29582 9422
rect 29610 9394 29634 9422
rect 29662 9394 29686 9422
rect 29714 9394 29738 9422
rect 29766 9394 29790 9422
rect 29818 9394 29842 9422
rect 29870 9394 29894 9422
rect 29922 9394 29946 9422
rect 29974 9394 29998 9422
rect 30026 9394 30031 9422
rect 34577 9394 34582 9422
rect 34610 9394 34634 9422
rect 34662 9394 34686 9422
rect 34714 9394 34738 9422
rect 34766 9394 34790 9422
rect 34818 9394 34842 9422
rect 34870 9394 34894 9422
rect 34922 9394 34946 9422
rect 34974 9394 34998 9422
rect 35026 9394 35031 9422
rect 1913 9310 1918 9338
rect 1946 9310 2478 9338
rect 2506 9310 2511 9338
rect 14009 9310 14014 9338
rect 14042 9310 15134 9338
rect 15162 9310 15167 9338
rect 2025 9254 2030 9282
rect 2058 9254 3374 9282
rect 3402 9254 3822 9282
rect 3850 9254 3855 9282
rect 10537 9254 10542 9282
rect 10570 9254 11774 9282
rect 11802 9254 11942 9282
rect 11970 9254 11975 9282
rect 13337 9254 13342 9282
rect 13370 9254 14462 9282
rect 14490 9254 14495 9282
rect 17985 9254 17990 9282
rect 18018 9254 19278 9282
rect 19306 9254 19311 9282
rect 34169 9254 34174 9282
rect 34202 9254 34678 9282
rect 34706 9254 34711 9282
rect 1633 9198 1638 9226
rect 1666 9198 1862 9226
rect 1890 9198 1895 9226
rect 4489 9198 4494 9226
rect 4522 9198 5110 9226
rect 5138 9198 5143 9226
rect 10313 9198 10318 9226
rect 10346 9198 10486 9226
rect 10514 9198 10519 9226
rect 29409 9198 29414 9226
rect 29442 9198 29526 9226
rect 29554 9198 30982 9226
rect 31010 9198 31015 9226
rect 27953 9142 27958 9170
rect 27986 9142 32830 9170
rect 32858 9142 36190 9170
rect 36218 9142 36223 9170
rect 2077 9002 2082 9030
rect 2110 9002 2134 9030
rect 2162 9002 2186 9030
rect 2214 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2394 9030
rect 2422 9002 2446 9030
rect 2474 9002 2498 9030
rect 2526 9002 2531 9030
rect 7077 9002 7082 9030
rect 7110 9002 7134 9030
rect 7162 9002 7186 9030
rect 7214 9002 7238 9030
rect 7266 9002 7290 9030
rect 7318 9002 7342 9030
rect 7370 9002 7394 9030
rect 7422 9002 7446 9030
rect 7474 9002 7498 9030
rect 7526 9002 7531 9030
rect 12077 9002 12082 9030
rect 12110 9002 12134 9030
rect 12162 9002 12186 9030
rect 12214 9002 12238 9030
rect 12266 9002 12290 9030
rect 12318 9002 12342 9030
rect 12370 9002 12394 9030
rect 12422 9002 12446 9030
rect 12474 9002 12498 9030
rect 12526 9002 12531 9030
rect 17077 9002 17082 9030
rect 17110 9002 17134 9030
rect 17162 9002 17186 9030
rect 17214 9002 17238 9030
rect 17266 9002 17290 9030
rect 17318 9002 17342 9030
rect 17370 9002 17394 9030
rect 17422 9002 17446 9030
rect 17474 9002 17498 9030
rect 17526 9002 17531 9030
rect 22077 9002 22082 9030
rect 22110 9002 22134 9030
rect 22162 9002 22186 9030
rect 22214 9002 22238 9030
rect 22266 9002 22290 9030
rect 22318 9002 22342 9030
rect 22370 9002 22394 9030
rect 22422 9002 22446 9030
rect 22474 9002 22498 9030
rect 22526 9002 22531 9030
rect 27077 9002 27082 9030
rect 27110 9002 27134 9030
rect 27162 9002 27186 9030
rect 27214 9002 27238 9030
rect 27266 9002 27290 9030
rect 27318 9002 27342 9030
rect 27370 9002 27394 9030
rect 27422 9002 27446 9030
rect 27474 9002 27498 9030
rect 27526 9002 27531 9030
rect 32077 9002 32082 9030
rect 32110 9002 32134 9030
rect 32162 9002 32186 9030
rect 32214 9002 32238 9030
rect 32266 9002 32290 9030
rect 32318 9002 32342 9030
rect 32370 9002 32394 9030
rect 32422 9002 32446 9030
rect 32474 9002 32498 9030
rect 32526 9002 32531 9030
rect 37077 9002 37082 9030
rect 37110 9002 37134 9030
rect 37162 9002 37186 9030
rect 37214 9002 37238 9030
rect 37266 9002 37290 9030
rect 37318 9002 37342 9030
rect 37370 9002 37394 9030
rect 37422 9002 37446 9030
rect 37474 9002 37498 9030
rect 37526 9002 37531 9030
rect 23417 8862 23422 8890
rect 23450 8862 23870 8890
rect 23898 8862 25214 8890
rect 25242 8862 27566 8890
rect 27594 8862 32886 8890
rect 32914 8862 32919 8890
rect 4993 8806 4998 8834
rect 5026 8806 5110 8834
rect 5138 8806 5558 8834
rect 5586 8806 5894 8834
rect 5922 8806 5927 8834
rect 28849 8806 28854 8834
rect 28882 8806 29414 8834
rect 29442 8806 29447 8834
rect 30193 8806 30198 8834
rect 30226 8806 31150 8834
rect 31178 8806 31374 8834
rect 31402 8806 31407 8834
rect 32825 8750 32830 8778
rect 32858 8750 33110 8778
rect 33138 8750 33143 8778
rect 35849 8750 35854 8778
rect 35882 8750 36974 8778
rect 37002 8750 37007 8778
rect 4577 8610 4582 8638
rect 4610 8610 4634 8638
rect 4662 8610 4686 8638
rect 4714 8610 4738 8638
rect 4766 8610 4790 8638
rect 4818 8610 4842 8638
rect 4870 8610 4894 8638
rect 4922 8610 4946 8638
rect 4974 8610 4998 8638
rect 5026 8610 5031 8638
rect 9577 8610 9582 8638
rect 9610 8610 9634 8638
rect 9662 8610 9686 8638
rect 9714 8610 9738 8638
rect 9766 8610 9790 8638
rect 9818 8610 9842 8638
rect 9870 8610 9894 8638
rect 9922 8610 9946 8638
rect 9974 8610 9998 8638
rect 10026 8610 10031 8638
rect 14577 8610 14582 8638
rect 14610 8610 14634 8638
rect 14662 8610 14686 8638
rect 14714 8610 14738 8638
rect 14766 8610 14790 8638
rect 14818 8610 14842 8638
rect 14870 8610 14894 8638
rect 14922 8610 14946 8638
rect 14974 8610 14998 8638
rect 15026 8610 15031 8638
rect 19577 8610 19582 8638
rect 19610 8610 19634 8638
rect 19662 8610 19686 8638
rect 19714 8610 19738 8638
rect 19766 8610 19790 8638
rect 19818 8610 19842 8638
rect 19870 8610 19894 8638
rect 19922 8610 19946 8638
rect 19974 8610 19998 8638
rect 20026 8610 20031 8638
rect 24577 8610 24582 8638
rect 24610 8610 24634 8638
rect 24662 8610 24686 8638
rect 24714 8610 24738 8638
rect 24766 8610 24790 8638
rect 24818 8610 24842 8638
rect 24870 8610 24894 8638
rect 24922 8610 24946 8638
rect 24974 8610 24998 8638
rect 25026 8610 25031 8638
rect 29577 8610 29582 8638
rect 29610 8610 29634 8638
rect 29662 8610 29686 8638
rect 29714 8610 29738 8638
rect 29766 8610 29790 8638
rect 29818 8610 29842 8638
rect 29870 8610 29894 8638
rect 29922 8610 29946 8638
rect 29974 8610 29998 8638
rect 30026 8610 30031 8638
rect 34577 8610 34582 8638
rect 34610 8610 34634 8638
rect 34662 8610 34686 8638
rect 34714 8610 34738 8638
rect 34766 8610 34790 8638
rect 34818 8610 34842 8638
rect 34870 8610 34894 8638
rect 34922 8610 34946 8638
rect 34974 8610 34998 8638
rect 35026 8610 35031 8638
rect 18774 8470 20230 8498
rect 20258 8470 20790 8498
rect 20818 8470 20823 8498
rect 31425 8470 31430 8498
rect 31458 8470 32830 8498
rect 32858 8470 32863 8498
rect 18774 8442 18802 8470
rect 1409 8414 1414 8442
rect 1442 8414 1862 8442
rect 1890 8414 4494 8442
rect 4522 8414 4527 8442
rect 6113 8414 6118 8442
rect 6146 8414 7014 8442
rect 7042 8414 7047 8442
rect 9809 8414 9814 8442
rect 9842 8414 10038 8442
rect 10066 8414 11438 8442
rect 11466 8414 11471 8442
rect 14401 8414 14406 8442
rect 14434 8414 14966 8442
rect 14994 8414 16254 8442
rect 16282 8414 16814 8442
rect 16842 8414 18270 8442
rect 18298 8414 18774 8442
rect 18802 8414 18807 8442
rect 19441 8414 19446 8442
rect 19474 8414 19950 8442
rect 19978 8414 21406 8442
rect 21434 8414 21439 8442
rect 31033 8414 31038 8442
rect 31066 8414 31934 8442
rect 31962 8414 31967 8442
rect 32153 8414 32158 8442
rect 32186 8414 32718 8442
rect 32746 8414 34398 8442
rect 34426 8414 34431 8442
rect 24425 8358 24430 8386
rect 24458 8358 25158 8386
rect 25186 8358 26222 8386
rect 26250 8358 26255 8386
rect 27393 8358 27398 8386
rect 27426 8358 27678 8386
rect 27706 8358 27711 8386
rect 33161 8358 33166 8386
rect 33194 8358 33614 8386
rect 33642 8358 33647 8386
rect 27398 8330 27426 8358
rect 21401 8302 21406 8330
rect 21434 8302 21798 8330
rect 21826 8302 23422 8330
rect 23450 8302 23455 8330
rect 25377 8302 25382 8330
rect 25410 8302 25942 8330
rect 25970 8302 27426 8330
rect 2077 8218 2082 8246
rect 2110 8218 2134 8246
rect 2162 8218 2186 8246
rect 2214 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2394 8246
rect 2422 8218 2446 8246
rect 2474 8218 2498 8246
rect 2526 8218 2531 8246
rect 7077 8218 7082 8246
rect 7110 8218 7134 8246
rect 7162 8218 7186 8246
rect 7214 8218 7238 8246
rect 7266 8218 7290 8246
rect 7318 8218 7342 8246
rect 7370 8218 7394 8246
rect 7422 8218 7446 8246
rect 7474 8218 7498 8246
rect 7526 8218 7531 8246
rect 12077 8218 12082 8246
rect 12110 8218 12134 8246
rect 12162 8218 12186 8246
rect 12214 8218 12238 8246
rect 12266 8218 12290 8246
rect 12318 8218 12342 8246
rect 12370 8218 12394 8246
rect 12422 8218 12446 8246
rect 12474 8218 12498 8246
rect 12526 8218 12531 8246
rect 17077 8218 17082 8246
rect 17110 8218 17134 8246
rect 17162 8218 17186 8246
rect 17214 8218 17238 8246
rect 17266 8218 17290 8246
rect 17318 8218 17342 8246
rect 17370 8218 17394 8246
rect 17422 8218 17446 8246
rect 17474 8218 17498 8246
rect 17526 8218 17531 8246
rect 22077 8218 22082 8246
rect 22110 8218 22134 8246
rect 22162 8218 22186 8246
rect 22214 8218 22238 8246
rect 22266 8218 22290 8246
rect 22318 8218 22342 8246
rect 22370 8218 22394 8246
rect 22422 8218 22446 8246
rect 22474 8218 22498 8246
rect 22526 8218 22531 8246
rect 27077 8218 27082 8246
rect 27110 8218 27134 8246
rect 27162 8218 27186 8246
rect 27214 8218 27238 8246
rect 27266 8218 27290 8246
rect 27318 8218 27342 8246
rect 27370 8218 27394 8246
rect 27422 8218 27446 8246
rect 27474 8218 27498 8246
rect 27526 8218 27531 8246
rect 32077 8218 32082 8246
rect 32110 8218 32134 8246
rect 32162 8218 32186 8246
rect 32214 8218 32238 8246
rect 32266 8218 32290 8246
rect 32318 8218 32342 8246
rect 32370 8218 32394 8246
rect 32422 8218 32446 8246
rect 32474 8218 32498 8246
rect 32526 8218 32531 8246
rect 37077 8218 37082 8246
rect 37110 8218 37134 8246
rect 37162 8218 37186 8246
rect 37214 8218 37238 8246
rect 37266 8218 37290 8246
rect 37318 8218 37342 8246
rect 37370 8218 37394 8246
rect 37422 8218 37446 8246
rect 37474 8218 37498 8246
rect 37526 8218 37531 8246
rect 8745 8022 8750 8050
rect 8778 8022 10150 8050
rect 10178 8022 10318 8050
rect 10346 8022 10351 8050
rect 26217 8022 26222 8050
rect 26250 8022 26726 8050
rect 26754 8022 26759 8050
rect 31929 8022 31934 8050
rect 31962 8022 32438 8050
rect 32466 8022 32471 8050
rect 34673 8022 34678 8050
rect 34706 8022 36134 8050
rect 36162 8022 36167 8050
rect 10537 7966 10542 7994
rect 10570 7966 32774 7994
rect 32802 7966 32807 7994
rect 4577 7826 4582 7854
rect 4610 7826 4634 7854
rect 4662 7826 4686 7854
rect 4714 7826 4738 7854
rect 4766 7826 4790 7854
rect 4818 7826 4842 7854
rect 4870 7826 4894 7854
rect 4922 7826 4946 7854
rect 4974 7826 4998 7854
rect 5026 7826 5031 7854
rect 9577 7826 9582 7854
rect 9610 7826 9634 7854
rect 9662 7826 9686 7854
rect 9714 7826 9738 7854
rect 9766 7826 9790 7854
rect 9818 7826 9842 7854
rect 9870 7826 9894 7854
rect 9922 7826 9946 7854
rect 9974 7826 9998 7854
rect 10026 7826 10031 7854
rect 14577 7826 14582 7854
rect 14610 7826 14634 7854
rect 14662 7826 14686 7854
rect 14714 7826 14738 7854
rect 14766 7826 14790 7854
rect 14818 7826 14842 7854
rect 14870 7826 14894 7854
rect 14922 7826 14946 7854
rect 14974 7826 14998 7854
rect 15026 7826 15031 7854
rect 19577 7826 19582 7854
rect 19610 7826 19634 7854
rect 19662 7826 19686 7854
rect 19714 7826 19738 7854
rect 19766 7826 19790 7854
rect 19818 7826 19842 7854
rect 19870 7826 19894 7854
rect 19922 7826 19946 7854
rect 19974 7826 19998 7854
rect 20026 7826 20031 7854
rect 24577 7826 24582 7854
rect 24610 7826 24634 7854
rect 24662 7826 24686 7854
rect 24714 7826 24738 7854
rect 24766 7826 24790 7854
rect 24818 7826 24842 7854
rect 24870 7826 24894 7854
rect 24922 7826 24946 7854
rect 24974 7826 24998 7854
rect 25026 7826 25031 7854
rect 29577 7826 29582 7854
rect 29610 7826 29634 7854
rect 29662 7826 29686 7854
rect 29714 7826 29738 7854
rect 29766 7826 29790 7854
rect 29818 7826 29842 7854
rect 29870 7826 29894 7854
rect 29922 7826 29946 7854
rect 29974 7826 29998 7854
rect 30026 7826 30031 7854
rect 34577 7826 34582 7854
rect 34610 7826 34634 7854
rect 34662 7826 34686 7854
rect 34714 7826 34738 7854
rect 34766 7826 34790 7854
rect 34818 7826 34842 7854
rect 34870 7826 34894 7854
rect 34922 7826 34946 7854
rect 34974 7826 34998 7854
rect 35026 7826 35031 7854
rect 6505 7686 6510 7714
rect 6538 7686 7742 7714
rect 7770 7686 7775 7714
rect 5553 7630 5558 7658
rect 5586 7630 6118 7658
rect 6146 7630 7574 7658
rect 7602 7630 7607 7658
rect 20001 7630 20006 7658
rect 20034 7630 21406 7658
rect 21434 7630 21798 7658
rect 21826 7630 21831 7658
rect 25153 7630 25158 7658
rect 25186 7630 25191 7658
rect 33385 7630 33390 7658
rect 33418 7630 35238 7658
rect 35266 7630 35798 7658
rect 35826 7630 35831 7658
rect 36129 7630 36134 7658
rect 36162 7630 36694 7658
rect 36722 7630 36727 7658
rect 25158 7602 25186 7630
rect 10201 7574 10206 7602
rect 10234 7574 10239 7602
rect 23529 7574 23534 7602
rect 23562 7574 23870 7602
rect 23898 7574 24654 7602
rect 24682 7574 25942 7602
rect 25970 7574 25975 7602
rect 32433 7574 32438 7602
rect 32466 7574 32606 7602
rect 32634 7574 32998 7602
rect 33026 7574 33031 7602
rect 10206 7546 10234 7574
rect 7289 7518 7294 7546
rect 7322 7518 7798 7546
rect 7826 7518 9254 7546
rect 9282 7518 9287 7546
rect 10066 7518 10234 7546
rect 24369 7518 24374 7546
rect 24402 7518 24766 7546
rect 24794 7518 24799 7546
rect 35345 7518 35350 7546
rect 35378 7518 35518 7546
rect 35546 7518 35854 7546
rect 35882 7518 35887 7546
rect 10066 7490 10094 7518
rect 8465 7462 8470 7490
rect 8498 7462 10094 7490
rect 2077 7434 2082 7462
rect 2110 7434 2134 7462
rect 2162 7434 2186 7462
rect 2214 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2394 7462
rect 2422 7434 2446 7462
rect 2474 7434 2498 7462
rect 2526 7434 2531 7462
rect 7077 7434 7082 7462
rect 7110 7434 7134 7462
rect 7162 7434 7186 7462
rect 7214 7434 7238 7462
rect 7266 7434 7290 7462
rect 7318 7434 7342 7462
rect 7370 7434 7394 7462
rect 7422 7434 7446 7462
rect 7474 7434 7498 7462
rect 7526 7434 7531 7462
rect 12077 7434 12082 7462
rect 12110 7434 12134 7462
rect 12162 7434 12186 7462
rect 12214 7434 12238 7462
rect 12266 7434 12290 7462
rect 12318 7434 12342 7462
rect 12370 7434 12394 7462
rect 12422 7434 12446 7462
rect 12474 7434 12498 7462
rect 12526 7434 12531 7462
rect 17077 7434 17082 7462
rect 17110 7434 17134 7462
rect 17162 7434 17186 7462
rect 17214 7434 17238 7462
rect 17266 7434 17290 7462
rect 17318 7434 17342 7462
rect 17370 7434 17394 7462
rect 17422 7434 17446 7462
rect 17474 7434 17498 7462
rect 17526 7434 17531 7462
rect 22077 7434 22082 7462
rect 22110 7434 22134 7462
rect 22162 7434 22186 7462
rect 22214 7434 22238 7462
rect 22266 7434 22290 7462
rect 22318 7434 22342 7462
rect 22370 7434 22394 7462
rect 22422 7434 22446 7462
rect 22474 7434 22498 7462
rect 22526 7434 22531 7462
rect 27077 7434 27082 7462
rect 27110 7434 27134 7462
rect 27162 7434 27186 7462
rect 27214 7434 27238 7462
rect 27266 7434 27290 7462
rect 27318 7434 27342 7462
rect 27370 7434 27394 7462
rect 27422 7434 27446 7462
rect 27474 7434 27498 7462
rect 27526 7434 27531 7462
rect 32077 7434 32082 7462
rect 32110 7434 32134 7462
rect 32162 7434 32186 7462
rect 32214 7434 32238 7462
rect 32266 7434 32290 7462
rect 32318 7434 32342 7462
rect 32370 7434 32394 7462
rect 32422 7434 32446 7462
rect 32474 7434 32498 7462
rect 32526 7434 32531 7462
rect 37077 7434 37082 7462
rect 37110 7434 37134 7462
rect 37162 7434 37186 7462
rect 37214 7434 37238 7462
rect 37266 7434 37290 7462
rect 37318 7434 37342 7462
rect 37370 7434 37394 7462
rect 37422 7434 37446 7462
rect 37474 7434 37498 7462
rect 37526 7434 37531 7462
rect 2473 7238 2478 7266
rect 2506 7238 2590 7266
rect 2618 7238 3038 7266
rect 3066 7238 3071 7266
rect 11993 7238 11998 7266
rect 12026 7238 13118 7266
rect 13146 7238 13454 7266
rect 13482 7238 13487 7266
rect 20505 7238 20510 7266
rect 20538 7238 20958 7266
rect 20986 7238 20991 7266
rect 22745 7238 22750 7266
rect 22778 7238 24374 7266
rect 24402 7238 24407 7266
rect 32825 7238 32830 7266
rect 32858 7238 33334 7266
rect 33362 7238 33367 7266
rect 34393 7238 34398 7266
rect 34426 7238 34958 7266
rect 34986 7238 36750 7266
rect 36778 7238 36783 7266
rect 4489 7182 4494 7210
rect 4522 7182 4998 7210
rect 5026 7182 6454 7210
rect 6482 7182 6958 7210
rect 6986 7182 6991 7210
rect 21345 7182 21350 7210
rect 21378 7182 21742 7210
rect 21770 7182 21775 7210
rect 35849 7182 35854 7210
rect 35882 7182 37310 7210
rect 37338 7182 37646 7210
rect 37674 7182 37679 7210
rect 4577 7042 4582 7070
rect 4610 7042 4634 7070
rect 4662 7042 4686 7070
rect 4714 7042 4738 7070
rect 4766 7042 4790 7070
rect 4818 7042 4842 7070
rect 4870 7042 4894 7070
rect 4922 7042 4946 7070
rect 4974 7042 4998 7070
rect 5026 7042 5031 7070
rect 9577 7042 9582 7070
rect 9610 7042 9634 7070
rect 9662 7042 9686 7070
rect 9714 7042 9738 7070
rect 9766 7042 9790 7070
rect 9818 7042 9842 7070
rect 9870 7042 9894 7070
rect 9922 7042 9946 7070
rect 9974 7042 9998 7070
rect 10026 7042 10031 7070
rect 14577 7042 14582 7070
rect 14610 7042 14634 7070
rect 14662 7042 14686 7070
rect 14714 7042 14738 7070
rect 14766 7042 14790 7070
rect 14818 7042 14842 7070
rect 14870 7042 14894 7070
rect 14922 7042 14946 7070
rect 14974 7042 14998 7070
rect 15026 7042 15031 7070
rect 19577 7042 19582 7070
rect 19610 7042 19634 7070
rect 19662 7042 19686 7070
rect 19714 7042 19738 7070
rect 19766 7042 19790 7070
rect 19818 7042 19842 7070
rect 19870 7042 19894 7070
rect 19922 7042 19946 7070
rect 19974 7042 19998 7070
rect 20026 7042 20031 7070
rect 24577 7042 24582 7070
rect 24610 7042 24634 7070
rect 24662 7042 24686 7070
rect 24714 7042 24738 7070
rect 24766 7042 24790 7070
rect 24818 7042 24842 7070
rect 24870 7042 24894 7070
rect 24922 7042 24946 7070
rect 24974 7042 24998 7070
rect 25026 7042 25031 7070
rect 29577 7042 29582 7070
rect 29610 7042 29634 7070
rect 29662 7042 29686 7070
rect 29714 7042 29738 7070
rect 29766 7042 29790 7070
rect 29818 7042 29842 7070
rect 29870 7042 29894 7070
rect 29922 7042 29946 7070
rect 29974 7042 29998 7070
rect 30026 7042 30031 7070
rect 34577 7042 34582 7070
rect 34610 7042 34634 7070
rect 34662 7042 34686 7070
rect 34714 7042 34738 7070
rect 34766 7042 34790 7070
rect 34818 7042 34842 7070
rect 34870 7042 34894 7070
rect 34922 7042 34946 7070
rect 34974 7042 34998 7070
rect 35026 7042 35031 7070
rect 13113 6902 13118 6930
rect 13146 6902 14406 6930
rect 14434 6902 14439 6930
rect 35177 6902 35182 6930
rect 35210 6902 35294 6930
rect 3033 6846 3038 6874
rect 3066 6846 3598 6874
rect 3626 6846 4102 6874
rect 4130 6846 4135 6874
rect 13505 6846 13510 6874
rect 13538 6846 15134 6874
rect 15162 6846 15246 6874
rect 15274 6846 15279 6874
rect 20953 6846 20958 6874
rect 20986 6846 22526 6874
rect 22554 6846 22559 6874
rect 27561 6846 27566 6874
rect 27594 6846 27678 6874
rect 27706 6846 27790 6874
rect 27818 6846 27823 6874
rect 35266 6846 35294 6902
rect 35322 6846 35630 6874
rect 35658 6846 35663 6874
rect 28345 6734 28350 6762
rect 28378 6734 28854 6762
rect 28882 6734 29358 6762
rect 29386 6734 29391 6762
rect 32993 6734 32998 6762
rect 33026 6734 33031 6762
rect 33329 6734 33334 6762
rect 33362 6734 33894 6762
rect 33922 6734 35350 6762
rect 35378 6734 35383 6762
rect 32998 6706 33026 6734
rect 10369 6678 10374 6706
rect 10402 6678 11830 6706
rect 11858 6678 11863 6706
rect 32998 6678 34398 6706
rect 34426 6678 34431 6706
rect 2077 6650 2082 6678
rect 2110 6650 2134 6678
rect 2162 6650 2186 6678
rect 2214 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2394 6678
rect 2422 6650 2446 6678
rect 2474 6650 2498 6678
rect 2526 6650 2531 6678
rect 7077 6650 7082 6678
rect 7110 6650 7134 6678
rect 7162 6650 7186 6678
rect 7214 6650 7238 6678
rect 7266 6650 7290 6678
rect 7318 6650 7342 6678
rect 7370 6650 7394 6678
rect 7422 6650 7446 6678
rect 7474 6650 7498 6678
rect 7526 6650 7531 6678
rect 12077 6650 12082 6678
rect 12110 6650 12134 6678
rect 12162 6650 12186 6678
rect 12214 6650 12238 6678
rect 12266 6650 12290 6678
rect 12318 6650 12342 6678
rect 12370 6650 12394 6678
rect 12422 6650 12446 6678
rect 12474 6650 12498 6678
rect 12526 6650 12531 6678
rect 17077 6650 17082 6678
rect 17110 6650 17134 6678
rect 17162 6650 17186 6678
rect 17214 6650 17238 6678
rect 17266 6650 17290 6678
rect 17318 6650 17342 6678
rect 17370 6650 17394 6678
rect 17422 6650 17446 6678
rect 17474 6650 17498 6678
rect 17526 6650 17531 6678
rect 22077 6650 22082 6678
rect 22110 6650 22134 6678
rect 22162 6650 22186 6678
rect 22214 6650 22238 6678
rect 22266 6650 22290 6678
rect 22318 6650 22342 6678
rect 22370 6650 22394 6678
rect 22422 6650 22446 6678
rect 22474 6650 22498 6678
rect 22526 6650 22531 6678
rect 27077 6650 27082 6678
rect 27110 6650 27134 6678
rect 27162 6650 27186 6678
rect 27214 6650 27238 6678
rect 27266 6650 27290 6678
rect 27318 6650 27342 6678
rect 27370 6650 27394 6678
rect 27422 6650 27446 6678
rect 27474 6650 27498 6678
rect 27526 6650 27531 6678
rect 32077 6650 32082 6678
rect 32110 6650 32134 6678
rect 32162 6650 32186 6678
rect 32214 6650 32238 6678
rect 32266 6650 32290 6678
rect 32318 6650 32342 6678
rect 32370 6650 32394 6678
rect 32422 6650 32446 6678
rect 32474 6650 32498 6678
rect 32526 6650 32531 6678
rect 37077 6650 37082 6678
rect 37110 6650 37134 6678
rect 37162 6650 37186 6678
rect 37214 6650 37238 6678
rect 37266 6650 37290 6678
rect 37318 6650 37342 6678
rect 37370 6650 37394 6678
rect 37422 6650 37446 6678
rect 37474 6650 37498 6678
rect 37526 6650 37531 6678
rect 3985 6510 3990 6538
rect 4018 6510 4270 6538
rect 4298 6510 4303 6538
rect 1913 6454 1918 6482
rect 1946 6454 2198 6482
rect 2226 6454 2758 6482
rect 2786 6454 2791 6482
rect 4097 6454 4102 6482
rect 4130 6454 5558 6482
rect 5586 6454 5591 6482
rect 15745 6454 15750 6482
rect 15778 6454 17486 6482
rect 17514 6454 17519 6482
rect 23193 6454 23198 6482
rect 23226 6454 23534 6482
rect 23562 6454 23567 6482
rect 33721 6454 33726 6482
rect 33754 6454 33894 6482
rect 33922 6454 35798 6482
rect 35826 6454 35831 6482
rect 4577 6258 4582 6286
rect 4610 6258 4634 6286
rect 4662 6258 4686 6286
rect 4714 6258 4738 6286
rect 4766 6258 4790 6286
rect 4818 6258 4842 6286
rect 4870 6258 4894 6286
rect 4922 6258 4946 6286
rect 4974 6258 4998 6286
rect 5026 6258 5031 6286
rect 9577 6258 9582 6286
rect 9610 6258 9634 6286
rect 9662 6258 9686 6286
rect 9714 6258 9738 6286
rect 9766 6258 9790 6286
rect 9818 6258 9842 6286
rect 9870 6258 9894 6286
rect 9922 6258 9946 6286
rect 9974 6258 9998 6286
rect 10026 6258 10031 6286
rect 14577 6258 14582 6286
rect 14610 6258 14634 6286
rect 14662 6258 14686 6286
rect 14714 6258 14738 6286
rect 14766 6258 14790 6286
rect 14818 6258 14842 6286
rect 14870 6258 14894 6286
rect 14922 6258 14946 6286
rect 14974 6258 14998 6286
rect 15026 6258 15031 6286
rect 19577 6258 19582 6286
rect 19610 6258 19634 6286
rect 19662 6258 19686 6286
rect 19714 6258 19738 6286
rect 19766 6258 19790 6286
rect 19818 6258 19842 6286
rect 19870 6258 19894 6286
rect 19922 6258 19946 6286
rect 19974 6258 19998 6286
rect 20026 6258 20031 6286
rect 24577 6258 24582 6286
rect 24610 6258 24634 6286
rect 24662 6258 24686 6286
rect 24714 6258 24738 6286
rect 24766 6258 24790 6286
rect 24818 6258 24842 6286
rect 24870 6258 24894 6286
rect 24922 6258 24946 6286
rect 24974 6258 24998 6286
rect 25026 6258 25031 6286
rect 29577 6258 29582 6286
rect 29610 6258 29634 6286
rect 29662 6258 29686 6286
rect 29714 6258 29738 6286
rect 29766 6258 29790 6286
rect 29818 6258 29842 6286
rect 29870 6258 29894 6286
rect 29922 6258 29946 6286
rect 29974 6258 29998 6286
rect 30026 6258 30031 6286
rect 34577 6258 34582 6286
rect 34610 6258 34634 6286
rect 34662 6258 34686 6286
rect 34714 6258 34738 6286
rect 34766 6258 34790 6286
rect 34818 6258 34842 6286
rect 34870 6258 34894 6286
rect 34922 6258 34946 6286
rect 34974 6258 34998 6286
rect 35026 6258 35031 6286
rect 7569 6062 7574 6090
rect 7602 6062 8078 6090
rect 8106 6062 8111 6090
rect 19105 6062 19110 6090
rect 19138 6062 20510 6090
rect 20538 6062 20543 6090
rect 37361 6062 37366 6090
rect 37394 6062 37646 6090
rect 37674 6062 37679 6090
rect 33665 5894 33670 5922
rect 33698 5894 35574 5922
rect 35602 5894 35607 5922
rect 2077 5866 2082 5894
rect 2110 5866 2134 5894
rect 2162 5866 2186 5894
rect 2214 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2394 5894
rect 2422 5866 2446 5894
rect 2474 5866 2498 5894
rect 2526 5866 2531 5894
rect 7077 5866 7082 5894
rect 7110 5866 7134 5894
rect 7162 5866 7186 5894
rect 7214 5866 7238 5894
rect 7266 5866 7290 5894
rect 7318 5866 7342 5894
rect 7370 5866 7394 5894
rect 7422 5866 7446 5894
rect 7474 5866 7498 5894
rect 7526 5866 7531 5894
rect 12077 5866 12082 5894
rect 12110 5866 12134 5894
rect 12162 5866 12186 5894
rect 12214 5866 12238 5894
rect 12266 5866 12290 5894
rect 12318 5866 12342 5894
rect 12370 5866 12394 5894
rect 12422 5866 12446 5894
rect 12474 5866 12498 5894
rect 12526 5866 12531 5894
rect 17077 5866 17082 5894
rect 17110 5866 17134 5894
rect 17162 5866 17186 5894
rect 17214 5866 17238 5894
rect 17266 5866 17290 5894
rect 17318 5866 17342 5894
rect 17370 5866 17394 5894
rect 17422 5866 17446 5894
rect 17474 5866 17498 5894
rect 17526 5866 17531 5894
rect 22077 5866 22082 5894
rect 22110 5866 22134 5894
rect 22162 5866 22186 5894
rect 22214 5866 22238 5894
rect 22266 5866 22290 5894
rect 22318 5866 22342 5894
rect 22370 5866 22394 5894
rect 22422 5866 22446 5894
rect 22474 5866 22498 5894
rect 22526 5866 22531 5894
rect 27077 5866 27082 5894
rect 27110 5866 27134 5894
rect 27162 5866 27186 5894
rect 27214 5866 27238 5894
rect 27266 5866 27290 5894
rect 27318 5866 27342 5894
rect 27370 5866 27394 5894
rect 27422 5866 27446 5894
rect 27474 5866 27498 5894
rect 27526 5866 27531 5894
rect 32077 5866 32082 5894
rect 32110 5866 32134 5894
rect 32162 5866 32186 5894
rect 32214 5866 32238 5894
rect 32266 5866 32290 5894
rect 32318 5866 32342 5894
rect 32370 5866 32394 5894
rect 32422 5866 32446 5894
rect 32474 5866 32498 5894
rect 32526 5866 32531 5894
rect 37077 5866 37082 5894
rect 37110 5866 37134 5894
rect 37162 5866 37186 5894
rect 37214 5866 37238 5894
rect 37266 5866 37290 5894
rect 37318 5866 37342 5894
rect 37370 5866 37394 5894
rect 37422 5866 37446 5894
rect 37474 5866 37498 5894
rect 37526 5866 37531 5894
rect 8073 5838 8078 5866
rect 8106 5838 9534 5866
rect 9562 5838 10038 5866
rect 10066 5838 11550 5866
rect 11578 5838 11583 5866
rect 30193 5838 30198 5866
rect 30226 5838 31822 5866
rect 31850 5838 31855 5866
rect 21793 5782 21798 5810
rect 21826 5782 21854 5810
rect 21882 5782 21887 5810
rect 23417 5782 23422 5810
rect 23450 5782 23870 5810
rect 23898 5782 25158 5810
rect 25186 5782 25191 5810
rect 35681 5726 35686 5754
rect 35714 5726 36974 5754
rect 11937 5670 11942 5698
rect 11970 5670 12502 5698
rect 12530 5670 12726 5698
rect 12754 5670 12759 5698
rect 32433 5670 32438 5698
rect 32466 5670 32718 5698
rect 32746 5670 32751 5698
rect 36946 5642 36974 5726
rect 11545 5614 11550 5642
rect 11578 5614 12334 5642
rect 12362 5614 12614 5642
rect 12642 5614 13118 5642
rect 13146 5614 13151 5642
rect 24481 5614 24486 5642
rect 24514 5614 25046 5642
rect 25074 5614 26502 5642
rect 26530 5614 26535 5642
rect 36946 5614 37590 5642
rect 37618 5614 38990 5642
rect 39018 5614 39023 5642
rect 16865 5558 16870 5586
rect 16898 5558 26894 5586
rect 26922 5558 27006 5586
rect 27034 5558 27039 5586
rect 4577 5474 4582 5502
rect 4610 5474 4634 5502
rect 4662 5474 4686 5502
rect 4714 5474 4738 5502
rect 4766 5474 4790 5502
rect 4818 5474 4842 5502
rect 4870 5474 4894 5502
rect 4922 5474 4946 5502
rect 4974 5474 4998 5502
rect 5026 5474 5031 5502
rect 9577 5474 9582 5502
rect 9610 5474 9634 5502
rect 9662 5474 9686 5502
rect 9714 5474 9738 5502
rect 9766 5474 9790 5502
rect 9818 5474 9842 5502
rect 9870 5474 9894 5502
rect 9922 5474 9946 5502
rect 9974 5474 9998 5502
rect 10026 5474 10031 5502
rect 14577 5474 14582 5502
rect 14610 5474 14634 5502
rect 14662 5474 14686 5502
rect 14714 5474 14738 5502
rect 14766 5474 14790 5502
rect 14818 5474 14842 5502
rect 14870 5474 14894 5502
rect 14922 5474 14946 5502
rect 14974 5474 14998 5502
rect 15026 5474 15031 5502
rect 19577 5474 19582 5502
rect 19610 5474 19634 5502
rect 19662 5474 19686 5502
rect 19714 5474 19738 5502
rect 19766 5474 19790 5502
rect 19818 5474 19842 5502
rect 19870 5474 19894 5502
rect 19922 5474 19946 5502
rect 19974 5474 19998 5502
rect 20026 5474 20031 5502
rect 24577 5474 24582 5502
rect 24610 5474 24634 5502
rect 24662 5474 24686 5502
rect 24714 5474 24738 5502
rect 24766 5474 24790 5502
rect 24818 5474 24842 5502
rect 24870 5474 24894 5502
rect 24922 5474 24946 5502
rect 24974 5474 24998 5502
rect 25026 5474 25031 5502
rect 29577 5474 29582 5502
rect 29610 5474 29634 5502
rect 29662 5474 29686 5502
rect 29714 5474 29738 5502
rect 29766 5474 29790 5502
rect 29818 5474 29842 5502
rect 29870 5474 29894 5502
rect 29922 5474 29946 5502
rect 29974 5474 29998 5502
rect 30026 5474 30031 5502
rect 34577 5474 34582 5502
rect 34610 5474 34634 5502
rect 34662 5474 34686 5502
rect 34714 5474 34738 5502
rect 34766 5474 34790 5502
rect 34818 5474 34842 5502
rect 34870 5474 34894 5502
rect 34922 5474 34946 5502
rect 34974 5474 34998 5502
rect 35026 5474 35031 5502
rect 22521 5390 22526 5418
rect 22554 5390 23030 5418
rect 23058 5390 24430 5418
rect 24458 5390 25046 5418
rect 25074 5390 25079 5418
rect 3593 5278 3598 5306
rect 3626 5278 4102 5306
rect 4130 5278 4135 5306
rect 6505 5278 6510 5306
rect 6538 5278 7742 5306
rect 7770 5278 7966 5306
rect 7994 5278 8246 5306
rect 8274 5278 8279 5306
rect 9529 5278 9534 5306
rect 9562 5278 9814 5306
rect 9842 5278 10094 5306
rect 12721 5278 12726 5306
rect 12754 5278 13286 5306
rect 13314 5278 13510 5306
rect 13538 5278 13543 5306
rect 20001 5278 20006 5306
rect 20034 5278 20118 5306
rect 20146 5278 21462 5306
rect 21490 5278 23422 5306
rect 23450 5278 23455 5306
rect 29353 5278 29358 5306
rect 29386 5278 30926 5306
rect 30954 5278 30959 5306
rect 32713 5278 32718 5306
rect 32746 5278 34174 5306
rect 34202 5278 34207 5306
rect 10066 5250 10094 5278
rect 10033 5222 10038 5250
rect 10066 5222 11550 5250
rect 11578 5222 11583 5250
rect 33385 5222 33390 5250
rect 33418 5222 34622 5250
rect 34650 5222 34846 5250
rect 34874 5222 34879 5250
rect 16417 5166 16422 5194
rect 16450 5166 16758 5194
rect 16786 5166 18438 5194
rect 18466 5166 18471 5194
rect 2077 5082 2082 5110
rect 2110 5082 2134 5110
rect 2162 5082 2186 5110
rect 2214 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2394 5110
rect 2422 5082 2446 5110
rect 2474 5082 2498 5110
rect 2526 5082 2531 5110
rect 7077 5082 7082 5110
rect 7110 5082 7134 5110
rect 7162 5082 7186 5110
rect 7214 5082 7238 5110
rect 7266 5082 7290 5110
rect 7318 5082 7342 5110
rect 7370 5082 7394 5110
rect 7422 5082 7446 5110
rect 7474 5082 7498 5110
rect 7526 5082 7531 5110
rect 12077 5082 12082 5110
rect 12110 5082 12134 5110
rect 12162 5082 12186 5110
rect 12214 5082 12238 5110
rect 12266 5082 12290 5110
rect 12318 5082 12342 5110
rect 12370 5082 12394 5110
rect 12422 5082 12446 5110
rect 12474 5082 12498 5110
rect 12526 5082 12531 5110
rect 17077 5082 17082 5110
rect 17110 5082 17134 5110
rect 17162 5082 17186 5110
rect 17214 5082 17238 5110
rect 17266 5082 17290 5110
rect 17318 5082 17342 5110
rect 17370 5082 17394 5110
rect 17422 5082 17446 5110
rect 17474 5082 17498 5110
rect 17526 5082 17531 5110
rect 22077 5082 22082 5110
rect 22110 5082 22134 5110
rect 22162 5082 22186 5110
rect 22214 5082 22238 5110
rect 22266 5082 22290 5110
rect 22318 5082 22342 5110
rect 22370 5082 22394 5110
rect 22422 5082 22446 5110
rect 22474 5082 22498 5110
rect 22526 5082 22531 5110
rect 27077 5082 27082 5110
rect 27110 5082 27134 5110
rect 27162 5082 27186 5110
rect 27214 5082 27238 5110
rect 27266 5082 27290 5110
rect 27318 5082 27342 5110
rect 27370 5082 27394 5110
rect 27422 5082 27446 5110
rect 27474 5082 27498 5110
rect 27526 5082 27531 5110
rect 32077 5082 32082 5110
rect 32110 5082 32134 5110
rect 32162 5082 32186 5110
rect 32214 5082 32238 5110
rect 32266 5082 32290 5110
rect 32318 5082 32342 5110
rect 32370 5082 32394 5110
rect 32422 5082 32446 5110
rect 32474 5082 32498 5110
rect 32526 5082 32531 5110
rect 37077 5082 37082 5110
rect 37110 5082 37134 5110
rect 37162 5082 37186 5110
rect 37214 5082 37238 5110
rect 37266 5082 37290 5110
rect 37318 5082 37342 5110
rect 37370 5082 37394 5110
rect 37422 5082 37446 5110
rect 37474 5082 37498 5110
rect 37526 5082 37531 5110
rect 4097 5054 4102 5082
rect 4130 5054 5558 5082
rect 5586 5054 5591 5082
rect 18433 5054 18438 5082
rect 18466 5054 19950 5082
rect 19978 5054 19983 5082
rect 33665 5054 33670 5082
rect 33698 5054 35630 5082
rect 35658 5054 35663 5082
rect 26889 4998 26894 5026
rect 26922 4998 27174 5026
rect 27202 4998 27207 5026
rect 28233 4998 28238 5026
rect 28266 4998 30142 5026
rect 30170 4998 30366 5026
rect 30394 4998 33782 5026
rect 33810 4998 35742 5026
rect 35770 4998 37702 5026
rect 37730 4998 37735 5026
rect 23193 4886 23198 4914
rect 23226 4886 24654 4914
rect 24682 4886 24878 4914
rect 24906 4886 25158 4914
rect 25186 4886 25191 4914
rect 27001 4886 27006 4914
rect 27034 4886 28462 4914
rect 28490 4886 28495 4914
rect 35569 4886 35574 4914
rect 35602 4886 37618 4914
rect 37590 4858 37618 4886
rect 28289 4830 28294 4858
rect 28322 4830 30030 4858
rect 30058 4830 31934 4858
rect 31962 4830 31967 4858
rect 37585 4830 37590 4858
rect 37618 4830 38206 4858
rect 38234 4830 38239 4858
rect 26497 4718 26502 4746
rect 26530 4718 26894 4746
rect 26922 4718 28182 4746
rect 28210 4718 28215 4746
rect 4577 4690 4582 4718
rect 4610 4690 4634 4718
rect 4662 4690 4686 4718
rect 4714 4690 4738 4718
rect 4766 4690 4790 4718
rect 4818 4690 4842 4718
rect 4870 4690 4894 4718
rect 4922 4690 4946 4718
rect 4974 4690 4998 4718
rect 5026 4690 5031 4718
rect 9577 4690 9582 4718
rect 9610 4690 9634 4718
rect 9662 4690 9686 4718
rect 9714 4690 9738 4718
rect 9766 4690 9790 4718
rect 9818 4690 9842 4718
rect 9870 4690 9894 4718
rect 9922 4690 9946 4718
rect 9974 4690 9998 4718
rect 10026 4690 10031 4718
rect 14577 4690 14582 4718
rect 14610 4690 14634 4718
rect 14662 4690 14686 4718
rect 14714 4690 14738 4718
rect 14766 4690 14790 4718
rect 14818 4690 14842 4718
rect 14870 4690 14894 4718
rect 14922 4690 14946 4718
rect 14974 4690 14998 4718
rect 15026 4690 15031 4718
rect 19577 4690 19582 4718
rect 19610 4690 19634 4718
rect 19662 4690 19686 4718
rect 19714 4690 19738 4718
rect 19766 4690 19790 4718
rect 19818 4690 19842 4718
rect 19870 4690 19894 4718
rect 19922 4690 19946 4718
rect 19974 4690 19998 4718
rect 20026 4690 20031 4718
rect 24577 4690 24582 4718
rect 24610 4690 24634 4718
rect 24662 4690 24686 4718
rect 24714 4690 24738 4718
rect 24766 4690 24790 4718
rect 24818 4690 24842 4718
rect 24870 4690 24894 4718
rect 24922 4690 24946 4718
rect 24974 4690 24998 4718
rect 25026 4690 25031 4718
rect 29577 4690 29582 4718
rect 29610 4690 29634 4718
rect 29662 4690 29686 4718
rect 29714 4690 29738 4718
rect 29766 4690 29790 4718
rect 29818 4690 29842 4718
rect 29870 4690 29894 4718
rect 29922 4690 29946 4718
rect 29974 4690 29998 4718
rect 30026 4690 30031 4718
rect 34577 4690 34582 4718
rect 34610 4690 34634 4718
rect 34662 4690 34686 4718
rect 34714 4690 34738 4718
rect 34766 4690 34790 4718
rect 34818 4690 34842 4718
rect 34870 4690 34894 4718
rect 34922 4690 34946 4718
rect 34974 4690 34998 4718
rect 35026 4690 35031 4718
rect 5777 4606 5782 4634
rect 5810 4606 16366 4634
rect 16394 4606 16399 4634
rect 21345 4550 21350 4578
rect 21378 4550 21798 4578
rect 2753 4494 2758 4522
rect 2786 4494 2982 4522
rect 3010 4494 3318 4522
rect 3346 4494 3598 4522
rect 3626 4494 3631 4522
rect 6001 4494 6006 4522
rect 6034 4494 7294 4522
rect 7322 4494 7574 4522
rect 7602 4494 7607 4522
rect 9025 4494 9030 4522
rect 9058 4494 10262 4522
rect 10290 4494 10486 4522
rect 10514 4494 11774 4522
rect 11802 4494 11942 4522
rect 11970 4494 11975 4522
rect 21826 4494 21854 4578
rect 28065 4550 28070 4578
rect 28098 4550 28238 4578
rect 28266 4550 28271 4578
rect 21882 4494 22694 4522
rect 22722 4494 22918 4522
rect 22946 4494 23198 4522
rect 23226 4494 23231 4522
rect 25433 4494 25438 4522
rect 25466 4494 26894 4522
rect 26922 4494 27174 4522
rect 27202 4494 27207 4522
rect 28457 4494 28462 4522
rect 28490 4494 28742 4522
rect 28770 4494 28775 4522
rect 31929 4494 31934 4522
rect 31962 4494 32046 4522
rect 32074 4494 32079 4522
rect 16977 4438 16982 4466
rect 17010 4438 28070 4466
rect 28098 4438 28103 4466
rect 31985 4438 31990 4466
rect 32018 4438 32158 4466
rect 32186 4438 32326 4466
rect 32354 4438 32359 4466
rect 2077 4298 2082 4326
rect 2110 4298 2134 4326
rect 2162 4298 2186 4326
rect 2214 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2394 4326
rect 2422 4298 2446 4326
rect 2474 4298 2498 4326
rect 2526 4298 2531 4326
rect 7077 4298 7082 4326
rect 7110 4298 7134 4326
rect 7162 4298 7186 4326
rect 7214 4298 7238 4326
rect 7266 4298 7290 4326
rect 7318 4298 7342 4326
rect 7370 4298 7394 4326
rect 7422 4298 7446 4326
rect 7474 4298 7498 4326
rect 7526 4298 7531 4326
rect 12077 4298 12082 4326
rect 12110 4298 12134 4326
rect 12162 4298 12186 4326
rect 12214 4298 12238 4326
rect 12266 4298 12290 4326
rect 12318 4298 12342 4326
rect 12370 4298 12394 4326
rect 12422 4298 12446 4326
rect 12474 4298 12498 4326
rect 12526 4298 12531 4326
rect 17077 4298 17082 4326
rect 17110 4298 17134 4326
rect 17162 4298 17186 4326
rect 17214 4298 17238 4326
rect 17266 4298 17290 4326
rect 17318 4298 17342 4326
rect 17370 4298 17394 4326
rect 17422 4298 17446 4326
rect 17474 4298 17498 4326
rect 17526 4298 17531 4326
rect 22077 4298 22082 4326
rect 22110 4298 22134 4326
rect 22162 4298 22186 4326
rect 22214 4298 22238 4326
rect 22266 4298 22290 4326
rect 22318 4298 22342 4326
rect 22370 4298 22394 4326
rect 22422 4298 22446 4326
rect 22474 4298 22498 4326
rect 22526 4298 22531 4326
rect 27077 4298 27082 4326
rect 27110 4298 27134 4326
rect 27162 4298 27186 4326
rect 27214 4298 27238 4326
rect 27266 4298 27290 4326
rect 27318 4298 27342 4326
rect 27370 4298 27394 4326
rect 27422 4298 27446 4326
rect 27474 4298 27498 4326
rect 27526 4298 27531 4326
rect 32077 4298 32082 4326
rect 32110 4298 32134 4326
rect 32162 4298 32186 4326
rect 32214 4298 32238 4326
rect 32266 4298 32290 4326
rect 32318 4298 32342 4326
rect 32370 4298 32394 4326
rect 32422 4298 32446 4326
rect 32474 4298 32498 4326
rect 32526 4298 32531 4326
rect 37077 4298 37082 4326
rect 37110 4298 37134 4326
rect 37162 4298 37186 4326
rect 37214 4298 37238 4326
rect 37266 4298 37290 4326
rect 37318 4298 37342 4326
rect 37370 4298 37394 4326
rect 37422 4298 37446 4326
rect 37474 4298 37498 4326
rect 37526 4298 37531 4326
rect 5273 4214 5278 4242
rect 5306 4214 6006 4242
rect 6034 4214 6039 4242
rect 11377 4214 11382 4242
rect 11410 4214 11998 4242
rect 12026 4214 12031 4242
rect 26889 4214 26894 4242
rect 26922 4214 27510 4242
rect 27538 4214 27678 4242
rect 27706 4214 28686 4242
rect 28714 4214 28910 4242
rect 28938 4214 29414 4242
rect 29442 4214 29447 4242
rect 30977 4214 30982 4242
rect 31010 4214 31990 4242
rect 32018 4214 32158 4242
rect 32186 4214 32718 4242
rect 32746 4214 32751 4242
rect 38593 4214 38598 4242
rect 38626 4214 38822 4242
rect 38850 4214 38855 4242
rect 4265 4158 4270 4186
rect 4298 4158 4494 4186
rect 4522 4158 4998 4186
rect 5026 4158 6454 4186
rect 6482 4158 7014 4186
rect 7042 4158 7047 4186
rect 28233 4158 28238 4186
rect 28266 4158 28271 4186
rect 35625 4158 35630 4186
rect 35658 4158 35854 4186
rect 35882 4158 36918 4186
rect 28238 4130 28266 4158
rect 36946 4130 36974 4186
rect 1801 4102 1806 4130
rect 1834 4102 1918 4130
rect 1946 4102 2030 4130
rect 2058 4102 2063 4130
rect 12945 4102 12950 4130
rect 12978 4102 13230 4130
rect 13258 4102 13263 4130
rect 20505 4102 20510 4130
rect 20538 4102 20958 4130
rect 20986 4102 20991 4130
rect 24481 4102 24486 4130
rect 24514 4102 25102 4130
rect 25130 4102 26502 4130
rect 26530 4102 26838 4130
rect 26866 4102 26871 4130
rect 28238 4102 28462 4130
rect 28490 4102 28495 4130
rect 36946 4102 37086 4130
rect 37114 4102 37119 4130
rect 30137 4046 30142 4074
rect 30170 4046 30310 4074
rect 30338 4046 30343 4074
rect 38649 3934 38654 3962
rect 38682 3934 38934 3962
rect 38962 3934 38967 3962
rect 4577 3906 4582 3934
rect 4610 3906 4634 3934
rect 4662 3906 4686 3934
rect 4714 3906 4738 3934
rect 4766 3906 4790 3934
rect 4818 3906 4842 3934
rect 4870 3906 4894 3934
rect 4922 3906 4946 3934
rect 4974 3906 4998 3934
rect 5026 3906 5031 3934
rect 9577 3906 9582 3934
rect 9610 3906 9634 3934
rect 9662 3906 9686 3934
rect 9714 3906 9738 3934
rect 9766 3906 9790 3934
rect 9818 3906 9842 3934
rect 9870 3906 9894 3934
rect 9922 3906 9946 3934
rect 9974 3906 9998 3934
rect 10026 3906 10031 3934
rect 14577 3906 14582 3934
rect 14610 3906 14634 3934
rect 14662 3906 14686 3934
rect 14714 3906 14738 3934
rect 14766 3906 14790 3934
rect 14818 3906 14842 3934
rect 14870 3906 14894 3934
rect 14922 3906 14946 3934
rect 14974 3906 14998 3934
rect 15026 3906 15031 3934
rect 19577 3906 19582 3934
rect 19610 3906 19634 3934
rect 19662 3906 19686 3934
rect 19714 3906 19738 3934
rect 19766 3906 19790 3934
rect 19818 3906 19842 3934
rect 19870 3906 19894 3934
rect 19922 3906 19946 3934
rect 19974 3906 19998 3934
rect 20026 3906 20031 3934
rect 24577 3906 24582 3934
rect 24610 3906 24634 3934
rect 24662 3906 24686 3934
rect 24714 3906 24738 3934
rect 24766 3906 24790 3934
rect 24818 3906 24842 3934
rect 24870 3906 24894 3934
rect 24922 3906 24946 3934
rect 24974 3906 24998 3934
rect 25026 3906 25031 3934
rect 29577 3906 29582 3934
rect 29610 3906 29634 3934
rect 29662 3906 29686 3934
rect 29714 3906 29738 3934
rect 29766 3906 29790 3934
rect 29818 3906 29842 3934
rect 29870 3906 29894 3934
rect 29922 3906 29946 3934
rect 29974 3906 29998 3934
rect 30026 3906 30031 3934
rect 34577 3906 34582 3934
rect 34610 3906 34634 3934
rect 34662 3906 34686 3934
rect 34714 3906 34738 3934
rect 34766 3906 34790 3934
rect 34818 3906 34842 3934
rect 34870 3906 34894 3934
rect 34922 3906 34946 3934
rect 34974 3906 34998 3934
rect 35026 3906 35031 3934
rect 26889 3878 26894 3906
rect 26922 3878 27174 3906
rect 27202 3878 27207 3906
rect 26161 3822 26166 3850
rect 26194 3822 30814 3850
rect 30842 3822 30847 3850
rect 3257 3766 3262 3794
rect 3290 3766 8806 3794
rect 8834 3766 8839 3794
rect 8465 3710 8470 3738
rect 8498 3710 8974 3738
rect 9002 3710 9007 3738
rect 9473 3710 9478 3738
rect 9506 3710 9814 3738
rect 9842 3710 9847 3738
rect 10481 3710 10486 3738
rect 10514 3710 10878 3738
rect 10906 3710 11774 3738
rect 11802 3710 11807 3738
rect 13225 3710 13230 3738
rect 13258 3710 13790 3738
rect 13818 3710 14070 3738
rect 14098 3710 14103 3738
rect 15241 3710 15246 3738
rect 15274 3710 15526 3738
rect 15554 3710 15559 3738
rect 20953 3710 20958 3738
rect 20986 3710 22526 3738
rect 22554 3710 23030 3738
rect 23058 3710 23063 3738
rect 31985 3710 31990 3738
rect 32018 3710 32158 3738
rect 32186 3710 32326 3738
rect 32354 3710 32359 3738
rect 33889 3710 33894 3738
rect 33922 3710 34454 3738
rect 34482 3710 35350 3738
rect 35378 3710 35630 3738
rect 35658 3710 35663 3738
rect 37585 3710 37590 3738
rect 37618 3710 38150 3738
rect 38178 3710 38183 3738
rect 38649 3710 38654 3738
rect 38682 3710 38822 3738
rect 38850 3710 38855 3738
rect 1913 3598 1918 3626
rect 1946 3598 2030 3626
rect 2058 3598 2478 3626
rect 2506 3598 4494 3626
rect 4522 3598 4527 3626
rect 2077 3514 2082 3542
rect 2110 3514 2134 3542
rect 2162 3514 2186 3542
rect 2214 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2394 3542
rect 2422 3514 2446 3542
rect 2474 3514 2498 3542
rect 2526 3514 2531 3542
rect 7077 3514 7082 3542
rect 7110 3514 7134 3542
rect 7162 3514 7186 3542
rect 7214 3514 7238 3542
rect 7266 3514 7290 3542
rect 7318 3514 7342 3542
rect 7370 3514 7394 3542
rect 7422 3514 7446 3542
rect 7474 3514 7498 3542
rect 7526 3514 7531 3542
rect 12077 3514 12082 3542
rect 12110 3514 12134 3542
rect 12162 3514 12186 3542
rect 12214 3514 12238 3542
rect 12266 3514 12290 3542
rect 12318 3514 12342 3542
rect 12370 3514 12394 3542
rect 12422 3514 12446 3542
rect 12474 3514 12498 3542
rect 12526 3514 12531 3542
rect 17077 3514 17082 3542
rect 17110 3514 17134 3542
rect 17162 3514 17186 3542
rect 17214 3514 17238 3542
rect 17266 3514 17290 3542
rect 17318 3514 17342 3542
rect 17370 3514 17394 3542
rect 17422 3514 17446 3542
rect 17474 3514 17498 3542
rect 17526 3514 17531 3542
rect 22077 3514 22082 3542
rect 22110 3514 22134 3542
rect 22162 3514 22186 3542
rect 22214 3514 22238 3542
rect 22266 3514 22290 3542
rect 22318 3514 22342 3542
rect 22370 3514 22394 3542
rect 22422 3514 22446 3542
rect 22474 3514 22498 3542
rect 22526 3514 22531 3542
rect 27077 3514 27082 3542
rect 27110 3514 27134 3542
rect 27162 3514 27186 3542
rect 27214 3514 27238 3542
rect 27266 3514 27290 3542
rect 27318 3514 27342 3542
rect 27370 3514 27394 3542
rect 27422 3514 27446 3542
rect 27474 3514 27498 3542
rect 27526 3514 27531 3542
rect 32077 3514 32082 3542
rect 32110 3514 32134 3542
rect 32162 3514 32186 3542
rect 32214 3514 32238 3542
rect 32266 3514 32290 3542
rect 32318 3514 32342 3542
rect 32370 3514 32394 3542
rect 32422 3514 32446 3542
rect 32474 3514 32498 3542
rect 32526 3514 32531 3542
rect 37077 3514 37082 3542
rect 37110 3514 37134 3542
rect 37162 3514 37186 3542
rect 37214 3514 37238 3542
rect 37266 3514 37290 3542
rect 37318 3514 37342 3542
rect 37370 3514 37394 3542
rect 37422 3514 37446 3542
rect 37474 3514 37498 3542
rect 37526 3514 37531 3542
rect 8017 3430 8022 3458
rect 8050 3430 8302 3458
rect 8330 3430 10486 3458
rect 10514 3430 10519 3458
rect 23865 3430 23870 3458
rect 23898 3430 25382 3458
rect 25410 3430 25415 3458
rect 8022 3346 8050 3430
rect 8969 3374 8974 3402
rect 9002 3374 9478 3402
rect 9506 3374 9511 3402
rect 14065 3374 14070 3402
rect 14098 3374 15246 3402
rect 15274 3374 15750 3402
rect 15778 3374 15783 3402
rect 17593 3374 17598 3402
rect 17626 3374 19110 3402
rect 19138 3374 20510 3402
rect 20538 3374 20543 3402
rect 24257 3374 24262 3402
rect 24290 3374 26166 3402
rect 26194 3374 26199 3402
rect 30473 3374 30478 3402
rect 30506 3374 30982 3402
rect 31010 3374 31015 3402
rect 36913 3374 36918 3402
rect 36946 3374 37142 3402
rect 37170 3374 37175 3402
rect 30982 3346 31010 3374
rect 5721 3318 5726 3346
rect 5754 3318 6006 3346
rect 6034 3318 8050 3346
rect 11937 3318 11942 3346
rect 11970 3318 12334 3346
rect 12362 3318 12367 3346
rect 25993 3318 25998 3346
rect 26026 3318 30702 3346
rect 30730 3318 30735 3346
rect 30982 3318 31598 3346
rect 31626 3318 31631 3346
rect 34169 3318 34174 3346
rect 34202 3318 34510 3346
rect 34538 3318 34678 3346
rect 34706 3318 36134 3346
rect 36162 3318 36694 3346
rect 36722 3318 36727 3346
rect 11769 3262 11774 3290
rect 11802 3262 14406 3290
rect 14434 3262 15078 3290
rect 15106 3262 15111 3290
rect 30025 3262 30030 3290
rect 30058 3262 35686 3290
rect 35714 3262 35719 3290
rect 4577 3122 4582 3150
rect 4610 3122 4634 3150
rect 4662 3122 4686 3150
rect 4714 3122 4738 3150
rect 4766 3122 4790 3150
rect 4818 3122 4842 3150
rect 4870 3122 4894 3150
rect 4922 3122 4946 3150
rect 4974 3122 4998 3150
rect 5026 3122 5031 3150
rect 9577 3122 9582 3150
rect 9610 3122 9634 3150
rect 9662 3122 9686 3150
rect 9714 3122 9738 3150
rect 9766 3122 9790 3150
rect 9818 3122 9842 3150
rect 9870 3122 9894 3150
rect 9922 3122 9946 3150
rect 9974 3122 9998 3150
rect 10026 3122 10031 3150
rect 14577 3122 14582 3150
rect 14610 3122 14634 3150
rect 14662 3122 14686 3150
rect 14714 3122 14738 3150
rect 14766 3122 14790 3150
rect 14818 3122 14842 3150
rect 14870 3122 14894 3150
rect 14922 3122 14946 3150
rect 14974 3122 14998 3150
rect 15026 3122 15031 3150
rect 19577 3122 19582 3150
rect 19610 3122 19634 3150
rect 19662 3122 19686 3150
rect 19714 3122 19738 3150
rect 19766 3122 19790 3150
rect 19818 3122 19842 3150
rect 19870 3122 19894 3150
rect 19922 3122 19946 3150
rect 19974 3122 19998 3150
rect 20026 3122 20031 3150
rect 24577 3122 24582 3150
rect 24610 3122 24634 3150
rect 24662 3122 24686 3150
rect 24714 3122 24738 3150
rect 24766 3122 24790 3150
rect 24818 3122 24842 3150
rect 24870 3122 24894 3150
rect 24922 3122 24946 3150
rect 24974 3122 24998 3150
rect 25026 3122 25031 3150
rect 29577 3122 29582 3150
rect 29610 3122 29634 3150
rect 29662 3122 29686 3150
rect 29714 3122 29738 3150
rect 29766 3122 29790 3150
rect 29818 3122 29842 3150
rect 29870 3122 29894 3150
rect 29922 3122 29946 3150
rect 29974 3122 29998 3150
rect 30026 3122 30031 3150
rect 34577 3122 34582 3150
rect 34610 3122 34634 3150
rect 34662 3122 34686 3150
rect 34714 3122 34738 3150
rect 34766 3122 34790 3150
rect 34818 3122 34842 3150
rect 34870 3122 34894 3150
rect 34922 3122 34946 3150
rect 34974 3122 34998 3150
rect 35026 3122 35031 3150
rect 37305 3038 37310 3066
rect 37338 3038 37646 3066
rect 37674 3038 37679 3066
rect 14401 2982 14406 3010
rect 14434 2982 18214 3010
rect 18242 2982 18247 3010
rect 28345 2982 28350 3010
rect 28378 2982 28518 3010
rect 28546 2982 30086 3010
rect 30114 2982 30119 3010
rect 30305 2982 30310 3010
rect 30338 2982 31990 3010
rect 32018 2982 32158 3010
rect 32186 2982 32326 3010
rect 32354 2982 32359 3010
rect 32881 2982 32886 3010
rect 32914 2982 34174 3010
rect 34202 2982 34678 3010
rect 34706 2982 34711 3010
rect 12441 2926 12446 2954
rect 12474 2926 13174 2954
rect 13202 2926 13207 2954
rect 14961 2926 14966 2954
rect 14994 2926 15078 2954
rect 15106 2926 15694 2954
rect 15722 2926 16422 2954
rect 16450 2926 16758 2954
rect 16786 2926 16791 2954
rect 20001 2926 20006 2954
rect 20034 2926 20118 2954
rect 20146 2926 21350 2954
rect 21378 2926 21383 2954
rect 29353 2926 29358 2954
rect 29386 2926 29470 2954
rect 29498 2926 29918 2954
rect 29946 2926 31318 2954
rect 31346 2926 32830 2954
rect 32858 2926 33166 2954
rect 33194 2926 33390 2954
rect 33418 2926 33423 2954
rect 15521 2870 15526 2898
rect 15554 2870 32438 2898
rect 32466 2870 32998 2898
rect 33026 2870 34230 2898
rect 34258 2870 34263 2898
rect 35905 2870 35910 2898
rect 35938 2870 38318 2898
rect 38346 2870 38654 2898
rect 38682 2870 38822 2898
rect 38850 2870 38855 2898
rect 2077 2730 2082 2758
rect 2110 2730 2134 2758
rect 2162 2730 2186 2758
rect 2214 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2394 2758
rect 2422 2730 2446 2758
rect 2474 2730 2498 2758
rect 2526 2730 2531 2758
rect 7077 2730 7082 2758
rect 7110 2730 7134 2758
rect 7162 2730 7186 2758
rect 7214 2730 7238 2758
rect 7266 2730 7290 2758
rect 7318 2730 7342 2758
rect 7370 2730 7394 2758
rect 7422 2730 7446 2758
rect 7474 2730 7498 2758
rect 7526 2730 7531 2758
rect 12077 2730 12082 2758
rect 12110 2730 12134 2758
rect 12162 2730 12186 2758
rect 12214 2730 12238 2758
rect 12266 2730 12290 2758
rect 12318 2730 12342 2758
rect 12370 2730 12394 2758
rect 12422 2730 12446 2758
rect 12474 2730 12498 2758
rect 12526 2730 12531 2758
rect 17077 2730 17082 2758
rect 17110 2730 17134 2758
rect 17162 2730 17186 2758
rect 17214 2730 17238 2758
rect 17266 2730 17290 2758
rect 17318 2730 17342 2758
rect 17370 2730 17394 2758
rect 17422 2730 17446 2758
rect 17474 2730 17498 2758
rect 17526 2730 17531 2758
rect 22077 2730 22082 2758
rect 22110 2730 22134 2758
rect 22162 2730 22186 2758
rect 22214 2730 22238 2758
rect 22266 2730 22290 2758
rect 22318 2730 22342 2758
rect 22370 2730 22394 2758
rect 22422 2730 22446 2758
rect 22474 2730 22498 2758
rect 22526 2730 22531 2758
rect 27077 2730 27082 2758
rect 27110 2730 27134 2758
rect 27162 2730 27186 2758
rect 27214 2730 27238 2758
rect 27266 2730 27290 2758
rect 27318 2730 27342 2758
rect 27370 2730 27394 2758
rect 27422 2730 27446 2758
rect 27474 2730 27498 2758
rect 27526 2730 27531 2758
rect 32077 2730 32082 2758
rect 32110 2730 32134 2758
rect 32162 2730 32186 2758
rect 32214 2730 32238 2758
rect 32266 2730 32290 2758
rect 32318 2730 32342 2758
rect 32370 2730 32394 2758
rect 32422 2730 32446 2758
rect 32474 2730 32498 2758
rect 32526 2730 32531 2758
rect 37077 2730 37082 2758
rect 37110 2730 37134 2758
rect 37162 2730 37186 2758
rect 37214 2730 37238 2758
rect 37266 2730 37290 2758
rect 37318 2730 37342 2758
rect 37370 2730 37394 2758
rect 37422 2730 37446 2758
rect 37474 2730 37498 2758
rect 37526 2730 37531 2758
rect 1185 2646 1190 2674
rect 1218 2646 5446 2674
rect 5474 2646 5479 2674
rect 25937 2646 25942 2674
rect 25970 2646 27622 2674
rect 27650 2646 29358 2674
rect 29386 2646 29391 2674
rect 2473 2590 2478 2618
rect 2506 2590 3038 2618
rect 3066 2590 3542 2618
rect 3570 2590 4046 2618
rect 4074 2590 16870 2618
rect 16898 2590 16903 2618
rect 23921 2590 23926 2618
rect 23954 2590 28070 2618
rect 28098 2590 30142 2618
rect 30170 2590 30310 2618
rect 30338 2590 30343 2618
rect 1969 2534 1974 2562
rect 2002 2534 2366 2562
rect 2394 2534 4998 2562
rect 5026 2534 5726 2562
rect 5754 2534 5838 2562
rect 5866 2534 5871 2562
rect 6449 2534 6454 2562
rect 6482 2534 7014 2562
rect 7042 2534 7047 2562
rect 7569 2534 7574 2562
rect 7602 2534 8078 2562
rect 8106 2534 9366 2562
rect 9394 2534 9399 2562
rect 16753 2534 16758 2562
rect 16786 2534 18270 2562
rect 18298 2534 19502 2562
rect 19530 2534 19950 2562
rect 19978 2534 19983 2562
rect 21793 2534 21798 2562
rect 21826 2534 23422 2562
rect 23450 2534 23455 2562
rect 26217 2534 26222 2562
rect 26250 2534 26726 2562
rect 26754 2534 26759 2562
rect 27706 2534 28462 2562
rect 28490 2534 28742 2562
rect 28770 2534 28775 2562
rect 30697 2534 30702 2562
rect 30730 2534 32158 2562
rect 32186 2534 32606 2562
rect 32634 2534 32639 2562
rect 27706 2506 27734 2534
rect 8465 2478 8470 2506
rect 8498 2478 8974 2506
rect 9002 2478 9007 2506
rect 24425 2478 24430 2506
rect 24458 2478 24766 2506
rect 24794 2478 24799 2506
rect 26385 2478 26390 2506
rect 26418 2478 27734 2506
rect 33329 2478 33334 2506
rect 33362 2478 33838 2506
rect 33866 2478 35854 2506
rect 35882 2478 37646 2506
rect 37674 2478 37679 2506
rect 38201 2478 38206 2506
rect 38234 2478 39046 2506
rect 39074 2478 39079 2506
rect 3593 2422 3598 2450
rect 3626 2422 4102 2450
rect 4130 2422 9422 2450
rect 9450 2422 9455 2450
rect 24369 2422 24374 2450
rect 24402 2422 28966 2450
rect 28994 2422 28999 2450
rect 33945 2422 33950 2450
rect 33978 2422 36582 2450
rect 36610 2422 38150 2450
rect 38178 2422 38183 2450
rect 37585 2366 37590 2394
rect 37618 2366 38206 2394
rect 38234 2366 38239 2394
rect 4577 2338 4582 2366
rect 4610 2338 4634 2366
rect 4662 2338 4686 2366
rect 4714 2338 4738 2366
rect 4766 2338 4790 2366
rect 4818 2338 4842 2366
rect 4870 2338 4894 2366
rect 4922 2338 4946 2366
rect 4974 2338 4998 2366
rect 5026 2338 5031 2366
rect 9577 2338 9582 2366
rect 9610 2338 9634 2366
rect 9662 2338 9686 2366
rect 9714 2338 9738 2366
rect 9766 2338 9790 2366
rect 9818 2338 9842 2366
rect 9870 2338 9894 2366
rect 9922 2338 9946 2366
rect 9974 2338 9998 2366
rect 10026 2338 10031 2366
rect 14577 2338 14582 2366
rect 14610 2338 14634 2366
rect 14662 2338 14686 2366
rect 14714 2338 14738 2366
rect 14766 2338 14790 2366
rect 14818 2338 14842 2366
rect 14870 2338 14894 2366
rect 14922 2338 14946 2366
rect 14974 2338 14998 2366
rect 15026 2338 15031 2366
rect 19577 2338 19582 2366
rect 19610 2338 19634 2366
rect 19662 2338 19686 2366
rect 19714 2338 19738 2366
rect 19766 2338 19790 2366
rect 19818 2338 19842 2366
rect 19870 2338 19894 2366
rect 19922 2338 19946 2366
rect 19974 2338 19998 2366
rect 20026 2338 20031 2366
rect 24577 2338 24582 2366
rect 24610 2338 24634 2366
rect 24662 2338 24686 2366
rect 24714 2338 24738 2366
rect 24766 2338 24790 2366
rect 24818 2338 24842 2366
rect 24870 2338 24894 2366
rect 24922 2338 24946 2366
rect 24974 2338 24998 2366
rect 25026 2338 25031 2366
rect 29577 2338 29582 2366
rect 29610 2338 29634 2366
rect 29662 2338 29686 2366
rect 29714 2338 29738 2366
rect 29766 2338 29790 2366
rect 29818 2338 29842 2366
rect 29870 2338 29894 2366
rect 29922 2338 29946 2366
rect 29974 2338 29998 2366
rect 30026 2338 30031 2366
rect 34577 2338 34582 2366
rect 34610 2338 34634 2366
rect 34662 2338 34686 2366
rect 34714 2338 34738 2366
rect 34766 2338 34790 2366
rect 34818 2338 34842 2366
rect 34870 2338 34894 2366
rect 34922 2338 34946 2366
rect 34974 2338 34998 2366
rect 35026 2338 35031 2366
rect 2585 2254 2590 2282
rect 2618 2254 8246 2282
rect 8274 2254 8279 2282
rect 18097 2254 18102 2282
rect 18130 2254 24374 2282
rect 24402 2254 24407 2282
rect 26721 2254 26726 2282
rect 26754 2254 26950 2282
rect 26978 2254 36134 2282
rect 36162 2254 36694 2282
rect 36722 2254 36727 2282
rect 1633 2198 1638 2226
rect 1666 2198 4494 2226
rect 4522 2198 6342 2226
rect 6370 2198 6375 2226
rect 9473 2198 9478 2226
rect 9506 2198 10038 2226
rect 10066 2198 13062 2226
rect 13090 2198 13790 2226
rect 13818 2198 13823 2226
rect 27393 2198 27398 2226
rect 27426 2198 27678 2226
rect 27706 2198 27711 2226
rect 31985 2198 31990 2226
rect 32018 2198 32158 2226
rect 32186 2198 32326 2226
rect 32354 2198 33726 2226
rect 33754 2198 33759 2226
rect 35737 2198 35742 2226
rect 35770 2198 35910 2226
rect 35938 2198 37702 2226
rect 37730 2198 38262 2226
rect 38290 2198 38710 2226
rect 38738 2198 38878 2226
rect 38906 2198 38911 2226
rect 3033 2142 3038 2170
rect 3066 2142 5502 2170
rect 5530 2142 5535 2170
rect 10873 2142 10878 2170
rect 10906 2142 11382 2170
rect 11410 2142 11415 2170
rect 11769 2142 11774 2170
rect 11802 2142 11942 2170
rect 11970 2142 11975 2170
rect 14233 2142 14238 2170
rect 14266 2142 14462 2170
rect 14490 2142 16254 2170
rect 16282 2142 16287 2170
rect 24761 2142 24766 2170
rect 24794 2142 26222 2170
rect 26250 2142 26255 2170
rect 29409 2142 29414 2170
rect 29442 2142 29918 2170
rect 29946 2142 31262 2170
rect 31290 2142 31486 2170
rect 31514 2142 31519 2170
rect 32097 2142 32102 2170
rect 32130 2142 33670 2170
rect 33698 2142 35686 2170
rect 35714 2142 37534 2170
rect 37562 2142 37814 2170
rect 37842 2142 37847 2170
rect 38145 2142 38150 2170
rect 38178 2142 38934 2170
rect 38962 2142 38967 2170
rect 11774 2114 11802 2142
rect 4489 2086 4494 2114
rect 4522 2086 10542 2114
rect 10570 2086 10575 2114
rect 10817 2086 10822 2114
rect 10850 2086 11802 2114
rect 13785 2086 13790 2114
rect 13818 2086 20510 2114
rect 20538 2086 20790 2114
rect 20818 2086 21630 2114
rect 21658 2086 22246 2114
rect 22274 2086 22582 2114
rect 22610 2086 22615 2114
rect 28345 2086 28350 2114
rect 28378 2086 34118 2114
rect 34146 2086 38822 2114
rect 38850 2086 38855 2114
rect 7009 2030 7014 2058
rect 7042 2030 7518 2058
rect 7546 2030 19334 2058
rect 19362 2030 19367 2058
rect 2077 1946 2082 1974
rect 2110 1946 2134 1974
rect 2162 1946 2186 1974
rect 2214 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2394 1974
rect 2422 1946 2446 1974
rect 2474 1946 2498 1974
rect 2526 1946 2531 1974
rect 7077 1946 7082 1974
rect 7110 1946 7134 1974
rect 7162 1946 7186 1974
rect 7214 1946 7238 1974
rect 7266 1946 7290 1974
rect 7318 1946 7342 1974
rect 7370 1946 7394 1974
rect 7422 1946 7446 1974
rect 7474 1946 7498 1974
rect 7526 1946 7531 1974
rect 7574 1890 7602 2030
rect 12077 1946 12082 1974
rect 12110 1946 12134 1974
rect 12162 1946 12186 1974
rect 12214 1946 12238 1974
rect 12266 1946 12290 1974
rect 12318 1946 12342 1974
rect 12370 1946 12394 1974
rect 12422 1946 12446 1974
rect 12474 1946 12498 1974
rect 12526 1946 12531 1974
rect 17077 1946 17082 1974
rect 17110 1946 17134 1974
rect 17162 1946 17186 1974
rect 17214 1946 17238 1974
rect 17266 1946 17290 1974
rect 17318 1946 17342 1974
rect 17370 1946 17394 1974
rect 17422 1946 17446 1974
rect 17474 1946 17498 1974
rect 17526 1946 17531 1974
rect 22077 1946 22082 1974
rect 22110 1946 22134 1974
rect 22162 1946 22186 1974
rect 22214 1946 22238 1974
rect 22266 1946 22290 1974
rect 22318 1946 22342 1974
rect 22370 1946 22394 1974
rect 22422 1946 22446 1974
rect 22474 1946 22498 1974
rect 22526 1946 22531 1974
rect 27077 1946 27082 1974
rect 27110 1946 27134 1974
rect 27162 1946 27186 1974
rect 27214 1946 27238 1974
rect 27266 1946 27290 1974
rect 27318 1946 27342 1974
rect 27370 1946 27394 1974
rect 27422 1946 27446 1974
rect 27474 1946 27498 1974
rect 27526 1946 27531 1974
rect 32077 1946 32082 1974
rect 32110 1946 32134 1974
rect 32162 1946 32186 1974
rect 32214 1946 32238 1974
rect 32266 1946 32290 1974
rect 32318 1946 32342 1974
rect 32370 1946 32394 1974
rect 32422 1946 32446 1974
rect 32474 1946 32498 1974
rect 32526 1946 32531 1974
rect 37077 1946 37082 1974
rect 37110 1946 37134 1974
rect 37162 1946 37186 1974
rect 37214 1946 37238 1974
rect 37266 1946 37290 1974
rect 37318 1946 37342 1974
rect 37370 1946 37394 1974
rect 37422 1946 37446 1974
rect 37474 1946 37498 1974
rect 37526 1946 37531 1974
rect 2081 1862 2086 1890
rect 2114 1862 3934 1890
rect 3962 1862 3967 1890
rect 7457 1862 7462 1890
rect 7490 1862 7602 1890
rect 9361 1806 9366 1834
rect 9394 1806 10094 1834
rect 11377 1806 11382 1834
rect 11410 1806 20566 1834
rect 20594 1806 22470 1834
rect 22498 1806 24430 1834
rect 24458 1806 24766 1834
rect 24794 1806 24799 1834
rect 10066 1778 10094 1806
rect 8969 1750 8974 1778
rect 9002 1750 9702 1778
rect 9730 1750 9735 1778
rect 10066 1750 10710 1778
rect 10738 1750 10743 1778
rect 15577 1750 15582 1778
rect 15610 1750 15694 1778
rect 15722 1750 15727 1778
rect 28513 1750 28518 1778
rect 28546 1750 28966 1778
rect 28994 1750 30310 1778
rect 30338 1750 30343 1778
rect 31873 1750 31878 1778
rect 31906 1750 33446 1778
rect 33474 1750 34454 1778
rect 34482 1750 34487 1778
rect 35345 1750 35350 1778
rect 35378 1750 38934 1778
rect 38962 1750 39102 1778
rect 39130 1750 39135 1778
rect 6393 1694 6398 1722
rect 6426 1694 8358 1722
rect 8386 1694 13510 1722
rect 13538 1694 13734 1722
rect 13762 1694 14238 1722
rect 14266 1694 14271 1722
rect 19329 1694 19334 1722
rect 19362 1694 26390 1722
rect 26418 1694 26423 1722
rect 31481 1694 31486 1722
rect 31514 1694 35182 1722
rect 35210 1694 35215 1722
rect 5497 1638 5502 1666
rect 5530 1638 18102 1666
rect 18130 1638 18135 1666
rect 4577 1554 4582 1582
rect 4610 1554 4634 1582
rect 4662 1554 4686 1582
rect 4714 1554 4738 1582
rect 4766 1554 4790 1582
rect 4818 1554 4842 1582
rect 4870 1554 4894 1582
rect 4922 1554 4946 1582
rect 4974 1554 4998 1582
rect 5026 1554 5031 1582
rect 9577 1554 9582 1582
rect 9610 1554 9634 1582
rect 9662 1554 9686 1582
rect 9714 1554 9738 1582
rect 9766 1554 9790 1582
rect 9818 1554 9842 1582
rect 9870 1554 9894 1582
rect 9922 1554 9946 1582
rect 9974 1554 9998 1582
rect 10026 1554 10031 1582
rect 14577 1554 14582 1582
rect 14610 1554 14634 1582
rect 14662 1554 14686 1582
rect 14714 1554 14738 1582
rect 14766 1554 14790 1582
rect 14818 1554 14842 1582
rect 14870 1554 14894 1582
rect 14922 1554 14946 1582
rect 14974 1554 14998 1582
rect 15026 1554 15031 1582
rect 19577 1554 19582 1582
rect 19610 1554 19634 1582
rect 19662 1554 19686 1582
rect 19714 1554 19738 1582
rect 19766 1554 19790 1582
rect 19818 1554 19842 1582
rect 19870 1554 19894 1582
rect 19922 1554 19946 1582
rect 19974 1554 19998 1582
rect 20026 1554 20031 1582
rect 24577 1554 24582 1582
rect 24610 1554 24634 1582
rect 24662 1554 24686 1582
rect 24714 1554 24738 1582
rect 24766 1554 24790 1582
rect 24818 1554 24842 1582
rect 24870 1554 24894 1582
rect 24922 1554 24946 1582
rect 24974 1554 24998 1582
rect 25026 1554 25031 1582
rect 29577 1554 29582 1582
rect 29610 1554 29634 1582
rect 29662 1554 29686 1582
rect 29714 1554 29738 1582
rect 29766 1554 29790 1582
rect 29818 1554 29842 1582
rect 29870 1554 29894 1582
rect 29922 1554 29946 1582
rect 29974 1554 29998 1582
rect 30026 1554 30031 1582
rect 34577 1554 34582 1582
rect 34610 1554 34634 1582
rect 34662 1554 34686 1582
rect 34714 1554 34738 1582
rect 34766 1554 34790 1582
rect 34818 1554 34842 1582
rect 34870 1554 34894 1582
rect 34922 1554 34946 1582
rect 34974 1554 34998 1582
rect 35026 1554 35031 1582
<< via3 >>
rect 2082 18410 2110 18438
rect 2134 18410 2162 18438
rect 2186 18410 2214 18438
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 2394 18410 2422 18438
rect 2446 18410 2474 18438
rect 2498 18410 2526 18438
rect 7082 18410 7110 18438
rect 7134 18410 7162 18438
rect 7186 18410 7214 18438
rect 7238 18410 7266 18438
rect 7290 18410 7318 18438
rect 7342 18410 7370 18438
rect 7394 18410 7422 18438
rect 7446 18410 7474 18438
rect 7498 18410 7526 18438
rect 12082 18410 12110 18438
rect 12134 18410 12162 18438
rect 12186 18410 12214 18438
rect 12238 18410 12266 18438
rect 12290 18410 12318 18438
rect 12342 18410 12370 18438
rect 12394 18410 12422 18438
rect 12446 18410 12474 18438
rect 12498 18410 12526 18438
rect 17082 18410 17110 18438
rect 17134 18410 17162 18438
rect 17186 18410 17214 18438
rect 17238 18410 17266 18438
rect 17290 18410 17318 18438
rect 17342 18410 17370 18438
rect 17394 18410 17422 18438
rect 17446 18410 17474 18438
rect 17498 18410 17526 18438
rect 22082 18410 22110 18438
rect 22134 18410 22162 18438
rect 22186 18410 22214 18438
rect 22238 18410 22266 18438
rect 22290 18410 22318 18438
rect 22342 18410 22370 18438
rect 22394 18410 22422 18438
rect 22446 18410 22474 18438
rect 22498 18410 22526 18438
rect 27082 18410 27110 18438
rect 27134 18410 27162 18438
rect 27186 18410 27214 18438
rect 27238 18410 27266 18438
rect 27290 18410 27318 18438
rect 27342 18410 27370 18438
rect 27394 18410 27422 18438
rect 27446 18410 27474 18438
rect 27498 18410 27526 18438
rect 32082 18410 32110 18438
rect 32134 18410 32162 18438
rect 32186 18410 32214 18438
rect 32238 18410 32266 18438
rect 32290 18410 32318 18438
rect 32342 18410 32370 18438
rect 32394 18410 32422 18438
rect 32446 18410 32474 18438
rect 32498 18410 32526 18438
rect 37082 18410 37110 18438
rect 37134 18410 37162 18438
rect 37186 18410 37214 18438
rect 37238 18410 37266 18438
rect 37290 18410 37318 18438
rect 37342 18410 37370 18438
rect 37394 18410 37422 18438
rect 37446 18410 37474 18438
rect 37498 18410 37526 18438
rect 4582 18018 4610 18046
rect 4634 18018 4662 18046
rect 4686 18018 4714 18046
rect 4738 18018 4766 18046
rect 4790 18018 4818 18046
rect 4842 18018 4870 18046
rect 4894 18018 4922 18046
rect 4946 18018 4974 18046
rect 4998 18018 5026 18046
rect 9582 18018 9610 18046
rect 9634 18018 9662 18046
rect 9686 18018 9714 18046
rect 9738 18018 9766 18046
rect 9790 18018 9818 18046
rect 9842 18018 9870 18046
rect 9894 18018 9922 18046
rect 9946 18018 9974 18046
rect 9998 18018 10026 18046
rect 14582 18018 14610 18046
rect 14634 18018 14662 18046
rect 14686 18018 14714 18046
rect 14738 18018 14766 18046
rect 14790 18018 14818 18046
rect 14842 18018 14870 18046
rect 14894 18018 14922 18046
rect 14946 18018 14974 18046
rect 14998 18018 15026 18046
rect 19582 18018 19610 18046
rect 19634 18018 19662 18046
rect 19686 18018 19714 18046
rect 19738 18018 19766 18046
rect 19790 18018 19818 18046
rect 19842 18018 19870 18046
rect 19894 18018 19922 18046
rect 19946 18018 19974 18046
rect 19998 18018 20026 18046
rect 24582 18018 24610 18046
rect 24634 18018 24662 18046
rect 24686 18018 24714 18046
rect 24738 18018 24766 18046
rect 24790 18018 24818 18046
rect 24842 18018 24870 18046
rect 24894 18018 24922 18046
rect 24946 18018 24974 18046
rect 24998 18018 25026 18046
rect 29582 18018 29610 18046
rect 29634 18018 29662 18046
rect 29686 18018 29714 18046
rect 29738 18018 29766 18046
rect 29790 18018 29818 18046
rect 29842 18018 29870 18046
rect 29894 18018 29922 18046
rect 29946 18018 29974 18046
rect 29998 18018 30026 18046
rect 34582 18018 34610 18046
rect 34634 18018 34662 18046
rect 34686 18018 34714 18046
rect 34738 18018 34766 18046
rect 34790 18018 34818 18046
rect 34842 18018 34870 18046
rect 34894 18018 34922 18046
rect 34946 18018 34974 18046
rect 34998 18018 35026 18046
rect 2082 17626 2110 17654
rect 2134 17626 2162 17654
rect 2186 17626 2214 17654
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 2394 17626 2422 17654
rect 2446 17626 2474 17654
rect 2498 17626 2526 17654
rect 7082 17626 7110 17654
rect 7134 17626 7162 17654
rect 7186 17626 7214 17654
rect 7238 17626 7266 17654
rect 7290 17626 7318 17654
rect 7342 17626 7370 17654
rect 7394 17626 7422 17654
rect 7446 17626 7474 17654
rect 7498 17626 7526 17654
rect 12082 17626 12110 17654
rect 12134 17626 12162 17654
rect 12186 17626 12214 17654
rect 12238 17626 12266 17654
rect 12290 17626 12318 17654
rect 12342 17626 12370 17654
rect 12394 17626 12422 17654
rect 12446 17626 12474 17654
rect 12498 17626 12526 17654
rect 17082 17626 17110 17654
rect 17134 17626 17162 17654
rect 17186 17626 17214 17654
rect 17238 17626 17266 17654
rect 17290 17626 17318 17654
rect 17342 17626 17370 17654
rect 17394 17626 17422 17654
rect 17446 17626 17474 17654
rect 17498 17626 17526 17654
rect 22082 17626 22110 17654
rect 22134 17626 22162 17654
rect 22186 17626 22214 17654
rect 22238 17626 22266 17654
rect 22290 17626 22318 17654
rect 22342 17626 22370 17654
rect 22394 17626 22422 17654
rect 22446 17626 22474 17654
rect 22498 17626 22526 17654
rect 27082 17626 27110 17654
rect 27134 17626 27162 17654
rect 27186 17626 27214 17654
rect 27238 17626 27266 17654
rect 27290 17626 27318 17654
rect 27342 17626 27370 17654
rect 27394 17626 27422 17654
rect 27446 17626 27474 17654
rect 27498 17626 27526 17654
rect 32082 17626 32110 17654
rect 32134 17626 32162 17654
rect 32186 17626 32214 17654
rect 32238 17626 32266 17654
rect 32290 17626 32318 17654
rect 32342 17626 32370 17654
rect 32394 17626 32422 17654
rect 32446 17626 32474 17654
rect 32498 17626 32526 17654
rect 37082 17626 37110 17654
rect 37134 17626 37162 17654
rect 37186 17626 37214 17654
rect 37238 17626 37266 17654
rect 37290 17626 37318 17654
rect 37342 17626 37370 17654
rect 37394 17626 37422 17654
rect 37446 17626 37474 17654
rect 37498 17626 37526 17654
rect 4582 17234 4610 17262
rect 4634 17234 4662 17262
rect 4686 17234 4714 17262
rect 4738 17234 4766 17262
rect 4790 17234 4818 17262
rect 4842 17234 4870 17262
rect 4894 17234 4922 17262
rect 4946 17234 4974 17262
rect 4998 17234 5026 17262
rect 9582 17234 9610 17262
rect 9634 17234 9662 17262
rect 9686 17234 9714 17262
rect 9738 17234 9766 17262
rect 9790 17234 9818 17262
rect 9842 17234 9870 17262
rect 9894 17234 9922 17262
rect 9946 17234 9974 17262
rect 9998 17234 10026 17262
rect 14582 17234 14610 17262
rect 14634 17234 14662 17262
rect 14686 17234 14714 17262
rect 14738 17234 14766 17262
rect 14790 17234 14818 17262
rect 14842 17234 14870 17262
rect 14894 17234 14922 17262
rect 14946 17234 14974 17262
rect 14998 17234 15026 17262
rect 19582 17234 19610 17262
rect 19634 17234 19662 17262
rect 19686 17234 19714 17262
rect 19738 17234 19766 17262
rect 19790 17234 19818 17262
rect 19842 17234 19870 17262
rect 19894 17234 19922 17262
rect 19946 17234 19974 17262
rect 19998 17234 20026 17262
rect 24582 17234 24610 17262
rect 24634 17234 24662 17262
rect 24686 17234 24714 17262
rect 24738 17234 24766 17262
rect 24790 17234 24818 17262
rect 24842 17234 24870 17262
rect 24894 17234 24922 17262
rect 24946 17234 24974 17262
rect 24998 17234 25026 17262
rect 29582 17234 29610 17262
rect 29634 17234 29662 17262
rect 29686 17234 29714 17262
rect 29738 17234 29766 17262
rect 29790 17234 29818 17262
rect 29842 17234 29870 17262
rect 29894 17234 29922 17262
rect 29946 17234 29974 17262
rect 29998 17234 30026 17262
rect 34582 17234 34610 17262
rect 34634 17234 34662 17262
rect 34686 17234 34714 17262
rect 34738 17234 34766 17262
rect 34790 17234 34818 17262
rect 34842 17234 34870 17262
rect 34894 17234 34922 17262
rect 34946 17234 34974 17262
rect 34998 17234 35026 17262
rect 2082 16842 2110 16870
rect 2134 16842 2162 16870
rect 2186 16842 2214 16870
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 2394 16842 2422 16870
rect 2446 16842 2474 16870
rect 2498 16842 2526 16870
rect 7082 16842 7110 16870
rect 7134 16842 7162 16870
rect 7186 16842 7214 16870
rect 7238 16842 7266 16870
rect 7290 16842 7318 16870
rect 7342 16842 7370 16870
rect 7394 16842 7422 16870
rect 7446 16842 7474 16870
rect 7498 16842 7526 16870
rect 12082 16842 12110 16870
rect 12134 16842 12162 16870
rect 12186 16842 12214 16870
rect 12238 16842 12266 16870
rect 12290 16842 12318 16870
rect 12342 16842 12370 16870
rect 12394 16842 12422 16870
rect 12446 16842 12474 16870
rect 12498 16842 12526 16870
rect 17082 16842 17110 16870
rect 17134 16842 17162 16870
rect 17186 16842 17214 16870
rect 17238 16842 17266 16870
rect 17290 16842 17318 16870
rect 17342 16842 17370 16870
rect 17394 16842 17422 16870
rect 17446 16842 17474 16870
rect 17498 16842 17526 16870
rect 22082 16842 22110 16870
rect 22134 16842 22162 16870
rect 22186 16842 22214 16870
rect 22238 16842 22266 16870
rect 22290 16842 22318 16870
rect 22342 16842 22370 16870
rect 22394 16842 22422 16870
rect 22446 16842 22474 16870
rect 22498 16842 22526 16870
rect 27082 16842 27110 16870
rect 27134 16842 27162 16870
rect 27186 16842 27214 16870
rect 27238 16842 27266 16870
rect 27290 16842 27318 16870
rect 27342 16842 27370 16870
rect 27394 16842 27422 16870
rect 27446 16842 27474 16870
rect 27498 16842 27526 16870
rect 32082 16842 32110 16870
rect 32134 16842 32162 16870
rect 32186 16842 32214 16870
rect 32238 16842 32266 16870
rect 32290 16842 32318 16870
rect 32342 16842 32370 16870
rect 32394 16842 32422 16870
rect 32446 16842 32474 16870
rect 32498 16842 32526 16870
rect 37082 16842 37110 16870
rect 37134 16842 37162 16870
rect 37186 16842 37214 16870
rect 37238 16842 37266 16870
rect 37290 16842 37318 16870
rect 37342 16842 37370 16870
rect 37394 16842 37422 16870
rect 37446 16842 37474 16870
rect 37498 16842 37526 16870
rect 4582 16450 4610 16478
rect 4634 16450 4662 16478
rect 4686 16450 4714 16478
rect 4738 16450 4766 16478
rect 4790 16450 4818 16478
rect 4842 16450 4870 16478
rect 4894 16450 4922 16478
rect 4946 16450 4974 16478
rect 4998 16450 5026 16478
rect 9582 16450 9610 16478
rect 9634 16450 9662 16478
rect 9686 16450 9714 16478
rect 9738 16450 9766 16478
rect 9790 16450 9818 16478
rect 9842 16450 9870 16478
rect 9894 16450 9922 16478
rect 9946 16450 9974 16478
rect 9998 16450 10026 16478
rect 14582 16450 14610 16478
rect 14634 16450 14662 16478
rect 14686 16450 14714 16478
rect 14738 16450 14766 16478
rect 14790 16450 14818 16478
rect 14842 16450 14870 16478
rect 14894 16450 14922 16478
rect 14946 16450 14974 16478
rect 14998 16450 15026 16478
rect 19582 16450 19610 16478
rect 19634 16450 19662 16478
rect 19686 16450 19714 16478
rect 19738 16450 19766 16478
rect 19790 16450 19818 16478
rect 19842 16450 19870 16478
rect 19894 16450 19922 16478
rect 19946 16450 19974 16478
rect 19998 16450 20026 16478
rect 24582 16450 24610 16478
rect 24634 16450 24662 16478
rect 24686 16450 24714 16478
rect 24738 16450 24766 16478
rect 24790 16450 24818 16478
rect 24842 16450 24870 16478
rect 24894 16450 24922 16478
rect 24946 16450 24974 16478
rect 24998 16450 25026 16478
rect 29582 16450 29610 16478
rect 29634 16450 29662 16478
rect 29686 16450 29714 16478
rect 29738 16450 29766 16478
rect 29790 16450 29818 16478
rect 29842 16450 29870 16478
rect 29894 16450 29922 16478
rect 29946 16450 29974 16478
rect 29998 16450 30026 16478
rect 34582 16450 34610 16478
rect 34634 16450 34662 16478
rect 34686 16450 34714 16478
rect 34738 16450 34766 16478
rect 34790 16450 34818 16478
rect 34842 16450 34870 16478
rect 34894 16450 34922 16478
rect 34946 16450 34974 16478
rect 34998 16450 35026 16478
rect 2082 16058 2110 16086
rect 2134 16058 2162 16086
rect 2186 16058 2214 16086
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 2394 16058 2422 16086
rect 2446 16058 2474 16086
rect 2498 16058 2526 16086
rect 7082 16058 7110 16086
rect 7134 16058 7162 16086
rect 7186 16058 7214 16086
rect 7238 16058 7266 16086
rect 7290 16058 7318 16086
rect 7342 16058 7370 16086
rect 7394 16058 7422 16086
rect 7446 16058 7474 16086
rect 7498 16058 7526 16086
rect 12082 16058 12110 16086
rect 12134 16058 12162 16086
rect 12186 16058 12214 16086
rect 12238 16058 12266 16086
rect 12290 16058 12318 16086
rect 12342 16058 12370 16086
rect 12394 16058 12422 16086
rect 12446 16058 12474 16086
rect 12498 16058 12526 16086
rect 17082 16058 17110 16086
rect 17134 16058 17162 16086
rect 17186 16058 17214 16086
rect 17238 16058 17266 16086
rect 17290 16058 17318 16086
rect 17342 16058 17370 16086
rect 17394 16058 17422 16086
rect 17446 16058 17474 16086
rect 17498 16058 17526 16086
rect 22082 16058 22110 16086
rect 22134 16058 22162 16086
rect 22186 16058 22214 16086
rect 22238 16058 22266 16086
rect 22290 16058 22318 16086
rect 22342 16058 22370 16086
rect 22394 16058 22422 16086
rect 22446 16058 22474 16086
rect 22498 16058 22526 16086
rect 27082 16058 27110 16086
rect 27134 16058 27162 16086
rect 27186 16058 27214 16086
rect 27238 16058 27266 16086
rect 27290 16058 27318 16086
rect 27342 16058 27370 16086
rect 27394 16058 27422 16086
rect 27446 16058 27474 16086
rect 27498 16058 27526 16086
rect 32082 16058 32110 16086
rect 32134 16058 32162 16086
rect 32186 16058 32214 16086
rect 32238 16058 32266 16086
rect 32290 16058 32318 16086
rect 32342 16058 32370 16086
rect 32394 16058 32422 16086
rect 32446 16058 32474 16086
rect 32498 16058 32526 16086
rect 37082 16058 37110 16086
rect 37134 16058 37162 16086
rect 37186 16058 37214 16086
rect 37238 16058 37266 16086
rect 37290 16058 37318 16086
rect 37342 16058 37370 16086
rect 37394 16058 37422 16086
rect 37446 16058 37474 16086
rect 37498 16058 37526 16086
rect 4582 15666 4610 15694
rect 4634 15666 4662 15694
rect 4686 15666 4714 15694
rect 4738 15666 4766 15694
rect 4790 15666 4818 15694
rect 4842 15666 4870 15694
rect 4894 15666 4922 15694
rect 4946 15666 4974 15694
rect 4998 15666 5026 15694
rect 9582 15666 9610 15694
rect 9634 15666 9662 15694
rect 9686 15666 9714 15694
rect 9738 15666 9766 15694
rect 9790 15666 9818 15694
rect 9842 15666 9870 15694
rect 9894 15666 9922 15694
rect 9946 15666 9974 15694
rect 9998 15666 10026 15694
rect 14582 15666 14610 15694
rect 14634 15666 14662 15694
rect 14686 15666 14714 15694
rect 14738 15666 14766 15694
rect 14790 15666 14818 15694
rect 14842 15666 14870 15694
rect 14894 15666 14922 15694
rect 14946 15666 14974 15694
rect 14998 15666 15026 15694
rect 19582 15666 19610 15694
rect 19634 15666 19662 15694
rect 19686 15666 19714 15694
rect 19738 15666 19766 15694
rect 19790 15666 19818 15694
rect 19842 15666 19870 15694
rect 19894 15666 19922 15694
rect 19946 15666 19974 15694
rect 19998 15666 20026 15694
rect 24582 15666 24610 15694
rect 24634 15666 24662 15694
rect 24686 15666 24714 15694
rect 24738 15666 24766 15694
rect 24790 15666 24818 15694
rect 24842 15666 24870 15694
rect 24894 15666 24922 15694
rect 24946 15666 24974 15694
rect 24998 15666 25026 15694
rect 29582 15666 29610 15694
rect 29634 15666 29662 15694
rect 29686 15666 29714 15694
rect 29738 15666 29766 15694
rect 29790 15666 29818 15694
rect 29842 15666 29870 15694
rect 29894 15666 29922 15694
rect 29946 15666 29974 15694
rect 29998 15666 30026 15694
rect 34582 15666 34610 15694
rect 34634 15666 34662 15694
rect 34686 15666 34714 15694
rect 34738 15666 34766 15694
rect 34790 15666 34818 15694
rect 34842 15666 34870 15694
rect 34894 15666 34922 15694
rect 34946 15666 34974 15694
rect 34998 15666 35026 15694
rect 2082 15274 2110 15302
rect 2134 15274 2162 15302
rect 2186 15274 2214 15302
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 2394 15274 2422 15302
rect 2446 15274 2474 15302
rect 2498 15274 2526 15302
rect 7082 15274 7110 15302
rect 7134 15274 7162 15302
rect 7186 15274 7214 15302
rect 7238 15274 7266 15302
rect 7290 15274 7318 15302
rect 7342 15274 7370 15302
rect 7394 15274 7422 15302
rect 7446 15274 7474 15302
rect 7498 15274 7526 15302
rect 12082 15274 12110 15302
rect 12134 15274 12162 15302
rect 12186 15274 12214 15302
rect 12238 15274 12266 15302
rect 12290 15274 12318 15302
rect 12342 15274 12370 15302
rect 12394 15274 12422 15302
rect 12446 15274 12474 15302
rect 12498 15274 12526 15302
rect 17082 15274 17110 15302
rect 17134 15274 17162 15302
rect 17186 15274 17214 15302
rect 17238 15274 17266 15302
rect 17290 15274 17318 15302
rect 17342 15274 17370 15302
rect 17394 15274 17422 15302
rect 17446 15274 17474 15302
rect 17498 15274 17526 15302
rect 22082 15274 22110 15302
rect 22134 15274 22162 15302
rect 22186 15274 22214 15302
rect 22238 15274 22266 15302
rect 22290 15274 22318 15302
rect 22342 15274 22370 15302
rect 22394 15274 22422 15302
rect 22446 15274 22474 15302
rect 22498 15274 22526 15302
rect 27082 15274 27110 15302
rect 27134 15274 27162 15302
rect 27186 15274 27214 15302
rect 27238 15274 27266 15302
rect 27290 15274 27318 15302
rect 27342 15274 27370 15302
rect 27394 15274 27422 15302
rect 27446 15274 27474 15302
rect 27498 15274 27526 15302
rect 32082 15274 32110 15302
rect 32134 15274 32162 15302
rect 32186 15274 32214 15302
rect 32238 15274 32266 15302
rect 32290 15274 32318 15302
rect 32342 15274 32370 15302
rect 32394 15274 32422 15302
rect 32446 15274 32474 15302
rect 32498 15274 32526 15302
rect 37082 15274 37110 15302
rect 37134 15274 37162 15302
rect 37186 15274 37214 15302
rect 37238 15274 37266 15302
rect 37290 15274 37318 15302
rect 37342 15274 37370 15302
rect 37394 15274 37422 15302
rect 37446 15274 37474 15302
rect 37498 15274 37526 15302
rect 4582 14882 4610 14910
rect 4634 14882 4662 14910
rect 4686 14882 4714 14910
rect 4738 14882 4766 14910
rect 4790 14882 4818 14910
rect 4842 14882 4870 14910
rect 4894 14882 4922 14910
rect 4946 14882 4974 14910
rect 4998 14882 5026 14910
rect 9582 14882 9610 14910
rect 9634 14882 9662 14910
rect 9686 14882 9714 14910
rect 9738 14882 9766 14910
rect 9790 14882 9818 14910
rect 9842 14882 9870 14910
rect 9894 14882 9922 14910
rect 9946 14882 9974 14910
rect 9998 14882 10026 14910
rect 14582 14882 14610 14910
rect 14634 14882 14662 14910
rect 14686 14882 14714 14910
rect 14738 14882 14766 14910
rect 14790 14882 14818 14910
rect 14842 14882 14870 14910
rect 14894 14882 14922 14910
rect 14946 14882 14974 14910
rect 14998 14882 15026 14910
rect 19582 14882 19610 14910
rect 19634 14882 19662 14910
rect 19686 14882 19714 14910
rect 19738 14882 19766 14910
rect 19790 14882 19818 14910
rect 19842 14882 19870 14910
rect 19894 14882 19922 14910
rect 19946 14882 19974 14910
rect 19998 14882 20026 14910
rect 24582 14882 24610 14910
rect 24634 14882 24662 14910
rect 24686 14882 24714 14910
rect 24738 14882 24766 14910
rect 24790 14882 24818 14910
rect 24842 14882 24870 14910
rect 24894 14882 24922 14910
rect 24946 14882 24974 14910
rect 24998 14882 25026 14910
rect 29582 14882 29610 14910
rect 29634 14882 29662 14910
rect 29686 14882 29714 14910
rect 29738 14882 29766 14910
rect 29790 14882 29818 14910
rect 29842 14882 29870 14910
rect 29894 14882 29922 14910
rect 29946 14882 29974 14910
rect 29998 14882 30026 14910
rect 34582 14882 34610 14910
rect 34634 14882 34662 14910
rect 34686 14882 34714 14910
rect 34738 14882 34766 14910
rect 34790 14882 34818 14910
rect 34842 14882 34870 14910
rect 34894 14882 34922 14910
rect 34946 14882 34974 14910
rect 34998 14882 35026 14910
rect 2082 14490 2110 14518
rect 2134 14490 2162 14518
rect 2186 14490 2214 14518
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 2394 14490 2422 14518
rect 2446 14490 2474 14518
rect 2498 14490 2526 14518
rect 7082 14490 7110 14518
rect 7134 14490 7162 14518
rect 7186 14490 7214 14518
rect 7238 14490 7266 14518
rect 7290 14490 7318 14518
rect 7342 14490 7370 14518
rect 7394 14490 7422 14518
rect 7446 14490 7474 14518
rect 7498 14490 7526 14518
rect 12082 14490 12110 14518
rect 12134 14490 12162 14518
rect 12186 14490 12214 14518
rect 12238 14490 12266 14518
rect 12290 14490 12318 14518
rect 12342 14490 12370 14518
rect 12394 14490 12422 14518
rect 12446 14490 12474 14518
rect 12498 14490 12526 14518
rect 17082 14490 17110 14518
rect 17134 14490 17162 14518
rect 17186 14490 17214 14518
rect 17238 14490 17266 14518
rect 17290 14490 17318 14518
rect 17342 14490 17370 14518
rect 17394 14490 17422 14518
rect 17446 14490 17474 14518
rect 17498 14490 17526 14518
rect 22082 14490 22110 14518
rect 22134 14490 22162 14518
rect 22186 14490 22214 14518
rect 22238 14490 22266 14518
rect 22290 14490 22318 14518
rect 22342 14490 22370 14518
rect 22394 14490 22422 14518
rect 22446 14490 22474 14518
rect 22498 14490 22526 14518
rect 27082 14490 27110 14518
rect 27134 14490 27162 14518
rect 27186 14490 27214 14518
rect 27238 14490 27266 14518
rect 27290 14490 27318 14518
rect 27342 14490 27370 14518
rect 27394 14490 27422 14518
rect 27446 14490 27474 14518
rect 27498 14490 27526 14518
rect 32082 14490 32110 14518
rect 32134 14490 32162 14518
rect 32186 14490 32214 14518
rect 32238 14490 32266 14518
rect 32290 14490 32318 14518
rect 32342 14490 32370 14518
rect 32394 14490 32422 14518
rect 32446 14490 32474 14518
rect 32498 14490 32526 14518
rect 37082 14490 37110 14518
rect 37134 14490 37162 14518
rect 37186 14490 37214 14518
rect 37238 14490 37266 14518
rect 37290 14490 37318 14518
rect 37342 14490 37370 14518
rect 37394 14490 37422 14518
rect 37446 14490 37474 14518
rect 37498 14490 37526 14518
rect 4582 14098 4610 14126
rect 4634 14098 4662 14126
rect 4686 14098 4714 14126
rect 4738 14098 4766 14126
rect 4790 14098 4818 14126
rect 4842 14098 4870 14126
rect 4894 14098 4922 14126
rect 4946 14098 4974 14126
rect 4998 14098 5026 14126
rect 9582 14098 9610 14126
rect 9634 14098 9662 14126
rect 9686 14098 9714 14126
rect 9738 14098 9766 14126
rect 9790 14098 9818 14126
rect 9842 14098 9870 14126
rect 9894 14098 9922 14126
rect 9946 14098 9974 14126
rect 9998 14098 10026 14126
rect 14582 14098 14610 14126
rect 14634 14098 14662 14126
rect 14686 14098 14714 14126
rect 14738 14098 14766 14126
rect 14790 14098 14818 14126
rect 14842 14098 14870 14126
rect 14894 14098 14922 14126
rect 14946 14098 14974 14126
rect 14998 14098 15026 14126
rect 19582 14098 19610 14126
rect 19634 14098 19662 14126
rect 19686 14098 19714 14126
rect 19738 14098 19766 14126
rect 19790 14098 19818 14126
rect 19842 14098 19870 14126
rect 19894 14098 19922 14126
rect 19946 14098 19974 14126
rect 19998 14098 20026 14126
rect 24582 14098 24610 14126
rect 24634 14098 24662 14126
rect 24686 14098 24714 14126
rect 24738 14098 24766 14126
rect 24790 14098 24818 14126
rect 24842 14098 24870 14126
rect 24894 14098 24922 14126
rect 24946 14098 24974 14126
rect 24998 14098 25026 14126
rect 29582 14098 29610 14126
rect 29634 14098 29662 14126
rect 29686 14098 29714 14126
rect 29738 14098 29766 14126
rect 29790 14098 29818 14126
rect 29842 14098 29870 14126
rect 29894 14098 29922 14126
rect 29946 14098 29974 14126
rect 29998 14098 30026 14126
rect 34582 14098 34610 14126
rect 34634 14098 34662 14126
rect 34686 14098 34714 14126
rect 34738 14098 34766 14126
rect 34790 14098 34818 14126
rect 34842 14098 34870 14126
rect 34894 14098 34922 14126
rect 34946 14098 34974 14126
rect 34998 14098 35026 14126
rect 2082 13706 2110 13734
rect 2134 13706 2162 13734
rect 2186 13706 2214 13734
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 2394 13706 2422 13734
rect 2446 13706 2474 13734
rect 2498 13706 2526 13734
rect 7082 13706 7110 13734
rect 7134 13706 7162 13734
rect 7186 13706 7214 13734
rect 7238 13706 7266 13734
rect 7290 13706 7318 13734
rect 7342 13706 7370 13734
rect 7394 13706 7422 13734
rect 7446 13706 7474 13734
rect 7498 13706 7526 13734
rect 12082 13706 12110 13734
rect 12134 13706 12162 13734
rect 12186 13706 12214 13734
rect 12238 13706 12266 13734
rect 12290 13706 12318 13734
rect 12342 13706 12370 13734
rect 12394 13706 12422 13734
rect 12446 13706 12474 13734
rect 12498 13706 12526 13734
rect 17082 13706 17110 13734
rect 17134 13706 17162 13734
rect 17186 13706 17214 13734
rect 17238 13706 17266 13734
rect 17290 13706 17318 13734
rect 17342 13706 17370 13734
rect 17394 13706 17422 13734
rect 17446 13706 17474 13734
rect 17498 13706 17526 13734
rect 22082 13706 22110 13734
rect 22134 13706 22162 13734
rect 22186 13706 22214 13734
rect 22238 13706 22266 13734
rect 22290 13706 22318 13734
rect 22342 13706 22370 13734
rect 22394 13706 22422 13734
rect 22446 13706 22474 13734
rect 22498 13706 22526 13734
rect 27082 13706 27110 13734
rect 27134 13706 27162 13734
rect 27186 13706 27214 13734
rect 27238 13706 27266 13734
rect 27290 13706 27318 13734
rect 27342 13706 27370 13734
rect 27394 13706 27422 13734
rect 27446 13706 27474 13734
rect 27498 13706 27526 13734
rect 32082 13706 32110 13734
rect 32134 13706 32162 13734
rect 32186 13706 32214 13734
rect 32238 13706 32266 13734
rect 32290 13706 32318 13734
rect 32342 13706 32370 13734
rect 32394 13706 32422 13734
rect 32446 13706 32474 13734
rect 32498 13706 32526 13734
rect 37082 13706 37110 13734
rect 37134 13706 37162 13734
rect 37186 13706 37214 13734
rect 37238 13706 37266 13734
rect 37290 13706 37318 13734
rect 37342 13706 37370 13734
rect 37394 13706 37422 13734
rect 37446 13706 37474 13734
rect 37498 13706 37526 13734
rect 4582 13314 4610 13342
rect 4634 13314 4662 13342
rect 4686 13314 4714 13342
rect 4738 13314 4766 13342
rect 4790 13314 4818 13342
rect 4842 13314 4870 13342
rect 4894 13314 4922 13342
rect 4946 13314 4974 13342
rect 4998 13314 5026 13342
rect 9582 13314 9610 13342
rect 9634 13314 9662 13342
rect 9686 13314 9714 13342
rect 9738 13314 9766 13342
rect 9790 13314 9818 13342
rect 9842 13314 9870 13342
rect 9894 13314 9922 13342
rect 9946 13314 9974 13342
rect 9998 13314 10026 13342
rect 14582 13314 14610 13342
rect 14634 13314 14662 13342
rect 14686 13314 14714 13342
rect 14738 13314 14766 13342
rect 14790 13314 14818 13342
rect 14842 13314 14870 13342
rect 14894 13314 14922 13342
rect 14946 13314 14974 13342
rect 14998 13314 15026 13342
rect 19582 13314 19610 13342
rect 19634 13314 19662 13342
rect 19686 13314 19714 13342
rect 19738 13314 19766 13342
rect 19790 13314 19818 13342
rect 19842 13314 19870 13342
rect 19894 13314 19922 13342
rect 19946 13314 19974 13342
rect 19998 13314 20026 13342
rect 24582 13314 24610 13342
rect 24634 13314 24662 13342
rect 24686 13314 24714 13342
rect 24738 13314 24766 13342
rect 24790 13314 24818 13342
rect 24842 13314 24870 13342
rect 24894 13314 24922 13342
rect 24946 13314 24974 13342
rect 24998 13314 25026 13342
rect 29582 13314 29610 13342
rect 29634 13314 29662 13342
rect 29686 13314 29714 13342
rect 29738 13314 29766 13342
rect 29790 13314 29818 13342
rect 29842 13314 29870 13342
rect 29894 13314 29922 13342
rect 29946 13314 29974 13342
rect 29998 13314 30026 13342
rect 34582 13314 34610 13342
rect 34634 13314 34662 13342
rect 34686 13314 34714 13342
rect 34738 13314 34766 13342
rect 34790 13314 34818 13342
rect 34842 13314 34870 13342
rect 34894 13314 34922 13342
rect 34946 13314 34974 13342
rect 34998 13314 35026 13342
rect 2082 12922 2110 12950
rect 2134 12922 2162 12950
rect 2186 12922 2214 12950
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 2394 12922 2422 12950
rect 2446 12922 2474 12950
rect 2498 12922 2526 12950
rect 7082 12922 7110 12950
rect 7134 12922 7162 12950
rect 7186 12922 7214 12950
rect 7238 12922 7266 12950
rect 7290 12922 7318 12950
rect 7342 12922 7370 12950
rect 7394 12922 7422 12950
rect 7446 12922 7474 12950
rect 7498 12922 7526 12950
rect 12082 12922 12110 12950
rect 12134 12922 12162 12950
rect 12186 12922 12214 12950
rect 12238 12922 12266 12950
rect 12290 12922 12318 12950
rect 12342 12922 12370 12950
rect 12394 12922 12422 12950
rect 12446 12922 12474 12950
rect 12498 12922 12526 12950
rect 17082 12922 17110 12950
rect 17134 12922 17162 12950
rect 17186 12922 17214 12950
rect 17238 12922 17266 12950
rect 17290 12922 17318 12950
rect 17342 12922 17370 12950
rect 17394 12922 17422 12950
rect 17446 12922 17474 12950
rect 17498 12922 17526 12950
rect 22082 12922 22110 12950
rect 22134 12922 22162 12950
rect 22186 12922 22214 12950
rect 22238 12922 22266 12950
rect 22290 12922 22318 12950
rect 22342 12922 22370 12950
rect 22394 12922 22422 12950
rect 22446 12922 22474 12950
rect 22498 12922 22526 12950
rect 27082 12922 27110 12950
rect 27134 12922 27162 12950
rect 27186 12922 27214 12950
rect 27238 12922 27266 12950
rect 27290 12922 27318 12950
rect 27342 12922 27370 12950
rect 27394 12922 27422 12950
rect 27446 12922 27474 12950
rect 27498 12922 27526 12950
rect 32082 12922 32110 12950
rect 32134 12922 32162 12950
rect 32186 12922 32214 12950
rect 32238 12922 32266 12950
rect 32290 12922 32318 12950
rect 32342 12922 32370 12950
rect 32394 12922 32422 12950
rect 32446 12922 32474 12950
rect 32498 12922 32526 12950
rect 37082 12922 37110 12950
rect 37134 12922 37162 12950
rect 37186 12922 37214 12950
rect 37238 12922 37266 12950
rect 37290 12922 37318 12950
rect 37342 12922 37370 12950
rect 37394 12922 37422 12950
rect 37446 12922 37474 12950
rect 37498 12922 37526 12950
rect 4582 12530 4610 12558
rect 4634 12530 4662 12558
rect 4686 12530 4714 12558
rect 4738 12530 4766 12558
rect 4790 12530 4818 12558
rect 4842 12530 4870 12558
rect 4894 12530 4922 12558
rect 4946 12530 4974 12558
rect 4998 12530 5026 12558
rect 9582 12530 9610 12558
rect 9634 12530 9662 12558
rect 9686 12530 9714 12558
rect 9738 12530 9766 12558
rect 9790 12530 9818 12558
rect 9842 12530 9870 12558
rect 9894 12530 9922 12558
rect 9946 12530 9974 12558
rect 9998 12530 10026 12558
rect 14582 12530 14610 12558
rect 14634 12530 14662 12558
rect 14686 12530 14714 12558
rect 14738 12530 14766 12558
rect 14790 12530 14818 12558
rect 14842 12530 14870 12558
rect 14894 12530 14922 12558
rect 14946 12530 14974 12558
rect 14998 12530 15026 12558
rect 19582 12530 19610 12558
rect 19634 12530 19662 12558
rect 19686 12530 19714 12558
rect 19738 12530 19766 12558
rect 19790 12530 19818 12558
rect 19842 12530 19870 12558
rect 19894 12530 19922 12558
rect 19946 12530 19974 12558
rect 19998 12530 20026 12558
rect 24582 12530 24610 12558
rect 24634 12530 24662 12558
rect 24686 12530 24714 12558
rect 24738 12530 24766 12558
rect 24790 12530 24818 12558
rect 24842 12530 24870 12558
rect 24894 12530 24922 12558
rect 24946 12530 24974 12558
rect 24998 12530 25026 12558
rect 29582 12530 29610 12558
rect 29634 12530 29662 12558
rect 29686 12530 29714 12558
rect 29738 12530 29766 12558
rect 29790 12530 29818 12558
rect 29842 12530 29870 12558
rect 29894 12530 29922 12558
rect 29946 12530 29974 12558
rect 29998 12530 30026 12558
rect 34582 12530 34610 12558
rect 34634 12530 34662 12558
rect 34686 12530 34714 12558
rect 34738 12530 34766 12558
rect 34790 12530 34818 12558
rect 34842 12530 34870 12558
rect 34894 12530 34922 12558
rect 34946 12530 34974 12558
rect 34998 12530 35026 12558
rect 2082 12138 2110 12166
rect 2134 12138 2162 12166
rect 2186 12138 2214 12166
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 2394 12138 2422 12166
rect 2446 12138 2474 12166
rect 2498 12138 2526 12166
rect 7082 12138 7110 12166
rect 7134 12138 7162 12166
rect 7186 12138 7214 12166
rect 7238 12138 7266 12166
rect 7290 12138 7318 12166
rect 7342 12138 7370 12166
rect 7394 12138 7422 12166
rect 7446 12138 7474 12166
rect 7498 12138 7526 12166
rect 12082 12138 12110 12166
rect 12134 12138 12162 12166
rect 12186 12138 12214 12166
rect 12238 12138 12266 12166
rect 12290 12138 12318 12166
rect 12342 12138 12370 12166
rect 12394 12138 12422 12166
rect 12446 12138 12474 12166
rect 12498 12138 12526 12166
rect 17082 12138 17110 12166
rect 17134 12138 17162 12166
rect 17186 12138 17214 12166
rect 17238 12138 17266 12166
rect 17290 12138 17318 12166
rect 17342 12138 17370 12166
rect 17394 12138 17422 12166
rect 17446 12138 17474 12166
rect 17498 12138 17526 12166
rect 22082 12138 22110 12166
rect 22134 12138 22162 12166
rect 22186 12138 22214 12166
rect 22238 12138 22266 12166
rect 22290 12138 22318 12166
rect 22342 12138 22370 12166
rect 22394 12138 22422 12166
rect 22446 12138 22474 12166
rect 22498 12138 22526 12166
rect 27082 12138 27110 12166
rect 27134 12138 27162 12166
rect 27186 12138 27214 12166
rect 27238 12138 27266 12166
rect 27290 12138 27318 12166
rect 27342 12138 27370 12166
rect 27394 12138 27422 12166
rect 27446 12138 27474 12166
rect 27498 12138 27526 12166
rect 32082 12138 32110 12166
rect 32134 12138 32162 12166
rect 32186 12138 32214 12166
rect 32238 12138 32266 12166
rect 32290 12138 32318 12166
rect 32342 12138 32370 12166
rect 32394 12138 32422 12166
rect 32446 12138 32474 12166
rect 32498 12138 32526 12166
rect 37082 12138 37110 12166
rect 37134 12138 37162 12166
rect 37186 12138 37214 12166
rect 37238 12138 37266 12166
rect 37290 12138 37318 12166
rect 37342 12138 37370 12166
rect 37394 12138 37422 12166
rect 37446 12138 37474 12166
rect 37498 12138 37526 12166
rect 4582 11746 4610 11774
rect 4634 11746 4662 11774
rect 4686 11746 4714 11774
rect 4738 11746 4766 11774
rect 4790 11746 4818 11774
rect 4842 11746 4870 11774
rect 4894 11746 4922 11774
rect 4946 11746 4974 11774
rect 4998 11746 5026 11774
rect 9582 11746 9610 11774
rect 9634 11746 9662 11774
rect 9686 11746 9714 11774
rect 9738 11746 9766 11774
rect 9790 11746 9818 11774
rect 9842 11746 9870 11774
rect 9894 11746 9922 11774
rect 9946 11746 9974 11774
rect 9998 11746 10026 11774
rect 14582 11746 14610 11774
rect 14634 11746 14662 11774
rect 14686 11746 14714 11774
rect 14738 11746 14766 11774
rect 14790 11746 14818 11774
rect 14842 11746 14870 11774
rect 14894 11746 14922 11774
rect 14946 11746 14974 11774
rect 14998 11746 15026 11774
rect 19582 11746 19610 11774
rect 19634 11746 19662 11774
rect 19686 11746 19714 11774
rect 19738 11746 19766 11774
rect 19790 11746 19818 11774
rect 19842 11746 19870 11774
rect 19894 11746 19922 11774
rect 19946 11746 19974 11774
rect 19998 11746 20026 11774
rect 24582 11746 24610 11774
rect 24634 11746 24662 11774
rect 24686 11746 24714 11774
rect 24738 11746 24766 11774
rect 24790 11746 24818 11774
rect 24842 11746 24870 11774
rect 24894 11746 24922 11774
rect 24946 11746 24974 11774
rect 24998 11746 25026 11774
rect 29582 11746 29610 11774
rect 29634 11746 29662 11774
rect 29686 11746 29714 11774
rect 29738 11746 29766 11774
rect 29790 11746 29818 11774
rect 29842 11746 29870 11774
rect 29894 11746 29922 11774
rect 29946 11746 29974 11774
rect 29998 11746 30026 11774
rect 34582 11746 34610 11774
rect 34634 11746 34662 11774
rect 34686 11746 34714 11774
rect 34738 11746 34766 11774
rect 34790 11746 34818 11774
rect 34842 11746 34870 11774
rect 34894 11746 34922 11774
rect 34946 11746 34974 11774
rect 34998 11746 35026 11774
rect 2082 11354 2110 11382
rect 2134 11354 2162 11382
rect 2186 11354 2214 11382
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 2394 11354 2422 11382
rect 2446 11354 2474 11382
rect 2498 11354 2526 11382
rect 7082 11354 7110 11382
rect 7134 11354 7162 11382
rect 7186 11354 7214 11382
rect 7238 11354 7266 11382
rect 7290 11354 7318 11382
rect 7342 11354 7370 11382
rect 7394 11354 7422 11382
rect 7446 11354 7474 11382
rect 7498 11354 7526 11382
rect 12082 11354 12110 11382
rect 12134 11354 12162 11382
rect 12186 11354 12214 11382
rect 12238 11354 12266 11382
rect 12290 11354 12318 11382
rect 12342 11354 12370 11382
rect 12394 11354 12422 11382
rect 12446 11354 12474 11382
rect 12498 11354 12526 11382
rect 17082 11354 17110 11382
rect 17134 11354 17162 11382
rect 17186 11354 17214 11382
rect 17238 11354 17266 11382
rect 17290 11354 17318 11382
rect 17342 11354 17370 11382
rect 17394 11354 17422 11382
rect 17446 11354 17474 11382
rect 17498 11354 17526 11382
rect 22082 11354 22110 11382
rect 22134 11354 22162 11382
rect 22186 11354 22214 11382
rect 22238 11354 22266 11382
rect 22290 11354 22318 11382
rect 22342 11354 22370 11382
rect 22394 11354 22422 11382
rect 22446 11354 22474 11382
rect 22498 11354 22526 11382
rect 27082 11354 27110 11382
rect 27134 11354 27162 11382
rect 27186 11354 27214 11382
rect 27238 11354 27266 11382
rect 27290 11354 27318 11382
rect 27342 11354 27370 11382
rect 27394 11354 27422 11382
rect 27446 11354 27474 11382
rect 27498 11354 27526 11382
rect 32082 11354 32110 11382
rect 32134 11354 32162 11382
rect 32186 11354 32214 11382
rect 32238 11354 32266 11382
rect 32290 11354 32318 11382
rect 32342 11354 32370 11382
rect 32394 11354 32422 11382
rect 32446 11354 32474 11382
rect 32498 11354 32526 11382
rect 37082 11354 37110 11382
rect 37134 11354 37162 11382
rect 37186 11354 37214 11382
rect 37238 11354 37266 11382
rect 37290 11354 37318 11382
rect 37342 11354 37370 11382
rect 37394 11354 37422 11382
rect 37446 11354 37474 11382
rect 37498 11354 37526 11382
rect 4582 10962 4610 10990
rect 4634 10962 4662 10990
rect 4686 10962 4714 10990
rect 4738 10962 4766 10990
rect 4790 10962 4818 10990
rect 4842 10962 4870 10990
rect 4894 10962 4922 10990
rect 4946 10962 4974 10990
rect 4998 10962 5026 10990
rect 9582 10962 9610 10990
rect 9634 10962 9662 10990
rect 9686 10962 9714 10990
rect 9738 10962 9766 10990
rect 9790 10962 9818 10990
rect 9842 10962 9870 10990
rect 9894 10962 9922 10990
rect 9946 10962 9974 10990
rect 9998 10962 10026 10990
rect 14582 10962 14610 10990
rect 14634 10962 14662 10990
rect 14686 10962 14714 10990
rect 14738 10962 14766 10990
rect 14790 10962 14818 10990
rect 14842 10962 14870 10990
rect 14894 10962 14922 10990
rect 14946 10962 14974 10990
rect 14998 10962 15026 10990
rect 19582 10962 19610 10990
rect 19634 10962 19662 10990
rect 19686 10962 19714 10990
rect 19738 10962 19766 10990
rect 19790 10962 19818 10990
rect 19842 10962 19870 10990
rect 19894 10962 19922 10990
rect 19946 10962 19974 10990
rect 19998 10962 20026 10990
rect 24582 10962 24610 10990
rect 24634 10962 24662 10990
rect 24686 10962 24714 10990
rect 24738 10962 24766 10990
rect 24790 10962 24818 10990
rect 24842 10962 24870 10990
rect 24894 10962 24922 10990
rect 24946 10962 24974 10990
rect 24998 10962 25026 10990
rect 29582 10962 29610 10990
rect 29634 10962 29662 10990
rect 29686 10962 29714 10990
rect 29738 10962 29766 10990
rect 29790 10962 29818 10990
rect 29842 10962 29870 10990
rect 29894 10962 29922 10990
rect 29946 10962 29974 10990
rect 29998 10962 30026 10990
rect 34582 10962 34610 10990
rect 34634 10962 34662 10990
rect 34686 10962 34714 10990
rect 34738 10962 34766 10990
rect 34790 10962 34818 10990
rect 34842 10962 34870 10990
rect 34894 10962 34922 10990
rect 34946 10962 34974 10990
rect 34998 10962 35026 10990
rect 2082 10570 2110 10598
rect 2134 10570 2162 10598
rect 2186 10570 2214 10598
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 2394 10570 2422 10598
rect 2446 10570 2474 10598
rect 2498 10570 2526 10598
rect 7082 10570 7110 10598
rect 7134 10570 7162 10598
rect 7186 10570 7214 10598
rect 7238 10570 7266 10598
rect 7290 10570 7318 10598
rect 7342 10570 7370 10598
rect 7394 10570 7422 10598
rect 7446 10570 7474 10598
rect 7498 10570 7526 10598
rect 12082 10570 12110 10598
rect 12134 10570 12162 10598
rect 12186 10570 12214 10598
rect 12238 10570 12266 10598
rect 12290 10570 12318 10598
rect 12342 10570 12370 10598
rect 12394 10570 12422 10598
rect 12446 10570 12474 10598
rect 12498 10570 12526 10598
rect 17082 10570 17110 10598
rect 17134 10570 17162 10598
rect 17186 10570 17214 10598
rect 17238 10570 17266 10598
rect 17290 10570 17318 10598
rect 17342 10570 17370 10598
rect 17394 10570 17422 10598
rect 17446 10570 17474 10598
rect 17498 10570 17526 10598
rect 22082 10570 22110 10598
rect 22134 10570 22162 10598
rect 22186 10570 22214 10598
rect 22238 10570 22266 10598
rect 22290 10570 22318 10598
rect 22342 10570 22370 10598
rect 22394 10570 22422 10598
rect 22446 10570 22474 10598
rect 22498 10570 22526 10598
rect 27082 10570 27110 10598
rect 27134 10570 27162 10598
rect 27186 10570 27214 10598
rect 27238 10570 27266 10598
rect 27290 10570 27318 10598
rect 27342 10570 27370 10598
rect 27394 10570 27422 10598
rect 27446 10570 27474 10598
rect 27498 10570 27526 10598
rect 32082 10570 32110 10598
rect 32134 10570 32162 10598
rect 32186 10570 32214 10598
rect 32238 10570 32266 10598
rect 32290 10570 32318 10598
rect 32342 10570 32370 10598
rect 32394 10570 32422 10598
rect 32446 10570 32474 10598
rect 32498 10570 32526 10598
rect 37082 10570 37110 10598
rect 37134 10570 37162 10598
rect 37186 10570 37214 10598
rect 37238 10570 37266 10598
rect 37290 10570 37318 10598
rect 37342 10570 37370 10598
rect 37394 10570 37422 10598
rect 37446 10570 37474 10598
rect 37498 10570 37526 10598
rect 4582 10178 4610 10206
rect 4634 10178 4662 10206
rect 4686 10178 4714 10206
rect 4738 10178 4766 10206
rect 4790 10178 4818 10206
rect 4842 10178 4870 10206
rect 4894 10178 4922 10206
rect 4946 10178 4974 10206
rect 4998 10178 5026 10206
rect 9582 10178 9610 10206
rect 9634 10178 9662 10206
rect 9686 10178 9714 10206
rect 9738 10178 9766 10206
rect 9790 10178 9818 10206
rect 9842 10178 9870 10206
rect 9894 10178 9922 10206
rect 9946 10178 9974 10206
rect 9998 10178 10026 10206
rect 14582 10178 14610 10206
rect 14634 10178 14662 10206
rect 14686 10178 14714 10206
rect 14738 10178 14766 10206
rect 14790 10178 14818 10206
rect 14842 10178 14870 10206
rect 14894 10178 14922 10206
rect 14946 10178 14974 10206
rect 14998 10178 15026 10206
rect 19582 10178 19610 10206
rect 19634 10178 19662 10206
rect 19686 10178 19714 10206
rect 19738 10178 19766 10206
rect 19790 10178 19818 10206
rect 19842 10178 19870 10206
rect 19894 10178 19922 10206
rect 19946 10178 19974 10206
rect 19998 10178 20026 10206
rect 24582 10178 24610 10206
rect 24634 10178 24662 10206
rect 24686 10178 24714 10206
rect 24738 10178 24766 10206
rect 24790 10178 24818 10206
rect 24842 10178 24870 10206
rect 24894 10178 24922 10206
rect 24946 10178 24974 10206
rect 24998 10178 25026 10206
rect 29582 10178 29610 10206
rect 29634 10178 29662 10206
rect 29686 10178 29714 10206
rect 29738 10178 29766 10206
rect 29790 10178 29818 10206
rect 29842 10178 29870 10206
rect 29894 10178 29922 10206
rect 29946 10178 29974 10206
rect 29998 10178 30026 10206
rect 34582 10178 34610 10206
rect 34634 10178 34662 10206
rect 34686 10178 34714 10206
rect 34738 10178 34766 10206
rect 34790 10178 34818 10206
rect 34842 10178 34870 10206
rect 34894 10178 34922 10206
rect 34946 10178 34974 10206
rect 34998 10178 35026 10206
rect 2082 9786 2110 9814
rect 2134 9786 2162 9814
rect 2186 9786 2214 9814
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 2394 9786 2422 9814
rect 2446 9786 2474 9814
rect 2498 9786 2526 9814
rect 7082 9786 7110 9814
rect 7134 9786 7162 9814
rect 7186 9786 7214 9814
rect 7238 9786 7266 9814
rect 7290 9786 7318 9814
rect 7342 9786 7370 9814
rect 7394 9786 7422 9814
rect 7446 9786 7474 9814
rect 7498 9786 7526 9814
rect 12082 9786 12110 9814
rect 12134 9786 12162 9814
rect 12186 9786 12214 9814
rect 12238 9786 12266 9814
rect 12290 9786 12318 9814
rect 12342 9786 12370 9814
rect 12394 9786 12422 9814
rect 12446 9786 12474 9814
rect 12498 9786 12526 9814
rect 17082 9786 17110 9814
rect 17134 9786 17162 9814
rect 17186 9786 17214 9814
rect 17238 9786 17266 9814
rect 17290 9786 17318 9814
rect 17342 9786 17370 9814
rect 17394 9786 17422 9814
rect 17446 9786 17474 9814
rect 17498 9786 17526 9814
rect 22082 9786 22110 9814
rect 22134 9786 22162 9814
rect 22186 9786 22214 9814
rect 22238 9786 22266 9814
rect 22290 9786 22318 9814
rect 22342 9786 22370 9814
rect 22394 9786 22422 9814
rect 22446 9786 22474 9814
rect 22498 9786 22526 9814
rect 27082 9786 27110 9814
rect 27134 9786 27162 9814
rect 27186 9786 27214 9814
rect 27238 9786 27266 9814
rect 27290 9786 27318 9814
rect 27342 9786 27370 9814
rect 27394 9786 27422 9814
rect 27446 9786 27474 9814
rect 27498 9786 27526 9814
rect 32082 9786 32110 9814
rect 32134 9786 32162 9814
rect 32186 9786 32214 9814
rect 32238 9786 32266 9814
rect 32290 9786 32318 9814
rect 32342 9786 32370 9814
rect 32394 9786 32422 9814
rect 32446 9786 32474 9814
rect 32498 9786 32526 9814
rect 37082 9786 37110 9814
rect 37134 9786 37162 9814
rect 37186 9786 37214 9814
rect 37238 9786 37266 9814
rect 37290 9786 37318 9814
rect 37342 9786 37370 9814
rect 37394 9786 37422 9814
rect 37446 9786 37474 9814
rect 37498 9786 37526 9814
rect 4582 9394 4610 9422
rect 4634 9394 4662 9422
rect 4686 9394 4714 9422
rect 4738 9394 4766 9422
rect 4790 9394 4818 9422
rect 4842 9394 4870 9422
rect 4894 9394 4922 9422
rect 4946 9394 4974 9422
rect 4998 9394 5026 9422
rect 9582 9394 9610 9422
rect 9634 9394 9662 9422
rect 9686 9394 9714 9422
rect 9738 9394 9766 9422
rect 9790 9394 9818 9422
rect 9842 9394 9870 9422
rect 9894 9394 9922 9422
rect 9946 9394 9974 9422
rect 9998 9394 10026 9422
rect 14582 9394 14610 9422
rect 14634 9394 14662 9422
rect 14686 9394 14714 9422
rect 14738 9394 14766 9422
rect 14790 9394 14818 9422
rect 14842 9394 14870 9422
rect 14894 9394 14922 9422
rect 14946 9394 14974 9422
rect 14998 9394 15026 9422
rect 19582 9394 19610 9422
rect 19634 9394 19662 9422
rect 19686 9394 19714 9422
rect 19738 9394 19766 9422
rect 19790 9394 19818 9422
rect 19842 9394 19870 9422
rect 19894 9394 19922 9422
rect 19946 9394 19974 9422
rect 19998 9394 20026 9422
rect 24582 9394 24610 9422
rect 24634 9394 24662 9422
rect 24686 9394 24714 9422
rect 24738 9394 24766 9422
rect 24790 9394 24818 9422
rect 24842 9394 24870 9422
rect 24894 9394 24922 9422
rect 24946 9394 24974 9422
rect 24998 9394 25026 9422
rect 29582 9394 29610 9422
rect 29634 9394 29662 9422
rect 29686 9394 29714 9422
rect 29738 9394 29766 9422
rect 29790 9394 29818 9422
rect 29842 9394 29870 9422
rect 29894 9394 29922 9422
rect 29946 9394 29974 9422
rect 29998 9394 30026 9422
rect 34582 9394 34610 9422
rect 34634 9394 34662 9422
rect 34686 9394 34714 9422
rect 34738 9394 34766 9422
rect 34790 9394 34818 9422
rect 34842 9394 34870 9422
rect 34894 9394 34922 9422
rect 34946 9394 34974 9422
rect 34998 9394 35026 9422
rect 2082 9002 2110 9030
rect 2134 9002 2162 9030
rect 2186 9002 2214 9030
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 2394 9002 2422 9030
rect 2446 9002 2474 9030
rect 2498 9002 2526 9030
rect 7082 9002 7110 9030
rect 7134 9002 7162 9030
rect 7186 9002 7214 9030
rect 7238 9002 7266 9030
rect 7290 9002 7318 9030
rect 7342 9002 7370 9030
rect 7394 9002 7422 9030
rect 7446 9002 7474 9030
rect 7498 9002 7526 9030
rect 12082 9002 12110 9030
rect 12134 9002 12162 9030
rect 12186 9002 12214 9030
rect 12238 9002 12266 9030
rect 12290 9002 12318 9030
rect 12342 9002 12370 9030
rect 12394 9002 12422 9030
rect 12446 9002 12474 9030
rect 12498 9002 12526 9030
rect 17082 9002 17110 9030
rect 17134 9002 17162 9030
rect 17186 9002 17214 9030
rect 17238 9002 17266 9030
rect 17290 9002 17318 9030
rect 17342 9002 17370 9030
rect 17394 9002 17422 9030
rect 17446 9002 17474 9030
rect 17498 9002 17526 9030
rect 22082 9002 22110 9030
rect 22134 9002 22162 9030
rect 22186 9002 22214 9030
rect 22238 9002 22266 9030
rect 22290 9002 22318 9030
rect 22342 9002 22370 9030
rect 22394 9002 22422 9030
rect 22446 9002 22474 9030
rect 22498 9002 22526 9030
rect 27082 9002 27110 9030
rect 27134 9002 27162 9030
rect 27186 9002 27214 9030
rect 27238 9002 27266 9030
rect 27290 9002 27318 9030
rect 27342 9002 27370 9030
rect 27394 9002 27422 9030
rect 27446 9002 27474 9030
rect 27498 9002 27526 9030
rect 32082 9002 32110 9030
rect 32134 9002 32162 9030
rect 32186 9002 32214 9030
rect 32238 9002 32266 9030
rect 32290 9002 32318 9030
rect 32342 9002 32370 9030
rect 32394 9002 32422 9030
rect 32446 9002 32474 9030
rect 32498 9002 32526 9030
rect 37082 9002 37110 9030
rect 37134 9002 37162 9030
rect 37186 9002 37214 9030
rect 37238 9002 37266 9030
rect 37290 9002 37318 9030
rect 37342 9002 37370 9030
rect 37394 9002 37422 9030
rect 37446 9002 37474 9030
rect 37498 9002 37526 9030
rect 4582 8610 4610 8638
rect 4634 8610 4662 8638
rect 4686 8610 4714 8638
rect 4738 8610 4766 8638
rect 4790 8610 4818 8638
rect 4842 8610 4870 8638
rect 4894 8610 4922 8638
rect 4946 8610 4974 8638
rect 4998 8610 5026 8638
rect 9582 8610 9610 8638
rect 9634 8610 9662 8638
rect 9686 8610 9714 8638
rect 9738 8610 9766 8638
rect 9790 8610 9818 8638
rect 9842 8610 9870 8638
rect 9894 8610 9922 8638
rect 9946 8610 9974 8638
rect 9998 8610 10026 8638
rect 14582 8610 14610 8638
rect 14634 8610 14662 8638
rect 14686 8610 14714 8638
rect 14738 8610 14766 8638
rect 14790 8610 14818 8638
rect 14842 8610 14870 8638
rect 14894 8610 14922 8638
rect 14946 8610 14974 8638
rect 14998 8610 15026 8638
rect 19582 8610 19610 8638
rect 19634 8610 19662 8638
rect 19686 8610 19714 8638
rect 19738 8610 19766 8638
rect 19790 8610 19818 8638
rect 19842 8610 19870 8638
rect 19894 8610 19922 8638
rect 19946 8610 19974 8638
rect 19998 8610 20026 8638
rect 24582 8610 24610 8638
rect 24634 8610 24662 8638
rect 24686 8610 24714 8638
rect 24738 8610 24766 8638
rect 24790 8610 24818 8638
rect 24842 8610 24870 8638
rect 24894 8610 24922 8638
rect 24946 8610 24974 8638
rect 24998 8610 25026 8638
rect 29582 8610 29610 8638
rect 29634 8610 29662 8638
rect 29686 8610 29714 8638
rect 29738 8610 29766 8638
rect 29790 8610 29818 8638
rect 29842 8610 29870 8638
rect 29894 8610 29922 8638
rect 29946 8610 29974 8638
rect 29998 8610 30026 8638
rect 34582 8610 34610 8638
rect 34634 8610 34662 8638
rect 34686 8610 34714 8638
rect 34738 8610 34766 8638
rect 34790 8610 34818 8638
rect 34842 8610 34870 8638
rect 34894 8610 34922 8638
rect 34946 8610 34974 8638
rect 34998 8610 35026 8638
rect 2082 8218 2110 8246
rect 2134 8218 2162 8246
rect 2186 8218 2214 8246
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 2394 8218 2422 8246
rect 2446 8218 2474 8246
rect 2498 8218 2526 8246
rect 7082 8218 7110 8246
rect 7134 8218 7162 8246
rect 7186 8218 7214 8246
rect 7238 8218 7266 8246
rect 7290 8218 7318 8246
rect 7342 8218 7370 8246
rect 7394 8218 7422 8246
rect 7446 8218 7474 8246
rect 7498 8218 7526 8246
rect 12082 8218 12110 8246
rect 12134 8218 12162 8246
rect 12186 8218 12214 8246
rect 12238 8218 12266 8246
rect 12290 8218 12318 8246
rect 12342 8218 12370 8246
rect 12394 8218 12422 8246
rect 12446 8218 12474 8246
rect 12498 8218 12526 8246
rect 17082 8218 17110 8246
rect 17134 8218 17162 8246
rect 17186 8218 17214 8246
rect 17238 8218 17266 8246
rect 17290 8218 17318 8246
rect 17342 8218 17370 8246
rect 17394 8218 17422 8246
rect 17446 8218 17474 8246
rect 17498 8218 17526 8246
rect 22082 8218 22110 8246
rect 22134 8218 22162 8246
rect 22186 8218 22214 8246
rect 22238 8218 22266 8246
rect 22290 8218 22318 8246
rect 22342 8218 22370 8246
rect 22394 8218 22422 8246
rect 22446 8218 22474 8246
rect 22498 8218 22526 8246
rect 27082 8218 27110 8246
rect 27134 8218 27162 8246
rect 27186 8218 27214 8246
rect 27238 8218 27266 8246
rect 27290 8218 27318 8246
rect 27342 8218 27370 8246
rect 27394 8218 27422 8246
rect 27446 8218 27474 8246
rect 27498 8218 27526 8246
rect 32082 8218 32110 8246
rect 32134 8218 32162 8246
rect 32186 8218 32214 8246
rect 32238 8218 32266 8246
rect 32290 8218 32318 8246
rect 32342 8218 32370 8246
rect 32394 8218 32422 8246
rect 32446 8218 32474 8246
rect 32498 8218 32526 8246
rect 37082 8218 37110 8246
rect 37134 8218 37162 8246
rect 37186 8218 37214 8246
rect 37238 8218 37266 8246
rect 37290 8218 37318 8246
rect 37342 8218 37370 8246
rect 37394 8218 37422 8246
rect 37446 8218 37474 8246
rect 37498 8218 37526 8246
rect 4582 7826 4610 7854
rect 4634 7826 4662 7854
rect 4686 7826 4714 7854
rect 4738 7826 4766 7854
rect 4790 7826 4818 7854
rect 4842 7826 4870 7854
rect 4894 7826 4922 7854
rect 4946 7826 4974 7854
rect 4998 7826 5026 7854
rect 9582 7826 9610 7854
rect 9634 7826 9662 7854
rect 9686 7826 9714 7854
rect 9738 7826 9766 7854
rect 9790 7826 9818 7854
rect 9842 7826 9870 7854
rect 9894 7826 9922 7854
rect 9946 7826 9974 7854
rect 9998 7826 10026 7854
rect 14582 7826 14610 7854
rect 14634 7826 14662 7854
rect 14686 7826 14714 7854
rect 14738 7826 14766 7854
rect 14790 7826 14818 7854
rect 14842 7826 14870 7854
rect 14894 7826 14922 7854
rect 14946 7826 14974 7854
rect 14998 7826 15026 7854
rect 19582 7826 19610 7854
rect 19634 7826 19662 7854
rect 19686 7826 19714 7854
rect 19738 7826 19766 7854
rect 19790 7826 19818 7854
rect 19842 7826 19870 7854
rect 19894 7826 19922 7854
rect 19946 7826 19974 7854
rect 19998 7826 20026 7854
rect 24582 7826 24610 7854
rect 24634 7826 24662 7854
rect 24686 7826 24714 7854
rect 24738 7826 24766 7854
rect 24790 7826 24818 7854
rect 24842 7826 24870 7854
rect 24894 7826 24922 7854
rect 24946 7826 24974 7854
rect 24998 7826 25026 7854
rect 29582 7826 29610 7854
rect 29634 7826 29662 7854
rect 29686 7826 29714 7854
rect 29738 7826 29766 7854
rect 29790 7826 29818 7854
rect 29842 7826 29870 7854
rect 29894 7826 29922 7854
rect 29946 7826 29974 7854
rect 29998 7826 30026 7854
rect 34582 7826 34610 7854
rect 34634 7826 34662 7854
rect 34686 7826 34714 7854
rect 34738 7826 34766 7854
rect 34790 7826 34818 7854
rect 34842 7826 34870 7854
rect 34894 7826 34922 7854
rect 34946 7826 34974 7854
rect 34998 7826 35026 7854
rect 2082 7434 2110 7462
rect 2134 7434 2162 7462
rect 2186 7434 2214 7462
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 2394 7434 2422 7462
rect 2446 7434 2474 7462
rect 2498 7434 2526 7462
rect 7082 7434 7110 7462
rect 7134 7434 7162 7462
rect 7186 7434 7214 7462
rect 7238 7434 7266 7462
rect 7290 7434 7318 7462
rect 7342 7434 7370 7462
rect 7394 7434 7422 7462
rect 7446 7434 7474 7462
rect 7498 7434 7526 7462
rect 12082 7434 12110 7462
rect 12134 7434 12162 7462
rect 12186 7434 12214 7462
rect 12238 7434 12266 7462
rect 12290 7434 12318 7462
rect 12342 7434 12370 7462
rect 12394 7434 12422 7462
rect 12446 7434 12474 7462
rect 12498 7434 12526 7462
rect 17082 7434 17110 7462
rect 17134 7434 17162 7462
rect 17186 7434 17214 7462
rect 17238 7434 17266 7462
rect 17290 7434 17318 7462
rect 17342 7434 17370 7462
rect 17394 7434 17422 7462
rect 17446 7434 17474 7462
rect 17498 7434 17526 7462
rect 22082 7434 22110 7462
rect 22134 7434 22162 7462
rect 22186 7434 22214 7462
rect 22238 7434 22266 7462
rect 22290 7434 22318 7462
rect 22342 7434 22370 7462
rect 22394 7434 22422 7462
rect 22446 7434 22474 7462
rect 22498 7434 22526 7462
rect 27082 7434 27110 7462
rect 27134 7434 27162 7462
rect 27186 7434 27214 7462
rect 27238 7434 27266 7462
rect 27290 7434 27318 7462
rect 27342 7434 27370 7462
rect 27394 7434 27422 7462
rect 27446 7434 27474 7462
rect 27498 7434 27526 7462
rect 32082 7434 32110 7462
rect 32134 7434 32162 7462
rect 32186 7434 32214 7462
rect 32238 7434 32266 7462
rect 32290 7434 32318 7462
rect 32342 7434 32370 7462
rect 32394 7434 32422 7462
rect 32446 7434 32474 7462
rect 32498 7434 32526 7462
rect 37082 7434 37110 7462
rect 37134 7434 37162 7462
rect 37186 7434 37214 7462
rect 37238 7434 37266 7462
rect 37290 7434 37318 7462
rect 37342 7434 37370 7462
rect 37394 7434 37422 7462
rect 37446 7434 37474 7462
rect 37498 7434 37526 7462
rect 4582 7042 4610 7070
rect 4634 7042 4662 7070
rect 4686 7042 4714 7070
rect 4738 7042 4766 7070
rect 4790 7042 4818 7070
rect 4842 7042 4870 7070
rect 4894 7042 4922 7070
rect 4946 7042 4974 7070
rect 4998 7042 5026 7070
rect 9582 7042 9610 7070
rect 9634 7042 9662 7070
rect 9686 7042 9714 7070
rect 9738 7042 9766 7070
rect 9790 7042 9818 7070
rect 9842 7042 9870 7070
rect 9894 7042 9922 7070
rect 9946 7042 9974 7070
rect 9998 7042 10026 7070
rect 14582 7042 14610 7070
rect 14634 7042 14662 7070
rect 14686 7042 14714 7070
rect 14738 7042 14766 7070
rect 14790 7042 14818 7070
rect 14842 7042 14870 7070
rect 14894 7042 14922 7070
rect 14946 7042 14974 7070
rect 14998 7042 15026 7070
rect 19582 7042 19610 7070
rect 19634 7042 19662 7070
rect 19686 7042 19714 7070
rect 19738 7042 19766 7070
rect 19790 7042 19818 7070
rect 19842 7042 19870 7070
rect 19894 7042 19922 7070
rect 19946 7042 19974 7070
rect 19998 7042 20026 7070
rect 24582 7042 24610 7070
rect 24634 7042 24662 7070
rect 24686 7042 24714 7070
rect 24738 7042 24766 7070
rect 24790 7042 24818 7070
rect 24842 7042 24870 7070
rect 24894 7042 24922 7070
rect 24946 7042 24974 7070
rect 24998 7042 25026 7070
rect 29582 7042 29610 7070
rect 29634 7042 29662 7070
rect 29686 7042 29714 7070
rect 29738 7042 29766 7070
rect 29790 7042 29818 7070
rect 29842 7042 29870 7070
rect 29894 7042 29922 7070
rect 29946 7042 29974 7070
rect 29998 7042 30026 7070
rect 34582 7042 34610 7070
rect 34634 7042 34662 7070
rect 34686 7042 34714 7070
rect 34738 7042 34766 7070
rect 34790 7042 34818 7070
rect 34842 7042 34870 7070
rect 34894 7042 34922 7070
rect 34946 7042 34974 7070
rect 34998 7042 35026 7070
rect 2082 6650 2110 6678
rect 2134 6650 2162 6678
rect 2186 6650 2214 6678
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 2394 6650 2422 6678
rect 2446 6650 2474 6678
rect 2498 6650 2526 6678
rect 7082 6650 7110 6678
rect 7134 6650 7162 6678
rect 7186 6650 7214 6678
rect 7238 6650 7266 6678
rect 7290 6650 7318 6678
rect 7342 6650 7370 6678
rect 7394 6650 7422 6678
rect 7446 6650 7474 6678
rect 7498 6650 7526 6678
rect 12082 6650 12110 6678
rect 12134 6650 12162 6678
rect 12186 6650 12214 6678
rect 12238 6650 12266 6678
rect 12290 6650 12318 6678
rect 12342 6650 12370 6678
rect 12394 6650 12422 6678
rect 12446 6650 12474 6678
rect 12498 6650 12526 6678
rect 17082 6650 17110 6678
rect 17134 6650 17162 6678
rect 17186 6650 17214 6678
rect 17238 6650 17266 6678
rect 17290 6650 17318 6678
rect 17342 6650 17370 6678
rect 17394 6650 17422 6678
rect 17446 6650 17474 6678
rect 17498 6650 17526 6678
rect 22082 6650 22110 6678
rect 22134 6650 22162 6678
rect 22186 6650 22214 6678
rect 22238 6650 22266 6678
rect 22290 6650 22318 6678
rect 22342 6650 22370 6678
rect 22394 6650 22422 6678
rect 22446 6650 22474 6678
rect 22498 6650 22526 6678
rect 27082 6650 27110 6678
rect 27134 6650 27162 6678
rect 27186 6650 27214 6678
rect 27238 6650 27266 6678
rect 27290 6650 27318 6678
rect 27342 6650 27370 6678
rect 27394 6650 27422 6678
rect 27446 6650 27474 6678
rect 27498 6650 27526 6678
rect 32082 6650 32110 6678
rect 32134 6650 32162 6678
rect 32186 6650 32214 6678
rect 32238 6650 32266 6678
rect 32290 6650 32318 6678
rect 32342 6650 32370 6678
rect 32394 6650 32422 6678
rect 32446 6650 32474 6678
rect 32498 6650 32526 6678
rect 37082 6650 37110 6678
rect 37134 6650 37162 6678
rect 37186 6650 37214 6678
rect 37238 6650 37266 6678
rect 37290 6650 37318 6678
rect 37342 6650 37370 6678
rect 37394 6650 37422 6678
rect 37446 6650 37474 6678
rect 37498 6650 37526 6678
rect 4582 6258 4610 6286
rect 4634 6258 4662 6286
rect 4686 6258 4714 6286
rect 4738 6258 4766 6286
rect 4790 6258 4818 6286
rect 4842 6258 4870 6286
rect 4894 6258 4922 6286
rect 4946 6258 4974 6286
rect 4998 6258 5026 6286
rect 9582 6258 9610 6286
rect 9634 6258 9662 6286
rect 9686 6258 9714 6286
rect 9738 6258 9766 6286
rect 9790 6258 9818 6286
rect 9842 6258 9870 6286
rect 9894 6258 9922 6286
rect 9946 6258 9974 6286
rect 9998 6258 10026 6286
rect 14582 6258 14610 6286
rect 14634 6258 14662 6286
rect 14686 6258 14714 6286
rect 14738 6258 14766 6286
rect 14790 6258 14818 6286
rect 14842 6258 14870 6286
rect 14894 6258 14922 6286
rect 14946 6258 14974 6286
rect 14998 6258 15026 6286
rect 19582 6258 19610 6286
rect 19634 6258 19662 6286
rect 19686 6258 19714 6286
rect 19738 6258 19766 6286
rect 19790 6258 19818 6286
rect 19842 6258 19870 6286
rect 19894 6258 19922 6286
rect 19946 6258 19974 6286
rect 19998 6258 20026 6286
rect 24582 6258 24610 6286
rect 24634 6258 24662 6286
rect 24686 6258 24714 6286
rect 24738 6258 24766 6286
rect 24790 6258 24818 6286
rect 24842 6258 24870 6286
rect 24894 6258 24922 6286
rect 24946 6258 24974 6286
rect 24998 6258 25026 6286
rect 29582 6258 29610 6286
rect 29634 6258 29662 6286
rect 29686 6258 29714 6286
rect 29738 6258 29766 6286
rect 29790 6258 29818 6286
rect 29842 6258 29870 6286
rect 29894 6258 29922 6286
rect 29946 6258 29974 6286
rect 29998 6258 30026 6286
rect 34582 6258 34610 6286
rect 34634 6258 34662 6286
rect 34686 6258 34714 6286
rect 34738 6258 34766 6286
rect 34790 6258 34818 6286
rect 34842 6258 34870 6286
rect 34894 6258 34922 6286
rect 34946 6258 34974 6286
rect 34998 6258 35026 6286
rect 2082 5866 2110 5894
rect 2134 5866 2162 5894
rect 2186 5866 2214 5894
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 2394 5866 2422 5894
rect 2446 5866 2474 5894
rect 2498 5866 2526 5894
rect 7082 5866 7110 5894
rect 7134 5866 7162 5894
rect 7186 5866 7214 5894
rect 7238 5866 7266 5894
rect 7290 5866 7318 5894
rect 7342 5866 7370 5894
rect 7394 5866 7422 5894
rect 7446 5866 7474 5894
rect 7498 5866 7526 5894
rect 12082 5866 12110 5894
rect 12134 5866 12162 5894
rect 12186 5866 12214 5894
rect 12238 5866 12266 5894
rect 12290 5866 12318 5894
rect 12342 5866 12370 5894
rect 12394 5866 12422 5894
rect 12446 5866 12474 5894
rect 12498 5866 12526 5894
rect 17082 5866 17110 5894
rect 17134 5866 17162 5894
rect 17186 5866 17214 5894
rect 17238 5866 17266 5894
rect 17290 5866 17318 5894
rect 17342 5866 17370 5894
rect 17394 5866 17422 5894
rect 17446 5866 17474 5894
rect 17498 5866 17526 5894
rect 22082 5866 22110 5894
rect 22134 5866 22162 5894
rect 22186 5866 22214 5894
rect 22238 5866 22266 5894
rect 22290 5866 22318 5894
rect 22342 5866 22370 5894
rect 22394 5866 22422 5894
rect 22446 5866 22474 5894
rect 22498 5866 22526 5894
rect 27082 5866 27110 5894
rect 27134 5866 27162 5894
rect 27186 5866 27214 5894
rect 27238 5866 27266 5894
rect 27290 5866 27318 5894
rect 27342 5866 27370 5894
rect 27394 5866 27422 5894
rect 27446 5866 27474 5894
rect 27498 5866 27526 5894
rect 32082 5866 32110 5894
rect 32134 5866 32162 5894
rect 32186 5866 32214 5894
rect 32238 5866 32266 5894
rect 32290 5866 32318 5894
rect 32342 5866 32370 5894
rect 32394 5866 32422 5894
rect 32446 5866 32474 5894
rect 32498 5866 32526 5894
rect 37082 5866 37110 5894
rect 37134 5866 37162 5894
rect 37186 5866 37214 5894
rect 37238 5866 37266 5894
rect 37290 5866 37318 5894
rect 37342 5866 37370 5894
rect 37394 5866 37422 5894
rect 37446 5866 37474 5894
rect 37498 5866 37526 5894
rect 4582 5474 4610 5502
rect 4634 5474 4662 5502
rect 4686 5474 4714 5502
rect 4738 5474 4766 5502
rect 4790 5474 4818 5502
rect 4842 5474 4870 5502
rect 4894 5474 4922 5502
rect 4946 5474 4974 5502
rect 4998 5474 5026 5502
rect 9582 5474 9610 5502
rect 9634 5474 9662 5502
rect 9686 5474 9714 5502
rect 9738 5474 9766 5502
rect 9790 5474 9818 5502
rect 9842 5474 9870 5502
rect 9894 5474 9922 5502
rect 9946 5474 9974 5502
rect 9998 5474 10026 5502
rect 14582 5474 14610 5502
rect 14634 5474 14662 5502
rect 14686 5474 14714 5502
rect 14738 5474 14766 5502
rect 14790 5474 14818 5502
rect 14842 5474 14870 5502
rect 14894 5474 14922 5502
rect 14946 5474 14974 5502
rect 14998 5474 15026 5502
rect 19582 5474 19610 5502
rect 19634 5474 19662 5502
rect 19686 5474 19714 5502
rect 19738 5474 19766 5502
rect 19790 5474 19818 5502
rect 19842 5474 19870 5502
rect 19894 5474 19922 5502
rect 19946 5474 19974 5502
rect 19998 5474 20026 5502
rect 24582 5474 24610 5502
rect 24634 5474 24662 5502
rect 24686 5474 24714 5502
rect 24738 5474 24766 5502
rect 24790 5474 24818 5502
rect 24842 5474 24870 5502
rect 24894 5474 24922 5502
rect 24946 5474 24974 5502
rect 24998 5474 25026 5502
rect 29582 5474 29610 5502
rect 29634 5474 29662 5502
rect 29686 5474 29714 5502
rect 29738 5474 29766 5502
rect 29790 5474 29818 5502
rect 29842 5474 29870 5502
rect 29894 5474 29922 5502
rect 29946 5474 29974 5502
rect 29998 5474 30026 5502
rect 34582 5474 34610 5502
rect 34634 5474 34662 5502
rect 34686 5474 34714 5502
rect 34738 5474 34766 5502
rect 34790 5474 34818 5502
rect 34842 5474 34870 5502
rect 34894 5474 34922 5502
rect 34946 5474 34974 5502
rect 34998 5474 35026 5502
rect 2082 5082 2110 5110
rect 2134 5082 2162 5110
rect 2186 5082 2214 5110
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 2394 5082 2422 5110
rect 2446 5082 2474 5110
rect 2498 5082 2526 5110
rect 7082 5082 7110 5110
rect 7134 5082 7162 5110
rect 7186 5082 7214 5110
rect 7238 5082 7266 5110
rect 7290 5082 7318 5110
rect 7342 5082 7370 5110
rect 7394 5082 7422 5110
rect 7446 5082 7474 5110
rect 7498 5082 7526 5110
rect 12082 5082 12110 5110
rect 12134 5082 12162 5110
rect 12186 5082 12214 5110
rect 12238 5082 12266 5110
rect 12290 5082 12318 5110
rect 12342 5082 12370 5110
rect 12394 5082 12422 5110
rect 12446 5082 12474 5110
rect 12498 5082 12526 5110
rect 17082 5082 17110 5110
rect 17134 5082 17162 5110
rect 17186 5082 17214 5110
rect 17238 5082 17266 5110
rect 17290 5082 17318 5110
rect 17342 5082 17370 5110
rect 17394 5082 17422 5110
rect 17446 5082 17474 5110
rect 17498 5082 17526 5110
rect 22082 5082 22110 5110
rect 22134 5082 22162 5110
rect 22186 5082 22214 5110
rect 22238 5082 22266 5110
rect 22290 5082 22318 5110
rect 22342 5082 22370 5110
rect 22394 5082 22422 5110
rect 22446 5082 22474 5110
rect 22498 5082 22526 5110
rect 27082 5082 27110 5110
rect 27134 5082 27162 5110
rect 27186 5082 27214 5110
rect 27238 5082 27266 5110
rect 27290 5082 27318 5110
rect 27342 5082 27370 5110
rect 27394 5082 27422 5110
rect 27446 5082 27474 5110
rect 27498 5082 27526 5110
rect 32082 5082 32110 5110
rect 32134 5082 32162 5110
rect 32186 5082 32214 5110
rect 32238 5082 32266 5110
rect 32290 5082 32318 5110
rect 32342 5082 32370 5110
rect 32394 5082 32422 5110
rect 32446 5082 32474 5110
rect 32498 5082 32526 5110
rect 37082 5082 37110 5110
rect 37134 5082 37162 5110
rect 37186 5082 37214 5110
rect 37238 5082 37266 5110
rect 37290 5082 37318 5110
rect 37342 5082 37370 5110
rect 37394 5082 37422 5110
rect 37446 5082 37474 5110
rect 37498 5082 37526 5110
rect 4582 4690 4610 4718
rect 4634 4690 4662 4718
rect 4686 4690 4714 4718
rect 4738 4690 4766 4718
rect 4790 4690 4818 4718
rect 4842 4690 4870 4718
rect 4894 4690 4922 4718
rect 4946 4690 4974 4718
rect 4998 4690 5026 4718
rect 9582 4690 9610 4718
rect 9634 4690 9662 4718
rect 9686 4690 9714 4718
rect 9738 4690 9766 4718
rect 9790 4690 9818 4718
rect 9842 4690 9870 4718
rect 9894 4690 9922 4718
rect 9946 4690 9974 4718
rect 9998 4690 10026 4718
rect 14582 4690 14610 4718
rect 14634 4690 14662 4718
rect 14686 4690 14714 4718
rect 14738 4690 14766 4718
rect 14790 4690 14818 4718
rect 14842 4690 14870 4718
rect 14894 4690 14922 4718
rect 14946 4690 14974 4718
rect 14998 4690 15026 4718
rect 19582 4690 19610 4718
rect 19634 4690 19662 4718
rect 19686 4690 19714 4718
rect 19738 4690 19766 4718
rect 19790 4690 19818 4718
rect 19842 4690 19870 4718
rect 19894 4690 19922 4718
rect 19946 4690 19974 4718
rect 19998 4690 20026 4718
rect 24582 4690 24610 4718
rect 24634 4690 24662 4718
rect 24686 4690 24714 4718
rect 24738 4690 24766 4718
rect 24790 4690 24818 4718
rect 24842 4690 24870 4718
rect 24894 4690 24922 4718
rect 24946 4690 24974 4718
rect 24998 4690 25026 4718
rect 29582 4690 29610 4718
rect 29634 4690 29662 4718
rect 29686 4690 29714 4718
rect 29738 4690 29766 4718
rect 29790 4690 29818 4718
rect 29842 4690 29870 4718
rect 29894 4690 29922 4718
rect 29946 4690 29974 4718
rect 29998 4690 30026 4718
rect 34582 4690 34610 4718
rect 34634 4690 34662 4718
rect 34686 4690 34714 4718
rect 34738 4690 34766 4718
rect 34790 4690 34818 4718
rect 34842 4690 34870 4718
rect 34894 4690 34922 4718
rect 34946 4690 34974 4718
rect 34998 4690 35026 4718
rect 31990 4438 32018 4466
rect 2082 4298 2110 4326
rect 2134 4298 2162 4326
rect 2186 4298 2214 4326
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 2394 4298 2422 4326
rect 2446 4298 2474 4326
rect 2498 4298 2526 4326
rect 7082 4298 7110 4326
rect 7134 4298 7162 4326
rect 7186 4298 7214 4326
rect 7238 4298 7266 4326
rect 7290 4298 7318 4326
rect 7342 4298 7370 4326
rect 7394 4298 7422 4326
rect 7446 4298 7474 4326
rect 7498 4298 7526 4326
rect 12082 4298 12110 4326
rect 12134 4298 12162 4326
rect 12186 4298 12214 4326
rect 12238 4298 12266 4326
rect 12290 4298 12318 4326
rect 12342 4298 12370 4326
rect 12394 4298 12422 4326
rect 12446 4298 12474 4326
rect 12498 4298 12526 4326
rect 17082 4298 17110 4326
rect 17134 4298 17162 4326
rect 17186 4298 17214 4326
rect 17238 4298 17266 4326
rect 17290 4298 17318 4326
rect 17342 4298 17370 4326
rect 17394 4298 17422 4326
rect 17446 4298 17474 4326
rect 17498 4298 17526 4326
rect 22082 4298 22110 4326
rect 22134 4298 22162 4326
rect 22186 4298 22214 4326
rect 22238 4298 22266 4326
rect 22290 4298 22318 4326
rect 22342 4298 22370 4326
rect 22394 4298 22422 4326
rect 22446 4298 22474 4326
rect 22498 4298 22526 4326
rect 27082 4298 27110 4326
rect 27134 4298 27162 4326
rect 27186 4298 27214 4326
rect 27238 4298 27266 4326
rect 27290 4298 27318 4326
rect 27342 4298 27370 4326
rect 27394 4298 27422 4326
rect 27446 4298 27474 4326
rect 27498 4298 27526 4326
rect 32082 4298 32110 4326
rect 32134 4298 32162 4326
rect 32186 4298 32214 4326
rect 32238 4298 32266 4326
rect 32290 4298 32318 4326
rect 32342 4298 32370 4326
rect 32394 4298 32422 4326
rect 32446 4298 32474 4326
rect 32498 4298 32526 4326
rect 37082 4298 37110 4326
rect 37134 4298 37162 4326
rect 37186 4298 37214 4326
rect 37238 4298 37266 4326
rect 37290 4298 37318 4326
rect 37342 4298 37370 4326
rect 37394 4298 37422 4326
rect 37446 4298 37474 4326
rect 37498 4298 37526 4326
rect 36918 4158 36946 4186
rect 4582 3906 4610 3934
rect 4634 3906 4662 3934
rect 4686 3906 4714 3934
rect 4738 3906 4766 3934
rect 4790 3906 4818 3934
rect 4842 3906 4870 3934
rect 4894 3906 4922 3934
rect 4946 3906 4974 3934
rect 4998 3906 5026 3934
rect 9582 3906 9610 3934
rect 9634 3906 9662 3934
rect 9686 3906 9714 3934
rect 9738 3906 9766 3934
rect 9790 3906 9818 3934
rect 9842 3906 9870 3934
rect 9894 3906 9922 3934
rect 9946 3906 9974 3934
rect 9998 3906 10026 3934
rect 14582 3906 14610 3934
rect 14634 3906 14662 3934
rect 14686 3906 14714 3934
rect 14738 3906 14766 3934
rect 14790 3906 14818 3934
rect 14842 3906 14870 3934
rect 14894 3906 14922 3934
rect 14946 3906 14974 3934
rect 14998 3906 15026 3934
rect 19582 3906 19610 3934
rect 19634 3906 19662 3934
rect 19686 3906 19714 3934
rect 19738 3906 19766 3934
rect 19790 3906 19818 3934
rect 19842 3906 19870 3934
rect 19894 3906 19922 3934
rect 19946 3906 19974 3934
rect 19998 3906 20026 3934
rect 24582 3906 24610 3934
rect 24634 3906 24662 3934
rect 24686 3906 24714 3934
rect 24738 3906 24766 3934
rect 24790 3906 24818 3934
rect 24842 3906 24870 3934
rect 24894 3906 24922 3934
rect 24946 3906 24974 3934
rect 24998 3906 25026 3934
rect 29582 3906 29610 3934
rect 29634 3906 29662 3934
rect 29686 3906 29714 3934
rect 29738 3906 29766 3934
rect 29790 3906 29818 3934
rect 29842 3906 29870 3934
rect 29894 3906 29922 3934
rect 29946 3906 29974 3934
rect 29998 3906 30026 3934
rect 34582 3906 34610 3934
rect 34634 3906 34662 3934
rect 34686 3906 34714 3934
rect 34738 3906 34766 3934
rect 34790 3906 34818 3934
rect 34842 3906 34870 3934
rect 34894 3906 34922 3934
rect 34946 3906 34974 3934
rect 34998 3906 35026 3934
rect 31990 3710 32018 3738
rect 2082 3514 2110 3542
rect 2134 3514 2162 3542
rect 2186 3514 2214 3542
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 2394 3514 2422 3542
rect 2446 3514 2474 3542
rect 2498 3514 2526 3542
rect 7082 3514 7110 3542
rect 7134 3514 7162 3542
rect 7186 3514 7214 3542
rect 7238 3514 7266 3542
rect 7290 3514 7318 3542
rect 7342 3514 7370 3542
rect 7394 3514 7422 3542
rect 7446 3514 7474 3542
rect 7498 3514 7526 3542
rect 12082 3514 12110 3542
rect 12134 3514 12162 3542
rect 12186 3514 12214 3542
rect 12238 3514 12266 3542
rect 12290 3514 12318 3542
rect 12342 3514 12370 3542
rect 12394 3514 12422 3542
rect 12446 3514 12474 3542
rect 12498 3514 12526 3542
rect 17082 3514 17110 3542
rect 17134 3514 17162 3542
rect 17186 3514 17214 3542
rect 17238 3514 17266 3542
rect 17290 3514 17318 3542
rect 17342 3514 17370 3542
rect 17394 3514 17422 3542
rect 17446 3514 17474 3542
rect 17498 3514 17526 3542
rect 22082 3514 22110 3542
rect 22134 3514 22162 3542
rect 22186 3514 22214 3542
rect 22238 3514 22266 3542
rect 22290 3514 22318 3542
rect 22342 3514 22370 3542
rect 22394 3514 22422 3542
rect 22446 3514 22474 3542
rect 22498 3514 22526 3542
rect 27082 3514 27110 3542
rect 27134 3514 27162 3542
rect 27186 3514 27214 3542
rect 27238 3514 27266 3542
rect 27290 3514 27318 3542
rect 27342 3514 27370 3542
rect 27394 3514 27422 3542
rect 27446 3514 27474 3542
rect 27498 3514 27526 3542
rect 32082 3514 32110 3542
rect 32134 3514 32162 3542
rect 32186 3514 32214 3542
rect 32238 3514 32266 3542
rect 32290 3514 32318 3542
rect 32342 3514 32370 3542
rect 32394 3514 32422 3542
rect 32446 3514 32474 3542
rect 32498 3514 32526 3542
rect 37082 3514 37110 3542
rect 37134 3514 37162 3542
rect 37186 3514 37214 3542
rect 37238 3514 37266 3542
rect 37290 3514 37318 3542
rect 37342 3514 37370 3542
rect 37394 3514 37422 3542
rect 37446 3514 37474 3542
rect 37498 3514 37526 3542
rect 36918 3374 36946 3402
rect 4582 3122 4610 3150
rect 4634 3122 4662 3150
rect 4686 3122 4714 3150
rect 4738 3122 4766 3150
rect 4790 3122 4818 3150
rect 4842 3122 4870 3150
rect 4894 3122 4922 3150
rect 4946 3122 4974 3150
rect 4998 3122 5026 3150
rect 9582 3122 9610 3150
rect 9634 3122 9662 3150
rect 9686 3122 9714 3150
rect 9738 3122 9766 3150
rect 9790 3122 9818 3150
rect 9842 3122 9870 3150
rect 9894 3122 9922 3150
rect 9946 3122 9974 3150
rect 9998 3122 10026 3150
rect 14582 3122 14610 3150
rect 14634 3122 14662 3150
rect 14686 3122 14714 3150
rect 14738 3122 14766 3150
rect 14790 3122 14818 3150
rect 14842 3122 14870 3150
rect 14894 3122 14922 3150
rect 14946 3122 14974 3150
rect 14998 3122 15026 3150
rect 19582 3122 19610 3150
rect 19634 3122 19662 3150
rect 19686 3122 19714 3150
rect 19738 3122 19766 3150
rect 19790 3122 19818 3150
rect 19842 3122 19870 3150
rect 19894 3122 19922 3150
rect 19946 3122 19974 3150
rect 19998 3122 20026 3150
rect 24582 3122 24610 3150
rect 24634 3122 24662 3150
rect 24686 3122 24714 3150
rect 24738 3122 24766 3150
rect 24790 3122 24818 3150
rect 24842 3122 24870 3150
rect 24894 3122 24922 3150
rect 24946 3122 24974 3150
rect 24998 3122 25026 3150
rect 29582 3122 29610 3150
rect 29634 3122 29662 3150
rect 29686 3122 29714 3150
rect 29738 3122 29766 3150
rect 29790 3122 29818 3150
rect 29842 3122 29870 3150
rect 29894 3122 29922 3150
rect 29946 3122 29974 3150
rect 29998 3122 30026 3150
rect 34582 3122 34610 3150
rect 34634 3122 34662 3150
rect 34686 3122 34714 3150
rect 34738 3122 34766 3150
rect 34790 3122 34818 3150
rect 34842 3122 34870 3150
rect 34894 3122 34922 3150
rect 34946 3122 34974 3150
rect 34998 3122 35026 3150
rect 31990 2982 32018 3010
rect 2082 2730 2110 2758
rect 2134 2730 2162 2758
rect 2186 2730 2214 2758
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 2394 2730 2422 2758
rect 2446 2730 2474 2758
rect 2498 2730 2526 2758
rect 7082 2730 7110 2758
rect 7134 2730 7162 2758
rect 7186 2730 7214 2758
rect 7238 2730 7266 2758
rect 7290 2730 7318 2758
rect 7342 2730 7370 2758
rect 7394 2730 7422 2758
rect 7446 2730 7474 2758
rect 7498 2730 7526 2758
rect 12082 2730 12110 2758
rect 12134 2730 12162 2758
rect 12186 2730 12214 2758
rect 12238 2730 12266 2758
rect 12290 2730 12318 2758
rect 12342 2730 12370 2758
rect 12394 2730 12422 2758
rect 12446 2730 12474 2758
rect 12498 2730 12526 2758
rect 17082 2730 17110 2758
rect 17134 2730 17162 2758
rect 17186 2730 17214 2758
rect 17238 2730 17266 2758
rect 17290 2730 17318 2758
rect 17342 2730 17370 2758
rect 17394 2730 17422 2758
rect 17446 2730 17474 2758
rect 17498 2730 17526 2758
rect 22082 2730 22110 2758
rect 22134 2730 22162 2758
rect 22186 2730 22214 2758
rect 22238 2730 22266 2758
rect 22290 2730 22318 2758
rect 22342 2730 22370 2758
rect 22394 2730 22422 2758
rect 22446 2730 22474 2758
rect 22498 2730 22526 2758
rect 27082 2730 27110 2758
rect 27134 2730 27162 2758
rect 27186 2730 27214 2758
rect 27238 2730 27266 2758
rect 27290 2730 27318 2758
rect 27342 2730 27370 2758
rect 27394 2730 27422 2758
rect 27446 2730 27474 2758
rect 27498 2730 27526 2758
rect 32082 2730 32110 2758
rect 32134 2730 32162 2758
rect 32186 2730 32214 2758
rect 32238 2730 32266 2758
rect 32290 2730 32318 2758
rect 32342 2730 32370 2758
rect 32394 2730 32422 2758
rect 32446 2730 32474 2758
rect 32498 2730 32526 2758
rect 37082 2730 37110 2758
rect 37134 2730 37162 2758
rect 37186 2730 37214 2758
rect 37238 2730 37266 2758
rect 37290 2730 37318 2758
rect 37342 2730 37370 2758
rect 37394 2730 37422 2758
rect 37446 2730 37474 2758
rect 37498 2730 37526 2758
rect 4582 2338 4610 2366
rect 4634 2338 4662 2366
rect 4686 2338 4714 2366
rect 4738 2338 4766 2366
rect 4790 2338 4818 2366
rect 4842 2338 4870 2366
rect 4894 2338 4922 2366
rect 4946 2338 4974 2366
rect 4998 2338 5026 2366
rect 9582 2338 9610 2366
rect 9634 2338 9662 2366
rect 9686 2338 9714 2366
rect 9738 2338 9766 2366
rect 9790 2338 9818 2366
rect 9842 2338 9870 2366
rect 9894 2338 9922 2366
rect 9946 2338 9974 2366
rect 9998 2338 10026 2366
rect 14582 2338 14610 2366
rect 14634 2338 14662 2366
rect 14686 2338 14714 2366
rect 14738 2338 14766 2366
rect 14790 2338 14818 2366
rect 14842 2338 14870 2366
rect 14894 2338 14922 2366
rect 14946 2338 14974 2366
rect 14998 2338 15026 2366
rect 19582 2338 19610 2366
rect 19634 2338 19662 2366
rect 19686 2338 19714 2366
rect 19738 2338 19766 2366
rect 19790 2338 19818 2366
rect 19842 2338 19870 2366
rect 19894 2338 19922 2366
rect 19946 2338 19974 2366
rect 19998 2338 20026 2366
rect 24582 2338 24610 2366
rect 24634 2338 24662 2366
rect 24686 2338 24714 2366
rect 24738 2338 24766 2366
rect 24790 2338 24818 2366
rect 24842 2338 24870 2366
rect 24894 2338 24922 2366
rect 24946 2338 24974 2366
rect 24998 2338 25026 2366
rect 29582 2338 29610 2366
rect 29634 2338 29662 2366
rect 29686 2338 29714 2366
rect 29738 2338 29766 2366
rect 29790 2338 29818 2366
rect 29842 2338 29870 2366
rect 29894 2338 29922 2366
rect 29946 2338 29974 2366
rect 29998 2338 30026 2366
rect 34582 2338 34610 2366
rect 34634 2338 34662 2366
rect 34686 2338 34714 2366
rect 34738 2338 34766 2366
rect 34790 2338 34818 2366
rect 34842 2338 34870 2366
rect 34894 2338 34922 2366
rect 34946 2338 34974 2366
rect 34998 2338 35026 2366
rect 31990 2198 32018 2226
rect 2082 1946 2110 1974
rect 2134 1946 2162 1974
rect 2186 1946 2214 1974
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 2394 1946 2422 1974
rect 2446 1946 2474 1974
rect 2498 1946 2526 1974
rect 7082 1946 7110 1974
rect 7134 1946 7162 1974
rect 7186 1946 7214 1974
rect 7238 1946 7266 1974
rect 7290 1946 7318 1974
rect 7342 1946 7370 1974
rect 7394 1946 7422 1974
rect 7446 1946 7474 1974
rect 7498 1946 7526 1974
rect 12082 1946 12110 1974
rect 12134 1946 12162 1974
rect 12186 1946 12214 1974
rect 12238 1946 12266 1974
rect 12290 1946 12318 1974
rect 12342 1946 12370 1974
rect 12394 1946 12422 1974
rect 12446 1946 12474 1974
rect 12498 1946 12526 1974
rect 17082 1946 17110 1974
rect 17134 1946 17162 1974
rect 17186 1946 17214 1974
rect 17238 1946 17266 1974
rect 17290 1946 17318 1974
rect 17342 1946 17370 1974
rect 17394 1946 17422 1974
rect 17446 1946 17474 1974
rect 17498 1946 17526 1974
rect 22082 1946 22110 1974
rect 22134 1946 22162 1974
rect 22186 1946 22214 1974
rect 22238 1946 22266 1974
rect 22290 1946 22318 1974
rect 22342 1946 22370 1974
rect 22394 1946 22422 1974
rect 22446 1946 22474 1974
rect 22498 1946 22526 1974
rect 27082 1946 27110 1974
rect 27134 1946 27162 1974
rect 27186 1946 27214 1974
rect 27238 1946 27266 1974
rect 27290 1946 27318 1974
rect 27342 1946 27370 1974
rect 27394 1946 27422 1974
rect 27446 1946 27474 1974
rect 27498 1946 27526 1974
rect 32082 1946 32110 1974
rect 32134 1946 32162 1974
rect 32186 1946 32214 1974
rect 32238 1946 32266 1974
rect 32290 1946 32318 1974
rect 32342 1946 32370 1974
rect 32394 1946 32422 1974
rect 32446 1946 32474 1974
rect 32498 1946 32526 1974
rect 37082 1946 37110 1974
rect 37134 1946 37162 1974
rect 37186 1946 37214 1974
rect 37238 1946 37266 1974
rect 37290 1946 37318 1974
rect 37342 1946 37370 1974
rect 37394 1946 37422 1974
rect 37446 1946 37474 1974
rect 37498 1946 37526 1974
rect 4582 1554 4610 1582
rect 4634 1554 4662 1582
rect 4686 1554 4714 1582
rect 4738 1554 4766 1582
rect 4790 1554 4818 1582
rect 4842 1554 4870 1582
rect 4894 1554 4922 1582
rect 4946 1554 4974 1582
rect 4998 1554 5026 1582
rect 9582 1554 9610 1582
rect 9634 1554 9662 1582
rect 9686 1554 9714 1582
rect 9738 1554 9766 1582
rect 9790 1554 9818 1582
rect 9842 1554 9870 1582
rect 9894 1554 9922 1582
rect 9946 1554 9974 1582
rect 9998 1554 10026 1582
rect 14582 1554 14610 1582
rect 14634 1554 14662 1582
rect 14686 1554 14714 1582
rect 14738 1554 14766 1582
rect 14790 1554 14818 1582
rect 14842 1554 14870 1582
rect 14894 1554 14922 1582
rect 14946 1554 14974 1582
rect 14998 1554 15026 1582
rect 19582 1554 19610 1582
rect 19634 1554 19662 1582
rect 19686 1554 19714 1582
rect 19738 1554 19766 1582
rect 19790 1554 19818 1582
rect 19842 1554 19870 1582
rect 19894 1554 19922 1582
rect 19946 1554 19974 1582
rect 19998 1554 20026 1582
rect 24582 1554 24610 1582
rect 24634 1554 24662 1582
rect 24686 1554 24714 1582
rect 24738 1554 24766 1582
rect 24790 1554 24818 1582
rect 24842 1554 24870 1582
rect 24894 1554 24922 1582
rect 24946 1554 24974 1582
rect 24998 1554 25026 1582
rect 29582 1554 29610 1582
rect 29634 1554 29662 1582
rect 29686 1554 29714 1582
rect 29738 1554 29766 1582
rect 29790 1554 29818 1582
rect 29842 1554 29870 1582
rect 29894 1554 29922 1582
rect 29946 1554 29974 1582
rect 29998 1554 30026 1582
rect 34582 1554 34610 1582
rect 34634 1554 34662 1582
rect 34686 1554 34714 1582
rect 34738 1554 34766 1582
rect 34790 1554 34818 1582
rect 34842 1554 34870 1582
rect 34894 1554 34922 1582
rect 34946 1554 34974 1582
rect 34998 1554 35026 1582
<< metal4 >>
rect 2054 18438 2554 18454
rect 2054 18410 2082 18438
rect 2110 18410 2134 18438
rect 2162 18410 2186 18438
rect 2214 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2394 18438
rect 2422 18410 2446 18438
rect 2474 18410 2498 18438
rect 2526 18410 2554 18438
rect 2054 17654 2554 18410
rect 2054 17626 2082 17654
rect 2110 17626 2134 17654
rect 2162 17626 2186 17654
rect 2214 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2394 17654
rect 2422 17626 2446 17654
rect 2474 17626 2498 17654
rect 2526 17626 2554 17654
rect 2054 16870 2554 17626
rect 2054 16842 2082 16870
rect 2110 16842 2134 16870
rect 2162 16842 2186 16870
rect 2214 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2394 16870
rect 2422 16842 2446 16870
rect 2474 16842 2498 16870
rect 2526 16842 2554 16870
rect 2054 16086 2554 16842
rect 2054 16058 2082 16086
rect 2110 16058 2134 16086
rect 2162 16058 2186 16086
rect 2214 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2394 16086
rect 2422 16058 2446 16086
rect 2474 16058 2498 16086
rect 2526 16058 2554 16086
rect 2054 15302 2554 16058
rect 2054 15274 2082 15302
rect 2110 15274 2134 15302
rect 2162 15274 2186 15302
rect 2214 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2394 15302
rect 2422 15274 2446 15302
rect 2474 15274 2498 15302
rect 2526 15274 2554 15302
rect 2054 14518 2554 15274
rect 2054 14490 2082 14518
rect 2110 14490 2134 14518
rect 2162 14490 2186 14518
rect 2214 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2394 14518
rect 2422 14490 2446 14518
rect 2474 14490 2498 14518
rect 2526 14490 2554 14518
rect 2054 13734 2554 14490
rect 2054 13706 2082 13734
rect 2110 13706 2134 13734
rect 2162 13706 2186 13734
rect 2214 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2394 13734
rect 2422 13706 2446 13734
rect 2474 13706 2498 13734
rect 2526 13706 2554 13734
rect 2054 12950 2554 13706
rect 2054 12922 2082 12950
rect 2110 12922 2134 12950
rect 2162 12922 2186 12950
rect 2214 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2394 12950
rect 2422 12922 2446 12950
rect 2474 12922 2498 12950
rect 2526 12922 2554 12950
rect 2054 12166 2554 12922
rect 2054 12138 2082 12166
rect 2110 12138 2134 12166
rect 2162 12138 2186 12166
rect 2214 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2394 12166
rect 2422 12138 2446 12166
rect 2474 12138 2498 12166
rect 2526 12138 2554 12166
rect 2054 11382 2554 12138
rect 2054 11354 2082 11382
rect 2110 11354 2134 11382
rect 2162 11354 2186 11382
rect 2214 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2394 11382
rect 2422 11354 2446 11382
rect 2474 11354 2498 11382
rect 2526 11354 2554 11382
rect 2054 10598 2554 11354
rect 2054 10570 2082 10598
rect 2110 10570 2134 10598
rect 2162 10570 2186 10598
rect 2214 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2394 10598
rect 2422 10570 2446 10598
rect 2474 10570 2498 10598
rect 2526 10570 2554 10598
rect 2054 9814 2554 10570
rect 2054 9786 2082 9814
rect 2110 9786 2134 9814
rect 2162 9786 2186 9814
rect 2214 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2394 9814
rect 2422 9786 2446 9814
rect 2474 9786 2498 9814
rect 2526 9786 2554 9814
rect 2054 9030 2554 9786
rect 2054 9002 2082 9030
rect 2110 9002 2134 9030
rect 2162 9002 2186 9030
rect 2214 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2394 9030
rect 2422 9002 2446 9030
rect 2474 9002 2498 9030
rect 2526 9002 2554 9030
rect 2054 8246 2554 9002
rect 2054 8218 2082 8246
rect 2110 8218 2134 8246
rect 2162 8218 2186 8246
rect 2214 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2394 8246
rect 2422 8218 2446 8246
rect 2474 8218 2498 8246
rect 2526 8218 2554 8246
rect 2054 7462 2554 8218
rect 2054 7434 2082 7462
rect 2110 7434 2134 7462
rect 2162 7434 2186 7462
rect 2214 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2394 7462
rect 2422 7434 2446 7462
rect 2474 7434 2498 7462
rect 2526 7434 2554 7462
rect 2054 6678 2554 7434
rect 2054 6650 2082 6678
rect 2110 6650 2134 6678
rect 2162 6650 2186 6678
rect 2214 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2394 6678
rect 2422 6650 2446 6678
rect 2474 6650 2498 6678
rect 2526 6650 2554 6678
rect 2054 5894 2554 6650
rect 2054 5866 2082 5894
rect 2110 5866 2134 5894
rect 2162 5866 2186 5894
rect 2214 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2394 5894
rect 2422 5866 2446 5894
rect 2474 5866 2498 5894
rect 2526 5866 2554 5894
rect 2054 5110 2554 5866
rect 2054 5082 2082 5110
rect 2110 5082 2134 5110
rect 2162 5082 2186 5110
rect 2214 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2394 5110
rect 2422 5082 2446 5110
rect 2474 5082 2498 5110
rect 2526 5082 2554 5110
rect 2054 4326 2554 5082
rect 2054 4298 2082 4326
rect 2110 4298 2134 4326
rect 2162 4298 2186 4326
rect 2214 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2394 4326
rect 2422 4298 2446 4326
rect 2474 4298 2498 4326
rect 2526 4298 2554 4326
rect 2054 3542 2554 4298
rect 2054 3514 2082 3542
rect 2110 3514 2134 3542
rect 2162 3514 2186 3542
rect 2214 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2394 3542
rect 2422 3514 2446 3542
rect 2474 3514 2498 3542
rect 2526 3514 2554 3542
rect 2054 2758 2554 3514
rect 2054 2730 2082 2758
rect 2110 2730 2134 2758
rect 2162 2730 2186 2758
rect 2214 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2394 2758
rect 2422 2730 2446 2758
rect 2474 2730 2498 2758
rect 2526 2730 2554 2758
rect 2054 1974 2554 2730
rect 2054 1946 2082 1974
rect 2110 1946 2134 1974
rect 2162 1946 2186 1974
rect 2214 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2394 1974
rect 2422 1946 2446 1974
rect 2474 1946 2498 1974
rect 2526 1946 2554 1974
rect 2054 1538 2554 1946
rect 4554 18046 5054 18454
rect 4554 18018 4582 18046
rect 4610 18018 4634 18046
rect 4662 18018 4686 18046
rect 4714 18018 4738 18046
rect 4766 18018 4790 18046
rect 4818 18018 4842 18046
rect 4870 18018 4894 18046
rect 4922 18018 4946 18046
rect 4974 18018 4998 18046
rect 5026 18018 5054 18046
rect 4554 17262 5054 18018
rect 4554 17234 4582 17262
rect 4610 17234 4634 17262
rect 4662 17234 4686 17262
rect 4714 17234 4738 17262
rect 4766 17234 4790 17262
rect 4818 17234 4842 17262
rect 4870 17234 4894 17262
rect 4922 17234 4946 17262
rect 4974 17234 4998 17262
rect 5026 17234 5054 17262
rect 4554 16478 5054 17234
rect 4554 16450 4582 16478
rect 4610 16450 4634 16478
rect 4662 16450 4686 16478
rect 4714 16450 4738 16478
rect 4766 16450 4790 16478
rect 4818 16450 4842 16478
rect 4870 16450 4894 16478
rect 4922 16450 4946 16478
rect 4974 16450 4998 16478
rect 5026 16450 5054 16478
rect 4554 15694 5054 16450
rect 4554 15666 4582 15694
rect 4610 15666 4634 15694
rect 4662 15666 4686 15694
rect 4714 15666 4738 15694
rect 4766 15666 4790 15694
rect 4818 15666 4842 15694
rect 4870 15666 4894 15694
rect 4922 15666 4946 15694
rect 4974 15666 4998 15694
rect 5026 15666 5054 15694
rect 4554 14910 5054 15666
rect 4554 14882 4582 14910
rect 4610 14882 4634 14910
rect 4662 14882 4686 14910
rect 4714 14882 4738 14910
rect 4766 14882 4790 14910
rect 4818 14882 4842 14910
rect 4870 14882 4894 14910
rect 4922 14882 4946 14910
rect 4974 14882 4998 14910
rect 5026 14882 5054 14910
rect 4554 14126 5054 14882
rect 4554 14098 4582 14126
rect 4610 14098 4634 14126
rect 4662 14098 4686 14126
rect 4714 14098 4738 14126
rect 4766 14098 4790 14126
rect 4818 14098 4842 14126
rect 4870 14098 4894 14126
rect 4922 14098 4946 14126
rect 4974 14098 4998 14126
rect 5026 14098 5054 14126
rect 4554 13342 5054 14098
rect 4554 13314 4582 13342
rect 4610 13314 4634 13342
rect 4662 13314 4686 13342
rect 4714 13314 4738 13342
rect 4766 13314 4790 13342
rect 4818 13314 4842 13342
rect 4870 13314 4894 13342
rect 4922 13314 4946 13342
rect 4974 13314 4998 13342
rect 5026 13314 5054 13342
rect 4554 12558 5054 13314
rect 4554 12530 4582 12558
rect 4610 12530 4634 12558
rect 4662 12530 4686 12558
rect 4714 12530 4738 12558
rect 4766 12530 4790 12558
rect 4818 12530 4842 12558
rect 4870 12530 4894 12558
rect 4922 12530 4946 12558
rect 4974 12530 4998 12558
rect 5026 12530 5054 12558
rect 4554 11774 5054 12530
rect 4554 11746 4582 11774
rect 4610 11746 4634 11774
rect 4662 11746 4686 11774
rect 4714 11746 4738 11774
rect 4766 11746 4790 11774
rect 4818 11746 4842 11774
rect 4870 11746 4894 11774
rect 4922 11746 4946 11774
rect 4974 11746 4998 11774
rect 5026 11746 5054 11774
rect 4554 10990 5054 11746
rect 4554 10962 4582 10990
rect 4610 10962 4634 10990
rect 4662 10962 4686 10990
rect 4714 10962 4738 10990
rect 4766 10962 4790 10990
rect 4818 10962 4842 10990
rect 4870 10962 4894 10990
rect 4922 10962 4946 10990
rect 4974 10962 4998 10990
rect 5026 10962 5054 10990
rect 4554 10206 5054 10962
rect 4554 10178 4582 10206
rect 4610 10178 4634 10206
rect 4662 10178 4686 10206
rect 4714 10178 4738 10206
rect 4766 10178 4790 10206
rect 4818 10178 4842 10206
rect 4870 10178 4894 10206
rect 4922 10178 4946 10206
rect 4974 10178 4998 10206
rect 5026 10178 5054 10206
rect 4554 9422 5054 10178
rect 4554 9394 4582 9422
rect 4610 9394 4634 9422
rect 4662 9394 4686 9422
rect 4714 9394 4738 9422
rect 4766 9394 4790 9422
rect 4818 9394 4842 9422
rect 4870 9394 4894 9422
rect 4922 9394 4946 9422
rect 4974 9394 4998 9422
rect 5026 9394 5054 9422
rect 4554 8638 5054 9394
rect 4554 8610 4582 8638
rect 4610 8610 4634 8638
rect 4662 8610 4686 8638
rect 4714 8610 4738 8638
rect 4766 8610 4790 8638
rect 4818 8610 4842 8638
rect 4870 8610 4894 8638
rect 4922 8610 4946 8638
rect 4974 8610 4998 8638
rect 5026 8610 5054 8638
rect 4554 7854 5054 8610
rect 4554 7826 4582 7854
rect 4610 7826 4634 7854
rect 4662 7826 4686 7854
rect 4714 7826 4738 7854
rect 4766 7826 4790 7854
rect 4818 7826 4842 7854
rect 4870 7826 4894 7854
rect 4922 7826 4946 7854
rect 4974 7826 4998 7854
rect 5026 7826 5054 7854
rect 4554 7070 5054 7826
rect 4554 7042 4582 7070
rect 4610 7042 4634 7070
rect 4662 7042 4686 7070
rect 4714 7042 4738 7070
rect 4766 7042 4790 7070
rect 4818 7042 4842 7070
rect 4870 7042 4894 7070
rect 4922 7042 4946 7070
rect 4974 7042 4998 7070
rect 5026 7042 5054 7070
rect 4554 6286 5054 7042
rect 4554 6258 4582 6286
rect 4610 6258 4634 6286
rect 4662 6258 4686 6286
rect 4714 6258 4738 6286
rect 4766 6258 4790 6286
rect 4818 6258 4842 6286
rect 4870 6258 4894 6286
rect 4922 6258 4946 6286
rect 4974 6258 4998 6286
rect 5026 6258 5054 6286
rect 4554 5502 5054 6258
rect 4554 5474 4582 5502
rect 4610 5474 4634 5502
rect 4662 5474 4686 5502
rect 4714 5474 4738 5502
rect 4766 5474 4790 5502
rect 4818 5474 4842 5502
rect 4870 5474 4894 5502
rect 4922 5474 4946 5502
rect 4974 5474 4998 5502
rect 5026 5474 5054 5502
rect 4554 4718 5054 5474
rect 4554 4690 4582 4718
rect 4610 4690 4634 4718
rect 4662 4690 4686 4718
rect 4714 4690 4738 4718
rect 4766 4690 4790 4718
rect 4818 4690 4842 4718
rect 4870 4690 4894 4718
rect 4922 4690 4946 4718
rect 4974 4690 4998 4718
rect 5026 4690 5054 4718
rect 4554 3934 5054 4690
rect 4554 3906 4582 3934
rect 4610 3906 4634 3934
rect 4662 3906 4686 3934
rect 4714 3906 4738 3934
rect 4766 3906 4790 3934
rect 4818 3906 4842 3934
rect 4870 3906 4894 3934
rect 4922 3906 4946 3934
rect 4974 3906 4998 3934
rect 5026 3906 5054 3934
rect 4554 3150 5054 3906
rect 4554 3122 4582 3150
rect 4610 3122 4634 3150
rect 4662 3122 4686 3150
rect 4714 3122 4738 3150
rect 4766 3122 4790 3150
rect 4818 3122 4842 3150
rect 4870 3122 4894 3150
rect 4922 3122 4946 3150
rect 4974 3122 4998 3150
rect 5026 3122 5054 3150
rect 4554 2366 5054 3122
rect 4554 2338 4582 2366
rect 4610 2338 4634 2366
rect 4662 2338 4686 2366
rect 4714 2338 4738 2366
rect 4766 2338 4790 2366
rect 4818 2338 4842 2366
rect 4870 2338 4894 2366
rect 4922 2338 4946 2366
rect 4974 2338 4998 2366
rect 5026 2338 5054 2366
rect 4554 1582 5054 2338
rect 4554 1554 4582 1582
rect 4610 1554 4634 1582
rect 4662 1554 4686 1582
rect 4714 1554 4738 1582
rect 4766 1554 4790 1582
rect 4818 1554 4842 1582
rect 4870 1554 4894 1582
rect 4922 1554 4946 1582
rect 4974 1554 4998 1582
rect 5026 1554 5054 1582
rect 4554 1538 5054 1554
rect 7054 18438 7554 18454
rect 7054 18410 7082 18438
rect 7110 18410 7134 18438
rect 7162 18410 7186 18438
rect 7214 18410 7238 18438
rect 7266 18410 7290 18438
rect 7318 18410 7342 18438
rect 7370 18410 7394 18438
rect 7422 18410 7446 18438
rect 7474 18410 7498 18438
rect 7526 18410 7554 18438
rect 7054 17654 7554 18410
rect 7054 17626 7082 17654
rect 7110 17626 7134 17654
rect 7162 17626 7186 17654
rect 7214 17626 7238 17654
rect 7266 17626 7290 17654
rect 7318 17626 7342 17654
rect 7370 17626 7394 17654
rect 7422 17626 7446 17654
rect 7474 17626 7498 17654
rect 7526 17626 7554 17654
rect 7054 16870 7554 17626
rect 7054 16842 7082 16870
rect 7110 16842 7134 16870
rect 7162 16842 7186 16870
rect 7214 16842 7238 16870
rect 7266 16842 7290 16870
rect 7318 16842 7342 16870
rect 7370 16842 7394 16870
rect 7422 16842 7446 16870
rect 7474 16842 7498 16870
rect 7526 16842 7554 16870
rect 7054 16086 7554 16842
rect 7054 16058 7082 16086
rect 7110 16058 7134 16086
rect 7162 16058 7186 16086
rect 7214 16058 7238 16086
rect 7266 16058 7290 16086
rect 7318 16058 7342 16086
rect 7370 16058 7394 16086
rect 7422 16058 7446 16086
rect 7474 16058 7498 16086
rect 7526 16058 7554 16086
rect 7054 15302 7554 16058
rect 7054 15274 7082 15302
rect 7110 15274 7134 15302
rect 7162 15274 7186 15302
rect 7214 15274 7238 15302
rect 7266 15274 7290 15302
rect 7318 15274 7342 15302
rect 7370 15274 7394 15302
rect 7422 15274 7446 15302
rect 7474 15274 7498 15302
rect 7526 15274 7554 15302
rect 7054 14518 7554 15274
rect 7054 14490 7082 14518
rect 7110 14490 7134 14518
rect 7162 14490 7186 14518
rect 7214 14490 7238 14518
rect 7266 14490 7290 14518
rect 7318 14490 7342 14518
rect 7370 14490 7394 14518
rect 7422 14490 7446 14518
rect 7474 14490 7498 14518
rect 7526 14490 7554 14518
rect 7054 13734 7554 14490
rect 7054 13706 7082 13734
rect 7110 13706 7134 13734
rect 7162 13706 7186 13734
rect 7214 13706 7238 13734
rect 7266 13706 7290 13734
rect 7318 13706 7342 13734
rect 7370 13706 7394 13734
rect 7422 13706 7446 13734
rect 7474 13706 7498 13734
rect 7526 13706 7554 13734
rect 7054 12950 7554 13706
rect 7054 12922 7082 12950
rect 7110 12922 7134 12950
rect 7162 12922 7186 12950
rect 7214 12922 7238 12950
rect 7266 12922 7290 12950
rect 7318 12922 7342 12950
rect 7370 12922 7394 12950
rect 7422 12922 7446 12950
rect 7474 12922 7498 12950
rect 7526 12922 7554 12950
rect 7054 12166 7554 12922
rect 7054 12138 7082 12166
rect 7110 12138 7134 12166
rect 7162 12138 7186 12166
rect 7214 12138 7238 12166
rect 7266 12138 7290 12166
rect 7318 12138 7342 12166
rect 7370 12138 7394 12166
rect 7422 12138 7446 12166
rect 7474 12138 7498 12166
rect 7526 12138 7554 12166
rect 7054 11382 7554 12138
rect 7054 11354 7082 11382
rect 7110 11354 7134 11382
rect 7162 11354 7186 11382
rect 7214 11354 7238 11382
rect 7266 11354 7290 11382
rect 7318 11354 7342 11382
rect 7370 11354 7394 11382
rect 7422 11354 7446 11382
rect 7474 11354 7498 11382
rect 7526 11354 7554 11382
rect 7054 10598 7554 11354
rect 7054 10570 7082 10598
rect 7110 10570 7134 10598
rect 7162 10570 7186 10598
rect 7214 10570 7238 10598
rect 7266 10570 7290 10598
rect 7318 10570 7342 10598
rect 7370 10570 7394 10598
rect 7422 10570 7446 10598
rect 7474 10570 7498 10598
rect 7526 10570 7554 10598
rect 7054 9814 7554 10570
rect 7054 9786 7082 9814
rect 7110 9786 7134 9814
rect 7162 9786 7186 9814
rect 7214 9786 7238 9814
rect 7266 9786 7290 9814
rect 7318 9786 7342 9814
rect 7370 9786 7394 9814
rect 7422 9786 7446 9814
rect 7474 9786 7498 9814
rect 7526 9786 7554 9814
rect 7054 9030 7554 9786
rect 7054 9002 7082 9030
rect 7110 9002 7134 9030
rect 7162 9002 7186 9030
rect 7214 9002 7238 9030
rect 7266 9002 7290 9030
rect 7318 9002 7342 9030
rect 7370 9002 7394 9030
rect 7422 9002 7446 9030
rect 7474 9002 7498 9030
rect 7526 9002 7554 9030
rect 7054 8246 7554 9002
rect 7054 8218 7082 8246
rect 7110 8218 7134 8246
rect 7162 8218 7186 8246
rect 7214 8218 7238 8246
rect 7266 8218 7290 8246
rect 7318 8218 7342 8246
rect 7370 8218 7394 8246
rect 7422 8218 7446 8246
rect 7474 8218 7498 8246
rect 7526 8218 7554 8246
rect 7054 7462 7554 8218
rect 7054 7434 7082 7462
rect 7110 7434 7134 7462
rect 7162 7434 7186 7462
rect 7214 7434 7238 7462
rect 7266 7434 7290 7462
rect 7318 7434 7342 7462
rect 7370 7434 7394 7462
rect 7422 7434 7446 7462
rect 7474 7434 7498 7462
rect 7526 7434 7554 7462
rect 7054 6678 7554 7434
rect 7054 6650 7082 6678
rect 7110 6650 7134 6678
rect 7162 6650 7186 6678
rect 7214 6650 7238 6678
rect 7266 6650 7290 6678
rect 7318 6650 7342 6678
rect 7370 6650 7394 6678
rect 7422 6650 7446 6678
rect 7474 6650 7498 6678
rect 7526 6650 7554 6678
rect 7054 5894 7554 6650
rect 7054 5866 7082 5894
rect 7110 5866 7134 5894
rect 7162 5866 7186 5894
rect 7214 5866 7238 5894
rect 7266 5866 7290 5894
rect 7318 5866 7342 5894
rect 7370 5866 7394 5894
rect 7422 5866 7446 5894
rect 7474 5866 7498 5894
rect 7526 5866 7554 5894
rect 7054 5110 7554 5866
rect 7054 5082 7082 5110
rect 7110 5082 7134 5110
rect 7162 5082 7186 5110
rect 7214 5082 7238 5110
rect 7266 5082 7290 5110
rect 7318 5082 7342 5110
rect 7370 5082 7394 5110
rect 7422 5082 7446 5110
rect 7474 5082 7498 5110
rect 7526 5082 7554 5110
rect 7054 4326 7554 5082
rect 7054 4298 7082 4326
rect 7110 4298 7134 4326
rect 7162 4298 7186 4326
rect 7214 4298 7238 4326
rect 7266 4298 7290 4326
rect 7318 4298 7342 4326
rect 7370 4298 7394 4326
rect 7422 4298 7446 4326
rect 7474 4298 7498 4326
rect 7526 4298 7554 4326
rect 7054 3542 7554 4298
rect 7054 3514 7082 3542
rect 7110 3514 7134 3542
rect 7162 3514 7186 3542
rect 7214 3514 7238 3542
rect 7266 3514 7290 3542
rect 7318 3514 7342 3542
rect 7370 3514 7394 3542
rect 7422 3514 7446 3542
rect 7474 3514 7498 3542
rect 7526 3514 7554 3542
rect 7054 2758 7554 3514
rect 7054 2730 7082 2758
rect 7110 2730 7134 2758
rect 7162 2730 7186 2758
rect 7214 2730 7238 2758
rect 7266 2730 7290 2758
rect 7318 2730 7342 2758
rect 7370 2730 7394 2758
rect 7422 2730 7446 2758
rect 7474 2730 7498 2758
rect 7526 2730 7554 2758
rect 7054 1974 7554 2730
rect 7054 1946 7082 1974
rect 7110 1946 7134 1974
rect 7162 1946 7186 1974
rect 7214 1946 7238 1974
rect 7266 1946 7290 1974
rect 7318 1946 7342 1974
rect 7370 1946 7394 1974
rect 7422 1946 7446 1974
rect 7474 1946 7498 1974
rect 7526 1946 7554 1974
rect 7054 1538 7554 1946
rect 9554 18046 10054 18454
rect 9554 18018 9582 18046
rect 9610 18018 9634 18046
rect 9662 18018 9686 18046
rect 9714 18018 9738 18046
rect 9766 18018 9790 18046
rect 9818 18018 9842 18046
rect 9870 18018 9894 18046
rect 9922 18018 9946 18046
rect 9974 18018 9998 18046
rect 10026 18018 10054 18046
rect 9554 17262 10054 18018
rect 9554 17234 9582 17262
rect 9610 17234 9634 17262
rect 9662 17234 9686 17262
rect 9714 17234 9738 17262
rect 9766 17234 9790 17262
rect 9818 17234 9842 17262
rect 9870 17234 9894 17262
rect 9922 17234 9946 17262
rect 9974 17234 9998 17262
rect 10026 17234 10054 17262
rect 9554 16478 10054 17234
rect 9554 16450 9582 16478
rect 9610 16450 9634 16478
rect 9662 16450 9686 16478
rect 9714 16450 9738 16478
rect 9766 16450 9790 16478
rect 9818 16450 9842 16478
rect 9870 16450 9894 16478
rect 9922 16450 9946 16478
rect 9974 16450 9998 16478
rect 10026 16450 10054 16478
rect 9554 15694 10054 16450
rect 9554 15666 9582 15694
rect 9610 15666 9634 15694
rect 9662 15666 9686 15694
rect 9714 15666 9738 15694
rect 9766 15666 9790 15694
rect 9818 15666 9842 15694
rect 9870 15666 9894 15694
rect 9922 15666 9946 15694
rect 9974 15666 9998 15694
rect 10026 15666 10054 15694
rect 9554 14910 10054 15666
rect 9554 14882 9582 14910
rect 9610 14882 9634 14910
rect 9662 14882 9686 14910
rect 9714 14882 9738 14910
rect 9766 14882 9790 14910
rect 9818 14882 9842 14910
rect 9870 14882 9894 14910
rect 9922 14882 9946 14910
rect 9974 14882 9998 14910
rect 10026 14882 10054 14910
rect 9554 14126 10054 14882
rect 9554 14098 9582 14126
rect 9610 14098 9634 14126
rect 9662 14098 9686 14126
rect 9714 14098 9738 14126
rect 9766 14098 9790 14126
rect 9818 14098 9842 14126
rect 9870 14098 9894 14126
rect 9922 14098 9946 14126
rect 9974 14098 9998 14126
rect 10026 14098 10054 14126
rect 9554 13342 10054 14098
rect 9554 13314 9582 13342
rect 9610 13314 9634 13342
rect 9662 13314 9686 13342
rect 9714 13314 9738 13342
rect 9766 13314 9790 13342
rect 9818 13314 9842 13342
rect 9870 13314 9894 13342
rect 9922 13314 9946 13342
rect 9974 13314 9998 13342
rect 10026 13314 10054 13342
rect 9554 12558 10054 13314
rect 9554 12530 9582 12558
rect 9610 12530 9634 12558
rect 9662 12530 9686 12558
rect 9714 12530 9738 12558
rect 9766 12530 9790 12558
rect 9818 12530 9842 12558
rect 9870 12530 9894 12558
rect 9922 12530 9946 12558
rect 9974 12530 9998 12558
rect 10026 12530 10054 12558
rect 9554 11774 10054 12530
rect 9554 11746 9582 11774
rect 9610 11746 9634 11774
rect 9662 11746 9686 11774
rect 9714 11746 9738 11774
rect 9766 11746 9790 11774
rect 9818 11746 9842 11774
rect 9870 11746 9894 11774
rect 9922 11746 9946 11774
rect 9974 11746 9998 11774
rect 10026 11746 10054 11774
rect 9554 10990 10054 11746
rect 9554 10962 9582 10990
rect 9610 10962 9634 10990
rect 9662 10962 9686 10990
rect 9714 10962 9738 10990
rect 9766 10962 9790 10990
rect 9818 10962 9842 10990
rect 9870 10962 9894 10990
rect 9922 10962 9946 10990
rect 9974 10962 9998 10990
rect 10026 10962 10054 10990
rect 9554 10206 10054 10962
rect 9554 10178 9582 10206
rect 9610 10178 9634 10206
rect 9662 10178 9686 10206
rect 9714 10178 9738 10206
rect 9766 10178 9790 10206
rect 9818 10178 9842 10206
rect 9870 10178 9894 10206
rect 9922 10178 9946 10206
rect 9974 10178 9998 10206
rect 10026 10178 10054 10206
rect 9554 9422 10054 10178
rect 9554 9394 9582 9422
rect 9610 9394 9634 9422
rect 9662 9394 9686 9422
rect 9714 9394 9738 9422
rect 9766 9394 9790 9422
rect 9818 9394 9842 9422
rect 9870 9394 9894 9422
rect 9922 9394 9946 9422
rect 9974 9394 9998 9422
rect 10026 9394 10054 9422
rect 9554 8638 10054 9394
rect 9554 8610 9582 8638
rect 9610 8610 9634 8638
rect 9662 8610 9686 8638
rect 9714 8610 9738 8638
rect 9766 8610 9790 8638
rect 9818 8610 9842 8638
rect 9870 8610 9894 8638
rect 9922 8610 9946 8638
rect 9974 8610 9998 8638
rect 10026 8610 10054 8638
rect 9554 7854 10054 8610
rect 9554 7826 9582 7854
rect 9610 7826 9634 7854
rect 9662 7826 9686 7854
rect 9714 7826 9738 7854
rect 9766 7826 9790 7854
rect 9818 7826 9842 7854
rect 9870 7826 9894 7854
rect 9922 7826 9946 7854
rect 9974 7826 9998 7854
rect 10026 7826 10054 7854
rect 9554 7070 10054 7826
rect 9554 7042 9582 7070
rect 9610 7042 9634 7070
rect 9662 7042 9686 7070
rect 9714 7042 9738 7070
rect 9766 7042 9790 7070
rect 9818 7042 9842 7070
rect 9870 7042 9894 7070
rect 9922 7042 9946 7070
rect 9974 7042 9998 7070
rect 10026 7042 10054 7070
rect 9554 6286 10054 7042
rect 9554 6258 9582 6286
rect 9610 6258 9634 6286
rect 9662 6258 9686 6286
rect 9714 6258 9738 6286
rect 9766 6258 9790 6286
rect 9818 6258 9842 6286
rect 9870 6258 9894 6286
rect 9922 6258 9946 6286
rect 9974 6258 9998 6286
rect 10026 6258 10054 6286
rect 9554 5502 10054 6258
rect 9554 5474 9582 5502
rect 9610 5474 9634 5502
rect 9662 5474 9686 5502
rect 9714 5474 9738 5502
rect 9766 5474 9790 5502
rect 9818 5474 9842 5502
rect 9870 5474 9894 5502
rect 9922 5474 9946 5502
rect 9974 5474 9998 5502
rect 10026 5474 10054 5502
rect 9554 4718 10054 5474
rect 9554 4690 9582 4718
rect 9610 4690 9634 4718
rect 9662 4690 9686 4718
rect 9714 4690 9738 4718
rect 9766 4690 9790 4718
rect 9818 4690 9842 4718
rect 9870 4690 9894 4718
rect 9922 4690 9946 4718
rect 9974 4690 9998 4718
rect 10026 4690 10054 4718
rect 9554 3934 10054 4690
rect 9554 3906 9582 3934
rect 9610 3906 9634 3934
rect 9662 3906 9686 3934
rect 9714 3906 9738 3934
rect 9766 3906 9790 3934
rect 9818 3906 9842 3934
rect 9870 3906 9894 3934
rect 9922 3906 9946 3934
rect 9974 3906 9998 3934
rect 10026 3906 10054 3934
rect 9554 3150 10054 3906
rect 9554 3122 9582 3150
rect 9610 3122 9634 3150
rect 9662 3122 9686 3150
rect 9714 3122 9738 3150
rect 9766 3122 9790 3150
rect 9818 3122 9842 3150
rect 9870 3122 9894 3150
rect 9922 3122 9946 3150
rect 9974 3122 9998 3150
rect 10026 3122 10054 3150
rect 9554 2366 10054 3122
rect 9554 2338 9582 2366
rect 9610 2338 9634 2366
rect 9662 2338 9686 2366
rect 9714 2338 9738 2366
rect 9766 2338 9790 2366
rect 9818 2338 9842 2366
rect 9870 2338 9894 2366
rect 9922 2338 9946 2366
rect 9974 2338 9998 2366
rect 10026 2338 10054 2366
rect 9554 1582 10054 2338
rect 9554 1554 9582 1582
rect 9610 1554 9634 1582
rect 9662 1554 9686 1582
rect 9714 1554 9738 1582
rect 9766 1554 9790 1582
rect 9818 1554 9842 1582
rect 9870 1554 9894 1582
rect 9922 1554 9946 1582
rect 9974 1554 9998 1582
rect 10026 1554 10054 1582
rect 9554 1538 10054 1554
rect 12054 18438 12554 18454
rect 12054 18410 12082 18438
rect 12110 18410 12134 18438
rect 12162 18410 12186 18438
rect 12214 18410 12238 18438
rect 12266 18410 12290 18438
rect 12318 18410 12342 18438
rect 12370 18410 12394 18438
rect 12422 18410 12446 18438
rect 12474 18410 12498 18438
rect 12526 18410 12554 18438
rect 12054 17654 12554 18410
rect 12054 17626 12082 17654
rect 12110 17626 12134 17654
rect 12162 17626 12186 17654
rect 12214 17626 12238 17654
rect 12266 17626 12290 17654
rect 12318 17626 12342 17654
rect 12370 17626 12394 17654
rect 12422 17626 12446 17654
rect 12474 17626 12498 17654
rect 12526 17626 12554 17654
rect 12054 16870 12554 17626
rect 12054 16842 12082 16870
rect 12110 16842 12134 16870
rect 12162 16842 12186 16870
rect 12214 16842 12238 16870
rect 12266 16842 12290 16870
rect 12318 16842 12342 16870
rect 12370 16842 12394 16870
rect 12422 16842 12446 16870
rect 12474 16842 12498 16870
rect 12526 16842 12554 16870
rect 12054 16086 12554 16842
rect 12054 16058 12082 16086
rect 12110 16058 12134 16086
rect 12162 16058 12186 16086
rect 12214 16058 12238 16086
rect 12266 16058 12290 16086
rect 12318 16058 12342 16086
rect 12370 16058 12394 16086
rect 12422 16058 12446 16086
rect 12474 16058 12498 16086
rect 12526 16058 12554 16086
rect 12054 15302 12554 16058
rect 12054 15274 12082 15302
rect 12110 15274 12134 15302
rect 12162 15274 12186 15302
rect 12214 15274 12238 15302
rect 12266 15274 12290 15302
rect 12318 15274 12342 15302
rect 12370 15274 12394 15302
rect 12422 15274 12446 15302
rect 12474 15274 12498 15302
rect 12526 15274 12554 15302
rect 12054 14518 12554 15274
rect 12054 14490 12082 14518
rect 12110 14490 12134 14518
rect 12162 14490 12186 14518
rect 12214 14490 12238 14518
rect 12266 14490 12290 14518
rect 12318 14490 12342 14518
rect 12370 14490 12394 14518
rect 12422 14490 12446 14518
rect 12474 14490 12498 14518
rect 12526 14490 12554 14518
rect 12054 13734 12554 14490
rect 12054 13706 12082 13734
rect 12110 13706 12134 13734
rect 12162 13706 12186 13734
rect 12214 13706 12238 13734
rect 12266 13706 12290 13734
rect 12318 13706 12342 13734
rect 12370 13706 12394 13734
rect 12422 13706 12446 13734
rect 12474 13706 12498 13734
rect 12526 13706 12554 13734
rect 12054 12950 12554 13706
rect 12054 12922 12082 12950
rect 12110 12922 12134 12950
rect 12162 12922 12186 12950
rect 12214 12922 12238 12950
rect 12266 12922 12290 12950
rect 12318 12922 12342 12950
rect 12370 12922 12394 12950
rect 12422 12922 12446 12950
rect 12474 12922 12498 12950
rect 12526 12922 12554 12950
rect 12054 12166 12554 12922
rect 12054 12138 12082 12166
rect 12110 12138 12134 12166
rect 12162 12138 12186 12166
rect 12214 12138 12238 12166
rect 12266 12138 12290 12166
rect 12318 12138 12342 12166
rect 12370 12138 12394 12166
rect 12422 12138 12446 12166
rect 12474 12138 12498 12166
rect 12526 12138 12554 12166
rect 12054 11382 12554 12138
rect 12054 11354 12082 11382
rect 12110 11354 12134 11382
rect 12162 11354 12186 11382
rect 12214 11354 12238 11382
rect 12266 11354 12290 11382
rect 12318 11354 12342 11382
rect 12370 11354 12394 11382
rect 12422 11354 12446 11382
rect 12474 11354 12498 11382
rect 12526 11354 12554 11382
rect 12054 10598 12554 11354
rect 12054 10570 12082 10598
rect 12110 10570 12134 10598
rect 12162 10570 12186 10598
rect 12214 10570 12238 10598
rect 12266 10570 12290 10598
rect 12318 10570 12342 10598
rect 12370 10570 12394 10598
rect 12422 10570 12446 10598
rect 12474 10570 12498 10598
rect 12526 10570 12554 10598
rect 12054 9814 12554 10570
rect 12054 9786 12082 9814
rect 12110 9786 12134 9814
rect 12162 9786 12186 9814
rect 12214 9786 12238 9814
rect 12266 9786 12290 9814
rect 12318 9786 12342 9814
rect 12370 9786 12394 9814
rect 12422 9786 12446 9814
rect 12474 9786 12498 9814
rect 12526 9786 12554 9814
rect 12054 9030 12554 9786
rect 12054 9002 12082 9030
rect 12110 9002 12134 9030
rect 12162 9002 12186 9030
rect 12214 9002 12238 9030
rect 12266 9002 12290 9030
rect 12318 9002 12342 9030
rect 12370 9002 12394 9030
rect 12422 9002 12446 9030
rect 12474 9002 12498 9030
rect 12526 9002 12554 9030
rect 12054 8246 12554 9002
rect 12054 8218 12082 8246
rect 12110 8218 12134 8246
rect 12162 8218 12186 8246
rect 12214 8218 12238 8246
rect 12266 8218 12290 8246
rect 12318 8218 12342 8246
rect 12370 8218 12394 8246
rect 12422 8218 12446 8246
rect 12474 8218 12498 8246
rect 12526 8218 12554 8246
rect 12054 7462 12554 8218
rect 12054 7434 12082 7462
rect 12110 7434 12134 7462
rect 12162 7434 12186 7462
rect 12214 7434 12238 7462
rect 12266 7434 12290 7462
rect 12318 7434 12342 7462
rect 12370 7434 12394 7462
rect 12422 7434 12446 7462
rect 12474 7434 12498 7462
rect 12526 7434 12554 7462
rect 12054 6678 12554 7434
rect 12054 6650 12082 6678
rect 12110 6650 12134 6678
rect 12162 6650 12186 6678
rect 12214 6650 12238 6678
rect 12266 6650 12290 6678
rect 12318 6650 12342 6678
rect 12370 6650 12394 6678
rect 12422 6650 12446 6678
rect 12474 6650 12498 6678
rect 12526 6650 12554 6678
rect 12054 5894 12554 6650
rect 12054 5866 12082 5894
rect 12110 5866 12134 5894
rect 12162 5866 12186 5894
rect 12214 5866 12238 5894
rect 12266 5866 12290 5894
rect 12318 5866 12342 5894
rect 12370 5866 12394 5894
rect 12422 5866 12446 5894
rect 12474 5866 12498 5894
rect 12526 5866 12554 5894
rect 12054 5110 12554 5866
rect 12054 5082 12082 5110
rect 12110 5082 12134 5110
rect 12162 5082 12186 5110
rect 12214 5082 12238 5110
rect 12266 5082 12290 5110
rect 12318 5082 12342 5110
rect 12370 5082 12394 5110
rect 12422 5082 12446 5110
rect 12474 5082 12498 5110
rect 12526 5082 12554 5110
rect 12054 4326 12554 5082
rect 12054 4298 12082 4326
rect 12110 4298 12134 4326
rect 12162 4298 12186 4326
rect 12214 4298 12238 4326
rect 12266 4298 12290 4326
rect 12318 4298 12342 4326
rect 12370 4298 12394 4326
rect 12422 4298 12446 4326
rect 12474 4298 12498 4326
rect 12526 4298 12554 4326
rect 12054 3542 12554 4298
rect 12054 3514 12082 3542
rect 12110 3514 12134 3542
rect 12162 3514 12186 3542
rect 12214 3514 12238 3542
rect 12266 3514 12290 3542
rect 12318 3514 12342 3542
rect 12370 3514 12394 3542
rect 12422 3514 12446 3542
rect 12474 3514 12498 3542
rect 12526 3514 12554 3542
rect 12054 2758 12554 3514
rect 12054 2730 12082 2758
rect 12110 2730 12134 2758
rect 12162 2730 12186 2758
rect 12214 2730 12238 2758
rect 12266 2730 12290 2758
rect 12318 2730 12342 2758
rect 12370 2730 12394 2758
rect 12422 2730 12446 2758
rect 12474 2730 12498 2758
rect 12526 2730 12554 2758
rect 12054 1974 12554 2730
rect 12054 1946 12082 1974
rect 12110 1946 12134 1974
rect 12162 1946 12186 1974
rect 12214 1946 12238 1974
rect 12266 1946 12290 1974
rect 12318 1946 12342 1974
rect 12370 1946 12394 1974
rect 12422 1946 12446 1974
rect 12474 1946 12498 1974
rect 12526 1946 12554 1974
rect 12054 1538 12554 1946
rect 14554 18046 15054 18454
rect 14554 18018 14582 18046
rect 14610 18018 14634 18046
rect 14662 18018 14686 18046
rect 14714 18018 14738 18046
rect 14766 18018 14790 18046
rect 14818 18018 14842 18046
rect 14870 18018 14894 18046
rect 14922 18018 14946 18046
rect 14974 18018 14998 18046
rect 15026 18018 15054 18046
rect 14554 17262 15054 18018
rect 14554 17234 14582 17262
rect 14610 17234 14634 17262
rect 14662 17234 14686 17262
rect 14714 17234 14738 17262
rect 14766 17234 14790 17262
rect 14818 17234 14842 17262
rect 14870 17234 14894 17262
rect 14922 17234 14946 17262
rect 14974 17234 14998 17262
rect 15026 17234 15054 17262
rect 14554 16478 15054 17234
rect 14554 16450 14582 16478
rect 14610 16450 14634 16478
rect 14662 16450 14686 16478
rect 14714 16450 14738 16478
rect 14766 16450 14790 16478
rect 14818 16450 14842 16478
rect 14870 16450 14894 16478
rect 14922 16450 14946 16478
rect 14974 16450 14998 16478
rect 15026 16450 15054 16478
rect 14554 15694 15054 16450
rect 14554 15666 14582 15694
rect 14610 15666 14634 15694
rect 14662 15666 14686 15694
rect 14714 15666 14738 15694
rect 14766 15666 14790 15694
rect 14818 15666 14842 15694
rect 14870 15666 14894 15694
rect 14922 15666 14946 15694
rect 14974 15666 14998 15694
rect 15026 15666 15054 15694
rect 14554 14910 15054 15666
rect 14554 14882 14582 14910
rect 14610 14882 14634 14910
rect 14662 14882 14686 14910
rect 14714 14882 14738 14910
rect 14766 14882 14790 14910
rect 14818 14882 14842 14910
rect 14870 14882 14894 14910
rect 14922 14882 14946 14910
rect 14974 14882 14998 14910
rect 15026 14882 15054 14910
rect 14554 14126 15054 14882
rect 14554 14098 14582 14126
rect 14610 14098 14634 14126
rect 14662 14098 14686 14126
rect 14714 14098 14738 14126
rect 14766 14098 14790 14126
rect 14818 14098 14842 14126
rect 14870 14098 14894 14126
rect 14922 14098 14946 14126
rect 14974 14098 14998 14126
rect 15026 14098 15054 14126
rect 14554 13342 15054 14098
rect 14554 13314 14582 13342
rect 14610 13314 14634 13342
rect 14662 13314 14686 13342
rect 14714 13314 14738 13342
rect 14766 13314 14790 13342
rect 14818 13314 14842 13342
rect 14870 13314 14894 13342
rect 14922 13314 14946 13342
rect 14974 13314 14998 13342
rect 15026 13314 15054 13342
rect 14554 12558 15054 13314
rect 14554 12530 14582 12558
rect 14610 12530 14634 12558
rect 14662 12530 14686 12558
rect 14714 12530 14738 12558
rect 14766 12530 14790 12558
rect 14818 12530 14842 12558
rect 14870 12530 14894 12558
rect 14922 12530 14946 12558
rect 14974 12530 14998 12558
rect 15026 12530 15054 12558
rect 14554 11774 15054 12530
rect 14554 11746 14582 11774
rect 14610 11746 14634 11774
rect 14662 11746 14686 11774
rect 14714 11746 14738 11774
rect 14766 11746 14790 11774
rect 14818 11746 14842 11774
rect 14870 11746 14894 11774
rect 14922 11746 14946 11774
rect 14974 11746 14998 11774
rect 15026 11746 15054 11774
rect 14554 10990 15054 11746
rect 14554 10962 14582 10990
rect 14610 10962 14634 10990
rect 14662 10962 14686 10990
rect 14714 10962 14738 10990
rect 14766 10962 14790 10990
rect 14818 10962 14842 10990
rect 14870 10962 14894 10990
rect 14922 10962 14946 10990
rect 14974 10962 14998 10990
rect 15026 10962 15054 10990
rect 14554 10206 15054 10962
rect 14554 10178 14582 10206
rect 14610 10178 14634 10206
rect 14662 10178 14686 10206
rect 14714 10178 14738 10206
rect 14766 10178 14790 10206
rect 14818 10178 14842 10206
rect 14870 10178 14894 10206
rect 14922 10178 14946 10206
rect 14974 10178 14998 10206
rect 15026 10178 15054 10206
rect 14554 9422 15054 10178
rect 14554 9394 14582 9422
rect 14610 9394 14634 9422
rect 14662 9394 14686 9422
rect 14714 9394 14738 9422
rect 14766 9394 14790 9422
rect 14818 9394 14842 9422
rect 14870 9394 14894 9422
rect 14922 9394 14946 9422
rect 14974 9394 14998 9422
rect 15026 9394 15054 9422
rect 14554 8638 15054 9394
rect 14554 8610 14582 8638
rect 14610 8610 14634 8638
rect 14662 8610 14686 8638
rect 14714 8610 14738 8638
rect 14766 8610 14790 8638
rect 14818 8610 14842 8638
rect 14870 8610 14894 8638
rect 14922 8610 14946 8638
rect 14974 8610 14998 8638
rect 15026 8610 15054 8638
rect 14554 7854 15054 8610
rect 14554 7826 14582 7854
rect 14610 7826 14634 7854
rect 14662 7826 14686 7854
rect 14714 7826 14738 7854
rect 14766 7826 14790 7854
rect 14818 7826 14842 7854
rect 14870 7826 14894 7854
rect 14922 7826 14946 7854
rect 14974 7826 14998 7854
rect 15026 7826 15054 7854
rect 14554 7070 15054 7826
rect 14554 7042 14582 7070
rect 14610 7042 14634 7070
rect 14662 7042 14686 7070
rect 14714 7042 14738 7070
rect 14766 7042 14790 7070
rect 14818 7042 14842 7070
rect 14870 7042 14894 7070
rect 14922 7042 14946 7070
rect 14974 7042 14998 7070
rect 15026 7042 15054 7070
rect 14554 6286 15054 7042
rect 14554 6258 14582 6286
rect 14610 6258 14634 6286
rect 14662 6258 14686 6286
rect 14714 6258 14738 6286
rect 14766 6258 14790 6286
rect 14818 6258 14842 6286
rect 14870 6258 14894 6286
rect 14922 6258 14946 6286
rect 14974 6258 14998 6286
rect 15026 6258 15054 6286
rect 14554 5502 15054 6258
rect 14554 5474 14582 5502
rect 14610 5474 14634 5502
rect 14662 5474 14686 5502
rect 14714 5474 14738 5502
rect 14766 5474 14790 5502
rect 14818 5474 14842 5502
rect 14870 5474 14894 5502
rect 14922 5474 14946 5502
rect 14974 5474 14998 5502
rect 15026 5474 15054 5502
rect 14554 4718 15054 5474
rect 14554 4690 14582 4718
rect 14610 4690 14634 4718
rect 14662 4690 14686 4718
rect 14714 4690 14738 4718
rect 14766 4690 14790 4718
rect 14818 4690 14842 4718
rect 14870 4690 14894 4718
rect 14922 4690 14946 4718
rect 14974 4690 14998 4718
rect 15026 4690 15054 4718
rect 14554 3934 15054 4690
rect 14554 3906 14582 3934
rect 14610 3906 14634 3934
rect 14662 3906 14686 3934
rect 14714 3906 14738 3934
rect 14766 3906 14790 3934
rect 14818 3906 14842 3934
rect 14870 3906 14894 3934
rect 14922 3906 14946 3934
rect 14974 3906 14998 3934
rect 15026 3906 15054 3934
rect 14554 3150 15054 3906
rect 14554 3122 14582 3150
rect 14610 3122 14634 3150
rect 14662 3122 14686 3150
rect 14714 3122 14738 3150
rect 14766 3122 14790 3150
rect 14818 3122 14842 3150
rect 14870 3122 14894 3150
rect 14922 3122 14946 3150
rect 14974 3122 14998 3150
rect 15026 3122 15054 3150
rect 14554 2366 15054 3122
rect 14554 2338 14582 2366
rect 14610 2338 14634 2366
rect 14662 2338 14686 2366
rect 14714 2338 14738 2366
rect 14766 2338 14790 2366
rect 14818 2338 14842 2366
rect 14870 2338 14894 2366
rect 14922 2338 14946 2366
rect 14974 2338 14998 2366
rect 15026 2338 15054 2366
rect 14554 1582 15054 2338
rect 14554 1554 14582 1582
rect 14610 1554 14634 1582
rect 14662 1554 14686 1582
rect 14714 1554 14738 1582
rect 14766 1554 14790 1582
rect 14818 1554 14842 1582
rect 14870 1554 14894 1582
rect 14922 1554 14946 1582
rect 14974 1554 14998 1582
rect 15026 1554 15054 1582
rect 14554 1538 15054 1554
rect 17054 18438 17554 18454
rect 17054 18410 17082 18438
rect 17110 18410 17134 18438
rect 17162 18410 17186 18438
rect 17214 18410 17238 18438
rect 17266 18410 17290 18438
rect 17318 18410 17342 18438
rect 17370 18410 17394 18438
rect 17422 18410 17446 18438
rect 17474 18410 17498 18438
rect 17526 18410 17554 18438
rect 17054 17654 17554 18410
rect 17054 17626 17082 17654
rect 17110 17626 17134 17654
rect 17162 17626 17186 17654
rect 17214 17626 17238 17654
rect 17266 17626 17290 17654
rect 17318 17626 17342 17654
rect 17370 17626 17394 17654
rect 17422 17626 17446 17654
rect 17474 17626 17498 17654
rect 17526 17626 17554 17654
rect 17054 16870 17554 17626
rect 17054 16842 17082 16870
rect 17110 16842 17134 16870
rect 17162 16842 17186 16870
rect 17214 16842 17238 16870
rect 17266 16842 17290 16870
rect 17318 16842 17342 16870
rect 17370 16842 17394 16870
rect 17422 16842 17446 16870
rect 17474 16842 17498 16870
rect 17526 16842 17554 16870
rect 17054 16086 17554 16842
rect 17054 16058 17082 16086
rect 17110 16058 17134 16086
rect 17162 16058 17186 16086
rect 17214 16058 17238 16086
rect 17266 16058 17290 16086
rect 17318 16058 17342 16086
rect 17370 16058 17394 16086
rect 17422 16058 17446 16086
rect 17474 16058 17498 16086
rect 17526 16058 17554 16086
rect 17054 15302 17554 16058
rect 17054 15274 17082 15302
rect 17110 15274 17134 15302
rect 17162 15274 17186 15302
rect 17214 15274 17238 15302
rect 17266 15274 17290 15302
rect 17318 15274 17342 15302
rect 17370 15274 17394 15302
rect 17422 15274 17446 15302
rect 17474 15274 17498 15302
rect 17526 15274 17554 15302
rect 17054 14518 17554 15274
rect 17054 14490 17082 14518
rect 17110 14490 17134 14518
rect 17162 14490 17186 14518
rect 17214 14490 17238 14518
rect 17266 14490 17290 14518
rect 17318 14490 17342 14518
rect 17370 14490 17394 14518
rect 17422 14490 17446 14518
rect 17474 14490 17498 14518
rect 17526 14490 17554 14518
rect 17054 13734 17554 14490
rect 17054 13706 17082 13734
rect 17110 13706 17134 13734
rect 17162 13706 17186 13734
rect 17214 13706 17238 13734
rect 17266 13706 17290 13734
rect 17318 13706 17342 13734
rect 17370 13706 17394 13734
rect 17422 13706 17446 13734
rect 17474 13706 17498 13734
rect 17526 13706 17554 13734
rect 17054 12950 17554 13706
rect 17054 12922 17082 12950
rect 17110 12922 17134 12950
rect 17162 12922 17186 12950
rect 17214 12922 17238 12950
rect 17266 12922 17290 12950
rect 17318 12922 17342 12950
rect 17370 12922 17394 12950
rect 17422 12922 17446 12950
rect 17474 12922 17498 12950
rect 17526 12922 17554 12950
rect 17054 12166 17554 12922
rect 17054 12138 17082 12166
rect 17110 12138 17134 12166
rect 17162 12138 17186 12166
rect 17214 12138 17238 12166
rect 17266 12138 17290 12166
rect 17318 12138 17342 12166
rect 17370 12138 17394 12166
rect 17422 12138 17446 12166
rect 17474 12138 17498 12166
rect 17526 12138 17554 12166
rect 17054 11382 17554 12138
rect 17054 11354 17082 11382
rect 17110 11354 17134 11382
rect 17162 11354 17186 11382
rect 17214 11354 17238 11382
rect 17266 11354 17290 11382
rect 17318 11354 17342 11382
rect 17370 11354 17394 11382
rect 17422 11354 17446 11382
rect 17474 11354 17498 11382
rect 17526 11354 17554 11382
rect 17054 10598 17554 11354
rect 17054 10570 17082 10598
rect 17110 10570 17134 10598
rect 17162 10570 17186 10598
rect 17214 10570 17238 10598
rect 17266 10570 17290 10598
rect 17318 10570 17342 10598
rect 17370 10570 17394 10598
rect 17422 10570 17446 10598
rect 17474 10570 17498 10598
rect 17526 10570 17554 10598
rect 17054 9814 17554 10570
rect 17054 9786 17082 9814
rect 17110 9786 17134 9814
rect 17162 9786 17186 9814
rect 17214 9786 17238 9814
rect 17266 9786 17290 9814
rect 17318 9786 17342 9814
rect 17370 9786 17394 9814
rect 17422 9786 17446 9814
rect 17474 9786 17498 9814
rect 17526 9786 17554 9814
rect 17054 9030 17554 9786
rect 17054 9002 17082 9030
rect 17110 9002 17134 9030
rect 17162 9002 17186 9030
rect 17214 9002 17238 9030
rect 17266 9002 17290 9030
rect 17318 9002 17342 9030
rect 17370 9002 17394 9030
rect 17422 9002 17446 9030
rect 17474 9002 17498 9030
rect 17526 9002 17554 9030
rect 17054 8246 17554 9002
rect 17054 8218 17082 8246
rect 17110 8218 17134 8246
rect 17162 8218 17186 8246
rect 17214 8218 17238 8246
rect 17266 8218 17290 8246
rect 17318 8218 17342 8246
rect 17370 8218 17394 8246
rect 17422 8218 17446 8246
rect 17474 8218 17498 8246
rect 17526 8218 17554 8246
rect 17054 7462 17554 8218
rect 17054 7434 17082 7462
rect 17110 7434 17134 7462
rect 17162 7434 17186 7462
rect 17214 7434 17238 7462
rect 17266 7434 17290 7462
rect 17318 7434 17342 7462
rect 17370 7434 17394 7462
rect 17422 7434 17446 7462
rect 17474 7434 17498 7462
rect 17526 7434 17554 7462
rect 17054 6678 17554 7434
rect 17054 6650 17082 6678
rect 17110 6650 17134 6678
rect 17162 6650 17186 6678
rect 17214 6650 17238 6678
rect 17266 6650 17290 6678
rect 17318 6650 17342 6678
rect 17370 6650 17394 6678
rect 17422 6650 17446 6678
rect 17474 6650 17498 6678
rect 17526 6650 17554 6678
rect 17054 5894 17554 6650
rect 17054 5866 17082 5894
rect 17110 5866 17134 5894
rect 17162 5866 17186 5894
rect 17214 5866 17238 5894
rect 17266 5866 17290 5894
rect 17318 5866 17342 5894
rect 17370 5866 17394 5894
rect 17422 5866 17446 5894
rect 17474 5866 17498 5894
rect 17526 5866 17554 5894
rect 17054 5110 17554 5866
rect 17054 5082 17082 5110
rect 17110 5082 17134 5110
rect 17162 5082 17186 5110
rect 17214 5082 17238 5110
rect 17266 5082 17290 5110
rect 17318 5082 17342 5110
rect 17370 5082 17394 5110
rect 17422 5082 17446 5110
rect 17474 5082 17498 5110
rect 17526 5082 17554 5110
rect 17054 4326 17554 5082
rect 17054 4298 17082 4326
rect 17110 4298 17134 4326
rect 17162 4298 17186 4326
rect 17214 4298 17238 4326
rect 17266 4298 17290 4326
rect 17318 4298 17342 4326
rect 17370 4298 17394 4326
rect 17422 4298 17446 4326
rect 17474 4298 17498 4326
rect 17526 4298 17554 4326
rect 17054 3542 17554 4298
rect 17054 3514 17082 3542
rect 17110 3514 17134 3542
rect 17162 3514 17186 3542
rect 17214 3514 17238 3542
rect 17266 3514 17290 3542
rect 17318 3514 17342 3542
rect 17370 3514 17394 3542
rect 17422 3514 17446 3542
rect 17474 3514 17498 3542
rect 17526 3514 17554 3542
rect 17054 2758 17554 3514
rect 17054 2730 17082 2758
rect 17110 2730 17134 2758
rect 17162 2730 17186 2758
rect 17214 2730 17238 2758
rect 17266 2730 17290 2758
rect 17318 2730 17342 2758
rect 17370 2730 17394 2758
rect 17422 2730 17446 2758
rect 17474 2730 17498 2758
rect 17526 2730 17554 2758
rect 17054 1974 17554 2730
rect 17054 1946 17082 1974
rect 17110 1946 17134 1974
rect 17162 1946 17186 1974
rect 17214 1946 17238 1974
rect 17266 1946 17290 1974
rect 17318 1946 17342 1974
rect 17370 1946 17394 1974
rect 17422 1946 17446 1974
rect 17474 1946 17498 1974
rect 17526 1946 17554 1974
rect 17054 1538 17554 1946
rect 19554 18046 20054 18454
rect 19554 18018 19582 18046
rect 19610 18018 19634 18046
rect 19662 18018 19686 18046
rect 19714 18018 19738 18046
rect 19766 18018 19790 18046
rect 19818 18018 19842 18046
rect 19870 18018 19894 18046
rect 19922 18018 19946 18046
rect 19974 18018 19998 18046
rect 20026 18018 20054 18046
rect 19554 17262 20054 18018
rect 19554 17234 19582 17262
rect 19610 17234 19634 17262
rect 19662 17234 19686 17262
rect 19714 17234 19738 17262
rect 19766 17234 19790 17262
rect 19818 17234 19842 17262
rect 19870 17234 19894 17262
rect 19922 17234 19946 17262
rect 19974 17234 19998 17262
rect 20026 17234 20054 17262
rect 19554 16478 20054 17234
rect 19554 16450 19582 16478
rect 19610 16450 19634 16478
rect 19662 16450 19686 16478
rect 19714 16450 19738 16478
rect 19766 16450 19790 16478
rect 19818 16450 19842 16478
rect 19870 16450 19894 16478
rect 19922 16450 19946 16478
rect 19974 16450 19998 16478
rect 20026 16450 20054 16478
rect 19554 15694 20054 16450
rect 19554 15666 19582 15694
rect 19610 15666 19634 15694
rect 19662 15666 19686 15694
rect 19714 15666 19738 15694
rect 19766 15666 19790 15694
rect 19818 15666 19842 15694
rect 19870 15666 19894 15694
rect 19922 15666 19946 15694
rect 19974 15666 19998 15694
rect 20026 15666 20054 15694
rect 19554 14910 20054 15666
rect 19554 14882 19582 14910
rect 19610 14882 19634 14910
rect 19662 14882 19686 14910
rect 19714 14882 19738 14910
rect 19766 14882 19790 14910
rect 19818 14882 19842 14910
rect 19870 14882 19894 14910
rect 19922 14882 19946 14910
rect 19974 14882 19998 14910
rect 20026 14882 20054 14910
rect 19554 14126 20054 14882
rect 19554 14098 19582 14126
rect 19610 14098 19634 14126
rect 19662 14098 19686 14126
rect 19714 14098 19738 14126
rect 19766 14098 19790 14126
rect 19818 14098 19842 14126
rect 19870 14098 19894 14126
rect 19922 14098 19946 14126
rect 19974 14098 19998 14126
rect 20026 14098 20054 14126
rect 19554 13342 20054 14098
rect 19554 13314 19582 13342
rect 19610 13314 19634 13342
rect 19662 13314 19686 13342
rect 19714 13314 19738 13342
rect 19766 13314 19790 13342
rect 19818 13314 19842 13342
rect 19870 13314 19894 13342
rect 19922 13314 19946 13342
rect 19974 13314 19998 13342
rect 20026 13314 20054 13342
rect 19554 12558 20054 13314
rect 19554 12530 19582 12558
rect 19610 12530 19634 12558
rect 19662 12530 19686 12558
rect 19714 12530 19738 12558
rect 19766 12530 19790 12558
rect 19818 12530 19842 12558
rect 19870 12530 19894 12558
rect 19922 12530 19946 12558
rect 19974 12530 19998 12558
rect 20026 12530 20054 12558
rect 19554 11774 20054 12530
rect 19554 11746 19582 11774
rect 19610 11746 19634 11774
rect 19662 11746 19686 11774
rect 19714 11746 19738 11774
rect 19766 11746 19790 11774
rect 19818 11746 19842 11774
rect 19870 11746 19894 11774
rect 19922 11746 19946 11774
rect 19974 11746 19998 11774
rect 20026 11746 20054 11774
rect 19554 10990 20054 11746
rect 19554 10962 19582 10990
rect 19610 10962 19634 10990
rect 19662 10962 19686 10990
rect 19714 10962 19738 10990
rect 19766 10962 19790 10990
rect 19818 10962 19842 10990
rect 19870 10962 19894 10990
rect 19922 10962 19946 10990
rect 19974 10962 19998 10990
rect 20026 10962 20054 10990
rect 19554 10206 20054 10962
rect 19554 10178 19582 10206
rect 19610 10178 19634 10206
rect 19662 10178 19686 10206
rect 19714 10178 19738 10206
rect 19766 10178 19790 10206
rect 19818 10178 19842 10206
rect 19870 10178 19894 10206
rect 19922 10178 19946 10206
rect 19974 10178 19998 10206
rect 20026 10178 20054 10206
rect 19554 9422 20054 10178
rect 19554 9394 19582 9422
rect 19610 9394 19634 9422
rect 19662 9394 19686 9422
rect 19714 9394 19738 9422
rect 19766 9394 19790 9422
rect 19818 9394 19842 9422
rect 19870 9394 19894 9422
rect 19922 9394 19946 9422
rect 19974 9394 19998 9422
rect 20026 9394 20054 9422
rect 19554 8638 20054 9394
rect 19554 8610 19582 8638
rect 19610 8610 19634 8638
rect 19662 8610 19686 8638
rect 19714 8610 19738 8638
rect 19766 8610 19790 8638
rect 19818 8610 19842 8638
rect 19870 8610 19894 8638
rect 19922 8610 19946 8638
rect 19974 8610 19998 8638
rect 20026 8610 20054 8638
rect 19554 7854 20054 8610
rect 19554 7826 19582 7854
rect 19610 7826 19634 7854
rect 19662 7826 19686 7854
rect 19714 7826 19738 7854
rect 19766 7826 19790 7854
rect 19818 7826 19842 7854
rect 19870 7826 19894 7854
rect 19922 7826 19946 7854
rect 19974 7826 19998 7854
rect 20026 7826 20054 7854
rect 19554 7070 20054 7826
rect 19554 7042 19582 7070
rect 19610 7042 19634 7070
rect 19662 7042 19686 7070
rect 19714 7042 19738 7070
rect 19766 7042 19790 7070
rect 19818 7042 19842 7070
rect 19870 7042 19894 7070
rect 19922 7042 19946 7070
rect 19974 7042 19998 7070
rect 20026 7042 20054 7070
rect 19554 6286 20054 7042
rect 19554 6258 19582 6286
rect 19610 6258 19634 6286
rect 19662 6258 19686 6286
rect 19714 6258 19738 6286
rect 19766 6258 19790 6286
rect 19818 6258 19842 6286
rect 19870 6258 19894 6286
rect 19922 6258 19946 6286
rect 19974 6258 19998 6286
rect 20026 6258 20054 6286
rect 19554 5502 20054 6258
rect 19554 5474 19582 5502
rect 19610 5474 19634 5502
rect 19662 5474 19686 5502
rect 19714 5474 19738 5502
rect 19766 5474 19790 5502
rect 19818 5474 19842 5502
rect 19870 5474 19894 5502
rect 19922 5474 19946 5502
rect 19974 5474 19998 5502
rect 20026 5474 20054 5502
rect 19554 4718 20054 5474
rect 19554 4690 19582 4718
rect 19610 4690 19634 4718
rect 19662 4690 19686 4718
rect 19714 4690 19738 4718
rect 19766 4690 19790 4718
rect 19818 4690 19842 4718
rect 19870 4690 19894 4718
rect 19922 4690 19946 4718
rect 19974 4690 19998 4718
rect 20026 4690 20054 4718
rect 19554 3934 20054 4690
rect 19554 3906 19582 3934
rect 19610 3906 19634 3934
rect 19662 3906 19686 3934
rect 19714 3906 19738 3934
rect 19766 3906 19790 3934
rect 19818 3906 19842 3934
rect 19870 3906 19894 3934
rect 19922 3906 19946 3934
rect 19974 3906 19998 3934
rect 20026 3906 20054 3934
rect 19554 3150 20054 3906
rect 19554 3122 19582 3150
rect 19610 3122 19634 3150
rect 19662 3122 19686 3150
rect 19714 3122 19738 3150
rect 19766 3122 19790 3150
rect 19818 3122 19842 3150
rect 19870 3122 19894 3150
rect 19922 3122 19946 3150
rect 19974 3122 19998 3150
rect 20026 3122 20054 3150
rect 19554 2366 20054 3122
rect 19554 2338 19582 2366
rect 19610 2338 19634 2366
rect 19662 2338 19686 2366
rect 19714 2338 19738 2366
rect 19766 2338 19790 2366
rect 19818 2338 19842 2366
rect 19870 2338 19894 2366
rect 19922 2338 19946 2366
rect 19974 2338 19998 2366
rect 20026 2338 20054 2366
rect 19554 1582 20054 2338
rect 19554 1554 19582 1582
rect 19610 1554 19634 1582
rect 19662 1554 19686 1582
rect 19714 1554 19738 1582
rect 19766 1554 19790 1582
rect 19818 1554 19842 1582
rect 19870 1554 19894 1582
rect 19922 1554 19946 1582
rect 19974 1554 19998 1582
rect 20026 1554 20054 1582
rect 19554 1538 20054 1554
rect 22054 18438 22554 18454
rect 22054 18410 22082 18438
rect 22110 18410 22134 18438
rect 22162 18410 22186 18438
rect 22214 18410 22238 18438
rect 22266 18410 22290 18438
rect 22318 18410 22342 18438
rect 22370 18410 22394 18438
rect 22422 18410 22446 18438
rect 22474 18410 22498 18438
rect 22526 18410 22554 18438
rect 22054 17654 22554 18410
rect 22054 17626 22082 17654
rect 22110 17626 22134 17654
rect 22162 17626 22186 17654
rect 22214 17626 22238 17654
rect 22266 17626 22290 17654
rect 22318 17626 22342 17654
rect 22370 17626 22394 17654
rect 22422 17626 22446 17654
rect 22474 17626 22498 17654
rect 22526 17626 22554 17654
rect 22054 16870 22554 17626
rect 22054 16842 22082 16870
rect 22110 16842 22134 16870
rect 22162 16842 22186 16870
rect 22214 16842 22238 16870
rect 22266 16842 22290 16870
rect 22318 16842 22342 16870
rect 22370 16842 22394 16870
rect 22422 16842 22446 16870
rect 22474 16842 22498 16870
rect 22526 16842 22554 16870
rect 22054 16086 22554 16842
rect 22054 16058 22082 16086
rect 22110 16058 22134 16086
rect 22162 16058 22186 16086
rect 22214 16058 22238 16086
rect 22266 16058 22290 16086
rect 22318 16058 22342 16086
rect 22370 16058 22394 16086
rect 22422 16058 22446 16086
rect 22474 16058 22498 16086
rect 22526 16058 22554 16086
rect 22054 15302 22554 16058
rect 22054 15274 22082 15302
rect 22110 15274 22134 15302
rect 22162 15274 22186 15302
rect 22214 15274 22238 15302
rect 22266 15274 22290 15302
rect 22318 15274 22342 15302
rect 22370 15274 22394 15302
rect 22422 15274 22446 15302
rect 22474 15274 22498 15302
rect 22526 15274 22554 15302
rect 22054 14518 22554 15274
rect 22054 14490 22082 14518
rect 22110 14490 22134 14518
rect 22162 14490 22186 14518
rect 22214 14490 22238 14518
rect 22266 14490 22290 14518
rect 22318 14490 22342 14518
rect 22370 14490 22394 14518
rect 22422 14490 22446 14518
rect 22474 14490 22498 14518
rect 22526 14490 22554 14518
rect 22054 13734 22554 14490
rect 22054 13706 22082 13734
rect 22110 13706 22134 13734
rect 22162 13706 22186 13734
rect 22214 13706 22238 13734
rect 22266 13706 22290 13734
rect 22318 13706 22342 13734
rect 22370 13706 22394 13734
rect 22422 13706 22446 13734
rect 22474 13706 22498 13734
rect 22526 13706 22554 13734
rect 22054 12950 22554 13706
rect 22054 12922 22082 12950
rect 22110 12922 22134 12950
rect 22162 12922 22186 12950
rect 22214 12922 22238 12950
rect 22266 12922 22290 12950
rect 22318 12922 22342 12950
rect 22370 12922 22394 12950
rect 22422 12922 22446 12950
rect 22474 12922 22498 12950
rect 22526 12922 22554 12950
rect 22054 12166 22554 12922
rect 22054 12138 22082 12166
rect 22110 12138 22134 12166
rect 22162 12138 22186 12166
rect 22214 12138 22238 12166
rect 22266 12138 22290 12166
rect 22318 12138 22342 12166
rect 22370 12138 22394 12166
rect 22422 12138 22446 12166
rect 22474 12138 22498 12166
rect 22526 12138 22554 12166
rect 22054 11382 22554 12138
rect 22054 11354 22082 11382
rect 22110 11354 22134 11382
rect 22162 11354 22186 11382
rect 22214 11354 22238 11382
rect 22266 11354 22290 11382
rect 22318 11354 22342 11382
rect 22370 11354 22394 11382
rect 22422 11354 22446 11382
rect 22474 11354 22498 11382
rect 22526 11354 22554 11382
rect 22054 10598 22554 11354
rect 22054 10570 22082 10598
rect 22110 10570 22134 10598
rect 22162 10570 22186 10598
rect 22214 10570 22238 10598
rect 22266 10570 22290 10598
rect 22318 10570 22342 10598
rect 22370 10570 22394 10598
rect 22422 10570 22446 10598
rect 22474 10570 22498 10598
rect 22526 10570 22554 10598
rect 22054 9814 22554 10570
rect 22054 9786 22082 9814
rect 22110 9786 22134 9814
rect 22162 9786 22186 9814
rect 22214 9786 22238 9814
rect 22266 9786 22290 9814
rect 22318 9786 22342 9814
rect 22370 9786 22394 9814
rect 22422 9786 22446 9814
rect 22474 9786 22498 9814
rect 22526 9786 22554 9814
rect 22054 9030 22554 9786
rect 22054 9002 22082 9030
rect 22110 9002 22134 9030
rect 22162 9002 22186 9030
rect 22214 9002 22238 9030
rect 22266 9002 22290 9030
rect 22318 9002 22342 9030
rect 22370 9002 22394 9030
rect 22422 9002 22446 9030
rect 22474 9002 22498 9030
rect 22526 9002 22554 9030
rect 22054 8246 22554 9002
rect 22054 8218 22082 8246
rect 22110 8218 22134 8246
rect 22162 8218 22186 8246
rect 22214 8218 22238 8246
rect 22266 8218 22290 8246
rect 22318 8218 22342 8246
rect 22370 8218 22394 8246
rect 22422 8218 22446 8246
rect 22474 8218 22498 8246
rect 22526 8218 22554 8246
rect 22054 7462 22554 8218
rect 22054 7434 22082 7462
rect 22110 7434 22134 7462
rect 22162 7434 22186 7462
rect 22214 7434 22238 7462
rect 22266 7434 22290 7462
rect 22318 7434 22342 7462
rect 22370 7434 22394 7462
rect 22422 7434 22446 7462
rect 22474 7434 22498 7462
rect 22526 7434 22554 7462
rect 22054 6678 22554 7434
rect 22054 6650 22082 6678
rect 22110 6650 22134 6678
rect 22162 6650 22186 6678
rect 22214 6650 22238 6678
rect 22266 6650 22290 6678
rect 22318 6650 22342 6678
rect 22370 6650 22394 6678
rect 22422 6650 22446 6678
rect 22474 6650 22498 6678
rect 22526 6650 22554 6678
rect 22054 5894 22554 6650
rect 22054 5866 22082 5894
rect 22110 5866 22134 5894
rect 22162 5866 22186 5894
rect 22214 5866 22238 5894
rect 22266 5866 22290 5894
rect 22318 5866 22342 5894
rect 22370 5866 22394 5894
rect 22422 5866 22446 5894
rect 22474 5866 22498 5894
rect 22526 5866 22554 5894
rect 22054 5110 22554 5866
rect 22054 5082 22082 5110
rect 22110 5082 22134 5110
rect 22162 5082 22186 5110
rect 22214 5082 22238 5110
rect 22266 5082 22290 5110
rect 22318 5082 22342 5110
rect 22370 5082 22394 5110
rect 22422 5082 22446 5110
rect 22474 5082 22498 5110
rect 22526 5082 22554 5110
rect 22054 4326 22554 5082
rect 22054 4298 22082 4326
rect 22110 4298 22134 4326
rect 22162 4298 22186 4326
rect 22214 4298 22238 4326
rect 22266 4298 22290 4326
rect 22318 4298 22342 4326
rect 22370 4298 22394 4326
rect 22422 4298 22446 4326
rect 22474 4298 22498 4326
rect 22526 4298 22554 4326
rect 22054 3542 22554 4298
rect 22054 3514 22082 3542
rect 22110 3514 22134 3542
rect 22162 3514 22186 3542
rect 22214 3514 22238 3542
rect 22266 3514 22290 3542
rect 22318 3514 22342 3542
rect 22370 3514 22394 3542
rect 22422 3514 22446 3542
rect 22474 3514 22498 3542
rect 22526 3514 22554 3542
rect 22054 2758 22554 3514
rect 22054 2730 22082 2758
rect 22110 2730 22134 2758
rect 22162 2730 22186 2758
rect 22214 2730 22238 2758
rect 22266 2730 22290 2758
rect 22318 2730 22342 2758
rect 22370 2730 22394 2758
rect 22422 2730 22446 2758
rect 22474 2730 22498 2758
rect 22526 2730 22554 2758
rect 22054 1974 22554 2730
rect 22054 1946 22082 1974
rect 22110 1946 22134 1974
rect 22162 1946 22186 1974
rect 22214 1946 22238 1974
rect 22266 1946 22290 1974
rect 22318 1946 22342 1974
rect 22370 1946 22394 1974
rect 22422 1946 22446 1974
rect 22474 1946 22498 1974
rect 22526 1946 22554 1974
rect 22054 1538 22554 1946
rect 24554 18046 25054 18454
rect 24554 18018 24582 18046
rect 24610 18018 24634 18046
rect 24662 18018 24686 18046
rect 24714 18018 24738 18046
rect 24766 18018 24790 18046
rect 24818 18018 24842 18046
rect 24870 18018 24894 18046
rect 24922 18018 24946 18046
rect 24974 18018 24998 18046
rect 25026 18018 25054 18046
rect 24554 17262 25054 18018
rect 24554 17234 24582 17262
rect 24610 17234 24634 17262
rect 24662 17234 24686 17262
rect 24714 17234 24738 17262
rect 24766 17234 24790 17262
rect 24818 17234 24842 17262
rect 24870 17234 24894 17262
rect 24922 17234 24946 17262
rect 24974 17234 24998 17262
rect 25026 17234 25054 17262
rect 24554 16478 25054 17234
rect 24554 16450 24582 16478
rect 24610 16450 24634 16478
rect 24662 16450 24686 16478
rect 24714 16450 24738 16478
rect 24766 16450 24790 16478
rect 24818 16450 24842 16478
rect 24870 16450 24894 16478
rect 24922 16450 24946 16478
rect 24974 16450 24998 16478
rect 25026 16450 25054 16478
rect 24554 15694 25054 16450
rect 24554 15666 24582 15694
rect 24610 15666 24634 15694
rect 24662 15666 24686 15694
rect 24714 15666 24738 15694
rect 24766 15666 24790 15694
rect 24818 15666 24842 15694
rect 24870 15666 24894 15694
rect 24922 15666 24946 15694
rect 24974 15666 24998 15694
rect 25026 15666 25054 15694
rect 24554 14910 25054 15666
rect 24554 14882 24582 14910
rect 24610 14882 24634 14910
rect 24662 14882 24686 14910
rect 24714 14882 24738 14910
rect 24766 14882 24790 14910
rect 24818 14882 24842 14910
rect 24870 14882 24894 14910
rect 24922 14882 24946 14910
rect 24974 14882 24998 14910
rect 25026 14882 25054 14910
rect 24554 14126 25054 14882
rect 24554 14098 24582 14126
rect 24610 14098 24634 14126
rect 24662 14098 24686 14126
rect 24714 14098 24738 14126
rect 24766 14098 24790 14126
rect 24818 14098 24842 14126
rect 24870 14098 24894 14126
rect 24922 14098 24946 14126
rect 24974 14098 24998 14126
rect 25026 14098 25054 14126
rect 24554 13342 25054 14098
rect 24554 13314 24582 13342
rect 24610 13314 24634 13342
rect 24662 13314 24686 13342
rect 24714 13314 24738 13342
rect 24766 13314 24790 13342
rect 24818 13314 24842 13342
rect 24870 13314 24894 13342
rect 24922 13314 24946 13342
rect 24974 13314 24998 13342
rect 25026 13314 25054 13342
rect 24554 12558 25054 13314
rect 24554 12530 24582 12558
rect 24610 12530 24634 12558
rect 24662 12530 24686 12558
rect 24714 12530 24738 12558
rect 24766 12530 24790 12558
rect 24818 12530 24842 12558
rect 24870 12530 24894 12558
rect 24922 12530 24946 12558
rect 24974 12530 24998 12558
rect 25026 12530 25054 12558
rect 24554 11774 25054 12530
rect 24554 11746 24582 11774
rect 24610 11746 24634 11774
rect 24662 11746 24686 11774
rect 24714 11746 24738 11774
rect 24766 11746 24790 11774
rect 24818 11746 24842 11774
rect 24870 11746 24894 11774
rect 24922 11746 24946 11774
rect 24974 11746 24998 11774
rect 25026 11746 25054 11774
rect 24554 10990 25054 11746
rect 24554 10962 24582 10990
rect 24610 10962 24634 10990
rect 24662 10962 24686 10990
rect 24714 10962 24738 10990
rect 24766 10962 24790 10990
rect 24818 10962 24842 10990
rect 24870 10962 24894 10990
rect 24922 10962 24946 10990
rect 24974 10962 24998 10990
rect 25026 10962 25054 10990
rect 24554 10206 25054 10962
rect 24554 10178 24582 10206
rect 24610 10178 24634 10206
rect 24662 10178 24686 10206
rect 24714 10178 24738 10206
rect 24766 10178 24790 10206
rect 24818 10178 24842 10206
rect 24870 10178 24894 10206
rect 24922 10178 24946 10206
rect 24974 10178 24998 10206
rect 25026 10178 25054 10206
rect 24554 9422 25054 10178
rect 24554 9394 24582 9422
rect 24610 9394 24634 9422
rect 24662 9394 24686 9422
rect 24714 9394 24738 9422
rect 24766 9394 24790 9422
rect 24818 9394 24842 9422
rect 24870 9394 24894 9422
rect 24922 9394 24946 9422
rect 24974 9394 24998 9422
rect 25026 9394 25054 9422
rect 24554 8638 25054 9394
rect 24554 8610 24582 8638
rect 24610 8610 24634 8638
rect 24662 8610 24686 8638
rect 24714 8610 24738 8638
rect 24766 8610 24790 8638
rect 24818 8610 24842 8638
rect 24870 8610 24894 8638
rect 24922 8610 24946 8638
rect 24974 8610 24998 8638
rect 25026 8610 25054 8638
rect 24554 7854 25054 8610
rect 24554 7826 24582 7854
rect 24610 7826 24634 7854
rect 24662 7826 24686 7854
rect 24714 7826 24738 7854
rect 24766 7826 24790 7854
rect 24818 7826 24842 7854
rect 24870 7826 24894 7854
rect 24922 7826 24946 7854
rect 24974 7826 24998 7854
rect 25026 7826 25054 7854
rect 24554 7070 25054 7826
rect 24554 7042 24582 7070
rect 24610 7042 24634 7070
rect 24662 7042 24686 7070
rect 24714 7042 24738 7070
rect 24766 7042 24790 7070
rect 24818 7042 24842 7070
rect 24870 7042 24894 7070
rect 24922 7042 24946 7070
rect 24974 7042 24998 7070
rect 25026 7042 25054 7070
rect 24554 6286 25054 7042
rect 24554 6258 24582 6286
rect 24610 6258 24634 6286
rect 24662 6258 24686 6286
rect 24714 6258 24738 6286
rect 24766 6258 24790 6286
rect 24818 6258 24842 6286
rect 24870 6258 24894 6286
rect 24922 6258 24946 6286
rect 24974 6258 24998 6286
rect 25026 6258 25054 6286
rect 24554 5502 25054 6258
rect 24554 5474 24582 5502
rect 24610 5474 24634 5502
rect 24662 5474 24686 5502
rect 24714 5474 24738 5502
rect 24766 5474 24790 5502
rect 24818 5474 24842 5502
rect 24870 5474 24894 5502
rect 24922 5474 24946 5502
rect 24974 5474 24998 5502
rect 25026 5474 25054 5502
rect 24554 4718 25054 5474
rect 24554 4690 24582 4718
rect 24610 4690 24634 4718
rect 24662 4690 24686 4718
rect 24714 4690 24738 4718
rect 24766 4690 24790 4718
rect 24818 4690 24842 4718
rect 24870 4690 24894 4718
rect 24922 4690 24946 4718
rect 24974 4690 24998 4718
rect 25026 4690 25054 4718
rect 24554 3934 25054 4690
rect 24554 3906 24582 3934
rect 24610 3906 24634 3934
rect 24662 3906 24686 3934
rect 24714 3906 24738 3934
rect 24766 3906 24790 3934
rect 24818 3906 24842 3934
rect 24870 3906 24894 3934
rect 24922 3906 24946 3934
rect 24974 3906 24998 3934
rect 25026 3906 25054 3934
rect 24554 3150 25054 3906
rect 24554 3122 24582 3150
rect 24610 3122 24634 3150
rect 24662 3122 24686 3150
rect 24714 3122 24738 3150
rect 24766 3122 24790 3150
rect 24818 3122 24842 3150
rect 24870 3122 24894 3150
rect 24922 3122 24946 3150
rect 24974 3122 24998 3150
rect 25026 3122 25054 3150
rect 24554 2366 25054 3122
rect 24554 2338 24582 2366
rect 24610 2338 24634 2366
rect 24662 2338 24686 2366
rect 24714 2338 24738 2366
rect 24766 2338 24790 2366
rect 24818 2338 24842 2366
rect 24870 2338 24894 2366
rect 24922 2338 24946 2366
rect 24974 2338 24998 2366
rect 25026 2338 25054 2366
rect 24554 1582 25054 2338
rect 24554 1554 24582 1582
rect 24610 1554 24634 1582
rect 24662 1554 24686 1582
rect 24714 1554 24738 1582
rect 24766 1554 24790 1582
rect 24818 1554 24842 1582
rect 24870 1554 24894 1582
rect 24922 1554 24946 1582
rect 24974 1554 24998 1582
rect 25026 1554 25054 1582
rect 24554 1538 25054 1554
rect 27054 18438 27554 18454
rect 27054 18410 27082 18438
rect 27110 18410 27134 18438
rect 27162 18410 27186 18438
rect 27214 18410 27238 18438
rect 27266 18410 27290 18438
rect 27318 18410 27342 18438
rect 27370 18410 27394 18438
rect 27422 18410 27446 18438
rect 27474 18410 27498 18438
rect 27526 18410 27554 18438
rect 27054 17654 27554 18410
rect 27054 17626 27082 17654
rect 27110 17626 27134 17654
rect 27162 17626 27186 17654
rect 27214 17626 27238 17654
rect 27266 17626 27290 17654
rect 27318 17626 27342 17654
rect 27370 17626 27394 17654
rect 27422 17626 27446 17654
rect 27474 17626 27498 17654
rect 27526 17626 27554 17654
rect 27054 16870 27554 17626
rect 27054 16842 27082 16870
rect 27110 16842 27134 16870
rect 27162 16842 27186 16870
rect 27214 16842 27238 16870
rect 27266 16842 27290 16870
rect 27318 16842 27342 16870
rect 27370 16842 27394 16870
rect 27422 16842 27446 16870
rect 27474 16842 27498 16870
rect 27526 16842 27554 16870
rect 27054 16086 27554 16842
rect 27054 16058 27082 16086
rect 27110 16058 27134 16086
rect 27162 16058 27186 16086
rect 27214 16058 27238 16086
rect 27266 16058 27290 16086
rect 27318 16058 27342 16086
rect 27370 16058 27394 16086
rect 27422 16058 27446 16086
rect 27474 16058 27498 16086
rect 27526 16058 27554 16086
rect 27054 15302 27554 16058
rect 27054 15274 27082 15302
rect 27110 15274 27134 15302
rect 27162 15274 27186 15302
rect 27214 15274 27238 15302
rect 27266 15274 27290 15302
rect 27318 15274 27342 15302
rect 27370 15274 27394 15302
rect 27422 15274 27446 15302
rect 27474 15274 27498 15302
rect 27526 15274 27554 15302
rect 27054 14518 27554 15274
rect 27054 14490 27082 14518
rect 27110 14490 27134 14518
rect 27162 14490 27186 14518
rect 27214 14490 27238 14518
rect 27266 14490 27290 14518
rect 27318 14490 27342 14518
rect 27370 14490 27394 14518
rect 27422 14490 27446 14518
rect 27474 14490 27498 14518
rect 27526 14490 27554 14518
rect 27054 13734 27554 14490
rect 27054 13706 27082 13734
rect 27110 13706 27134 13734
rect 27162 13706 27186 13734
rect 27214 13706 27238 13734
rect 27266 13706 27290 13734
rect 27318 13706 27342 13734
rect 27370 13706 27394 13734
rect 27422 13706 27446 13734
rect 27474 13706 27498 13734
rect 27526 13706 27554 13734
rect 27054 12950 27554 13706
rect 27054 12922 27082 12950
rect 27110 12922 27134 12950
rect 27162 12922 27186 12950
rect 27214 12922 27238 12950
rect 27266 12922 27290 12950
rect 27318 12922 27342 12950
rect 27370 12922 27394 12950
rect 27422 12922 27446 12950
rect 27474 12922 27498 12950
rect 27526 12922 27554 12950
rect 27054 12166 27554 12922
rect 27054 12138 27082 12166
rect 27110 12138 27134 12166
rect 27162 12138 27186 12166
rect 27214 12138 27238 12166
rect 27266 12138 27290 12166
rect 27318 12138 27342 12166
rect 27370 12138 27394 12166
rect 27422 12138 27446 12166
rect 27474 12138 27498 12166
rect 27526 12138 27554 12166
rect 27054 11382 27554 12138
rect 27054 11354 27082 11382
rect 27110 11354 27134 11382
rect 27162 11354 27186 11382
rect 27214 11354 27238 11382
rect 27266 11354 27290 11382
rect 27318 11354 27342 11382
rect 27370 11354 27394 11382
rect 27422 11354 27446 11382
rect 27474 11354 27498 11382
rect 27526 11354 27554 11382
rect 27054 10598 27554 11354
rect 27054 10570 27082 10598
rect 27110 10570 27134 10598
rect 27162 10570 27186 10598
rect 27214 10570 27238 10598
rect 27266 10570 27290 10598
rect 27318 10570 27342 10598
rect 27370 10570 27394 10598
rect 27422 10570 27446 10598
rect 27474 10570 27498 10598
rect 27526 10570 27554 10598
rect 27054 9814 27554 10570
rect 27054 9786 27082 9814
rect 27110 9786 27134 9814
rect 27162 9786 27186 9814
rect 27214 9786 27238 9814
rect 27266 9786 27290 9814
rect 27318 9786 27342 9814
rect 27370 9786 27394 9814
rect 27422 9786 27446 9814
rect 27474 9786 27498 9814
rect 27526 9786 27554 9814
rect 27054 9030 27554 9786
rect 27054 9002 27082 9030
rect 27110 9002 27134 9030
rect 27162 9002 27186 9030
rect 27214 9002 27238 9030
rect 27266 9002 27290 9030
rect 27318 9002 27342 9030
rect 27370 9002 27394 9030
rect 27422 9002 27446 9030
rect 27474 9002 27498 9030
rect 27526 9002 27554 9030
rect 27054 8246 27554 9002
rect 27054 8218 27082 8246
rect 27110 8218 27134 8246
rect 27162 8218 27186 8246
rect 27214 8218 27238 8246
rect 27266 8218 27290 8246
rect 27318 8218 27342 8246
rect 27370 8218 27394 8246
rect 27422 8218 27446 8246
rect 27474 8218 27498 8246
rect 27526 8218 27554 8246
rect 27054 7462 27554 8218
rect 27054 7434 27082 7462
rect 27110 7434 27134 7462
rect 27162 7434 27186 7462
rect 27214 7434 27238 7462
rect 27266 7434 27290 7462
rect 27318 7434 27342 7462
rect 27370 7434 27394 7462
rect 27422 7434 27446 7462
rect 27474 7434 27498 7462
rect 27526 7434 27554 7462
rect 27054 6678 27554 7434
rect 27054 6650 27082 6678
rect 27110 6650 27134 6678
rect 27162 6650 27186 6678
rect 27214 6650 27238 6678
rect 27266 6650 27290 6678
rect 27318 6650 27342 6678
rect 27370 6650 27394 6678
rect 27422 6650 27446 6678
rect 27474 6650 27498 6678
rect 27526 6650 27554 6678
rect 27054 5894 27554 6650
rect 27054 5866 27082 5894
rect 27110 5866 27134 5894
rect 27162 5866 27186 5894
rect 27214 5866 27238 5894
rect 27266 5866 27290 5894
rect 27318 5866 27342 5894
rect 27370 5866 27394 5894
rect 27422 5866 27446 5894
rect 27474 5866 27498 5894
rect 27526 5866 27554 5894
rect 27054 5110 27554 5866
rect 27054 5082 27082 5110
rect 27110 5082 27134 5110
rect 27162 5082 27186 5110
rect 27214 5082 27238 5110
rect 27266 5082 27290 5110
rect 27318 5082 27342 5110
rect 27370 5082 27394 5110
rect 27422 5082 27446 5110
rect 27474 5082 27498 5110
rect 27526 5082 27554 5110
rect 27054 4326 27554 5082
rect 27054 4298 27082 4326
rect 27110 4298 27134 4326
rect 27162 4298 27186 4326
rect 27214 4298 27238 4326
rect 27266 4298 27290 4326
rect 27318 4298 27342 4326
rect 27370 4298 27394 4326
rect 27422 4298 27446 4326
rect 27474 4298 27498 4326
rect 27526 4298 27554 4326
rect 27054 3542 27554 4298
rect 27054 3514 27082 3542
rect 27110 3514 27134 3542
rect 27162 3514 27186 3542
rect 27214 3514 27238 3542
rect 27266 3514 27290 3542
rect 27318 3514 27342 3542
rect 27370 3514 27394 3542
rect 27422 3514 27446 3542
rect 27474 3514 27498 3542
rect 27526 3514 27554 3542
rect 27054 2758 27554 3514
rect 27054 2730 27082 2758
rect 27110 2730 27134 2758
rect 27162 2730 27186 2758
rect 27214 2730 27238 2758
rect 27266 2730 27290 2758
rect 27318 2730 27342 2758
rect 27370 2730 27394 2758
rect 27422 2730 27446 2758
rect 27474 2730 27498 2758
rect 27526 2730 27554 2758
rect 27054 1974 27554 2730
rect 27054 1946 27082 1974
rect 27110 1946 27134 1974
rect 27162 1946 27186 1974
rect 27214 1946 27238 1974
rect 27266 1946 27290 1974
rect 27318 1946 27342 1974
rect 27370 1946 27394 1974
rect 27422 1946 27446 1974
rect 27474 1946 27498 1974
rect 27526 1946 27554 1974
rect 27054 1538 27554 1946
rect 29554 18046 30054 18454
rect 29554 18018 29582 18046
rect 29610 18018 29634 18046
rect 29662 18018 29686 18046
rect 29714 18018 29738 18046
rect 29766 18018 29790 18046
rect 29818 18018 29842 18046
rect 29870 18018 29894 18046
rect 29922 18018 29946 18046
rect 29974 18018 29998 18046
rect 30026 18018 30054 18046
rect 29554 17262 30054 18018
rect 29554 17234 29582 17262
rect 29610 17234 29634 17262
rect 29662 17234 29686 17262
rect 29714 17234 29738 17262
rect 29766 17234 29790 17262
rect 29818 17234 29842 17262
rect 29870 17234 29894 17262
rect 29922 17234 29946 17262
rect 29974 17234 29998 17262
rect 30026 17234 30054 17262
rect 29554 16478 30054 17234
rect 29554 16450 29582 16478
rect 29610 16450 29634 16478
rect 29662 16450 29686 16478
rect 29714 16450 29738 16478
rect 29766 16450 29790 16478
rect 29818 16450 29842 16478
rect 29870 16450 29894 16478
rect 29922 16450 29946 16478
rect 29974 16450 29998 16478
rect 30026 16450 30054 16478
rect 29554 15694 30054 16450
rect 29554 15666 29582 15694
rect 29610 15666 29634 15694
rect 29662 15666 29686 15694
rect 29714 15666 29738 15694
rect 29766 15666 29790 15694
rect 29818 15666 29842 15694
rect 29870 15666 29894 15694
rect 29922 15666 29946 15694
rect 29974 15666 29998 15694
rect 30026 15666 30054 15694
rect 29554 14910 30054 15666
rect 29554 14882 29582 14910
rect 29610 14882 29634 14910
rect 29662 14882 29686 14910
rect 29714 14882 29738 14910
rect 29766 14882 29790 14910
rect 29818 14882 29842 14910
rect 29870 14882 29894 14910
rect 29922 14882 29946 14910
rect 29974 14882 29998 14910
rect 30026 14882 30054 14910
rect 29554 14126 30054 14882
rect 29554 14098 29582 14126
rect 29610 14098 29634 14126
rect 29662 14098 29686 14126
rect 29714 14098 29738 14126
rect 29766 14098 29790 14126
rect 29818 14098 29842 14126
rect 29870 14098 29894 14126
rect 29922 14098 29946 14126
rect 29974 14098 29998 14126
rect 30026 14098 30054 14126
rect 29554 13342 30054 14098
rect 29554 13314 29582 13342
rect 29610 13314 29634 13342
rect 29662 13314 29686 13342
rect 29714 13314 29738 13342
rect 29766 13314 29790 13342
rect 29818 13314 29842 13342
rect 29870 13314 29894 13342
rect 29922 13314 29946 13342
rect 29974 13314 29998 13342
rect 30026 13314 30054 13342
rect 29554 12558 30054 13314
rect 29554 12530 29582 12558
rect 29610 12530 29634 12558
rect 29662 12530 29686 12558
rect 29714 12530 29738 12558
rect 29766 12530 29790 12558
rect 29818 12530 29842 12558
rect 29870 12530 29894 12558
rect 29922 12530 29946 12558
rect 29974 12530 29998 12558
rect 30026 12530 30054 12558
rect 29554 11774 30054 12530
rect 29554 11746 29582 11774
rect 29610 11746 29634 11774
rect 29662 11746 29686 11774
rect 29714 11746 29738 11774
rect 29766 11746 29790 11774
rect 29818 11746 29842 11774
rect 29870 11746 29894 11774
rect 29922 11746 29946 11774
rect 29974 11746 29998 11774
rect 30026 11746 30054 11774
rect 29554 10990 30054 11746
rect 29554 10962 29582 10990
rect 29610 10962 29634 10990
rect 29662 10962 29686 10990
rect 29714 10962 29738 10990
rect 29766 10962 29790 10990
rect 29818 10962 29842 10990
rect 29870 10962 29894 10990
rect 29922 10962 29946 10990
rect 29974 10962 29998 10990
rect 30026 10962 30054 10990
rect 29554 10206 30054 10962
rect 29554 10178 29582 10206
rect 29610 10178 29634 10206
rect 29662 10178 29686 10206
rect 29714 10178 29738 10206
rect 29766 10178 29790 10206
rect 29818 10178 29842 10206
rect 29870 10178 29894 10206
rect 29922 10178 29946 10206
rect 29974 10178 29998 10206
rect 30026 10178 30054 10206
rect 29554 9422 30054 10178
rect 29554 9394 29582 9422
rect 29610 9394 29634 9422
rect 29662 9394 29686 9422
rect 29714 9394 29738 9422
rect 29766 9394 29790 9422
rect 29818 9394 29842 9422
rect 29870 9394 29894 9422
rect 29922 9394 29946 9422
rect 29974 9394 29998 9422
rect 30026 9394 30054 9422
rect 29554 8638 30054 9394
rect 29554 8610 29582 8638
rect 29610 8610 29634 8638
rect 29662 8610 29686 8638
rect 29714 8610 29738 8638
rect 29766 8610 29790 8638
rect 29818 8610 29842 8638
rect 29870 8610 29894 8638
rect 29922 8610 29946 8638
rect 29974 8610 29998 8638
rect 30026 8610 30054 8638
rect 29554 7854 30054 8610
rect 29554 7826 29582 7854
rect 29610 7826 29634 7854
rect 29662 7826 29686 7854
rect 29714 7826 29738 7854
rect 29766 7826 29790 7854
rect 29818 7826 29842 7854
rect 29870 7826 29894 7854
rect 29922 7826 29946 7854
rect 29974 7826 29998 7854
rect 30026 7826 30054 7854
rect 29554 7070 30054 7826
rect 29554 7042 29582 7070
rect 29610 7042 29634 7070
rect 29662 7042 29686 7070
rect 29714 7042 29738 7070
rect 29766 7042 29790 7070
rect 29818 7042 29842 7070
rect 29870 7042 29894 7070
rect 29922 7042 29946 7070
rect 29974 7042 29998 7070
rect 30026 7042 30054 7070
rect 29554 6286 30054 7042
rect 29554 6258 29582 6286
rect 29610 6258 29634 6286
rect 29662 6258 29686 6286
rect 29714 6258 29738 6286
rect 29766 6258 29790 6286
rect 29818 6258 29842 6286
rect 29870 6258 29894 6286
rect 29922 6258 29946 6286
rect 29974 6258 29998 6286
rect 30026 6258 30054 6286
rect 29554 5502 30054 6258
rect 29554 5474 29582 5502
rect 29610 5474 29634 5502
rect 29662 5474 29686 5502
rect 29714 5474 29738 5502
rect 29766 5474 29790 5502
rect 29818 5474 29842 5502
rect 29870 5474 29894 5502
rect 29922 5474 29946 5502
rect 29974 5474 29998 5502
rect 30026 5474 30054 5502
rect 29554 4718 30054 5474
rect 29554 4690 29582 4718
rect 29610 4690 29634 4718
rect 29662 4690 29686 4718
rect 29714 4690 29738 4718
rect 29766 4690 29790 4718
rect 29818 4690 29842 4718
rect 29870 4690 29894 4718
rect 29922 4690 29946 4718
rect 29974 4690 29998 4718
rect 30026 4690 30054 4718
rect 29554 3934 30054 4690
rect 32054 18438 32554 18454
rect 32054 18410 32082 18438
rect 32110 18410 32134 18438
rect 32162 18410 32186 18438
rect 32214 18410 32238 18438
rect 32266 18410 32290 18438
rect 32318 18410 32342 18438
rect 32370 18410 32394 18438
rect 32422 18410 32446 18438
rect 32474 18410 32498 18438
rect 32526 18410 32554 18438
rect 32054 17654 32554 18410
rect 32054 17626 32082 17654
rect 32110 17626 32134 17654
rect 32162 17626 32186 17654
rect 32214 17626 32238 17654
rect 32266 17626 32290 17654
rect 32318 17626 32342 17654
rect 32370 17626 32394 17654
rect 32422 17626 32446 17654
rect 32474 17626 32498 17654
rect 32526 17626 32554 17654
rect 32054 16870 32554 17626
rect 32054 16842 32082 16870
rect 32110 16842 32134 16870
rect 32162 16842 32186 16870
rect 32214 16842 32238 16870
rect 32266 16842 32290 16870
rect 32318 16842 32342 16870
rect 32370 16842 32394 16870
rect 32422 16842 32446 16870
rect 32474 16842 32498 16870
rect 32526 16842 32554 16870
rect 32054 16086 32554 16842
rect 32054 16058 32082 16086
rect 32110 16058 32134 16086
rect 32162 16058 32186 16086
rect 32214 16058 32238 16086
rect 32266 16058 32290 16086
rect 32318 16058 32342 16086
rect 32370 16058 32394 16086
rect 32422 16058 32446 16086
rect 32474 16058 32498 16086
rect 32526 16058 32554 16086
rect 32054 15302 32554 16058
rect 32054 15274 32082 15302
rect 32110 15274 32134 15302
rect 32162 15274 32186 15302
rect 32214 15274 32238 15302
rect 32266 15274 32290 15302
rect 32318 15274 32342 15302
rect 32370 15274 32394 15302
rect 32422 15274 32446 15302
rect 32474 15274 32498 15302
rect 32526 15274 32554 15302
rect 32054 14518 32554 15274
rect 32054 14490 32082 14518
rect 32110 14490 32134 14518
rect 32162 14490 32186 14518
rect 32214 14490 32238 14518
rect 32266 14490 32290 14518
rect 32318 14490 32342 14518
rect 32370 14490 32394 14518
rect 32422 14490 32446 14518
rect 32474 14490 32498 14518
rect 32526 14490 32554 14518
rect 32054 13734 32554 14490
rect 32054 13706 32082 13734
rect 32110 13706 32134 13734
rect 32162 13706 32186 13734
rect 32214 13706 32238 13734
rect 32266 13706 32290 13734
rect 32318 13706 32342 13734
rect 32370 13706 32394 13734
rect 32422 13706 32446 13734
rect 32474 13706 32498 13734
rect 32526 13706 32554 13734
rect 32054 12950 32554 13706
rect 32054 12922 32082 12950
rect 32110 12922 32134 12950
rect 32162 12922 32186 12950
rect 32214 12922 32238 12950
rect 32266 12922 32290 12950
rect 32318 12922 32342 12950
rect 32370 12922 32394 12950
rect 32422 12922 32446 12950
rect 32474 12922 32498 12950
rect 32526 12922 32554 12950
rect 32054 12166 32554 12922
rect 32054 12138 32082 12166
rect 32110 12138 32134 12166
rect 32162 12138 32186 12166
rect 32214 12138 32238 12166
rect 32266 12138 32290 12166
rect 32318 12138 32342 12166
rect 32370 12138 32394 12166
rect 32422 12138 32446 12166
rect 32474 12138 32498 12166
rect 32526 12138 32554 12166
rect 32054 11382 32554 12138
rect 32054 11354 32082 11382
rect 32110 11354 32134 11382
rect 32162 11354 32186 11382
rect 32214 11354 32238 11382
rect 32266 11354 32290 11382
rect 32318 11354 32342 11382
rect 32370 11354 32394 11382
rect 32422 11354 32446 11382
rect 32474 11354 32498 11382
rect 32526 11354 32554 11382
rect 32054 10598 32554 11354
rect 32054 10570 32082 10598
rect 32110 10570 32134 10598
rect 32162 10570 32186 10598
rect 32214 10570 32238 10598
rect 32266 10570 32290 10598
rect 32318 10570 32342 10598
rect 32370 10570 32394 10598
rect 32422 10570 32446 10598
rect 32474 10570 32498 10598
rect 32526 10570 32554 10598
rect 32054 9814 32554 10570
rect 32054 9786 32082 9814
rect 32110 9786 32134 9814
rect 32162 9786 32186 9814
rect 32214 9786 32238 9814
rect 32266 9786 32290 9814
rect 32318 9786 32342 9814
rect 32370 9786 32394 9814
rect 32422 9786 32446 9814
rect 32474 9786 32498 9814
rect 32526 9786 32554 9814
rect 32054 9030 32554 9786
rect 32054 9002 32082 9030
rect 32110 9002 32134 9030
rect 32162 9002 32186 9030
rect 32214 9002 32238 9030
rect 32266 9002 32290 9030
rect 32318 9002 32342 9030
rect 32370 9002 32394 9030
rect 32422 9002 32446 9030
rect 32474 9002 32498 9030
rect 32526 9002 32554 9030
rect 32054 8246 32554 9002
rect 32054 8218 32082 8246
rect 32110 8218 32134 8246
rect 32162 8218 32186 8246
rect 32214 8218 32238 8246
rect 32266 8218 32290 8246
rect 32318 8218 32342 8246
rect 32370 8218 32394 8246
rect 32422 8218 32446 8246
rect 32474 8218 32498 8246
rect 32526 8218 32554 8246
rect 32054 7462 32554 8218
rect 32054 7434 32082 7462
rect 32110 7434 32134 7462
rect 32162 7434 32186 7462
rect 32214 7434 32238 7462
rect 32266 7434 32290 7462
rect 32318 7434 32342 7462
rect 32370 7434 32394 7462
rect 32422 7434 32446 7462
rect 32474 7434 32498 7462
rect 32526 7434 32554 7462
rect 32054 6678 32554 7434
rect 32054 6650 32082 6678
rect 32110 6650 32134 6678
rect 32162 6650 32186 6678
rect 32214 6650 32238 6678
rect 32266 6650 32290 6678
rect 32318 6650 32342 6678
rect 32370 6650 32394 6678
rect 32422 6650 32446 6678
rect 32474 6650 32498 6678
rect 32526 6650 32554 6678
rect 32054 5894 32554 6650
rect 32054 5866 32082 5894
rect 32110 5866 32134 5894
rect 32162 5866 32186 5894
rect 32214 5866 32238 5894
rect 32266 5866 32290 5894
rect 32318 5866 32342 5894
rect 32370 5866 32394 5894
rect 32422 5866 32446 5894
rect 32474 5866 32498 5894
rect 32526 5866 32554 5894
rect 32054 5110 32554 5866
rect 32054 5082 32082 5110
rect 32110 5082 32134 5110
rect 32162 5082 32186 5110
rect 32214 5082 32238 5110
rect 32266 5082 32290 5110
rect 32318 5082 32342 5110
rect 32370 5082 32394 5110
rect 32422 5082 32446 5110
rect 32474 5082 32498 5110
rect 32526 5082 32554 5110
rect 29554 3906 29582 3934
rect 29610 3906 29634 3934
rect 29662 3906 29686 3934
rect 29714 3906 29738 3934
rect 29766 3906 29790 3934
rect 29818 3906 29842 3934
rect 29870 3906 29894 3934
rect 29922 3906 29946 3934
rect 29974 3906 29998 3934
rect 30026 3906 30054 3934
rect 29554 3150 30054 3906
rect 29554 3122 29582 3150
rect 29610 3122 29634 3150
rect 29662 3122 29686 3150
rect 29714 3122 29738 3150
rect 29766 3122 29790 3150
rect 29818 3122 29842 3150
rect 29870 3122 29894 3150
rect 29922 3122 29946 3150
rect 29974 3122 29998 3150
rect 30026 3122 30054 3150
rect 29554 2366 30054 3122
rect 29554 2338 29582 2366
rect 29610 2338 29634 2366
rect 29662 2338 29686 2366
rect 29714 2338 29738 2366
rect 29766 2338 29790 2366
rect 29818 2338 29842 2366
rect 29870 2338 29894 2366
rect 29922 2338 29946 2366
rect 29974 2338 29998 2366
rect 30026 2338 30054 2366
rect 29554 1582 30054 2338
rect 31990 4466 32018 4471
rect 31990 3738 32018 4438
rect 31990 3010 32018 3710
rect 31990 2226 32018 2982
rect 31990 2193 32018 2198
rect 32054 4326 32554 5082
rect 32054 4298 32082 4326
rect 32110 4298 32134 4326
rect 32162 4298 32186 4326
rect 32214 4298 32238 4326
rect 32266 4298 32290 4326
rect 32318 4298 32342 4326
rect 32370 4298 32394 4326
rect 32422 4298 32446 4326
rect 32474 4298 32498 4326
rect 32526 4298 32554 4326
rect 32054 3542 32554 4298
rect 32054 3514 32082 3542
rect 32110 3514 32134 3542
rect 32162 3514 32186 3542
rect 32214 3514 32238 3542
rect 32266 3514 32290 3542
rect 32318 3514 32342 3542
rect 32370 3514 32394 3542
rect 32422 3514 32446 3542
rect 32474 3514 32498 3542
rect 32526 3514 32554 3542
rect 32054 2758 32554 3514
rect 32054 2730 32082 2758
rect 32110 2730 32134 2758
rect 32162 2730 32186 2758
rect 32214 2730 32238 2758
rect 32266 2730 32290 2758
rect 32318 2730 32342 2758
rect 32370 2730 32394 2758
rect 32422 2730 32446 2758
rect 32474 2730 32498 2758
rect 32526 2730 32554 2758
rect 29554 1554 29582 1582
rect 29610 1554 29634 1582
rect 29662 1554 29686 1582
rect 29714 1554 29738 1582
rect 29766 1554 29790 1582
rect 29818 1554 29842 1582
rect 29870 1554 29894 1582
rect 29922 1554 29946 1582
rect 29974 1554 29998 1582
rect 30026 1554 30054 1582
rect 29554 1538 30054 1554
rect 32054 1974 32554 2730
rect 32054 1946 32082 1974
rect 32110 1946 32134 1974
rect 32162 1946 32186 1974
rect 32214 1946 32238 1974
rect 32266 1946 32290 1974
rect 32318 1946 32342 1974
rect 32370 1946 32394 1974
rect 32422 1946 32446 1974
rect 32474 1946 32498 1974
rect 32526 1946 32554 1974
rect 32054 1538 32554 1946
rect 34554 18046 35054 18454
rect 34554 18018 34582 18046
rect 34610 18018 34634 18046
rect 34662 18018 34686 18046
rect 34714 18018 34738 18046
rect 34766 18018 34790 18046
rect 34818 18018 34842 18046
rect 34870 18018 34894 18046
rect 34922 18018 34946 18046
rect 34974 18018 34998 18046
rect 35026 18018 35054 18046
rect 34554 17262 35054 18018
rect 34554 17234 34582 17262
rect 34610 17234 34634 17262
rect 34662 17234 34686 17262
rect 34714 17234 34738 17262
rect 34766 17234 34790 17262
rect 34818 17234 34842 17262
rect 34870 17234 34894 17262
rect 34922 17234 34946 17262
rect 34974 17234 34998 17262
rect 35026 17234 35054 17262
rect 34554 16478 35054 17234
rect 34554 16450 34582 16478
rect 34610 16450 34634 16478
rect 34662 16450 34686 16478
rect 34714 16450 34738 16478
rect 34766 16450 34790 16478
rect 34818 16450 34842 16478
rect 34870 16450 34894 16478
rect 34922 16450 34946 16478
rect 34974 16450 34998 16478
rect 35026 16450 35054 16478
rect 34554 15694 35054 16450
rect 34554 15666 34582 15694
rect 34610 15666 34634 15694
rect 34662 15666 34686 15694
rect 34714 15666 34738 15694
rect 34766 15666 34790 15694
rect 34818 15666 34842 15694
rect 34870 15666 34894 15694
rect 34922 15666 34946 15694
rect 34974 15666 34998 15694
rect 35026 15666 35054 15694
rect 34554 14910 35054 15666
rect 34554 14882 34582 14910
rect 34610 14882 34634 14910
rect 34662 14882 34686 14910
rect 34714 14882 34738 14910
rect 34766 14882 34790 14910
rect 34818 14882 34842 14910
rect 34870 14882 34894 14910
rect 34922 14882 34946 14910
rect 34974 14882 34998 14910
rect 35026 14882 35054 14910
rect 34554 14126 35054 14882
rect 34554 14098 34582 14126
rect 34610 14098 34634 14126
rect 34662 14098 34686 14126
rect 34714 14098 34738 14126
rect 34766 14098 34790 14126
rect 34818 14098 34842 14126
rect 34870 14098 34894 14126
rect 34922 14098 34946 14126
rect 34974 14098 34998 14126
rect 35026 14098 35054 14126
rect 34554 13342 35054 14098
rect 34554 13314 34582 13342
rect 34610 13314 34634 13342
rect 34662 13314 34686 13342
rect 34714 13314 34738 13342
rect 34766 13314 34790 13342
rect 34818 13314 34842 13342
rect 34870 13314 34894 13342
rect 34922 13314 34946 13342
rect 34974 13314 34998 13342
rect 35026 13314 35054 13342
rect 34554 12558 35054 13314
rect 34554 12530 34582 12558
rect 34610 12530 34634 12558
rect 34662 12530 34686 12558
rect 34714 12530 34738 12558
rect 34766 12530 34790 12558
rect 34818 12530 34842 12558
rect 34870 12530 34894 12558
rect 34922 12530 34946 12558
rect 34974 12530 34998 12558
rect 35026 12530 35054 12558
rect 34554 11774 35054 12530
rect 34554 11746 34582 11774
rect 34610 11746 34634 11774
rect 34662 11746 34686 11774
rect 34714 11746 34738 11774
rect 34766 11746 34790 11774
rect 34818 11746 34842 11774
rect 34870 11746 34894 11774
rect 34922 11746 34946 11774
rect 34974 11746 34998 11774
rect 35026 11746 35054 11774
rect 34554 10990 35054 11746
rect 34554 10962 34582 10990
rect 34610 10962 34634 10990
rect 34662 10962 34686 10990
rect 34714 10962 34738 10990
rect 34766 10962 34790 10990
rect 34818 10962 34842 10990
rect 34870 10962 34894 10990
rect 34922 10962 34946 10990
rect 34974 10962 34998 10990
rect 35026 10962 35054 10990
rect 34554 10206 35054 10962
rect 34554 10178 34582 10206
rect 34610 10178 34634 10206
rect 34662 10178 34686 10206
rect 34714 10178 34738 10206
rect 34766 10178 34790 10206
rect 34818 10178 34842 10206
rect 34870 10178 34894 10206
rect 34922 10178 34946 10206
rect 34974 10178 34998 10206
rect 35026 10178 35054 10206
rect 34554 9422 35054 10178
rect 34554 9394 34582 9422
rect 34610 9394 34634 9422
rect 34662 9394 34686 9422
rect 34714 9394 34738 9422
rect 34766 9394 34790 9422
rect 34818 9394 34842 9422
rect 34870 9394 34894 9422
rect 34922 9394 34946 9422
rect 34974 9394 34998 9422
rect 35026 9394 35054 9422
rect 34554 8638 35054 9394
rect 34554 8610 34582 8638
rect 34610 8610 34634 8638
rect 34662 8610 34686 8638
rect 34714 8610 34738 8638
rect 34766 8610 34790 8638
rect 34818 8610 34842 8638
rect 34870 8610 34894 8638
rect 34922 8610 34946 8638
rect 34974 8610 34998 8638
rect 35026 8610 35054 8638
rect 34554 7854 35054 8610
rect 34554 7826 34582 7854
rect 34610 7826 34634 7854
rect 34662 7826 34686 7854
rect 34714 7826 34738 7854
rect 34766 7826 34790 7854
rect 34818 7826 34842 7854
rect 34870 7826 34894 7854
rect 34922 7826 34946 7854
rect 34974 7826 34998 7854
rect 35026 7826 35054 7854
rect 34554 7070 35054 7826
rect 34554 7042 34582 7070
rect 34610 7042 34634 7070
rect 34662 7042 34686 7070
rect 34714 7042 34738 7070
rect 34766 7042 34790 7070
rect 34818 7042 34842 7070
rect 34870 7042 34894 7070
rect 34922 7042 34946 7070
rect 34974 7042 34998 7070
rect 35026 7042 35054 7070
rect 34554 6286 35054 7042
rect 34554 6258 34582 6286
rect 34610 6258 34634 6286
rect 34662 6258 34686 6286
rect 34714 6258 34738 6286
rect 34766 6258 34790 6286
rect 34818 6258 34842 6286
rect 34870 6258 34894 6286
rect 34922 6258 34946 6286
rect 34974 6258 34998 6286
rect 35026 6258 35054 6286
rect 34554 5502 35054 6258
rect 34554 5474 34582 5502
rect 34610 5474 34634 5502
rect 34662 5474 34686 5502
rect 34714 5474 34738 5502
rect 34766 5474 34790 5502
rect 34818 5474 34842 5502
rect 34870 5474 34894 5502
rect 34922 5474 34946 5502
rect 34974 5474 34998 5502
rect 35026 5474 35054 5502
rect 34554 4718 35054 5474
rect 34554 4690 34582 4718
rect 34610 4690 34634 4718
rect 34662 4690 34686 4718
rect 34714 4690 34738 4718
rect 34766 4690 34790 4718
rect 34818 4690 34842 4718
rect 34870 4690 34894 4718
rect 34922 4690 34946 4718
rect 34974 4690 34998 4718
rect 35026 4690 35054 4718
rect 34554 3934 35054 4690
rect 37054 18438 37554 18454
rect 37054 18410 37082 18438
rect 37110 18410 37134 18438
rect 37162 18410 37186 18438
rect 37214 18410 37238 18438
rect 37266 18410 37290 18438
rect 37318 18410 37342 18438
rect 37370 18410 37394 18438
rect 37422 18410 37446 18438
rect 37474 18410 37498 18438
rect 37526 18410 37554 18438
rect 37054 17654 37554 18410
rect 37054 17626 37082 17654
rect 37110 17626 37134 17654
rect 37162 17626 37186 17654
rect 37214 17626 37238 17654
rect 37266 17626 37290 17654
rect 37318 17626 37342 17654
rect 37370 17626 37394 17654
rect 37422 17626 37446 17654
rect 37474 17626 37498 17654
rect 37526 17626 37554 17654
rect 37054 16870 37554 17626
rect 37054 16842 37082 16870
rect 37110 16842 37134 16870
rect 37162 16842 37186 16870
rect 37214 16842 37238 16870
rect 37266 16842 37290 16870
rect 37318 16842 37342 16870
rect 37370 16842 37394 16870
rect 37422 16842 37446 16870
rect 37474 16842 37498 16870
rect 37526 16842 37554 16870
rect 37054 16086 37554 16842
rect 37054 16058 37082 16086
rect 37110 16058 37134 16086
rect 37162 16058 37186 16086
rect 37214 16058 37238 16086
rect 37266 16058 37290 16086
rect 37318 16058 37342 16086
rect 37370 16058 37394 16086
rect 37422 16058 37446 16086
rect 37474 16058 37498 16086
rect 37526 16058 37554 16086
rect 37054 15302 37554 16058
rect 37054 15274 37082 15302
rect 37110 15274 37134 15302
rect 37162 15274 37186 15302
rect 37214 15274 37238 15302
rect 37266 15274 37290 15302
rect 37318 15274 37342 15302
rect 37370 15274 37394 15302
rect 37422 15274 37446 15302
rect 37474 15274 37498 15302
rect 37526 15274 37554 15302
rect 37054 14518 37554 15274
rect 37054 14490 37082 14518
rect 37110 14490 37134 14518
rect 37162 14490 37186 14518
rect 37214 14490 37238 14518
rect 37266 14490 37290 14518
rect 37318 14490 37342 14518
rect 37370 14490 37394 14518
rect 37422 14490 37446 14518
rect 37474 14490 37498 14518
rect 37526 14490 37554 14518
rect 37054 13734 37554 14490
rect 37054 13706 37082 13734
rect 37110 13706 37134 13734
rect 37162 13706 37186 13734
rect 37214 13706 37238 13734
rect 37266 13706 37290 13734
rect 37318 13706 37342 13734
rect 37370 13706 37394 13734
rect 37422 13706 37446 13734
rect 37474 13706 37498 13734
rect 37526 13706 37554 13734
rect 37054 12950 37554 13706
rect 37054 12922 37082 12950
rect 37110 12922 37134 12950
rect 37162 12922 37186 12950
rect 37214 12922 37238 12950
rect 37266 12922 37290 12950
rect 37318 12922 37342 12950
rect 37370 12922 37394 12950
rect 37422 12922 37446 12950
rect 37474 12922 37498 12950
rect 37526 12922 37554 12950
rect 37054 12166 37554 12922
rect 37054 12138 37082 12166
rect 37110 12138 37134 12166
rect 37162 12138 37186 12166
rect 37214 12138 37238 12166
rect 37266 12138 37290 12166
rect 37318 12138 37342 12166
rect 37370 12138 37394 12166
rect 37422 12138 37446 12166
rect 37474 12138 37498 12166
rect 37526 12138 37554 12166
rect 37054 11382 37554 12138
rect 37054 11354 37082 11382
rect 37110 11354 37134 11382
rect 37162 11354 37186 11382
rect 37214 11354 37238 11382
rect 37266 11354 37290 11382
rect 37318 11354 37342 11382
rect 37370 11354 37394 11382
rect 37422 11354 37446 11382
rect 37474 11354 37498 11382
rect 37526 11354 37554 11382
rect 37054 10598 37554 11354
rect 37054 10570 37082 10598
rect 37110 10570 37134 10598
rect 37162 10570 37186 10598
rect 37214 10570 37238 10598
rect 37266 10570 37290 10598
rect 37318 10570 37342 10598
rect 37370 10570 37394 10598
rect 37422 10570 37446 10598
rect 37474 10570 37498 10598
rect 37526 10570 37554 10598
rect 37054 9814 37554 10570
rect 37054 9786 37082 9814
rect 37110 9786 37134 9814
rect 37162 9786 37186 9814
rect 37214 9786 37238 9814
rect 37266 9786 37290 9814
rect 37318 9786 37342 9814
rect 37370 9786 37394 9814
rect 37422 9786 37446 9814
rect 37474 9786 37498 9814
rect 37526 9786 37554 9814
rect 37054 9030 37554 9786
rect 37054 9002 37082 9030
rect 37110 9002 37134 9030
rect 37162 9002 37186 9030
rect 37214 9002 37238 9030
rect 37266 9002 37290 9030
rect 37318 9002 37342 9030
rect 37370 9002 37394 9030
rect 37422 9002 37446 9030
rect 37474 9002 37498 9030
rect 37526 9002 37554 9030
rect 37054 8246 37554 9002
rect 37054 8218 37082 8246
rect 37110 8218 37134 8246
rect 37162 8218 37186 8246
rect 37214 8218 37238 8246
rect 37266 8218 37290 8246
rect 37318 8218 37342 8246
rect 37370 8218 37394 8246
rect 37422 8218 37446 8246
rect 37474 8218 37498 8246
rect 37526 8218 37554 8246
rect 37054 7462 37554 8218
rect 37054 7434 37082 7462
rect 37110 7434 37134 7462
rect 37162 7434 37186 7462
rect 37214 7434 37238 7462
rect 37266 7434 37290 7462
rect 37318 7434 37342 7462
rect 37370 7434 37394 7462
rect 37422 7434 37446 7462
rect 37474 7434 37498 7462
rect 37526 7434 37554 7462
rect 37054 6678 37554 7434
rect 37054 6650 37082 6678
rect 37110 6650 37134 6678
rect 37162 6650 37186 6678
rect 37214 6650 37238 6678
rect 37266 6650 37290 6678
rect 37318 6650 37342 6678
rect 37370 6650 37394 6678
rect 37422 6650 37446 6678
rect 37474 6650 37498 6678
rect 37526 6650 37554 6678
rect 37054 5894 37554 6650
rect 37054 5866 37082 5894
rect 37110 5866 37134 5894
rect 37162 5866 37186 5894
rect 37214 5866 37238 5894
rect 37266 5866 37290 5894
rect 37318 5866 37342 5894
rect 37370 5866 37394 5894
rect 37422 5866 37446 5894
rect 37474 5866 37498 5894
rect 37526 5866 37554 5894
rect 37054 5110 37554 5866
rect 37054 5082 37082 5110
rect 37110 5082 37134 5110
rect 37162 5082 37186 5110
rect 37214 5082 37238 5110
rect 37266 5082 37290 5110
rect 37318 5082 37342 5110
rect 37370 5082 37394 5110
rect 37422 5082 37446 5110
rect 37474 5082 37498 5110
rect 37526 5082 37554 5110
rect 37054 4326 37554 5082
rect 37054 4298 37082 4326
rect 37110 4298 37134 4326
rect 37162 4298 37186 4326
rect 37214 4298 37238 4326
rect 37266 4298 37290 4326
rect 37318 4298 37342 4326
rect 37370 4298 37394 4326
rect 37422 4298 37446 4326
rect 37474 4298 37498 4326
rect 37526 4298 37554 4326
rect 34554 3906 34582 3934
rect 34610 3906 34634 3934
rect 34662 3906 34686 3934
rect 34714 3906 34738 3934
rect 34766 3906 34790 3934
rect 34818 3906 34842 3934
rect 34870 3906 34894 3934
rect 34922 3906 34946 3934
rect 34974 3906 34998 3934
rect 35026 3906 35054 3934
rect 34554 3150 35054 3906
rect 36918 4186 36946 4191
rect 36918 3402 36946 4158
rect 36918 3369 36946 3374
rect 37054 3542 37554 4298
rect 37054 3514 37082 3542
rect 37110 3514 37134 3542
rect 37162 3514 37186 3542
rect 37214 3514 37238 3542
rect 37266 3514 37290 3542
rect 37318 3514 37342 3542
rect 37370 3514 37394 3542
rect 37422 3514 37446 3542
rect 37474 3514 37498 3542
rect 37526 3514 37554 3542
rect 34554 3122 34582 3150
rect 34610 3122 34634 3150
rect 34662 3122 34686 3150
rect 34714 3122 34738 3150
rect 34766 3122 34790 3150
rect 34818 3122 34842 3150
rect 34870 3122 34894 3150
rect 34922 3122 34946 3150
rect 34974 3122 34998 3150
rect 35026 3122 35054 3150
rect 34554 2366 35054 3122
rect 34554 2338 34582 2366
rect 34610 2338 34634 2366
rect 34662 2338 34686 2366
rect 34714 2338 34738 2366
rect 34766 2338 34790 2366
rect 34818 2338 34842 2366
rect 34870 2338 34894 2366
rect 34922 2338 34946 2366
rect 34974 2338 34998 2366
rect 35026 2338 35054 2366
rect 34554 1582 35054 2338
rect 34554 1554 34582 1582
rect 34610 1554 34634 1582
rect 34662 1554 34686 1582
rect 34714 1554 34738 1582
rect 34766 1554 34790 1582
rect 34818 1554 34842 1582
rect 34870 1554 34894 1582
rect 34922 1554 34946 1582
rect 34974 1554 34998 1582
rect 35026 1554 35054 1582
rect 34554 1538 35054 1554
rect 37054 2758 37554 3514
rect 37054 2730 37082 2758
rect 37110 2730 37134 2758
rect 37162 2730 37186 2758
rect 37214 2730 37238 2758
rect 37266 2730 37290 2758
rect 37318 2730 37342 2758
rect 37370 2730 37394 2758
rect 37422 2730 37446 2758
rect 37474 2730 37498 2758
rect 37526 2730 37554 2758
rect 37054 1974 37554 2730
rect 37054 1946 37082 1974
rect 37110 1946 37134 1974
rect 37162 1946 37186 1974
rect 37214 1946 37238 1974
rect 37266 1946 37290 1974
rect 37318 1946 37342 1974
rect 37370 1946 37394 1974
rect 37422 1946 37446 1974
rect 37474 1946 37498 1974
rect 37526 1946 37554 1974
rect 37054 1538 37554 1946
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2184 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 4536 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1667941163
transform 1 0 6664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 8456 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142
timestamp 1667941163
transform 1 0 8624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 10416 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_177
timestamp 1667941163
transform 1 0 10584 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1667941163
transform 1 0 12376 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_212
timestamp 1667941163
transform 1 0 12544 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1667941163
transform 1 0 14336 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_247
timestamp 1667941163
transform 1 0 14504 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 16296 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_282
timestamp 1667941163
transform 1 0 16464 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1667941163
transform 1 0 18256 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1667941163
transform 1 0 18424 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_342
timestamp 1667941163
transform 1 0 19824 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1667941163
transform 1 0 20384 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_377
timestamp 1667941163
transform 1 0 21784 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1667941163
transform 1 0 22344 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_412
timestamp 1667941163
transform 1 0 23744 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1667941163
transform 1 0 24304 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_447
timestamp 1667941163
transform 1 0 25704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1667941163
transform 1 0 26264 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_482
timestamp 1667941163
transform 1 0 27664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1667941163
transform 1 0 28224 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_517
timestamp 1667941163
transform 1 0 29624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1667941163
transform 1 0 30184 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_552
timestamp 1667941163
transform 1 0 31584 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1667941163
transform 1 0 32144 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_587
timestamp 1667941163
transform 1 0 33544 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1667941163
transform 1 0 34104 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_622
timestamp 1667941163
transform 1 0 35504 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1667941163
transform 1 0 36064 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_657
timestamp 1667941163
transform 1 0 37464 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1667941163
transform 1 0 38024 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_676 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 38528 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_686
timestamp 1667941163
transform 1 0 39088 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_18
timestamp 1667941163
transform 1 0 1680 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_44
timestamp 1667941163
transform 1 0 3136 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_89
timestamp 1667941163
transform 1 0 5656 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_115
timestamp 1667941163
transform 1 0 7112 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 8568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_144
timestamp 1667941163
transform 1 0 8736 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_160
timestamp 1667941163
transform 1 0 9632 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_186
timestamp 1667941163
transform 1 0 11088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 12544 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_215
timestamp 1667941163
transform 1 0 12712 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_231
timestamp 1667941163
transform 1 0 13608 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_257
timestamp 1667941163
transform 1 0 15064 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1667941163
transform 1 0 16520 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_286 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 16688 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_290
timestamp 1667941163
transform 1 0 16912 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_316
timestamp 1667941163
transform 1 0 18368 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_342
timestamp 1667941163
transform 1 0 19824 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1667941163
transform 1 0 20272 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1667941163
transform 1 0 20496 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1667941163
transform 1 0 20664 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_382
timestamp 1667941163
transform 1 0 22064 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_408
timestamp 1667941163
transform 1 0 23520 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_424
timestamp 1667941163
transform 1 0 24416 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1667941163
transform 1 0 24640 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_453
timestamp 1667941163
transform 1 0 26040 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_479
timestamp 1667941163
transform 1 0 27496 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_487
timestamp 1667941163
transform 1 0 27944 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1667941163
transform 1 0 28448 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1667941163
transform 1 0 28616 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_524
timestamp 1667941163
transform 1 0 30016 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_550
timestamp 1667941163
transform 1 0 31472 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_558
timestamp 1667941163
transform 1 0 31920 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1667941163
transform 1 0 32424 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1667941163
transform 1 0 32592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_595
timestamp 1667941163
transform 1 0 33992 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_621
timestamp 1667941163
transform 1 0 35448 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_631
timestamp 1667941163
transform 1 0 36008 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1667941163
transform 1 0 36568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_666
timestamp 1667941163
transform 1 0 37968 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_676
timestamp 1667941163
transform 1 0 38528 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_686
timestamp 1667941163
transform 1 0 39088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_53
timestamp 1667941163
transform 1 0 3640 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_79
timestamp 1667941163
transform 1 0 5096 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_108
timestamp 1667941163
transform 1 0 6720 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_124
timestamp 1667941163
transform 1 0 7616 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_150
timestamp 1667941163
transform 1 0 9072 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 10528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_179
timestamp 1667941163
transform 1 0 10696 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_195
timestamp 1667941163
transform 1 0 11592 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_203
timestamp 1667941163
transform 1 0 12040 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_229
timestamp 1667941163
transform 1 0 13496 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_245
timestamp 1667941163
transform 1 0 14392 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1667941163
transform 1 0 14504 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_250
timestamp 1667941163
transform 1 0 14672 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_290
timestamp 1667941163
transform 1 0 16912 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_316
timestamp 1667941163
transform 1 0 18368 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1667941163
transform 1 0 18480 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1667941163
transform 1 0 18648 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_346
timestamp 1667941163
transform 1 0 20048 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_372
timestamp 1667941163
transform 1 0 21504 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_388
timestamp 1667941163
transform 1 0 22400 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1667941163
transform 1 0 22624 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_417
timestamp 1667941163
transform 1 0 24024 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_443
timestamp 1667941163
transform 1 0 25480 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_459
timestamp 1667941163
transform 1 0 26376 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1667941163
transform 1 0 26600 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_488
timestamp 1667941163
transform 1 0 28000 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_514
timestamp 1667941163
transform 1 0 29456 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_522
timestamp 1667941163
transform 1 0 29904 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1667941163
transform 1 0 30408 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1667941163
transform 1 0 30576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_559
timestamp 1667941163
transform 1 0 31976 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_585
timestamp 1667941163
transform 1 0 33432 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_595
timestamp 1667941163
transform 1 0 33992 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1667941163
transform 1 0 34552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_630
timestamp 1667941163
transform 1 0 35952 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_656
timestamp 1667941163
transform 1 0 37408 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_666
timestamp 1667941163
transform 1 0 37968 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_676
timestamp 1667941163
transform 1 0 38528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_685
timestamp 1667941163
transform 1 0 39032 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_687
timestamp 1667941163
transform 1 0 39144 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_18
timestamp 1667941163
transform 1 0 1680 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_44
timestamp 1667941163
transform 1 0 3136 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_89
timestamp 1667941163
transform 1 0 5656 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_115
timestamp 1667941163
transform 1 0 7112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 8568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_144
timestamp 1667941163
transform 1 0 8736 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_160
timestamp 1667941163
transform 1 0 9632 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_186
timestamp 1667941163
transform 1 0 11088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1667941163
transform 1 0 12544 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_215
timestamp 1667941163
transform 1 0 12712 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_231
timestamp 1667941163
transform 1 0 13608 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_257
timestamp 1667941163
transform 1 0 15064 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1667941163
transform 1 0 16520 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_286
timestamp 1667941163
transform 1 0 16688 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_294
timestamp 1667941163
transform 1 0 17136 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_296
timestamp 1667941163
transform 1 0 17248 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_321
timestamp 1667941163
transform 1 0 18648 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_347
timestamp 1667941163
transform 1 0 20104 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1667941163
transform 1 0 20664 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_382
timestamp 1667941163
transform 1 0 22064 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_408
timestamp 1667941163
transform 1 0 23520 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_424
timestamp 1667941163
transform 1 0 24416 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1667941163
transform 1 0 24640 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_453
timestamp 1667941163
transform 1 0 26040 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_479
timestamp 1667941163
transform 1 0 27496 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_487
timestamp 1667941163
transform 1 0 27944 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1667941163
transform 1 0 28448 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1667941163
transform 1 0 28616 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_524
timestamp 1667941163
transform 1 0 30016 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_550
timestamp 1667941163
transform 1 0 31472 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_558
timestamp 1667941163
transform 1 0 31920 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1667941163
transform 1 0 32424 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1667941163
transform 1 0 32592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_595
timestamp 1667941163
transform 1 0 33992 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_621
timestamp 1667941163
transform 1 0 35448 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_631
timestamp 1667941163
transform 1 0 36008 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_641
timestamp 1667941163
transform 1 0 36568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_666
timestamp 1667941163
transform 1 0 37968 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_676
timestamp 1667941163
transform 1 0 38528 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_686
timestamp 1667941163
transform 1 0 39088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_53
timestamp 1667941163
transform 1 0 3640 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_79
timestamp 1667941163
transform 1 0 5096 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_108
timestamp 1667941163
transform 1 0 6720 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_124
timestamp 1667941163
transform 1 0 7616 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_150
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 10528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_179
timestamp 1667941163
transform 1 0 10696 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_195
timestamp 1667941163
transform 1 0 11592 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_221
timestamp 1667941163
transform 1 0 13048 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1667941163
transform 1 0 14504 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_250
timestamp 1667941163
transform 1 0 14672 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_266
timestamp 1667941163
transform 1 0 15568 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_292
timestamp 1667941163
transform 1 0 17024 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1667941163
transform 1 0 18480 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1667941163
transform 1 0 18648 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_346
timestamp 1667941163
transform 1 0 20048 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_372
timestamp 1667941163
transform 1 0 21504 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_388
timestamp 1667941163
transform 1 0 22400 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1667941163
transform 1 0 22624 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_417
timestamp 1667941163
transform 1 0 24024 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_443
timestamp 1667941163
transform 1 0 25480 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_459
timestamp 1667941163
transform 1 0 26376 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1667941163
transform 1 0 26600 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_488
timestamp 1667941163
transform 1 0 28000 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_514
timestamp 1667941163
transform 1 0 29456 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_522
timestamp 1667941163
transform 1 0 29904 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1667941163
transform 1 0 30408 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_534
timestamp 1667941163
transform 1 0 30576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_559
timestamp 1667941163
transform 1 0 31976 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_585
timestamp 1667941163
transform 1 0 33432 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_595
timestamp 1667941163
transform 1 0 33992 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1667941163
transform 1 0 34552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_630
timestamp 1667941163
transform 1 0 35952 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_656
timestamp 1667941163
transform 1 0 37408 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_666
timestamp 1667941163
transform 1 0 37968 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1667941163
transform 1 0 38528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_685
timestamp 1667941163
transform 1 0 39032 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_687
timestamp 1667941163
transform 1 0 39144 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_18
timestamp 1667941163
transform 1 0 1680 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_44
timestamp 1667941163
transform 1 0 3136 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_89
timestamp 1667941163
transform 1 0 5656 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_115
timestamp 1667941163
transform 1 0 7112 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 8568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_144
timestamp 1667941163
transform 1 0 8736 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_160
timestamp 1667941163
transform 1 0 9632 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_186
timestamp 1667941163
transform 1 0 11088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1667941163
transform 1 0 12544 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_215
timestamp 1667941163
transform 1 0 12712 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_231
timestamp 1667941163
transform 1 0 13608 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_257
timestamp 1667941163
transform 1 0 15064 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1667941163
transform 1 0 16520 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_286
timestamp 1667941163
transform 1 0 16688 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_294
timestamp 1667941163
transform 1 0 17136 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_296
timestamp 1667941163
transform 1 0 17248 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_321
timestamp 1667941163
transform 1 0 18648 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_347
timestamp 1667941163
transform 1 0 20104 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1667941163
transform 1 0 20664 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_382
timestamp 1667941163
transform 1 0 22064 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_408
timestamp 1667941163
transform 1 0 23520 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_424
timestamp 1667941163
transform 1 0 24416 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1667941163
transform 1 0 24640 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_453
timestamp 1667941163
transform 1 0 26040 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_479
timestamp 1667941163
transform 1 0 27496 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_487
timestamp 1667941163
transform 1 0 27944 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1667941163
transform 1 0 28448 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_499
timestamp 1667941163
transform 1 0 28616 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_524
timestamp 1667941163
transform 1 0 30016 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_550
timestamp 1667941163
transform 1 0 31472 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_558
timestamp 1667941163
transform 1 0 31920 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1667941163
transform 1 0 32424 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1667941163
transform 1 0 32592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_595
timestamp 1667941163
transform 1 0 33992 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_621
timestamp 1667941163
transform 1 0 35448 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_631
timestamp 1667941163
transform 1 0 36008 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_641
timestamp 1667941163
transform 1 0 36568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_666
timestamp 1667941163
transform 1 0 37968 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_676
timestamp 1667941163
transform 1 0 38528 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_686
timestamp 1667941163
transform 1 0 39088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_53
timestamp 1667941163
transform 1 0 3640 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_79
timestamp 1667941163
transform 1 0 5096 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 6552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_108
timestamp 1667941163
transform 1 0 6720 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_124
timestamp 1667941163
transform 1 0 7616 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_150
timestamp 1667941163
transform 1 0 9072 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 10528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_179
timestamp 1667941163
transform 1 0 10696 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_195
timestamp 1667941163
transform 1 0 11592 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_221
timestamp 1667941163
transform 1 0 13048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1667941163
transform 1 0 14504 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_250
timestamp 1667941163
transform 1 0 14672 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_266
timestamp 1667941163
transform 1 0 15568 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_292
timestamp 1667941163
transform 1 0 17024 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1667941163
transform 1 0 18480 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1667941163
transform 1 0 18648 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_346
timestamp 1667941163
transform 1 0 20048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_372
timestamp 1667941163
transform 1 0 21504 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_388
timestamp 1667941163
transform 1 0 22400 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_392
timestamp 1667941163
transform 1 0 22624 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_417
timestamp 1667941163
transform 1 0 24024 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_443
timestamp 1667941163
transform 1 0 25480 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_459
timestamp 1667941163
transform 1 0 26376 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1667941163
transform 1 0 26600 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_488
timestamp 1667941163
transform 1 0 28000 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_514
timestamp 1667941163
transform 1 0 29456 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_522
timestamp 1667941163
transform 1 0 29904 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1667941163
transform 1 0 30408 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_534
timestamp 1667941163
transform 1 0 30576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_559
timestamp 1667941163
transform 1 0 31976 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_585
timestamp 1667941163
transform 1 0 33432 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_595
timestamp 1667941163
transform 1 0 33992 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_605
timestamp 1667941163
transform 1 0 34552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_630
timestamp 1667941163
transform 1 0 35952 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_656
timestamp 1667941163
transform 1 0 37408 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_666
timestamp 1667941163
transform 1 0 37968 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_676
timestamp 1667941163
transform 1 0 38528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_685
timestamp 1667941163
transform 1 0 39032 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_687
timestamp 1667941163
transform 1 0 39144 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_2
timestamp 1667941163
transform 1 0 784 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_18
timestamp 1667941163
transform 1 0 1680 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_44
timestamp 1667941163
transform 1 0 3136 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 4592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1667941163
transform 1 0 4760 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_89
timestamp 1667941163
transform 1 0 5656 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_115
timestamp 1667941163
transform 1 0 7112 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 8568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_144
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1667941163
transform 1 0 9632 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_186
timestamp 1667941163
transform 1 0 11088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1667941163
transform 1 0 12544 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_215
timestamp 1667941163
transform 1 0 12712 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_231
timestamp 1667941163
transform 1 0 13608 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_257
timestamp 1667941163
transform 1 0 15064 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1667941163
transform 1 0 16520 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_286
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_294
timestamp 1667941163
transform 1 0 17136 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_296
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_321
timestamp 1667941163
transform 1 0 18648 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_347
timestamp 1667941163
transform 1 0 20104 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_357
timestamp 1667941163
transform 1 0 20664 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_382
timestamp 1667941163
transform 1 0 22064 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_408
timestamp 1667941163
transform 1 0 23520 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_424
timestamp 1667941163
transform 1 0 24416 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1667941163
transform 1 0 24640 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_453
timestamp 1667941163
transform 1 0 26040 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_479
timestamp 1667941163
transform 1 0 27496 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_487
timestamp 1667941163
transform 1 0 27944 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1667941163
transform 1 0 28448 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_499
timestamp 1667941163
transform 1 0 28616 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_524
timestamp 1667941163
transform 1 0 30016 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_550
timestamp 1667941163
transform 1 0 31472 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_558
timestamp 1667941163
transform 1 0 31920 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1667941163
transform 1 0 32424 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_570
timestamp 1667941163
transform 1 0 32592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_595
timestamp 1667941163
transform 1 0 33992 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_621
timestamp 1667941163
transform 1 0 35448 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_631
timestamp 1667941163
transform 1 0 36008 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_641
timestamp 1667941163
transform 1 0 36568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_666
timestamp 1667941163
transform 1 0 37968 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_676
timestamp 1667941163
transform 1 0 38528 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_686
timestamp 1667941163
transform 1 0 39088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_2
timestamp 1667941163
transform 1 0 784 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1667941163
transform 1 0 2744 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_53
timestamp 1667941163
transform 1 0 3640 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_79
timestamp 1667941163
transform 1 0 5096 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 6552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_108
timestamp 1667941163
transform 1 0 6720 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_124
timestamp 1667941163
transform 1 0 7616 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_150
timestamp 1667941163
transform 1 0 9072 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 10528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_179
timestamp 1667941163
transform 1 0 10696 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_195
timestamp 1667941163
transform 1 0 11592 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_199
timestamp 1667941163
transform 1 0 11816 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_201
timestamp 1667941163
transform 1 0 11928 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_226
timestamp 1667941163
transform 1 0 13328 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_242
timestamp 1667941163
transform 1 0 14224 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_246
timestamp 1667941163
transform 1 0 14448 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_250
timestamp 1667941163
transform 1 0 14672 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_266
timestamp 1667941163
transform 1 0 15568 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_292
timestamp 1667941163
transform 1 0 17024 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1667941163
transform 1 0 18480 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1667941163
transform 1 0 18648 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_346
timestamp 1667941163
transform 1 0 20048 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_372
timestamp 1667941163
transform 1 0 21504 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_388
timestamp 1667941163
transform 1 0 22400 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1667941163
transform 1 0 22624 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_417
timestamp 1667941163
transform 1 0 24024 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_443
timestamp 1667941163
transform 1 0 25480 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_459
timestamp 1667941163
transform 1 0 26376 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_463
timestamp 1667941163
transform 1 0 26600 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_488
timestamp 1667941163
transform 1 0 28000 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_514
timestamp 1667941163
transform 1 0 29456 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_522
timestamp 1667941163
transform 1 0 29904 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1667941163
transform 1 0 30408 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_534
timestamp 1667941163
transform 1 0 30576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_559
timestamp 1667941163
transform 1 0 31976 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_585
timestamp 1667941163
transform 1 0 33432 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_595
timestamp 1667941163
transform 1 0 33992 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_605
timestamp 1667941163
transform 1 0 34552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_630
timestamp 1667941163
transform 1 0 35952 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_656
timestamp 1667941163
transform 1 0 37408 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_666
timestamp 1667941163
transform 1 0 37968 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_676
timestamp 1667941163
transform 1 0 38528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_685
timestamp 1667941163
transform 1 0 39032 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_687
timestamp 1667941163
transform 1 0 39144 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_2
timestamp 1667941163
transform 1 0 784 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_18
timestamp 1667941163
transform 1 0 1680 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_44
timestamp 1667941163
transform 1 0 3136 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 4592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_73
timestamp 1667941163
transform 1 0 4760 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_89
timestamp 1667941163
transform 1 0 5656 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_115
timestamp 1667941163
transform 1 0 7112 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 8568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_144
timestamp 1667941163
transform 1 0 8736 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_160
timestamp 1667941163
transform 1 0 9632 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_186
timestamp 1667941163
transform 1 0 11088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1667941163
transform 1 0 12544 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1667941163
transform 1 0 12712 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_240
timestamp 1667941163
transform 1 0 14112 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_256
timestamp 1667941163
transform 1 0 15008 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_258
timestamp 1667941163
transform 1 0 15120 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1667941163
transform 1 0 16520 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_286
timestamp 1667941163
transform 1 0 16688 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_294
timestamp 1667941163
transform 1 0 17136 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_296
timestamp 1667941163
transform 1 0 17248 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_321
timestamp 1667941163
transform 1 0 18648 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_347
timestamp 1667941163
transform 1 0 20104 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1667941163
transform 1 0 20664 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_382
timestamp 1667941163
transform 1 0 22064 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_408
timestamp 1667941163
transform 1 0 23520 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_424
timestamp 1667941163
transform 1 0 24416 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_428
timestamp 1667941163
transform 1 0 24640 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_453
timestamp 1667941163
transform 1 0 26040 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_479
timestamp 1667941163
transform 1 0 27496 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_495
timestamp 1667941163
transform 1 0 28392 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_499
timestamp 1667941163
transform 1 0 28616 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_507
timestamp 1667941163
transform 1 0 29064 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_532
timestamp 1667941163
transform 1 0 30464 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_558
timestamp 1667941163
transform 1 0 31920 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_566
timestamp 1667941163
transform 1 0 32368 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_570
timestamp 1667941163
transform 1 0 32592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_595
timestamp 1667941163
transform 1 0 33992 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_621
timestamp 1667941163
transform 1 0 35448 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_631
timestamp 1667941163
transform 1 0 36008 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_641
timestamp 1667941163
transform 1 0 36568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_666
timestamp 1667941163
transform 1 0 37968 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_682
timestamp 1667941163
transform 1 0 38864 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_686
timestamp 1667941163
transform 1 0 39088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1667941163
transform 1 0 784 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 2576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1667941163
transform 1 0 2744 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1667941163
transform 1 0 3640 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_79
timestamp 1667941163
transform 1 0 5096 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 6552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_108
timestamp 1667941163
transform 1 0 6720 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_124
timestamp 1667941163
transform 1 0 7616 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_150
timestamp 1667941163
transform 1 0 9072 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 10528 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_179
timestamp 1667941163
transform 1 0 10696 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_195
timestamp 1667941163
transform 1 0 11592 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_199
timestamp 1667941163
transform 1 0 11816 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_201
timestamp 1667941163
transform 1 0 11928 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_226
timestamp 1667941163
transform 1 0 13328 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_242
timestamp 1667941163
transform 1 0 14224 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_246
timestamp 1667941163
transform 1 0 14448 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_250
timestamp 1667941163
transform 1 0 14672 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_266
timestamp 1667941163
transform 1 0 15568 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_292
timestamp 1667941163
transform 1 0 17024 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1667941163
transform 1 0 18480 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1667941163
transform 1 0 18648 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_346
timestamp 1667941163
transform 1 0 20048 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_372
timestamp 1667941163
transform 1 0 21504 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_388
timestamp 1667941163
transform 1 0 22400 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_392
timestamp 1667941163
transform 1 0 22624 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_417
timestamp 1667941163
transform 1 0 24024 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_443
timestamp 1667941163
transform 1 0 25480 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_459
timestamp 1667941163
transform 1 0 26376 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1667941163
transform 1 0 26600 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_488
timestamp 1667941163
transform 1 0 28000 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_504
timestamp 1667941163
transform 1 0 28896 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_506
timestamp 1667941163
transform 1 0 29008 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1667941163
transform 1 0 30408 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_534
timestamp 1667941163
transform 1 0 30576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_559
timestamp 1667941163
transform 1 0 31976 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_585
timestamp 1667941163
transform 1 0 33432 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_595
timestamp 1667941163
transform 1 0 33992 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_605
timestamp 1667941163
transform 1 0 34552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_630
timestamp 1667941163
transform 1 0 35952 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_656
timestamp 1667941163
transform 1 0 37408 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_666
timestamp 1667941163
transform 1 0 37968 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_676
timestamp 1667941163
transform 1 0 38528 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_684
timestamp 1667941163
transform 1 0 38976 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1667941163
transform 1 0 784 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_18
timestamp 1667941163
transform 1 0 1680 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_44
timestamp 1667941163
transform 1 0 3136 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 4592 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_73
timestamp 1667941163
transform 1 0 4760 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_89
timestamp 1667941163
transform 1 0 5656 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_115
timestamp 1667941163
transform 1 0 7112 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 8568 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_144
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_160
timestamp 1667941163
transform 1 0 9632 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_186
timestamp 1667941163
transform 1 0 11088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1667941163
transform 1 0 12544 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1667941163
transform 1 0 12712 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_240
timestamp 1667941163
transform 1 0 14112 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_256
timestamp 1667941163
transform 1 0 15008 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_258
timestamp 1667941163
transform 1 0 15120 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1667941163
transform 1 0 16520 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_286
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_294
timestamp 1667941163
transform 1 0 17136 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_296
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_321
timestamp 1667941163
transform 1 0 18648 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_347
timestamp 1667941163
transform 1 0 20104 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1667941163
transform 1 0 20664 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_382
timestamp 1667941163
transform 1 0 22064 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_408
timestamp 1667941163
transform 1 0 23520 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_424
timestamp 1667941163
transform 1 0 24416 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1667941163
transform 1 0 24640 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_453
timestamp 1667941163
transform 1 0 26040 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_479
timestamp 1667941163
transform 1 0 27496 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_495
timestamp 1667941163
transform 1 0 28392 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_499
timestamp 1667941163
transform 1 0 28616 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_507
timestamp 1667941163
transform 1 0 29064 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_532
timestamp 1667941163
transform 1 0 30464 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_558
timestamp 1667941163
transform 1 0 31920 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_566
timestamp 1667941163
transform 1 0 32368 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_570
timestamp 1667941163
transform 1 0 32592 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_595
timestamp 1667941163
transform 1 0 33992 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_621
timestamp 1667941163
transform 1 0 35448 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_631
timestamp 1667941163
transform 1 0 36008 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_641
timestamp 1667941163
transform 1 0 36568 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_666
timestamp 1667941163
transform 1 0 37968 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_682
timestamp 1667941163
transform 1 0 38864 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_686
timestamp 1667941163
transform 1 0 39088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_2
timestamp 1667941163
transform 1 0 784 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 2576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_37
timestamp 1667941163
transform 1 0 2744 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_53
timestamp 1667941163
transform 1 0 3640 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_79
timestamp 1667941163
transform 1 0 5096 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 6552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_108
timestamp 1667941163
transform 1 0 6720 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_124
timestamp 1667941163
transform 1 0 7616 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_150
timestamp 1667941163
transform 1 0 9072 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 10528 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_179
timestamp 1667941163
transform 1 0 10696 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_187
timestamp 1667941163
transform 1 0 11144 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_191
timestamp 1667941163
transform 1 0 11368 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_216
timestamp 1667941163
transform 1 0 12768 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_242
timestamp 1667941163
transform 1 0 14224 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_246
timestamp 1667941163
transform 1 0 14448 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_250
timestamp 1667941163
transform 1 0 14672 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_266
timestamp 1667941163
transform 1 0 15568 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_292
timestamp 1667941163
transform 1 0 17024 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1667941163
transform 1 0 18480 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1667941163
transform 1 0 18648 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_346
timestamp 1667941163
transform 1 0 20048 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_372
timestamp 1667941163
transform 1 0 21504 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_388
timestamp 1667941163
transform 1 0 22400 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1667941163
transform 1 0 22624 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_417
timestamp 1667941163
transform 1 0 24024 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_443
timestamp 1667941163
transform 1 0 25480 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_459
timestamp 1667941163
transform 1 0 26376 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_463
timestamp 1667941163
transform 1 0 26600 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_479
timestamp 1667941163
transform 1 0 27496 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_505
timestamp 1667941163
transform 1 0 28952 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1667941163
transform 1 0 30408 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_534
timestamp 1667941163
transform 1 0 30576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_559
timestamp 1667941163
transform 1 0 31976 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_585
timestamp 1667941163
transform 1 0 33432 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_595
timestamp 1667941163
transform 1 0 33992 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_605
timestamp 1667941163
transform 1 0 34552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_630
timestamp 1667941163
transform 1 0 35952 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_656
timestamp 1667941163
transform 1 0 37408 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_672
timestamp 1667941163
transform 1 0 38304 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_676
timestamp 1667941163
transform 1 0 38528 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_684
timestamp 1667941163
transform 1 0 38976 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1667941163
transform 1 0 784 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_18
timestamp 1667941163
transform 1 0 1680 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_44
timestamp 1667941163
transform 1 0 3136 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 4592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_73
timestamp 1667941163
transform 1 0 4760 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_89
timestamp 1667941163
transform 1 0 5656 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_115
timestamp 1667941163
transform 1 0 7112 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 8568 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_144
timestamp 1667941163
transform 1 0 8736 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_184
timestamp 1667941163
transform 1 0 10976 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_210
timestamp 1667941163
transform 1 0 12432 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 12544 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1667941163
transform 1 0 12712 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_240
timestamp 1667941163
transform 1 0 14112 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_266
timestamp 1667941163
transform 1 0 15568 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_282
timestamp 1667941163
transform 1 0 16464 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_286
timestamp 1667941163
transform 1 0 16688 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_294
timestamp 1667941163
transform 1 0 17136 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_296
timestamp 1667941163
transform 1 0 17248 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_321
timestamp 1667941163
transform 1 0 18648 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_347
timestamp 1667941163
transform 1 0 20104 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_357
timestamp 1667941163
transform 1 0 20664 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_382
timestamp 1667941163
transform 1 0 22064 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_408
timestamp 1667941163
transform 1 0 23520 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_424
timestamp 1667941163
transform 1 0 24416 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1667941163
transform 1 0 24640 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_453
timestamp 1667941163
transform 1 0 26040 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_469
timestamp 1667941163
transform 1 0 26936 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_471
timestamp 1667941163
transform 1 0 27048 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1667941163
transform 1 0 28448 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_499
timestamp 1667941163
transform 1 0 28616 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_507
timestamp 1667941163
transform 1 0 29064 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_532
timestamp 1667941163
transform 1 0 30464 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_558
timestamp 1667941163
transform 1 0 31920 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_566
timestamp 1667941163
transform 1 0 32368 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_570
timestamp 1667941163
transform 1 0 32592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_595
timestamp 1667941163
transform 1 0 33992 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_621
timestamp 1667941163
transform 1 0 35448 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_631
timestamp 1667941163
transform 1 0 36008 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_641
timestamp 1667941163
transform 1 0 36568 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_666
timestamp 1667941163
transform 1 0 37968 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_682
timestamp 1667941163
transform 1 0 38864 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_686
timestamp 1667941163
transform 1 0 39088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1667941163
transform 1 0 784 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 2576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_37
timestamp 1667941163
transform 1 0 2744 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_53
timestamp 1667941163
transform 1 0 3640 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_79
timestamp 1667941163
transform 1 0 5096 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 6552 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_108
timestamp 1667941163
transform 1 0 6720 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_124
timestamp 1667941163
transform 1 0 7616 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_150
timestamp 1667941163
transform 1 0 9072 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1667941163
transform 1 0 10528 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_179
timestamp 1667941163
transform 1 0 10696 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_211
timestamp 1667941163
transform 1 0 12488 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_237
timestamp 1667941163
transform 1 0 13944 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_245
timestamp 1667941163
transform 1 0 14392 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1667941163
transform 1 0 14504 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1667941163
transform 1 0 14672 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_275
timestamp 1667941163
transform 1 0 16072 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_291
timestamp 1667941163
transform 1 0 16968 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_293
timestamp 1667941163
transform 1 0 17080 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1667941163
transform 1 0 18480 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1667941163
transform 1 0 18648 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_346
timestamp 1667941163
transform 1 0 20048 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_372
timestamp 1667941163
transform 1 0 21504 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_388
timestamp 1667941163
transform 1 0 22400 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_392
timestamp 1667941163
transform 1 0 22624 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_417
timestamp 1667941163
transform 1 0 24024 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_443
timestamp 1667941163
transform 1 0 25480 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_459
timestamp 1667941163
transform 1 0 26376 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_463
timestamp 1667941163
transform 1 0 26600 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_479
timestamp 1667941163
transform 1 0 27496 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_505
timestamp 1667941163
transform 1 0 28952 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1667941163
transform 1 0 30408 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_534
timestamp 1667941163
transform 1 0 30576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_559
timestamp 1667941163
transform 1 0 31976 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_585
timestamp 1667941163
transform 1 0 33432 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_595
timestamp 1667941163
transform 1 0 33992 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_605
timestamp 1667941163
transform 1 0 34552 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_630
timestamp 1667941163
transform 1 0 35952 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_656
timestamp 1667941163
transform 1 0 37408 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_672
timestamp 1667941163
transform 1 0 38304 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_676
timestamp 1667941163
transform 1 0 38528 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_684
timestamp 1667941163
transform 1 0 38976 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_2
timestamp 1667941163
transform 1 0 784 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_18
timestamp 1667941163
transform 1 0 1680 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_44
timestamp 1667941163
transform 1 0 3136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 4592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_73
timestamp 1667941163
transform 1 0 4760 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_89
timestamp 1667941163
transform 1 0 5656 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_115
timestamp 1667941163
transform 1 0 7112 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 8568 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_144
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_160
timestamp 1667941163
transform 1 0 9632 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_185
timestamp 1667941163
transform 1 0 11032 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_211
timestamp 1667941163
transform 1 0 12488 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_215
timestamp 1667941163
transform 1 0 12712 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_240
timestamp 1667941163
transform 1 0 14112 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_266
timestamp 1667941163
transform 1 0 15568 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_282
timestamp 1667941163
transform 1 0 16464 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_286
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_294
timestamp 1667941163
transform 1 0 17136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_296
timestamp 1667941163
transform 1 0 17248 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_321
timestamp 1667941163
transform 1 0 18648 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_347
timestamp 1667941163
transform 1 0 20104 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_357
timestamp 1667941163
transform 1 0 20664 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_382
timestamp 1667941163
transform 1 0 22064 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_408
timestamp 1667941163
transform 1 0 23520 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_424
timestamp 1667941163
transform 1 0 24416 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_428
timestamp 1667941163
transform 1 0 24640 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_453
timestamp 1667941163
transform 1 0 26040 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_479
timestamp 1667941163
transform 1 0 27496 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_495
timestamp 1667941163
transform 1 0 28392 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_499
timestamp 1667941163
transform 1 0 28616 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_507
timestamp 1667941163
transform 1 0 29064 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_532
timestamp 1667941163
transform 1 0 30464 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_558
timestamp 1667941163
transform 1 0 31920 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_566
timestamp 1667941163
transform 1 0 32368 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_570
timestamp 1667941163
transform 1 0 32592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_595
timestamp 1667941163
transform 1 0 33992 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_621
timestamp 1667941163
transform 1 0 35448 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_637
timestamp 1667941163
transform 1 0 36344 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_641
timestamp 1667941163
transform 1 0 36568 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_666
timestamp 1667941163
transform 1 0 37968 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_682
timestamp 1667941163
transform 1 0 38864 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_686
timestamp 1667941163
transform 1 0 39088 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_2
timestamp 1667941163
transform 1 0 784 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1667941163
transform 1 0 2576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_37
timestamp 1667941163
transform 1 0 2744 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_53
timestamp 1667941163
transform 1 0 3640 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_79
timestamp 1667941163
transform 1 0 5096 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1667941163
transform 1 0 6552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_108
timestamp 1667941163
transform 1 0 6720 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_124
timestamp 1667941163
transform 1 0 7616 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_150
timestamp 1667941163
transform 1 0 9072 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1667941163
transform 1 0 10528 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_179
timestamp 1667941163
transform 1 0 10696 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_211
timestamp 1667941163
transform 1 0 12488 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_215
timestamp 1667941163
transform 1 0 12712 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_241
timestamp 1667941163
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_245
timestamp 1667941163
transform 1 0 14392 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1667941163
transform 1 0 14504 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1667941163
transform 1 0 14672 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_275
timestamp 1667941163
transform 1 0 16072 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_301
timestamp 1667941163
transform 1 0 17528 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_317
timestamp 1667941163
transform 1 0 18424 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_321
timestamp 1667941163
transform 1 0 18648 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_346
timestamp 1667941163
transform 1 0 20048 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_372
timestamp 1667941163
transform 1 0 21504 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_388
timestamp 1667941163
transform 1 0 22400 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_392
timestamp 1667941163
transform 1 0 22624 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_417
timestamp 1667941163
transform 1 0 24024 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_443
timestamp 1667941163
transform 1 0 25480 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_459
timestamp 1667941163
transform 1 0 26376 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_463
timestamp 1667941163
transform 1 0 26600 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_488
timestamp 1667941163
transform 1 0 28000 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_504
timestamp 1667941163
transform 1 0 28896 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_506
timestamp 1667941163
transform 1 0 29008 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1667941163
transform 1 0 30408 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_534
timestamp 1667941163
transform 1 0 30576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_559
timestamp 1667941163
transform 1 0 31976 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_585
timestamp 1667941163
transform 1 0 33432 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_595
timestamp 1667941163
transform 1 0 33992 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_605
timestamp 1667941163
transform 1 0 34552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_630
timestamp 1667941163
transform 1 0 35952 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_656
timestamp 1667941163
transform 1 0 37408 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_672
timestamp 1667941163
transform 1 0 38304 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_676
timestamp 1667941163
transform 1 0 38528 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_684
timestamp 1667941163
transform 1 0 38976 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_2
timestamp 1667941163
transform 1 0 784 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_18
timestamp 1667941163
transform 1 0 1680 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_44
timestamp 1667941163
transform 1 0 3136 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1667941163
transform 1 0 4592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_73
timestamp 1667941163
transform 1 0 4760 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_89
timestamp 1667941163
transform 1 0 5656 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_115
timestamp 1667941163
transform 1 0 7112 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1667941163
transform 1 0 8568 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_144
timestamp 1667941163
transform 1 0 8736 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_160
timestamp 1667941163
transform 1 0 9632 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_186
timestamp 1667941163
transform 1 0 11088 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1667941163
transform 1 0 12544 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_215
timestamp 1667941163
transform 1 0 12712 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_243
timestamp 1667941163
transform 1 0 14280 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_269
timestamp 1667941163
transform 1 0 15736 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_277
timestamp 1667941163
transform 1 0 16184 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 16408 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1667941163
transform 1 0 16520 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1667941163
transform 1 0 16688 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_311
timestamp 1667941163
transform 1 0 18088 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_337
timestamp 1667941163
transform 1 0 19544 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_353
timestamp 1667941163
transform 1 0 20440 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_357
timestamp 1667941163
transform 1 0 20664 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_382
timestamp 1667941163
transform 1 0 22064 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_408
timestamp 1667941163
transform 1 0 23520 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_424
timestamp 1667941163
transform 1 0 24416 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_428
timestamp 1667941163
transform 1 0 24640 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_453
timestamp 1667941163
transform 1 0 26040 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_479
timestamp 1667941163
transform 1 0 27496 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_495
timestamp 1667941163
transform 1 0 28392 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_499
timestamp 1667941163
transform 1 0 28616 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_507
timestamp 1667941163
transform 1 0 29064 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_509
timestamp 1667941163
transform 1 0 29176 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_534
timestamp 1667941163
transform 1 0 30576 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_560
timestamp 1667941163
transform 1 0 32032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_570
timestamp 1667941163
transform 1 0 32592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_595
timestamp 1667941163
transform 1 0 33992 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_621
timestamp 1667941163
transform 1 0 35448 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_637
timestamp 1667941163
transform 1 0 36344 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_641
timestamp 1667941163
transform 1 0 36568 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_666
timestamp 1667941163
transform 1 0 37968 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_682
timestamp 1667941163
transform 1 0 38864 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_686
timestamp 1667941163
transform 1 0 39088 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_2
timestamp 1667941163
transform 1 0 784 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1667941163
transform 1 0 2576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_37
timestamp 1667941163
transform 1 0 2744 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_53
timestamp 1667941163
transform 1 0 3640 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_79
timestamp 1667941163
transform 1 0 5096 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1667941163
transform 1 0 6552 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_108
timestamp 1667941163
transform 1 0 6720 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_124
timestamp 1667941163
transform 1 0 7616 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_150
timestamp 1667941163
transform 1 0 9072 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1667941163
transform 1 0 10528 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_179
timestamp 1667941163
transform 1 0 10696 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_187
timestamp 1667941163
transform 1 0 11144 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_191
timestamp 1667941163
transform 1 0 11368 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_193
timestamp 1667941163
transform 1 0 11480 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_218
timestamp 1667941163
transform 1 0 12880 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_244
timestamp 1667941163
transform 1 0 14336 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1667941163
transform 1 0 14672 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_275
timestamp 1667941163
transform 1 0 16072 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_301
timestamp 1667941163
transform 1 0 17528 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_317
timestamp 1667941163
transform 1 0 18424 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1667941163
transform 1 0 18648 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_346
timestamp 1667941163
transform 1 0 20048 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_372
timestamp 1667941163
transform 1 0 21504 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_388
timestamp 1667941163
transform 1 0 22400 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_392
timestamp 1667941163
transform 1 0 22624 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_417
timestamp 1667941163
transform 1 0 24024 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_443
timestamp 1667941163
transform 1 0 25480 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_459
timestamp 1667941163
transform 1 0 26376 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_463
timestamp 1667941163
transform 1 0 26600 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_479
timestamp 1667941163
transform 1 0 27496 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_505
timestamp 1667941163
transform 1 0 28952 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1667941163
transform 1 0 30408 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_534
timestamp 1667941163
transform 1 0 30576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_559
timestamp 1667941163
transform 1 0 31976 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_585
timestamp 1667941163
transform 1 0 33432 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_601
timestamp 1667941163
transform 1 0 34328 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_605
timestamp 1667941163
transform 1 0 34552 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_630
timestamp 1667941163
transform 1 0 35952 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_656
timestamp 1667941163
transform 1 0 37408 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_672
timestamp 1667941163
transform 1 0 38304 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_676
timestamp 1667941163
transform 1 0 38528 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_684
timestamp 1667941163
transform 1 0 38976 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_2
timestamp 1667941163
transform 1 0 784 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_18
timestamp 1667941163
transform 1 0 1680 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_44
timestamp 1667941163
transform 1 0 3136 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1667941163
transform 1 0 4592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_73
timestamp 1667941163
transform 1 0 4760 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_89
timestamp 1667941163
transform 1 0 5656 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_115
timestamp 1667941163
transform 1 0 7112 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1667941163
transform 1 0 8568 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_144
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_160
timestamp 1667941163
transform 1 0 9632 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_186
timestamp 1667941163
transform 1 0 11088 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1667941163
transform 1 0 12544 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_215
timestamp 1667941163
transform 1 0 12712 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_223
timestamp 1667941163
transform 1 0 13160 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_249
timestamp 1667941163
transform 1 0 14616 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_275
timestamp 1667941163
transform 1 0 16072 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1667941163
transform 1 0 16520 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_286
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_311
timestamp 1667941163
transform 1 0 18088 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_337
timestamp 1667941163
transform 1 0 19544 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_353
timestamp 1667941163
transform 1 0 20440 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_357
timestamp 1667941163
transform 1 0 20664 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_382
timestamp 1667941163
transform 1 0 22064 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_408
timestamp 1667941163
transform 1 0 23520 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_424
timestamp 1667941163
transform 1 0 24416 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1667941163
transform 1 0 24640 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_453
timestamp 1667941163
transform 1 0 26040 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_461
timestamp 1667941163
transform 1 0 26488 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_489
timestamp 1667941163
transform 1 0 28056 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_499
timestamp 1667941163
transform 1 0 28616 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_507
timestamp 1667941163
transform 1 0 29064 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_533
timestamp 1667941163
transform 1 0 30520 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_559
timestamp 1667941163
transform 1 0 31976 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1667941163
transform 1 0 32424 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_570
timestamp 1667941163
transform 1 0 32592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_595
timestamp 1667941163
transform 1 0 33992 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_621
timestamp 1667941163
transform 1 0 35448 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_637
timestamp 1667941163
transform 1 0 36344 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_641
timestamp 1667941163
transform 1 0 36568 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_666
timestamp 1667941163
transform 1 0 37968 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_682
timestamp 1667941163
transform 1 0 38864 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_686
timestamp 1667941163
transform 1 0 39088 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_2
timestamp 1667941163
transform 1 0 784 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1667941163
transform 1 0 2576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_37
timestamp 1667941163
transform 1 0 2744 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_53
timestamp 1667941163
transform 1 0 3640 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_79
timestamp 1667941163
transform 1 0 5096 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1667941163
transform 1 0 6552 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_108
timestamp 1667941163
transform 1 0 6720 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_124
timestamp 1667941163
transform 1 0 7616 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_150
timestamp 1667941163
transform 1 0 9072 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1667941163
transform 1 0 10528 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_179
timestamp 1667941163
transform 1 0 10696 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_187
timestamp 1667941163
transform 1 0 11144 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_191
timestamp 1667941163
transform 1 0 11368 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_193
timestamp 1667941163
transform 1 0 11480 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_218
timestamp 1667941163
transform 1 0 12880 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_244
timestamp 1667941163
transform 1 0 14336 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_250
timestamp 1667941163
transform 1 0 14672 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_275
timestamp 1667941163
transform 1 0 16072 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_301
timestamp 1667941163
transform 1 0 17528 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_317
timestamp 1667941163
transform 1 0 18424 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_321
timestamp 1667941163
transform 1 0 18648 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_346
timestamp 1667941163
transform 1 0 20048 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_372
timestamp 1667941163
transform 1 0 21504 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_388
timestamp 1667941163
transform 1 0 22400 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_392
timestamp 1667941163
transform 1 0 22624 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_417
timestamp 1667941163
transform 1 0 24024 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_443
timestamp 1667941163
transform 1 0 25480 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_459
timestamp 1667941163
transform 1 0 26376 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_463
timestamp 1667941163
transform 1 0 26600 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_479
timestamp 1667941163
transform 1 0 27496 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_505
timestamp 1667941163
transform 1 0 28952 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1667941163
transform 1 0 30408 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_534
timestamp 1667941163
transform 1 0 30576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_559
timestamp 1667941163
transform 1 0 31976 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_585
timestamp 1667941163
transform 1 0 33432 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_601
timestamp 1667941163
transform 1 0 34328 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_605
timestamp 1667941163
transform 1 0 34552 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_630
timestamp 1667941163
transform 1 0 35952 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_656
timestamp 1667941163
transform 1 0 37408 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_672
timestamp 1667941163
transform 1 0 38304 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_676
timestamp 1667941163
transform 1 0 38528 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_684
timestamp 1667941163
transform 1 0 38976 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_2
timestamp 1667941163
transform 1 0 784 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_18
timestamp 1667941163
transform 1 0 1680 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_44
timestamp 1667941163
transform 1 0 3136 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1667941163
transform 1 0 4592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_73
timestamp 1667941163
transform 1 0 4760 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_89
timestamp 1667941163
transform 1 0 5656 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_115
timestamp 1667941163
transform 1 0 7112 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1667941163
transform 1 0 8568 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_144
timestamp 1667941163
transform 1 0 8736 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_160
timestamp 1667941163
transform 1 0 9632 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_186
timestamp 1667941163
transform 1 0 11088 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1667941163
transform 1 0 12544 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_215
timestamp 1667941163
transform 1 0 12712 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_223
timestamp 1667941163
transform 1 0 13160 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_227
timestamp 1667941163
transform 1 0 13384 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_229
timestamp 1667941163
transform 1 0 13496 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_254
timestamp 1667941163
transform 1 0 14896 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_280
timestamp 1667941163
transform 1 0 16352 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1667941163
transform 1 0 16688 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_311
timestamp 1667941163
transform 1 0 18088 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_337
timestamp 1667941163
transform 1 0 19544 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_353
timestamp 1667941163
transform 1 0 20440 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_357
timestamp 1667941163
transform 1 0 20664 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_382
timestamp 1667941163
transform 1 0 22064 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_408
timestamp 1667941163
transform 1 0 23520 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_424
timestamp 1667941163
transform 1 0 24416 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_428
timestamp 1667941163
transform 1 0 24640 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_444
timestamp 1667941163
transform 1 0 25536 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_470
timestamp 1667941163
transform 1 0 26992 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1667941163
transform 1 0 28448 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_499
timestamp 1667941163
transform 1 0 28616 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_507
timestamp 1667941163
transform 1 0 29064 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_535
timestamp 1667941163
transform 1 0 30632 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_561
timestamp 1667941163
transform 1 0 32088 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_565
timestamp 1667941163
transform 1 0 32312 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1667941163
transform 1 0 32424 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_570
timestamp 1667941163
transform 1 0 32592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_595
timestamp 1667941163
transform 1 0 33992 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_621
timestamp 1667941163
transform 1 0 35448 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_637
timestamp 1667941163
transform 1 0 36344 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_641
timestamp 1667941163
transform 1 0 36568 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_666
timestamp 1667941163
transform 1 0 37968 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_682
timestamp 1667941163
transform 1 0 38864 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_686
timestamp 1667941163
transform 1 0 39088 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_2
timestamp 1667941163
transform 1 0 784 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1667941163
transform 1 0 2576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_37
timestamp 1667941163
transform 1 0 2744 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_53
timestamp 1667941163
transform 1 0 3640 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_79
timestamp 1667941163
transform 1 0 5096 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1667941163
transform 1 0 6552 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_108
timestamp 1667941163
transform 1 0 6720 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_124
timestamp 1667941163
transform 1 0 7616 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_150
timestamp 1667941163
transform 1 0 9072 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1667941163
transform 1 0 10528 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_179
timestamp 1667941163
transform 1 0 10696 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 11592 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_220
timestamp 1667941163
transform 1 0 12992 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_246
timestamp 1667941163
transform 1 0 14448 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1667941163
transform 1 0 14672 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_275
timestamp 1667941163
transform 1 0 16072 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_301
timestamp 1667941163
transform 1 0 17528 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1667941163
transform 1 0 18424 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1667941163
transform 1 0 18648 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_346
timestamp 1667941163
transform 1 0 20048 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_372
timestamp 1667941163
transform 1 0 21504 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_388
timestamp 1667941163
transform 1 0 22400 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1667941163
transform 1 0 22624 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_417
timestamp 1667941163
transform 1 0 24024 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_443
timestamp 1667941163
transform 1 0 25480 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_459
timestamp 1667941163
transform 1 0 26376 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_463
timestamp 1667941163
transform 1 0 26600 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_471
timestamp 1667941163
transform 1 0 27048 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_499
timestamp 1667941163
transform 1 0 28616 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_525
timestamp 1667941163
transform 1 0 30072 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_529
timestamp 1667941163
transform 1 0 30296 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1667941163
transform 1 0 30408 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_534
timestamp 1667941163
transform 1 0 30576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_559
timestamp 1667941163
transform 1 0 31976 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_585
timestamp 1667941163
transform 1 0 33432 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_601
timestamp 1667941163
transform 1 0 34328 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_605
timestamp 1667941163
transform 1 0 34552 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_630
timestamp 1667941163
transform 1 0 35952 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_656
timestamp 1667941163
transform 1 0 37408 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_672
timestamp 1667941163
transform 1 0 38304 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_676
timestamp 1667941163
transform 1 0 38528 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_684
timestamp 1667941163
transform 1 0 38976 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_2
timestamp 1667941163
transform 1 0 784 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_18
timestamp 1667941163
transform 1 0 1680 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_44
timestamp 1667941163
transform 1 0 3136 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1667941163
transform 1 0 4592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_73
timestamp 1667941163
transform 1 0 4760 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_89
timestamp 1667941163
transform 1 0 5656 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_115
timestamp 1667941163
transform 1 0 7112 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1667941163
transform 1 0 8568 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_144
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_160
timestamp 1667941163
transform 1 0 9632 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_186
timestamp 1667941163
transform 1 0 11088 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1667941163
transform 1 0 12544 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_215
timestamp 1667941163
transform 1 0 12712 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_223
timestamp 1667941163
transform 1 0 13160 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_251
timestamp 1667941163
transform 1 0 14728 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_277
timestamp 1667941163
transform 1 0 16184 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 16408 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1667941163
transform 1 0 16520 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_311
timestamp 1667941163
transform 1 0 18088 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_337
timestamp 1667941163
transform 1 0 19544 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_353
timestamp 1667941163
transform 1 0 20440 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_357
timestamp 1667941163
transform 1 0 20664 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_382
timestamp 1667941163
transform 1 0 22064 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_408
timestamp 1667941163
transform 1 0 23520 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_424
timestamp 1667941163
transform 1 0 24416 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1667941163
transform 1 0 24640 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_453
timestamp 1667941163
transform 1 0 26040 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_469
timestamp 1667941163
transform 1 0 26936 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_471
timestamp 1667941163
transform 1 0 27048 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1667941163
transform 1 0 28448 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_499
timestamp 1667941163
transform 1 0 28616 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_525
timestamp 1667941163
transform 1 0 30072 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_551
timestamp 1667941163
transform 1 0 31528 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1667941163
transform 1 0 32424 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_570
timestamp 1667941163
transform 1 0 32592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_595
timestamp 1667941163
transform 1 0 33992 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_621
timestamp 1667941163
transform 1 0 35448 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_637
timestamp 1667941163
transform 1 0 36344 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_641
timestamp 1667941163
transform 1 0 36568 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_666
timestamp 1667941163
transform 1 0 37968 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_682
timestamp 1667941163
transform 1 0 38864 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_686
timestamp 1667941163
transform 1 0 39088 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_2
timestamp 1667941163
transform 1 0 784 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1667941163
transform 1 0 2576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_37
timestamp 1667941163
transform 1 0 2744 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_53
timestamp 1667941163
transform 1 0 3640 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_79
timestamp 1667941163
transform 1 0 5096 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1667941163
transform 1 0 6552 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_108
timestamp 1667941163
transform 1 0 6720 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_124
timestamp 1667941163
transform 1 0 7616 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_150
timestamp 1667941163
transform 1 0 9072 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1667941163
transform 1 0 10528 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_179
timestamp 1667941163
transform 1 0 10696 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_195
timestamp 1667941163
transform 1 0 11592 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_221
timestamp 1667941163
transform 1 0 13048 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1667941163
transform 1 0 14504 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_250
timestamp 1667941163
transform 1 0 14672 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_275
timestamp 1667941163
transform 1 0 16072 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_301
timestamp 1667941163
transform 1 0 17528 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_317
timestamp 1667941163
transform 1 0 18424 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1667941163
transform 1 0 18648 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_346
timestamp 1667941163
transform 1 0 20048 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_372
timestamp 1667941163
transform 1 0 21504 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_388
timestamp 1667941163
transform 1 0 22400 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_392
timestamp 1667941163
transform 1 0 22624 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_417
timestamp 1667941163
transform 1 0 24024 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_443
timestamp 1667941163
transform 1 0 25480 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_459
timestamp 1667941163
transform 1 0 26376 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_463
timestamp 1667941163
transform 1 0 26600 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_471
timestamp 1667941163
transform 1 0 27048 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_499
timestamp 1667941163
transform 1 0 28616 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_525
timestamp 1667941163
transform 1 0 30072 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_529
timestamp 1667941163
transform 1 0 30296 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1667941163
transform 1 0 30408 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_534
timestamp 1667941163
transform 1 0 30576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_559
timestamp 1667941163
transform 1 0 31976 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_585
timestamp 1667941163
transform 1 0 33432 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_601
timestamp 1667941163
transform 1 0 34328 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_605
timestamp 1667941163
transform 1 0 34552 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_630
timestamp 1667941163
transform 1 0 35952 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_656
timestamp 1667941163
transform 1 0 37408 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_672
timestamp 1667941163
transform 1 0 38304 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_676
timestamp 1667941163
transform 1 0 38528 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_684
timestamp 1667941163
transform 1 0 38976 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_2
timestamp 1667941163
transform 1 0 784 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_18
timestamp 1667941163
transform 1 0 1680 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_44
timestamp 1667941163
transform 1 0 3136 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1667941163
transform 1 0 4592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_73
timestamp 1667941163
transform 1 0 4760 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_89
timestamp 1667941163
transform 1 0 5656 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_115
timestamp 1667941163
transform 1 0 7112 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1667941163
transform 1 0 8568 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_144
timestamp 1667941163
transform 1 0 8736 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_160
timestamp 1667941163
transform 1 0 9632 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_186
timestamp 1667941163
transform 1 0 11088 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1667941163
transform 1 0 12544 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_215
timestamp 1667941163
transform 1 0 12712 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_223
timestamp 1667941163
transform 1 0 13160 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_251
timestamp 1667941163
transform 1 0 14728 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_277
timestamp 1667941163
transform 1 0 16184 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 16408 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1667941163
transform 1 0 16520 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1667941163
transform 1 0 16688 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_311
timestamp 1667941163
transform 1 0 18088 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_337
timestamp 1667941163
transform 1 0 19544 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_353
timestamp 1667941163
transform 1 0 20440 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1667941163
transform 1 0 20664 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_382
timestamp 1667941163
transform 1 0 22064 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_408
timestamp 1667941163
transform 1 0 23520 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_424
timestamp 1667941163
transform 1 0 24416 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_428
timestamp 1667941163
transform 1 0 24640 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_453
timestamp 1667941163
transform 1 0 26040 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_469
timestamp 1667941163
transform 1 0 26936 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_471
timestamp 1667941163
transform 1 0 27048 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1667941163
transform 1 0 28448 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_499
timestamp 1667941163
transform 1 0 28616 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_501
timestamp 1667941163
transform 1 0 28728 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_526
timestamp 1667941163
transform 1 0 30128 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_552
timestamp 1667941163
transform 1 0 31584 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_570
timestamp 1667941163
transform 1 0 32592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_595 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 33992 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_627
timestamp 1667941163
transform 1 0 35784 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_635
timestamp 1667941163
transform 1 0 36232 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_641
timestamp 1667941163
transform 1 0 36568 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_673
timestamp 1667941163
transform 1 0 38360 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_681
timestamp 1667941163
transform 1 0 38808 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_685
timestamp 1667941163
transform 1 0 39032 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_687
timestamp 1667941163
transform 1 0 39144 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_2
timestamp 1667941163
transform 1 0 784 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1667941163
transform 1 0 2576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_37
timestamp 1667941163
transform 1 0 2744 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_53
timestamp 1667941163
transform 1 0 3640 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_79
timestamp 1667941163
transform 1 0 5096 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1667941163
transform 1 0 6552 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_108
timestamp 1667941163
transform 1 0 6720 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_124
timestamp 1667941163
transform 1 0 7616 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_150
timestamp 1667941163
transform 1 0 9072 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1667941163
transform 1 0 10528 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_179
timestamp 1667941163
transform 1 0 10696 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_195
timestamp 1667941163
transform 1 0 11592 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_221
timestamp 1667941163
transform 1 0 13048 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1667941163
transform 1 0 14504 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1667941163
transform 1 0 14672 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_275
timestamp 1667941163
transform 1 0 16072 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_301
timestamp 1667941163
transform 1 0 17528 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_317
timestamp 1667941163
transform 1 0 18424 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1667941163
transform 1 0 18648 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_346
timestamp 1667941163
transform 1 0 20048 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_372
timestamp 1667941163
transform 1 0 21504 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_388
timestamp 1667941163
transform 1 0 22400 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_392
timestamp 1667941163
transform 1 0 22624 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_417
timestamp 1667941163
transform 1 0 24024 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_443
timestamp 1667941163
transform 1 0 25480 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_459
timestamp 1667941163
transform 1 0 26376 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_463
timestamp 1667941163
transform 1 0 26600 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_488
timestamp 1667941163
transform 1 0 28000 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_490
timestamp 1667941163
transform 1 0 28112 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_515
timestamp 1667941163
transform 1 0 29512 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1667941163
transform 1 0 30408 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_534
timestamp 1667941163
transform 1 0 30576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_559
timestamp 1667941163
transform 1 0 31976 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_585
timestamp 1667941163
transform 1 0 33432 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_601
timestamp 1667941163
transform 1 0 34328 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 34552 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1667941163
transform 1 0 38136 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1667941163
transform 1 0 38360 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_676
timestamp 1667941163
transform 1 0 38528 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_684
timestamp 1667941163
transform 1 0 38976 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_2
timestamp 1667941163
transform 1 0 784 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_18
timestamp 1667941163
transform 1 0 1680 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_44
timestamp 1667941163
transform 1 0 3136 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1667941163
transform 1 0 4592 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_73
timestamp 1667941163
transform 1 0 4760 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_89
timestamp 1667941163
transform 1 0 5656 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_115
timestamp 1667941163
transform 1 0 7112 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1667941163
transform 1 0 8568 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_144
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_160
timestamp 1667941163
transform 1 0 9632 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_186
timestamp 1667941163
transform 1 0 11088 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1667941163
transform 1 0 12544 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_215
timestamp 1667941163
transform 1 0 12712 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 13160 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_248
timestamp 1667941163
transform 1 0 14560 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_274
timestamp 1667941163
transform 1 0 16016 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_282
timestamp 1667941163
transform 1 0 16464 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_311
timestamp 1667941163
transform 1 0 18088 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_337
timestamp 1667941163
transform 1 0 19544 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_353
timestamp 1667941163
transform 1 0 20440 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_357
timestamp 1667941163
transform 1 0 20664 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_382
timestamp 1667941163
transform 1 0 22064 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_408
timestamp 1667941163
transform 1 0 23520 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_424
timestamp 1667941163
transform 1 0 24416 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_428
timestamp 1667941163
transform 1 0 24640 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_453
timestamp 1667941163
transform 1 0 26040 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_479
timestamp 1667941163
transform 1 0 27496 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_495
timestamp 1667941163
transform 1 0 28392 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_499
timestamp 1667941163
transform 1 0 28616 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_507
timestamp 1667941163
transform 1 0 29064 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_532
timestamp 1667941163
transform 1 0 30464 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_558
timestamp 1667941163
transform 1 0 31920 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_566
timestamp 1667941163
transform 1 0 32368 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1667941163
transform 1 0 32592 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1667941163
transform 1 0 36176 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1667941163
transform 1 0 36400 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_641
timestamp 1667941163
transform 1 0 36568 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_673
timestamp 1667941163
transform 1 0 38360 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_681
timestamp 1667941163
transform 1 0 38808 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_685
timestamp 1667941163
transform 1 0 39032 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1667941163
transform 1 0 39144 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_2
timestamp 1667941163
transform 1 0 784 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1667941163
transform 1 0 2576 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_37
timestamp 1667941163
transform 1 0 2744 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_53
timestamp 1667941163
transform 1 0 3640 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_79
timestamp 1667941163
transform 1 0 5096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1667941163
transform 1 0 6552 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_108
timestamp 1667941163
transform 1 0 6720 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_124
timestamp 1667941163
transform 1 0 7616 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_150
timestamp 1667941163
transform 1 0 9072 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1667941163
transform 1 0 10528 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_179
timestamp 1667941163
transform 1 0 10696 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 11592 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_220
timestamp 1667941163
transform 1 0 12992 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_246
timestamp 1667941163
transform 1 0 14448 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_250
timestamp 1667941163
transform 1 0 14672 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_275
timestamp 1667941163
transform 1 0 16072 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_301
timestamp 1667941163
transform 1 0 17528 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_317
timestamp 1667941163
transform 1 0 18424 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1667941163
transform 1 0 18648 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_346
timestamp 1667941163
transform 1 0 20048 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_372
timestamp 1667941163
transform 1 0 21504 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_388
timestamp 1667941163
transform 1 0 22400 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1667941163
transform 1 0 22624 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_417
timestamp 1667941163
transform 1 0 24024 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_443
timestamp 1667941163
transform 1 0 25480 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_459
timestamp 1667941163
transform 1 0 26376 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_463
timestamp 1667941163
transform 1 0 26600 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_495
timestamp 1667941163
transform 1 0 28392 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_503
timestamp 1667941163
transform 1 0 28840 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1667941163
transform 1 0 30408 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1667941163
transform 1 0 30576 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1667941163
transform 1 0 34160 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1667941163
transform 1 0 34384 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1667941163
transform 1 0 34552 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1667941163
transform 1 0 38136 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1667941163
transform 1 0 38360 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_676
timestamp 1667941163
transform 1 0 38528 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_684
timestamp 1667941163
transform 1 0 38976 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_2
timestamp 1667941163
transform 1 0 784 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_18
timestamp 1667941163
transform 1 0 1680 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_44
timestamp 1667941163
transform 1 0 3136 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1667941163
transform 1 0 4592 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_73
timestamp 1667941163
transform 1 0 4760 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_89
timestamp 1667941163
transform 1 0 5656 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_115
timestamp 1667941163
transform 1 0 7112 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1667941163
transform 1 0 8568 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_144
timestamp 1667941163
transform 1 0 8736 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_160
timestamp 1667941163
transform 1 0 9632 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_186
timestamp 1667941163
transform 1 0 11088 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1667941163
transform 1 0 12544 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1667941163
transform 1 0 12712 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_240
timestamp 1667941163
transform 1 0 14112 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_266
timestamp 1667941163
transform 1 0 15568 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_282
timestamp 1667941163
transform 1 0 16464 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1667941163
transform 1 0 16688 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_311
timestamp 1667941163
transform 1 0 18088 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_337
timestamp 1667941163
transform 1 0 19544 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_353
timestamp 1667941163
transform 1 0 20440 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1667941163
transform 1 0 20664 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_382
timestamp 1667941163
transform 1 0 22064 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_408
timestamp 1667941163
transform 1 0 23520 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_424
timestamp 1667941163
transform 1 0 24416 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_428
timestamp 1667941163
transform 1 0 24640 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_453
timestamp 1667941163
transform 1 0 26040 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_485
timestamp 1667941163
transform 1 0 27832 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_493
timestamp 1667941163
transform 1 0 28280 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1667941163
transform 1 0 28616 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1667941163
transform 1 0 32200 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1667941163
transform 1 0 32424 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1667941163
transform 1 0 32592 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1667941163
transform 1 0 36176 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1667941163
transform 1 0 36400 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_641
timestamp 1667941163
transform 1 0 36568 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_673
timestamp 1667941163
transform 1 0 38360 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_681
timestamp 1667941163
transform 1 0 38808 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_685
timestamp 1667941163
transform 1 0 39032 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1667941163
transform 1 0 39144 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_2
timestamp 1667941163
transform 1 0 784 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1667941163
transform 1 0 2576 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_37
timestamp 1667941163
transform 1 0 2744 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_53
timestamp 1667941163
transform 1 0 3640 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_79
timestamp 1667941163
transform 1 0 5096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1667941163
transform 1 0 6552 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_108
timestamp 1667941163
transform 1 0 6720 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_124
timestamp 1667941163
transform 1 0 7616 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_150
timestamp 1667941163
transform 1 0 9072 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1667941163
transform 1 0 10528 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_179
timestamp 1667941163
transform 1 0 10696 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_181
timestamp 1667941163
transform 1 0 10808 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_206
timestamp 1667941163
transform 1 0 12208 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_232
timestamp 1667941163
transform 1 0 13664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_250
timestamp 1667941163
transform 1 0 14672 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_275
timestamp 1667941163
transform 1 0 16072 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_301
timestamp 1667941163
transform 1 0 17528 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_317
timestamp 1667941163
transform 1 0 18424 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1667941163
transform 1 0 18648 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_346
timestamp 1667941163
transform 1 0 20048 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_372
timestamp 1667941163
transform 1 0 21504 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_388
timestamp 1667941163
transform 1 0 22400 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_392
timestamp 1667941163
transform 1 0 22624 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_417
timestamp 1667941163
transform 1 0 24024 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_443
timestamp 1667941163
transform 1 0 25480 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_459
timestamp 1667941163
transform 1 0 26376 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1667941163
transform 1 0 26600 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1667941163
transform 1 0 30184 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1667941163
transform 1 0 30408 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1667941163
transform 1 0 30576 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1667941163
transform 1 0 34160 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1667941163
transform 1 0 34384 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1667941163
transform 1 0 34552 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1667941163
transform 1 0 38136 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1667941163
transform 1 0 38360 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_676
timestamp 1667941163
transform 1 0 38528 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_684
timestamp 1667941163
transform 1 0 38976 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_2
timestamp 1667941163
transform 1 0 784 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_18
timestamp 1667941163
transform 1 0 1680 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_44
timestamp 1667941163
transform 1 0 3136 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1667941163
transform 1 0 4592 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_73
timestamp 1667941163
transform 1 0 4760 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_89
timestamp 1667941163
transform 1 0 5656 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_115
timestamp 1667941163
transform 1 0 7112 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1667941163
transform 1 0 8568 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_144
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_160
timestamp 1667941163
transform 1 0 9632 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_186
timestamp 1667941163
transform 1 0 11088 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1667941163
transform 1 0 12544 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1667941163
transform 1 0 12712 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_240
timestamp 1667941163
transform 1 0 14112 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_266
timestamp 1667941163
transform 1 0 15568 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_282
timestamp 1667941163
transform 1 0 16464 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_286
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_311
timestamp 1667941163
transform 1 0 18088 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_337
timestamp 1667941163
transform 1 0 19544 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_353
timestamp 1667941163
transform 1 0 20440 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1667941163
transform 1 0 20664 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_382
timestamp 1667941163
transform 1 0 22064 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_408
timestamp 1667941163
transform 1 0 23520 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_424
timestamp 1667941163
transform 1 0 24416 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1667941163
transform 1 0 24640 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_453
timestamp 1667941163
transform 1 0 26040 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_485
timestamp 1667941163
transform 1 0 27832 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_493
timestamp 1667941163
transform 1 0 28280 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1667941163
transform 1 0 28616 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1667941163
transform 1 0 32200 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1667941163
transform 1 0 32424 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1667941163
transform 1 0 32592 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1667941163
transform 1 0 36176 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1667941163
transform 1 0 36400 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_641
timestamp 1667941163
transform 1 0 36568 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_673
timestamp 1667941163
transform 1 0 38360 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_681
timestamp 1667941163
transform 1 0 38808 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_685
timestamp 1667941163
transform 1 0 39032 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1667941163
transform 1 0 39144 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_2
timestamp 1667941163
transform 1 0 784 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1667941163
transform 1 0 2576 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_37
timestamp 1667941163
transform 1 0 2744 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_53
timestamp 1667941163
transform 1 0 3640 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_79
timestamp 1667941163
transform 1 0 5096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1667941163
transform 1 0 6552 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_108
timestamp 1667941163
transform 1 0 6720 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_124
timestamp 1667941163
transform 1 0 7616 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_150
timestamp 1667941163
transform 1 0 9072 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1667941163
transform 1 0 10528 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_179
timestamp 1667941163
transform 1 0 10696 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_195
timestamp 1667941163
transform 1 0 11592 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_221
timestamp 1667941163
transform 1 0 13048 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1667941163
transform 1 0 14504 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1667941163
transform 1 0 14672 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_275
timestamp 1667941163
transform 1 0 16072 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_301
timestamp 1667941163
transform 1 0 17528 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1667941163
transform 1 0 18424 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1667941163
transform 1 0 18648 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_346
timestamp 1667941163
transform 1 0 20048 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_372
timestamp 1667941163
transform 1 0 21504 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_388
timestamp 1667941163
transform 1 0 22400 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1667941163
transform 1 0 22624 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_417
timestamp 1667941163
transform 1 0 24024 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_443
timestamp 1667941163
transform 1 0 25480 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_459
timestamp 1667941163
transform 1 0 26376 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1667941163
transform 1 0 26600 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1667941163
transform 1 0 30184 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1667941163
transform 1 0 30408 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1667941163
transform 1 0 30576 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1667941163
transform 1 0 34160 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1667941163
transform 1 0 34384 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1667941163
transform 1 0 34552 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1667941163
transform 1 0 38136 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1667941163
transform 1 0 38360 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_676
timestamp 1667941163
transform 1 0 38528 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_684
timestamp 1667941163
transform 1 0 38976 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_2
timestamp 1667941163
transform 1 0 784 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_18
timestamp 1667941163
transform 1 0 1680 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_44
timestamp 1667941163
transform 1 0 3136 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1667941163
transform 1 0 4592 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_73
timestamp 1667941163
transform 1 0 4760 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_89
timestamp 1667941163
transform 1 0 5656 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_115
timestamp 1667941163
transform 1 0 7112 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1667941163
transform 1 0 8568 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_144
timestamp 1667941163
transform 1 0 8736 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_160
timestamp 1667941163
transform 1 0 9632 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_186
timestamp 1667941163
transform 1 0 11088 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1667941163
transform 1 0 12544 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1667941163
transform 1 0 12712 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_240
timestamp 1667941163
transform 1 0 14112 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_266
timestamp 1667941163
transform 1 0 15568 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_282
timestamp 1667941163
transform 1 0 16464 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1667941163
transform 1 0 16688 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_311
timestamp 1667941163
transform 1 0 18088 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_337
timestamp 1667941163
transform 1 0 19544 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_353
timestamp 1667941163
transform 1 0 20440 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1667941163
transform 1 0 20664 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1667941163
transform 1 0 24248 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1667941163
transform 1 0 24472 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1667941163
transform 1 0 24640 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1667941163
transform 1 0 28224 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1667941163
transform 1 0 28448 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1667941163
transform 1 0 28616 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1667941163
transform 1 0 32200 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1667941163
transform 1 0 32424 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1667941163
transform 1 0 32592 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1667941163
transform 1 0 36176 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1667941163
transform 1 0 36400 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_641
timestamp 1667941163
transform 1 0 36568 0 -1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_673
timestamp 1667941163
transform 1 0 38360 0 -1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_681
timestamp 1667941163
transform 1 0 38808 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_685
timestamp 1667941163
transform 1 0 39032 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_687
timestamp 1667941163
transform 1 0 39144 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_2
timestamp 1667941163
transform 1 0 784 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1667941163
transform 1 0 2576 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_37
timestamp 1667941163
transform 1 0 2744 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_53
timestamp 1667941163
transform 1 0 3640 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_79
timestamp 1667941163
transform 1 0 5096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1667941163
transform 1 0 6552 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_108
timestamp 1667941163
transform 1 0 6720 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_124
timestamp 1667941163
transform 1 0 7616 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_150
timestamp 1667941163
transform 1 0 9072 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1667941163
transform 1 0 10528 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_179
timestamp 1667941163
transform 1 0 10696 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_219
timestamp 1667941163
transform 1 0 12936 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_245
timestamp 1667941163
transform 1 0 14392 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1667941163
transform 1 0 14504 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1667941163
transform 1 0 14672 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_275
timestamp 1667941163
transform 1 0 16072 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_301
timestamp 1667941163
transform 1 0 17528 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1667941163
transform 1 0 18424 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1667941163
transform 1 0 18648 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_346
timestamp 1667941163
transform 1 0 20048 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_378
timestamp 1667941163
transform 1 0 21840 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_386
timestamp 1667941163
transform 1 0 22288 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1667941163
transform 1 0 22624 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1667941163
transform 1 0 26208 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1667941163
transform 1 0 26432 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1667941163
transform 1 0 26600 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1667941163
transform 1 0 30184 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1667941163
transform 1 0 30408 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1667941163
transform 1 0 30576 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1667941163
transform 1 0 34160 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1667941163
transform 1 0 34384 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1667941163
transform 1 0 34552 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1667941163
transform 1 0 38136 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1667941163
transform 1 0 38360 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_676
timestamp 1667941163
transform 1 0 38528 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_684
timestamp 1667941163
transform 1 0 38976 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1667941163
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1667941163
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1667941163
transform 1 0 4592 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_73
timestamp 1667941163
transform 1 0 4760 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_89
timestamp 1667941163
transform 1 0 5656 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_115
timestamp 1667941163
transform 1 0 7112 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1667941163
transform 1 0 8568 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_144
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_160
timestamp 1667941163
transform 1 0 9632 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_186
timestamp 1667941163
transform 1 0 11088 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1667941163
transform 1 0 12544 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1667941163
transform 1 0 12712 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_240
timestamp 1667941163
transform 1 0 14112 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_266
timestamp 1667941163
transform 1 0 15568 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1667941163
transform 1 0 16464 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1667941163
transform 1 0 20272 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1667941163
transform 1 0 20496 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_357
timestamp 1667941163
transform 1 0 20664 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_373
timestamp 1667941163
transform 1 0 21560 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_377
timestamp 1667941163
transform 1 0 21784 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_382
timestamp 1667941163
transform 1 0 22064 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_388
timestamp 1667941163
transform 1 0 22400 0 -1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_420
timestamp 1667941163
transform 1 0 24192 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_424
timestamp 1667941163
transform 1 0 24416 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1667941163
transform 1 0 24640 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1667941163
transform 1 0 28224 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1667941163
transform 1 0 28448 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1667941163
transform 1 0 28616 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1667941163
transform 1 0 32200 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1667941163
transform 1 0 32424 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1667941163
transform 1 0 32592 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1667941163
transform 1 0 36176 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1667941163
transform 1 0 36400 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_641
timestamp 1667941163
transform 1 0 36568 0 -1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_673
timestamp 1667941163
transform 1 0 38360 0 -1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_681
timestamp 1667941163
transform 1 0 38808 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_685
timestamp 1667941163
transform 1 0 39032 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1667941163
transform 1 0 39144 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1667941163
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1667941163
transform 1 0 2576 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_37
timestamp 1667941163
transform 1 0 2744 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_69
timestamp 1667941163
transform 1 0 4536 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_77
timestamp 1667941163
transform 1 0 4984 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1667941163
transform 1 0 6552 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_108
timestamp 1667941163
transform 1 0 6720 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_124
timestamp 1667941163
transform 1 0 7616 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_150
timestamp 1667941163
transform 1 0 9072 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1667941163
transform 1 0 10528 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_179
timestamp 1667941163
transform 1 0 10696 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_219
timestamp 1667941163
transform 1 0 12936 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_245
timestamp 1667941163
transform 1 0 14392 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1667941163
transform 1 0 14504 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_250
timestamp 1667941163
transform 1 0 14672 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_275
timestamp 1667941163
transform 1 0 16072 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_301
timestamp 1667941163
transform 1 0 17528 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_317
timestamp 1667941163
transform 1 0 18424 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_321
timestamp 1667941163
transform 1 0 18648 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_353
timestamp 1667941163
transform 1 0 20440 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_361
timestamp 1667941163
transform 1 0 20888 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_369
timestamp 1667941163
transform 1 0 21336 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_375
timestamp 1667941163
transform 1 0 21672 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_381
timestamp 1667941163
transform 1 0 22008 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_387
timestamp 1667941163
transform 1 0 22344 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1667941163
transform 1 0 22456 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1667941163
transform 1 0 22624 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1667941163
transform 1 0 26208 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1667941163
transform 1 0 26432 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1667941163
transform 1 0 26600 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1667941163
transform 1 0 30184 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1667941163
transform 1 0 30408 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1667941163
transform 1 0 30576 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1667941163
transform 1 0 34160 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1667941163
transform 1 0 34384 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1667941163
transform 1 0 34552 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1667941163
transform 1 0 38136 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1667941163
transform 1 0 38360 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_676
timestamp 1667941163
transform 1 0 38528 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_684
timestamp 1667941163
transform 1 0 38976 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1667941163
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1667941163
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1667941163
transform 1 0 4592 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_73
timestamp 1667941163
transform 1 0 4760 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_89
timestamp 1667941163
transform 1 0 5656 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_115
timestamp 1667941163
transform 1 0 7112 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1667941163
transform 1 0 8568 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_144
timestamp 1667941163
transform 1 0 8736 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_184
timestamp 1667941163
transform 1 0 10976 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_210
timestamp 1667941163
transform 1 0 12432 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1667941163
transform 1 0 12544 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_215
timestamp 1667941163
transform 1 0 12712 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_240
timestamp 1667941163
transform 1 0 14112 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_266
timestamp 1667941163
transform 1 0 15568 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1667941163
transform 1 0 16464 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1667941163
transform 1 0 16688 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1667941163
transform 1 0 20272 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1667941163
transform 1 0 20496 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_357
timestamp 1667941163
transform 1 0 20664 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_373
timestamp 1667941163
transform 1 0 21560 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_377
timestamp 1667941163
transform 1 0 21784 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_382
timestamp 1667941163
transform 1 0 22064 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_388
timestamp 1667941163
transform 1 0 22400 0 -1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_420
timestamp 1667941163
transform 1 0 24192 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_424
timestamp 1667941163
transform 1 0 24416 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1667941163
transform 1 0 24640 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1667941163
transform 1 0 28224 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1667941163
transform 1 0 28448 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1667941163
transform 1 0 28616 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1667941163
transform 1 0 32200 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1667941163
transform 1 0 32424 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1667941163
transform 1 0 32592 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1667941163
transform 1 0 36176 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1667941163
transform 1 0 36400 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_641
timestamp 1667941163
transform 1 0 36568 0 -1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_673
timestamp 1667941163
transform 1 0 38360 0 -1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_681
timestamp 1667941163
transform 1 0 38808 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_685
timestamp 1667941163
transform 1 0 39032 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_687
timestamp 1667941163
transform 1 0 39144 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1667941163
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1667941163
transform 1 0 2576 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1667941163
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1667941163
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1667941163
transform 1 0 6552 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_108
timestamp 1667941163
transform 1 0 6720 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_140
timestamp 1667941163
transform 1 0 8512 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_148
timestamp 1667941163
transform 1 0 8960 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1667941163
transform 1 0 10528 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1667941163
transform 1 0 10696 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_204
timestamp 1667941163
transform 1 0 12096 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_230
timestamp 1667941163
transform 1 0 13552 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_246
timestamp 1667941163
transform 1 0 14448 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1667941163
transform 1 0 14672 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1667941163
transform 1 0 18256 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1667941163
transform 1 0 18480 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1667941163
transform 1 0 18648 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1667941163
transform 1 0 22232 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1667941163
transform 1 0 22456 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1667941163
transform 1 0 22624 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1667941163
transform 1 0 26208 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1667941163
transform 1 0 26432 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1667941163
transform 1 0 26600 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1667941163
transform 1 0 30184 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1667941163
transform 1 0 30408 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1667941163
transform 1 0 30576 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1667941163
transform 1 0 34160 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1667941163
transform 1 0 34384 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1667941163
transform 1 0 34552 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1667941163
transform 1 0 38136 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1667941163
transform 1 0 38360 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_676
timestamp 1667941163
transform 1 0 38528 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_684
timestamp 1667941163
transform 1 0 38976 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1667941163
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1667941163
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1667941163
transform 1 0 4592 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1667941163
transform 1 0 4760 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1667941163
transform 1 0 8344 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1667941163
transform 1 0 8568 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_144
timestamp 1667941163
transform 1 0 8736 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_152
timestamp 1667941163
transform 1 0 9184 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_156
timestamp 1667941163
transform 1 0 9408 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_158
timestamp 1667941163
transform 1 0 9520 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_183
timestamp 1667941163
transform 1 0 10920 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_209
timestamp 1667941163
transform 1 0 12376 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1667941163
transform 1 0 12712 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_240
timestamp 1667941163
transform 1 0 14112 0 -1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_272
timestamp 1667941163
transform 1 0 15904 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_280
timestamp 1667941163
transform 1 0 16352 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1667941163
transform 1 0 16688 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1667941163
transform 1 0 20272 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1667941163
transform 1 0 20496 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1667941163
transform 1 0 20664 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1667941163
transform 1 0 24248 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1667941163
transform 1 0 24472 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1667941163
transform 1 0 24640 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1667941163
transform 1 0 28224 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1667941163
transform 1 0 28448 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1667941163
transform 1 0 28616 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1667941163
transform 1 0 32200 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1667941163
transform 1 0 32424 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1667941163
transform 1 0 32592 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1667941163
transform 1 0 36176 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1667941163
transform 1 0 36400 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_641
timestamp 1667941163
transform 1 0 36568 0 -1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_673
timestamp 1667941163
transform 1 0 38360 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_681
timestamp 1667941163
transform 1 0 38808 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_685
timestamp 1667941163
transform 1 0 39032 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_687
timestamp 1667941163
transform 1 0 39144 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1667941163
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1667941163
transform 1 0 2576 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1667941163
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1667941163
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1667941163
transform 1 0 6552 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1667941163
transform 1 0 6720 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1667941163
transform 1 0 10304 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1667941163
transform 1 0 10528 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_179
timestamp 1667941163
transform 1 0 10696 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_195
timestamp 1667941163
transform 1 0 11592 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_203
timestamp 1667941163
transform 1 0 12040 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_229
timestamp 1667941163
transform 1 0 13496 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_245
timestamp 1667941163
transform 1 0 14392 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1667941163
transform 1 0 14504 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1667941163
transform 1 0 14672 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1667941163
transform 1 0 18256 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1667941163
transform 1 0 18480 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1667941163
transform 1 0 18648 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1667941163
transform 1 0 22232 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1667941163
transform 1 0 22456 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1667941163
transform 1 0 22624 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1667941163
transform 1 0 26208 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1667941163
transform 1 0 26432 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1667941163
transform 1 0 26600 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1667941163
transform 1 0 30184 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1667941163
transform 1 0 30408 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1667941163
transform 1 0 30576 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1667941163
transform 1 0 34160 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1667941163
transform 1 0 34384 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1667941163
transform 1 0 34552 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1667941163
transform 1 0 38136 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1667941163
transform 1 0 38360 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_676
timestamp 1667941163
transform 1 0 38528 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_684
timestamp 1667941163
transform 1 0 38976 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1667941163
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1667941163
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1667941163
transform 1 0 4592 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1667941163
transform 1 0 4760 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1667941163
transform 1 0 8344 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1667941163
transform 1 0 8568 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1667941163
transform 1 0 8736 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1667941163
transform 1 0 12320 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1667941163
transform 1 0 12544 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1667941163
transform 1 0 12712 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1667941163
transform 1 0 16296 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1667941163
transform 1 0 16520 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1667941163
transform 1 0 16688 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1667941163
transform 1 0 20272 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1667941163
transform 1 0 20496 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1667941163
transform 1 0 20664 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1667941163
transform 1 0 24248 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1667941163
transform 1 0 24472 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1667941163
transform 1 0 24640 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1667941163
transform 1 0 28224 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1667941163
transform 1 0 28448 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1667941163
transform 1 0 28616 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1667941163
transform 1 0 32200 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1667941163
transform 1 0 32424 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1667941163
transform 1 0 32592 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1667941163
transform 1 0 36176 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1667941163
transform 1 0 36400 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_641
timestamp 1667941163
transform 1 0 36568 0 -1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_673
timestamp 1667941163
transform 1 0 38360 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_681
timestamp 1667941163
transform 1 0 38808 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_685
timestamp 1667941163
transform 1 0 39032 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_687
timestamp 1667941163
transform 1 0 39144 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1667941163
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1667941163
transform 1 0 2576 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_37
timestamp 1667941163
transform 1 0 2744 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_69
timestamp 1667941163
transform 1 0 4536 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_72
timestamp 1667941163
transform 1 0 4704 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1667941163
transform 1 0 6496 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_107
timestamp 1667941163
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 8456 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_142
timestamp 1667941163
transform 1 0 8624 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1667941163
transform 1 0 10416 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1667941163
transform 1 0 10584 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1667941163
transform 1 0 12376 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_212
timestamp 1667941163
transform 1 0 12544 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1667941163
transform 1 0 14336 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_247
timestamp 1667941163
transform 1 0 14504 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_279
timestamp 1667941163
transform 1 0 16296 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_282
timestamp 1667941163
transform 1 0 16464 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1667941163
transform 1 0 18256 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_317
timestamp 1667941163
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_349
timestamp 1667941163
transform 1 0 20216 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_352
timestamp 1667941163
transform 1 0 20384 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1667941163
transform 1 0 22176 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_387
timestamp 1667941163
transform 1 0 22344 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1667941163
transform 1 0 24136 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_422
timestamp 1667941163
transform 1 0 24304 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1667941163
transform 1 0 26096 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_457
timestamp 1667941163
transform 1 0 26264 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_489
timestamp 1667941163
transform 1 0 28056 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_492
timestamp 1667941163
transform 1 0 28224 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1667941163
transform 1 0 30016 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_527
timestamp 1667941163
transform 1 0 30184 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_559
timestamp 1667941163
transform 1 0 31976 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_562
timestamp 1667941163
transform 1 0 32144 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_594
timestamp 1667941163
transform 1 0 33936 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_597
timestamp 1667941163
transform 1 0 34104 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_629
timestamp 1667941163
transform 1 0 35896 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_632
timestamp 1667941163
transform 1 0 36064 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1667941163
transform 1 0 37856 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_667
timestamp 1667941163
transform 1 0 38024 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_683
timestamp 1667941163
transform 1 0 38920 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_687
timestamp 1667941163
transform 1 0 39144 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 39312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 39312 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 39312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 39312 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 39312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 39312 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 39312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 39312 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 39312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 39312 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 39312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 39312 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 39312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 39312 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 39312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 39312 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 39312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1667941163
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1667941163
transform -1 0 39312 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1667941163
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1667941163
transform -1 0 39312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1667941163
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1667941163
transform -1 0 39312 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1667941163
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1667941163
transform -1 0 39312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1667941163
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1667941163
transform -1 0 39312 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1667941163
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1667941163
transform -1 0 39312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1667941163
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1667941163
transform -1 0 39312 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1667941163
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1667941163
transform -1 0 39312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1667941163
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1667941163
transform -1 0 39312 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1667941163
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1667941163
transform -1 0 39312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1667941163
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1667941163
transform -1 0 39312 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1667941163
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1667941163
transform -1 0 39312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1667941163
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1667941163
transform -1 0 39312 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1667941163
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1667941163
transform -1 0 39312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1667941163
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1667941163
transform -1 0 39312 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1667941163
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1667941163
transform -1 0 39312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1667941163
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1667941163
transform -1 0 39312 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1667941163
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1667941163
transform -1 0 39312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1667941163
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1667941163
transform -1 0 39312 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1667941163
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1667941163
transform -1 0 39312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1667941163
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1667941163
transform -1 0 39312 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1667941163
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1667941163
transform -1 0 39312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1667941163
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1667941163
transform -1 0 39312 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1667941163
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1667941163
transform -1 0 39312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1667941163
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1667941163
transform -1 0 39312 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1667941163
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1667941163
transform -1 0 39312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1667941163
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1667941163
transform 1 0 8512 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1667941163
transform 1 0 10472 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1667941163
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1667941163
transform 1 0 14392 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1667941163
transform 1 0 16352 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1667941163
transform 1 0 18312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1667941163
transform 1 0 20272 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1667941163
transform 1 0 22232 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1667941163
transform 1 0 24192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1667941163
transform 1 0 26152 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1667941163
transform 1 0 28112 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1667941163
transform 1 0 30072 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1667941163
transform 1 0 32032 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1667941163
transform 1 0 33992 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1667941163
transform 1 0 35952 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1667941163
transform 1 0 37912 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1667941163
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1667941163
transform 1 0 12600 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1667941163
transform 1 0 16576 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1667941163
transform 1 0 20552 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1667941163
transform 1 0 24528 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1667941163
transform 1 0 28504 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1667941163
transform 1 0 32480 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1667941163
transform 1 0 36456 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1667941163
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1667941163
transform 1 0 10584 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1667941163
transform 1 0 14560 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1667941163
transform 1 0 18536 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1667941163
transform 1 0 22512 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1667941163
transform 1 0 26488 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1667941163
transform 1 0 30464 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1667941163
transform 1 0 34440 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1667941163
transform 1 0 38416 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1667941163
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1667941163
transform 1 0 12600 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1667941163
transform 1 0 16576 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1667941163
transform 1 0 20552 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1667941163
transform 1 0 24528 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1667941163
transform 1 0 28504 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1667941163
transform 1 0 32480 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1667941163
transform 1 0 36456 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1667941163
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1667941163
transform 1 0 10584 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1667941163
transform 1 0 14560 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1667941163
transform 1 0 18536 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1667941163
transform 1 0 22512 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1667941163
transform 1 0 26488 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1667941163
transform 1 0 30464 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1667941163
transform 1 0 34440 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1667941163
transform 1 0 38416 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1667941163
transform 1 0 8624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1667941163
transform 1 0 12600 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1667941163
transform 1 0 16576 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1667941163
transform 1 0 20552 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1667941163
transform 1 0 24528 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1667941163
transform 1 0 28504 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1667941163
transform 1 0 32480 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1667941163
transform 1 0 36456 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1667941163
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1667941163
transform 1 0 10584 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1667941163
transform 1 0 14560 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1667941163
transform 1 0 18536 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1667941163
transform 1 0 22512 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1667941163
transform 1 0 26488 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1667941163
transform 1 0 30464 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1667941163
transform 1 0 34440 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1667941163
transform 1 0 38416 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1667941163
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 8624 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 12600 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 16576 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 20552 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 24528 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 28504 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 32480 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 36456 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 10584 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 14560 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 18536 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 22512 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 26488 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 30464 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 34440 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 38416 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 8624 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 12600 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 16576 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 20552 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 24528 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 28504 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 32480 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 36456 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 10584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 14560 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 18536 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 22512 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 26488 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 30464 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 34440 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 38416 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 4648 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 12600 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 16576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 20552 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 24528 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 28504 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 32480 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 36456 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 6608 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 14560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 18536 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 22512 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 26488 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 30464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 34440 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 38416 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 4648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 12600 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 16576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 20552 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 24528 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 28504 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 32480 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 36456 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 6608 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 14560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 18536 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 22512 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 26488 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 30464 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 34440 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 38416 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 4648 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 12600 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 16576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 20552 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 24528 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 28504 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 32480 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 36456 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 6608 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 14560 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 18536 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 22512 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 26488 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 30464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 34440 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 38416 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 4648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 12600 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 16576 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 20552 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 24528 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 28504 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 32480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 36456 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 6608 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 14560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 18536 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 22512 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 26488 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 30464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 34440 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 38416 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 4648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 12600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 16576 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 20552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 24528 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 28504 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 32480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 36456 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 6608 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1667941163
transform 1 0 14560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1667941163
transform 1 0 18536 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1667941163
transform 1 0 22512 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1667941163
transform 1 0 26488 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1667941163
transform 1 0 30464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1667941163
transform 1 0 34440 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1667941163
transform 1 0 38416 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1667941163
transform 1 0 4648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1667941163
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1667941163
transform 1 0 12600 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1667941163
transform 1 0 16576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1667941163
transform 1 0 20552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1667941163
transform 1 0 24528 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1667941163
transform 1 0 28504 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1667941163
transform 1 0 32480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1667941163
transform 1 0 36456 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1667941163
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1667941163
transform 1 0 6608 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1667941163
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1667941163
transform 1 0 14560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1667941163
transform 1 0 18536 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1667941163
transform 1 0 22512 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1667941163
transform 1 0 26488 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1667941163
transform 1 0 30464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1667941163
transform 1 0 34440 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1667941163
transform 1 0 38416 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1667941163
transform 1 0 4648 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1667941163
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1667941163
transform 1 0 12600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1667941163
transform 1 0 16576 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1667941163
transform 1 0 20552 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1667941163
transform 1 0 24528 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1667941163
transform 1 0 28504 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1667941163
transform 1 0 32480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1667941163
transform 1 0 36456 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1667941163
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1667941163
transform 1 0 6608 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1667941163
transform 1 0 10584 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1667941163
transform 1 0 14560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1667941163
transform 1 0 18536 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1667941163
transform 1 0 22512 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1667941163
transform 1 0 26488 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1667941163
transform 1 0 30464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1667941163
transform 1 0 34440 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1667941163
transform 1 0 38416 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1667941163
transform 1 0 4648 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1667941163
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1667941163
transform 1 0 12600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1667941163
transform 1 0 16576 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1667941163
transform 1 0 20552 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1667941163
transform 1 0 24528 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1667941163
transform 1 0 28504 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1667941163
transform 1 0 32480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1667941163
transform 1 0 36456 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1667941163
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1667941163
transform 1 0 6608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1667941163
transform 1 0 10584 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1667941163
transform 1 0 14560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1667941163
transform 1 0 18536 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1667941163
transform 1 0 22512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1667941163
transform 1 0 26488 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1667941163
transform 1 0 30464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1667941163
transform 1 0 34440 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1667941163
transform 1 0 38416 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1667941163
transform 1 0 4648 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1667941163
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1667941163
transform 1 0 12600 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1667941163
transform 1 0 16576 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1667941163
transform 1 0 20552 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1667941163
transform 1 0 24528 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1667941163
transform 1 0 28504 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1667941163
transform 1 0 32480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1667941163
transform 1 0 36456 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1667941163
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1667941163
transform 1 0 6608 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1667941163
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1667941163
transform 1 0 14560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1667941163
transform 1 0 18536 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1667941163
transform 1 0 22512 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1667941163
transform 1 0 26488 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1667941163
transform 1 0 30464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1667941163
transform 1 0 34440 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1667941163
transform 1 0 38416 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1667941163
transform 1 0 4648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1667941163
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1667941163
transform 1 0 12600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1667941163
transform 1 0 16576 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1667941163
transform 1 0 20552 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1667941163
transform 1 0 24528 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1667941163
transform 1 0 28504 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1667941163
transform 1 0 32480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1667941163
transform 1 0 36456 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1667941163
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1667941163
transform 1 0 6608 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1667941163
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1667941163
transform 1 0 14560 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1667941163
transform 1 0 18536 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1667941163
transform 1 0 22512 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1667941163
transform 1 0 26488 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1667941163
transform 1 0 30464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1667941163
transform 1 0 34440 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1667941163
transform 1 0 38416 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1667941163
transform 1 0 4648 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1667941163
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1667941163
transform 1 0 12600 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1667941163
transform 1 0 16576 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1667941163
transform 1 0 20552 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1667941163
transform 1 0 24528 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1667941163
transform 1 0 28504 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1667941163
transform 1 0 32480 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1667941163
transform 1 0 36456 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1667941163
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1667941163
transform 1 0 6608 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1667941163
transform 1 0 10584 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1667941163
transform 1 0 14560 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1667941163
transform 1 0 18536 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1667941163
transform 1 0 22512 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1667941163
transform 1 0 26488 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1667941163
transform 1 0 30464 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1667941163
transform 1 0 34440 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1667941163
transform 1 0 38416 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1667941163
transform 1 0 4648 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1667941163
transform 1 0 8624 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1667941163
transform 1 0 12600 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1667941163
transform 1 0 16576 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1667941163
transform 1 0 20552 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1667941163
transform 1 0 24528 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1667941163
transform 1 0 28504 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1667941163
transform 1 0 32480 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1667941163
transform 1 0 36456 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1667941163
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1667941163
transform 1 0 6608 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1667941163
transform 1 0 10584 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1667941163
transform 1 0 14560 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1667941163
transform 1 0 18536 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1667941163
transform 1 0 22512 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1667941163
transform 1 0 26488 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1667941163
transform 1 0 30464 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1667941163
transform 1 0 34440 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1667941163
transform 1 0 38416 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1667941163
transform 1 0 4648 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1667941163
transform 1 0 8624 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1667941163
transform 1 0 12600 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1667941163
transform 1 0 16576 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1667941163
transform 1 0 20552 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1667941163
transform 1 0 24528 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1667941163
transform 1 0 28504 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1667941163
transform 1 0 32480 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1667941163
transform 1 0 36456 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1667941163
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1667941163
transform 1 0 6608 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1667941163
transform 1 0 10584 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1667941163
transform 1 0 14560 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1667941163
transform 1 0 18536 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1667941163
transform 1 0 22512 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1667941163
transform 1 0 26488 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1667941163
transform 1 0 30464 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1667941163
transform 1 0 34440 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1667941163
transform 1 0 38416 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1667941163
transform 1 0 4648 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1667941163
transform 1 0 8624 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1667941163
transform 1 0 12600 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1667941163
transform 1 0 16576 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1667941163
transform 1 0 20552 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1667941163
transform 1 0 24528 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1667941163
transform 1 0 28504 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1667941163
transform 1 0 32480 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1667941163
transform 1 0 36456 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1667941163
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1667941163
transform 1 0 6608 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1667941163
transform 1 0 10584 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1667941163
transform 1 0 14560 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1667941163
transform 1 0 18536 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1667941163
transform 1 0 22512 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1667941163
transform 1 0 26488 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1667941163
transform 1 0 30464 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1667941163
transform 1 0 34440 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1667941163
transform 1 0 38416 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1667941163
transform 1 0 4648 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1667941163
transform 1 0 8624 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1667941163
transform 1 0 12600 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1667941163
transform 1 0 16576 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1667941163
transform 1 0 20552 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1667941163
transform 1 0 24528 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1667941163
transform 1 0 28504 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1667941163
transform 1 0 32480 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1667941163
transform 1 0 36456 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1667941163
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1667941163
transform 1 0 6608 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1667941163
transform 1 0 10584 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1667941163
transform 1 0 14560 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1667941163
transform 1 0 18536 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1667941163
transform 1 0 22512 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1667941163
transform 1 0 26488 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1667941163
transform 1 0 30464 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1667941163
transform 1 0 34440 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1667941163
transform 1 0 38416 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1667941163
transform 1 0 4648 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1667941163
transform 1 0 8624 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1667941163
transform 1 0 12600 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1667941163
transform 1 0 16576 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1667941163
transform 1 0 20552 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1667941163
transform 1 0 24528 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1667941163
transform 1 0 28504 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1667941163
transform 1 0 32480 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1667941163
transform 1 0 36456 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1667941163
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1667941163
transform 1 0 4592 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1667941163
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1667941163
transform 1 0 8512 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1667941163
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1667941163
transform 1 0 12432 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1667941163
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1667941163
transform 1 0 16352 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1667941163
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1667941163
transform 1 0 20272 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1667941163
transform 1 0 22232 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1667941163
transform 1 0 24192 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1667941163
transform 1 0 26152 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1667941163
transform 1 0 28112 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1667941163
transform 1 0 30072 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1667941163
transform 1 0 32032 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1667941163
transform 1 0 33992 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1667941163
transform 1 0 35952 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1667941163
transform 1 0 37912 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 21672 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1_
timestamp 1667941163
transform -1 0 21336 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _2_
timestamp 1667941163
transform -1 0 22064 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _3_
timestamp 1667941163
transform -1 0 22064 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _4_
timestamp 1667941163
transform -1 0 22008 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _5_
timestamp 1667941163
transform -1 0 22400 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _6_
timestamp 1667941163
transform -1 0 22400 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  _7_
timestamp 1667941163
transform -1 0 22344 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 22064 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 18256 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 20048 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 20048 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 21504 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 20104 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 16520 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 16912 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 16520 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 15064 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 20104 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 19824 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 20104 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyp1
timestamp 1667941163
transform -1 0 23520 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 18368 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyp1
timestamp 1667941163
transform -1 0 22064 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyp1
timestamp 1667941163
transform -1 0 20048 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 20048 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyp1
timestamp 1667941163
transform -1 0 22064 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 22064 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 20048 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyp1
timestamp 1667941163
transform -1 0 16520 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 20104 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyp1
timestamp 1667941163
transform -1 0 22064 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[16\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[16\].u_series_gyp1
timestamp 1667941163
transform -1 0 16296 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[17\].u_series_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[17\].u_series_gyp1
timestamp 1667941163
transform 1 0 11704 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[18\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[18\].u_series_gyp1
timestamp 1667941163
transform -1 0 20104 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[19\].u_series_gyn1
timestamp 1667941163
transform -1 0 20104 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[19\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[20\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[20\].u_series_gyp1
timestamp 1667941163
transform -1 0 17024 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[21\].u_series_gyn1
timestamp 1667941163
transform -1 0 16520 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[21\].u_series_gyp1
timestamp 1667941163
transform -1 0 19824 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[22\].u_series_gyn1
timestamp 1667941163
transform -1 0 21504 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[22\].u_series_gyp1
timestamp 1667941163
transform -1 0 16520 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[23\].u_series_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[23\].u_series_gyp1
timestamp 1667941163
transform -1 0 20048 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[24\].u_series_gyn1
timestamp 1667941163
transform -1 0 18648 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[24\].u_series_gyp1
timestamp 1667941163
transform -1 0 14504 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[25\].u_series_gyn1
timestamp 1667941163
transform -1 0 17024 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[25\].u_series_gyp1
timestamp 1667941163
transform -1 0 15064 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[26\].u_series_gyn1
timestamp 1667941163
transform -1 0 17024 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[26\].u_series_gyp1
timestamp 1667941163
transform -1 0 16520 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[27\].u_series_gyn1
timestamp 1667941163
transform -1 0 20104 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[27\].u_series_gyp1
timestamp 1667941163
transform -1 0 15064 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[28\].u_series_gyn1
timestamp 1667941163
transform -1 0 17024 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[28\].u_series_gyp1
timestamp 1667941163
transform -1 0 23520 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[29\].u_series_gyn1
timestamp 1667941163
transform -1 0 20048 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[29\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[30\].u_series_gyn1
timestamp 1667941163
transform -1 0 18480 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[30\].u_series_gyp1
timestamp 1667941163
transform -1 0 14504 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[31\].u_series_gyn1
timestamp 1667941163
transform -1 0 17024 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[31\].u_series_gyp1
timestamp 1667941163
transform -1 0 18368 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyp1
timestamp 1667941163
transform 1 0 7728 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 22064 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 22064 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 23520 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 24024 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 14336 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 15064 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 23520 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 25480 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 23520 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[8\].u_series_gyp1
timestamp 1667941163
transform -1 0 26040 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 23520 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 28000 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[10\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 21504 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[11\].u_series_gyp1
timestamp 1667941163
transform 1 0 7728 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[12\].u_series_gyp1
timestamp 1667941163
transform 1 0 7224 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 22064 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 23520 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[14\].u_series_gyp1
timestamp 1667941163
transform -1 0 27496 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 21784 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[15\].u_series_gyp1
timestamp 1667941163
transform -1 0 28000 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyn2
timestamp 1667941163
transform 1 0 5768 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 12544 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyp2
timestamp 1667941163
transform -1 0 26040 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 27496 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyn2
timestamp 1667941163
transform -1 0 27664 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyp1
timestamp 1667941163
transform 1 0 9744 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyp2
timestamp 1667941163
transform 1 0 5208 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyn2
timestamp 1667941163
transform -1 0 29456 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 12376 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyp2
timestamp 1667941163
transform -1 0 29456 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyn2
timestamp 1667941163
transform -1 0 29456 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 25480 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyp2
timestamp 1667941163
transform 1 0 5768 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[4\].u_series_gyn2
timestamp 1667941163
transform -1 0 8568 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 26040 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[4\].u_series_gyp2
timestamp 1667941163
transform 1 0 5208 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 25704 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[5\].u_series_gyn2
timestamp 1667941163
transform -1 0 30016 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 27496 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[5\].u_series_gyp2
timestamp 1667941163
transform -1 0 27496 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[6\].u_series_gyn2
timestamp 1667941163
transform -1 0 8456 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 27496 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[6\].u_series_gyp2
timestamp 1667941163
transform -1 0 30016 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 23744 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[7\].u_series_gyn2
timestamp 1667941163
transform -1 0 25480 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 28000 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[7\].u_series_gyp2
timestamp 1667941163
transform -1 0 28000 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 29624 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyn2
timestamp 1667941163
transform -1 0 4592 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 31584 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyp2
timestamp 1667941163
transform -1 0 5096 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 30016 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyn2
timestamp 1667941163
transform -1 0 4536 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 26040 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyp2
timestamp 1667941163
transform -1 0 29456 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 6496 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[2\].u_series_gyn2
timestamp 1667941163
transform -1 0 28000 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[2\].u_series_gyp1
timestamp 1667941163
transform 1 0 1792 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[2\].u_series_gyp2
timestamp 1667941163
transform -1 0 30016 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 31472 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[3\].u_series_gyn2
timestamp 1667941163
transform 1 0 1232 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[3\].u_series_gyp2
timestamp 1667941163
transform 1 0 1792 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 33432 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 35504 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 35448 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g6\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g6\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 25480 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 10976 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 14336 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 12880 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 14728 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 12880 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 16352 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 15736 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 14448 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 14168 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 12432 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 14616 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 12992 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 14560 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 14336 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 12488 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 12488 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 14896 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 16016 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 14448 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 12432 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 12488 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 13664 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 12208 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 12936 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 13944 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 12992 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 16184 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 12936 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_p
timestamp 1667941163
transform -1 0 11032 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_n
timestamp 1667941163
transform -1 0 16184 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_n
timestamp 1667941163
transform -1 0 14392 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_n
timestamp 1667941163
transform -1 0 14728 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_p
timestamp 1667941163
transform -1 0 14280 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_p
timestamp 1667941163
transform -1 0 12768 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_n1
timestamp 1667941163
transform -1 0 19544 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_n2
timestamp 1667941163
transform -1 0 8568 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_p1
timestamp 1667941163
transform -1 0 22064 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_p2
timestamp 1667941163
transform -1 0 15568 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_n1
timestamp 1667941163
transform -1 0 14112 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_n2
timestamp 1667941163
transform -1 0 6552 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_p1
timestamp 1667941163
transform -1 0 19544 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_p2
timestamp 1667941163
transform -1 0 19544 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_n1
timestamp 1667941163
transform -1 0 17528 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_n2
timestamp 1667941163
transform 1 0 1232 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_p1
timestamp 1667941163
transform -1 0 10528 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_p2
timestamp 1667941163
transform -1 0 7112 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_n1
timestamp 1667941163
transform -1 0 9072 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_n2
timestamp 1667941163
transform -1 0 8568 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_p1
timestamp 1667941163
transform -1 0 19544 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_p2
timestamp 1667941163
transform -1 0 10416 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_n1
timestamp 1667941163
transform -1 0 20048 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_n2
timestamp 1667941163
transform -1 0 14392 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_p1
timestamp 1667941163
transform -1 0 9072 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_p2
timestamp 1667941163
transform -1 0 26040 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_n1
timestamp 1667941163
transform -1 0 15568 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_n2
timestamp 1667941163
transform -1 0 15568 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_p1
timestamp 1667941163
transform -1 0 11088 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_p2
timestamp 1667941163
transform -1 0 14112 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_n1
timestamp 1667941163
transform -1 0 15568 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_n2
timestamp 1667941163
transform -1 0 21504 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_p1
timestamp 1667941163
transform -1 0 6552 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_p2
timestamp 1667941163
transform -1 0 4592 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_n1
timestamp 1667941163
transform -1 0 13328 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_n2
timestamp 1667941163
transform -1 0 20048 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_p1
timestamp 1667941163
transform -1 0 10528 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_p2
timestamp 1667941163
transform -1 0 13496 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_n1
timestamp 1667941163
transform -1 0 7112 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_n2
timestamp 1667941163
transform -1 0 23520 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_p1
timestamp 1667941163
transform -1 0 21504 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_p2
timestamp 1667941163
transform -1 0 6552 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_n1
timestamp 1667941163
transform -1 0 17528 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_n2
timestamp 1667941163
transform -1 0 5096 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_p1
timestamp 1667941163
transform -1 0 6552 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_p2
timestamp 1667941163
transform -1 0 9072 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_n1
timestamp 1667941163
transform -1 0 14224 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_n2
timestamp 1667941163
transform -1 0 17528 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_p1
timestamp 1667941163
transform -1 0 7112 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_p2
timestamp 1667941163
transform -1 0 8568 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_n1
timestamp 1667941163
transform -1 0 8568 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_n2
timestamp 1667941163
transform 1 0 1792 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_p1
timestamp 1667941163
transform -1 0 20048 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_p2
timestamp 1667941163
transform 1 0 1232 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_n1
timestamp 1667941163
transform -1 0 17528 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_n2
timestamp 1667941163
transform -1 0 7112 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_p1
timestamp 1667941163
transform -1 0 20048 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_p2
timestamp 1667941163
transform -1 0 25480 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_n1
timestamp 1667941163
transform -1 0 13328 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_n2
timestamp 1667941163
transform -1 0 13552 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_p1
timestamp 1667941163
transform 1 0 3248 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_p2
timestamp 1667941163
transform -1 0 24024 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_n1
timestamp 1667941163
transform -1 0 14112 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_n2
timestamp 1667941163
transform -1 0 16072 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_p1
timestamp 1667941163
transform -1 0 16072 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_p2
timestamp 1667941163
transform -1 0 5096 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_n1
timestamp 1667941163
transform -1 0 16072 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_n2
timestamp 1667941163
transform -1 0 23520 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_p1
timestamp 1667941163
transform -1 0 8568 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_p2
timestamp 1667941163
transform -1 0 23520 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_n1
timestamp 1667941163
transform -1 0 10528 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_n2
timestamp 1667941163
transform -1 0 22064 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_p1
timestamp 1667941163
transform -1 0 9072 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_p2
timestamp 1667941163
transform -1 0 4592 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_n1
timestamp 1667941163
transform -1 0 10528 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_n2
timestamp 1667941163
transform -1 0 6552 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_p1
timestamp 1667941163
transform -1 0 8568 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_p2
timestamp 1667941163
transform -1 0 6552 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_n1
timestamp 1667941163
transform -1 0 18088 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_n2
timestamp 1667941163
transform -1 0 17528 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_p1
timestamp 1667941163
transform -1 0 20048 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_p2
timestamp 1667941163
transform 1 0 1792 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_n1
timestamp 1667941163
transform -1 0 16072 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_n2
timestamp 1667941163
transform -1 0 18088 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_p1
timestamp 1667941163
transform -1 0 11088 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_p2
timestamp 1667941163
transform 1 0 1232 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_n1
timestamp 1667941163
transform -1 0 19544 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_n2
timestamp 1667941163
transform -1 0 7112 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_p1
timestamp 1667941163
transform -1 0 15568 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_p2
timestamp 1667941163
transform 1 0 1792 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_n1
timestamp 1667941163
transform -1 0 12544 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_n2
timestamp 1667941163
transform -1 0 4592 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_p1
timestamp 1667941163
transform 1 0 3752 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_p2
timestamp 1667941163
transform -1 0 5096 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_n1
timestamp 1667941163
transform -1 0 20048 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_n2
timestamp 1667941163
transform -1 0 18088 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_p1
timestamp 1667941163
transform -1 0 21504 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_p2
timestamp 1667941163
transform -1 0 25480 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_n1
timestamp 1667941163
transform -1 0 9072 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_n2
timestamp 1667941163
transform -1 0 6552 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_p1
timestamp 1667941163
transform -1 0 12544 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_p2
timestamp 1667941163
transform -1 0 25480 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_n1
timestamp 1667941163
transform -1 0 12544 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_n2
timestamp 1667941163
transform -1 0 5096 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_p1
timestamp 1667941163
transform -1 0 22064 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_p2
timestamp 1667941163
transform -1 0 7112 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_n1
timestamp 1667941163
transform -1 0 14112 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_n2
timestamp 1667941163
transform -1 0 4592 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_p1
timestamp 1667941163
transform -1 0 13496 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_p2
timestamp 1667941163
transform -1 0 26040 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_n1
timestamp 1667941163
transform -1 0 8568 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_n2
timestamp 1667941163
transform -1 0 14112 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_p1
timestamp 1667941163
transform -1 0 13048 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_p2
timestamp 1667941163
transform -1 0 23520 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_n1
timestamp 1667941163
transform -1 0 19544 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_n2
timestamp 1667941163
transform -1 0 19544 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_p1
timestamp 1667941163
transform -1 0 21504 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_p2
timestamp 1667941163
transform -1 0 24024 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_n1
timestamp 1667941163
transform -1 0 18088 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_n2
timestamp 1667941163
transform -1 0 9072 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_p1
timestamp 1667941163
transform 1 0 3752 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_p2
timestamp 1667941163
transform -1 0 20048 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_n1
timestamp 1667941163
transform -1 0 11088 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_n2
timestamp 1667941163
transform 1 0 1792 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_p1
timestamp 1667941163
transform -1 0 12544 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_p2
timestamp 1667941163
transform -1 0 24024 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_n1
timestamp 1667941163
transform -1 0 10976 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_n2
timestamp 1667941163
transform -1 0 7112 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_p1
timestamp 1667941163
transform -1 0 21504 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_p2
timestamp 1667941163
transform -1 0 5096 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_n1
timestamp 1667941163
transform -1 0 18088 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_n2
timestamp 1667941163
transform -1 0 24024 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_p1
timestamp 1667941163
transform -1 0 22064 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_p2
timestamp 1667941163
transform -1 0 4592 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_n1
timestamp 1667941163
transform -1 0 16072 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_n2
timestamp 1667941163
transform 1 0 1232 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_p1
timestamp 1667941163
transform -1 0 4592 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_p2
timestamp 1667941163
transform -1 0 28000 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_n1
timestamp 1667941163
transform -1 0 10920 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_n2
timestamp 1667941163
transform -1 0 4592 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_p1
timestamp 1667941163
transform 1 0 1792 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_p2
timestamp 1667941163
transform -1 0 23520 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_n1
timestamp 1667941163
transform -1 0 8568 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_n2
timestamp 1667941163
transform -1 0 6552 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_p1
timestamp 1667941163
transform 1 0 1232 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_p2
timestamp 1667941163
transform -1 0 20048 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_n1
timestamp 1667941163
transform 1 0 1232 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_n2
timestamp 1667941163
transform -1 0 7112 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_p1
timestamp 1667941163
transform -1 0 5096 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_p2
timestamp 1667941163
transform -1 0 25480 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_n1
timestamp 1667941163
transform -1 0 10528 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_n2
timestamp 1667941163
transform -1 0 5096 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_p1
timestamp 1667941163
transform 1 0 1792 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_p2
timestamp 1667941163
transform -1 0 24024 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_n1
timestamp 1667941163
transform -1 0 21504 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_n2
timestamp 1667941163
transform -1 0 17528 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_p1
timestamp 1667941163
transform 1 0 1232 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_p2
timestamp 1667941163
transform -1 0 27496 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_n1
timestamp 1667941163
transform -1 0 7112 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_n2
timestamp 1667941163
transform -1 0 8568 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_p1
timestamp 1667941163
transform 1 0 1792 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_p2
timestamp 1667941163
transform -1 0 6552 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_n1
timestamp 1667941163
transform -1 0 22064 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_n2
timestamp 1667941163
transform -1 0 6552 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_p1
timestamp 1667941163
transform 1 0 1232 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_p2
timestamp 1667941163
transform -1 0 17528 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_n1
timestamp 1667941163
transform -1 0 12376 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_n2
timestamp 1667941163
transform 1 0 1792 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_p1
timestamp 1667941163
transform -1 0 5096 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_p2
timestamp 1667941163
transform 1 0 1232 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_n1
timestamp 1667941163
transform -1 0 9072 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_n2
timestamp 1667941163
transform -1 0 18088 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_p1
timestamp 1667941163
transform -1 0 4592 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_p2
timestamp 1667941163
transform -1 0 26040 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_n1
timestamp 1667941163
transform 1 0 1792 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_n2
timestamp 1667941163
transform -1 0 27496 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_p1
timestamp 1667941163
transform -1 0 4592 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_p2
timestamp 1667941163
transform 1 0 1792 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_n1
timestamp 1667941163
transform 1 0 1232 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_n2
timestamp 1667941163
transform 1 0 1232 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_p1
timestamp 1667941163
transform 1 0 1792 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_p2
timestamp 1667941163
transform -1 0 24024 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_n1
timestamp 1667941163
transform -1 0 5096 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_n2
timestamp 1667941163
transform -1 0 4592 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_p1
timestamp 1667941163
transform 1 0 1792 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_p2
timestamp 1667941163
transform -1 0 21504 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_n1
timestamp 1667941163
transform -1 0 8568 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_n2
timestamp 1667941163
transform -1 0 7112 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_p1
timestamp 1667941163
transform 1 0 1232 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_p2
timestamp 1667941163
transform -1 0 19544 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_n1
timestamp 1667941163
transform -1 0 4592 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_n2
timestamp 1667941163
transform -1 0 5096 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_p1
timestamp 1667941163
transform 1 0 1232 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_p2
timestamp 1667941163
transform -1 0 22064 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_n1
timestamp 1667941163
transform -1 0 6552 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_n2
timestamp 1667941163
transform -1 0 7112 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_p1
timestamp 1667941163
transform 1 0 1792 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_p2
timestamp 1667941163
transform -1 0 23520 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_n1
timestamp 1667941163
transform -1 0 5096 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_n2
timestamp 1667941163
transform -1 0 23520 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_p1
timestamp 1667941163
transform -1 0 20048 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_p2
timestamp 1667941163
transform -1 0 26040 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_n1
timestamp 1667941163
transform -1 0 4592 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_n2
timestamp 1667941163
transform -1 0 24024 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_p1
timestamp 1667941163
transform -1 0 21504 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_p2
timestamp 1667941163
transform -1 0 27496 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_n1
timestamp 1667941163
transform 1 0 1792 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_n2
timestamp 1667941163
transform -1 0 22064 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_p1
timestamp 1667941163
transform -1 0 22064 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_p2
timestamp 1667941163
transform -1 0 28000 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_n1
timestamp 1667941163
transform 1 0 1232 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_n2
timestamp 1667941163
transform -1 0 25480 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_p1
timestamp 1667941163
transform -1 0 23520 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_p2
timestamp 1667941163
transform -1 0 26040 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_n1
timestamp 1667941163
transform 1 0 1232 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_n2
timestamp 1667941163
transform -1 0 26040 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_p1
timestamp 1667941163
transform -1 0 24024 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_p2
timestamp 1667941163
transform -1 0 25480 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_n1
timestamp 1667941163
transform 1 0 1792 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_n2
timestamp 1667941163
transform -1 0 24024 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_p1
timestamp 1667941163
transform -1 0 20048 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_p2
timestamp 1667941163
transform -1 0 26040 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_n1
timestamp 1667941163
transform 1 0 1232 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_n2
timestamp 1667941163
transform -1 0 23520 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_p1
timestamp 1667941163
transform -1 0 26040 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_p2
timestamp 1667941163
transform -1 0 24024 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_n1
timestamp 1667941163
transform -1 0 19544 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_n2
timestamp 1667941163
transform -1 0 25480 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_p1
timestamp 1667941163
transform -1 0 21504 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_p2
timestamp 1667941163
transform -1 0 25480 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 33992 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 37408 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 35952 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 33432 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 35448 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 33992 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 33432 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 37968 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_n1
timestamp 1667941163
transform -1 0 37408 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_n2
timestamp 1667941163
transform -1 0 37968 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_p1
timestamp 1667941163
transform -1 0 35448 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_p2
timestamp 1667941163
transform -1 0 35952 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_n1
timestamp 1667941163
transform -1 0 37968 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_n2
timestamp 1667941163
transform -1 0 37408 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_p1
timestamp 1667941163
transform -1 0 35952 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_p2
timestamp 1667941163
transform -1 0 37408 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 37968 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 36008 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 28000 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33992 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 38640 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 37968 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 36008 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 28000 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 30408 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 30408 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 28000 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 37968 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 30408 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 37968 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 38528 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 36008 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 37968 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 36008 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 36008 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 38528 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 36008 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33992 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 38528 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 33992 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 30408 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 39032 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 38640 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 33544 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 38528 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 38528 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 38584 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 38640 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 38584 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 37968 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 38640 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 38640 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 36008 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 39032 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_p
timestamp 1667941163
transform 1 0 28000 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_series_gygyn1
timestamp 1667941163
transform -1 0 30408 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_series_gygyn2
timestamp 1667941163
transform -1 0 35448 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_series_gygyp1
timestamp 1667941163
transform -1 0 32032 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31976 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37408 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_series_gygyn2
timestamp 1667941163
transform -1 0 30408 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35448 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30408 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37408 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_series_gygyn2
timestamp 1667941163
transform -1 0 30576 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_series_gygyp1
timestamp 1667941163
transform -1 0 33992 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31976 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37408 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33992 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35952 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31472 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_series_gygyn1
timestamp 1667941163
transform -1 0 35952 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_series_gygyn2
timestamp 1667941163
transform -1 0 31920 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35448 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31976 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37968 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33432 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_series_gygyp1
timestamp 1667941163
transform -1 0 37408 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30464 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_series_gygyn1
timestamp 1667941163
transform -1 0 30632 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_series_gygyn2
timestamp 1667941163
transform 1 0 27608 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35952 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30408 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37968 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_series_gygyn2
timestamp 1667941163
transform 1 0 27104 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35952 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30464 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[8\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37968 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[8\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33432 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[8\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35952 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[8\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31920 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[9\].u_series_gygyn1
timestamp 1667941163
transform -1 0 35952 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[9\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33992 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[9\].u_series_gygyp1
timestamp 1667941163
transform -1 0 30408 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[9\].u_series_gygyp2
timestamp 1667941163
transform 1 0 27608 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[10\].u_series_gygyn1
timestamp 1667941163
transform -1 0 31976 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[10\].u_series_gygyn2
timestamp 1667941163
transform -1 0 31920 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[10\].u_series_gygyp1
timestamp 1667941163
transform -1 0 33432 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[10\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30464 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[11\].u_series_gygyn1
timestamp 1667941163
transform -1 0 33432 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[11\].u_series_gygyn2
timestamp 1667941163
transform -1 0 31976 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[11\].u_series_gygyp1
timestamp 1667941163
transform -1 0 31976 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[11\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30408 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[12\].u_series_gygyn1
timestamp 1667941163
transform -1 0 31976 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[12\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33432 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[12\].u_series_gygyp1
timestamp 1667941163
transform -1 0 33992 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[12\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30464 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[13\].u_series_gygyn1
timestamp 1667941163
transform -1 0 33992 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[13\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33432 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[13\].u_series_gygyp1
timestamp 1667941163
transform -1 0 30520 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[13\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31920 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[14\].u_series_gygyn1
timestamp 1667941163
transform 1 0 27608 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[14\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33992 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[14\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35448 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[14\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31976 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[15\].u_series_gygyn1
timestamp 1667941163
transform -1 0 35448 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[15\].u_series_gygyn2
timestamp 1667941163
transform -1 0 31976 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[15\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35448 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[15\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31472 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_series_gygyn1
timestamp 1667941163
transform -1 0 33992 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_series_gygyn2
timestamp 1667941163
transform -1 0 31528 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_series_gygyp1
timestamp 1667941163
transform -1 0 31976 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_series_gygyp2
timestamp 1667941163
transform -1 0 37968 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_series_gygyn1
timestamp 1667941163
transform -1 0 31976 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33992 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_series_gygyp1
timestamp 1667941163
transform -1 0 37968 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30072 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37408 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_series_gygyn2
timestamp 1667941163
transform -1 0 35448 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_series_gygyp1
timestamp 1667941163
transform -1 0 37408 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_series_gygyp2
timestamp 1667941163
transform 1 0 27608 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37968 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_series_gygyn2
timestamp 1667941163
transform -1 0 35952 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_series_gygyp1
timestamp 1667941163
transform 1 0 29120 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30072 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[4\].u_series_gygyn1
timestamp 1667941163
transform 1 0 29064 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[4\].u_series_gygyn2
timestamp 1667941163
transform -1 0 30128 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[4\].u_series_gygyp1
timestamp 1667941163
transform -1 0 31584 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[4\].u_series_gygyp2
timestamp 1667941163
transform -1 0 30072 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[5\].u_series_gygyn1
timestamp 1667941163
transform -1 0 35448 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[5\].u_series_gygyn2
timestamp 1667941163
transform -1 0 31976 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[5\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35448 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[5\].u_series_gygyp2
timestamp 1667941163
transform 1 0 27104 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[6\].u_series_gygyn1
timestamp 1667941163
transform -1 0 35952 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[6\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33432 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[6\].u_series_gygyp1
timestamp 1667941163
transform -1 0 33432 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[6\].u_series_gygyp2
timestamp 1667941163
transform -1 0 32088 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[7\].u_series_gygyn1
timestamp 1667941163
transform -1 0 31920 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[7\].u_series_gygyn2
timestamp 1667941163
transform 1 0 27272 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[7\].u_series_gygyp1
timestamp 1667941163
transform -1 0 35952 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[7\].u_series_gygyp2
timestamp 1667941163
transform -1 0 33432 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37408 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_series_gygyp1
timestamp 1667941163
transform -1 0 29512 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37968 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_series_gygyp1
timestamp 1667941163
transform -1 0 28448 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[2\].u_series_gygyn1
timestamp 1667941163
transform -1 0 28448 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[2\].u_series_gygyp1
timestamp 1667941163
transform -1 0 28616 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[3\].u_series_gygyn1
timestamp 1667941163
transform -1 0 33992 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[3\].u_series_gygyp1
timestamp 1667941163
transform 1 0 25648 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[0\].u_series_gygyn1
timestamp 1667941163
transform -1 0 37968 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[0\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33432 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[0\].u_series_gygyp1
timestamp 1667941163
transform -1 0 37464 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[0\].u_series_gygyp2
timestamp 1667941163
transform -1 0 31976 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[1\].u_series_gygyn1
timestamp 1667941163
transform -1 0 28056 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[1\].u_series_gygyn2
timestamp 1667941163
transform -1 0 33992 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[1\].u_series_gygyp1
timestamp 1667941163
transform -1 0 37408 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g4\[1\].u_series_gygyp2
timestamp 1667941163
transform -1 0 33544 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g5\[0\].u_series_gygyn1
timestamp 1667941163
transform -1 0 27496 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g5\[0\].u_series_gygyp1
timestamp 1667941163
transform -1 0 31976 0 1 2352
box -43 -43 1387 435
<< labels >>
flabel metal2 s 37408 19600 37464 20000 0 FreeSans 224 90 0 0 cap_series_gygyn
port 0 nsew signal bidirectional
flabel metal2 s 32424 19600 32480 20000 0 FreeSans 224 90 0 0 cap_series_gygyp
port 1 nsew signal bidirectional
flabel metal2 s 27440 19600 27496 20000 0 FreeSans 224 90 0 0 cap_series_gyn
port 2 nsew signal bidirectional
flabel metal2 s 22456 19600 22512 20000 0 FreeSans 224 90 0 0 cap_series_gyp
port 3 nsew signal bidirectional
flabel metal2 s 17472 19600 17528 20000 0 FreeSans 224 90 0 0 cap_shunt_gyn
port 4 nsew signal bidirectional
flabel metal2 s 12488 19600 12544 20000 0 FreeSans 224 90 0 0 cap_shunt_gyp
port 5 nsew signal bidirectional
flabel metal2 s 7504 19600 7560 20000 0 FreeSans 224 90 0 0 cap_shunt_n
port 6 nsew signal bidirectional
flabel metal2 s 2520 19600 2576 20000 0 FreeSans 224 90 0 0 cap_shunt_p
port 7 nsew signal bidirectional
flabel metal2 s 14392 0 14448 400 0 FreeSans 224 90 0 0 tune_series_gy[0]
port 8 nsew signal input
flabel metal2 s 15624 0 15680 400 0 FreeSans 224 90 0 0 tune_series_gy[1]
port 9 nsew signal input
flabel metal2 s 16856 0 16912 400 0 FreeSans 224 90 0 0 tune_series_gy[2]
port 10 nsew signal input
flabel metal2 s 18088 0 18144 400 0 FreeSans 224 90 0 0 tune_series_gy[3]
port 11 nsew signal input
flabel metal2 s 19320 0 19376 400 0 FreeSans 224 90 0 0 tune_series_gy[4]
port 12 nsew signal input
flabel metal2 s 20552 0 20608 400 0 FreeSans 224 90 0 0 tune_series_gy[5]
port 13 nsew signal input
flabel metal2 s 21784 0 21840 400 0 FreeSans 224 90 0 0 tune_series_gy[6]
port 14 nsew signal input
flabel metal2 s 23016 0 23072 400 0 FreeSans 224 90 0 0 tune_series_gy[7]
port 15 nsew signal input
flabel metal2 s 24248 0 24304 400 0 FreeSans 224 90 0 0 tune_series_gygy[0]
port 16 nsew signal input
flabel metal2 s 25480 0 25536 400 0 FreeSans 224 90 0 0 tune_series_gygy[1]
port 17 nsew signal input
flabel metal2 s 26712 0 26768 400 0 FreeSans 224 90 0 0 tune_series_gygy[2]
port 18 nsew signal input
flabel metal2 s 27944 0 28000 400 0 FreeSans 224 90 0 0 tune_series_gygy[3]
port 19 nsew signal input
flabel metal2 s 29176 0 29232 400 0 FreeSans 224 90 0 0 tune_series_gygy[4]
port 20 nsew signal input
flabel metal2 s 30408 0 30464 400 0 FreeSans 224 90 0 0 tune_series_gygy[5]
port 21 nsew signal input
flabel metal2 s 31640 0 31696 400 0 FreeSans 224 90 0 0 tune_series_gygy[6]
port 22 nsew signal input
flabel metal2 s 32872 0 32928 400 0 FreeSans 224 90 0 0 tune_series_gygy[7]
port 23 nsew signal input
flabel metal2 s 840 0 896 400 0 FreeSans 224 90 0 0 tune_shunt[0]
port 24 nsew signal input
flabel metal2 s 13160 0 13216 400 0 FreeSans 224 90 0 0 tune_shunt[10]
port 25 nsew signal input
flabel metal2 s 2072 0 2128 400 0 FreeSans 224 90 0 0 tune_shunt[1]
port 26 nsew signal input
flabel metal2 s 3304 0 3360 400 0 FreeSans 224 90 0 0 tune_shunt[2]
port 27 nsew signal input
flabel metal2 s 4536 0 4592 400 0 FreeSans 224 90 0 0 tune_shunt[3]
port 28 nsew signal input
flabel metal2 s 5768 0 5824 400 0 FreeSans 224 90 0 0 tune_shunt[4]
port 29 nsew signal input
flabel metal2 s 7000 0 7056 400 0 FreeSans 224 90 0 0 tune_shunt[5]
port 30 nsew signal input
flabel metal2 s 8232 0 8288 400 0 FreeSans 224 90 0 0 tune_shunt[6]
port 31 nsew signal input
flabel metal2 s 9464 0 9520 400 0 FreeSans 224 90 0 0 tune_shunt[7]
port 32 nsew signal input
flabel metal2 s 10696 0 10752 400 0 FreeSans 224 90 0 0 tune_shunt[8]
port 33 nsew signal input
flabel metal2 s 11928 0 11984 400 0 FreeSans 224 90 0 0 tune_shunt[9]
port 34 nsew signal input
flabel metal2 s 34104 0 34160 400 0 FreeSans 224 90 0 0 tune_shunt_gy[0]
port 35 nsew signal input
flabel metal2 s 35336 0 35392 400 0 FreeSans 224 90 0 0 tune_shunt_gy[1]
port 36 nsew signal input
flabel metal2 s 36568 0 36624 400 0 FreeSans 224 90 0 0 tune_shunt_gy[2]
port 37 nsew signal input
flabel metal2 s 37800 0 37856 400 0 FreeSans 224 90 0 0 tune_shunt_gy[3]
port 38 nsew signal input
flabel metal2 s 39032 0 39088 400 0 FreeSans 224 90 0 0 tune_shunt_gy[4]
port 39 nsew signal input
flabel metal4 s 2054 1538 2554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 7054 1538 7554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 12054 1538 12554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 17054 1538 17554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 22054 1538 22554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 27054 1538 27554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 32054 1538 32554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 37054 1538 37554 18454 0 FreeSans 2560 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 4554 1538 5054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 9554 1538 10054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 14554 1538 15054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 19554 1538 20054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 24554 1538 25054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 29554 1538 30054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 34554 1538 35054 18454 0 FreeSans 2560 90 0 0 vss
port 41 nsew ground bidirectional
rlabel metal1 19992 18424 19992 18424 0 vdd
rlabel metal1 19992 18032 19992 18032 0 vss
rlabel metal2 27412 6104 27412 6104 0 cap_series_gygyn
rlabel metal2 35868 8008 35868 8008 0 cap_series_gygyp
rlabel metal2 1652 2380 1652 2380 0 cap_series_gyn
rlabel metal2 2380 2352 2380 2352 0 cap_series_gyp
rlabel metal2 33684 8036 33684 8036 0 cap_shunt_gyn
rlabel metal2 12628 17528 12628 17528 0 cap_shunt_gyp
rlabel metal2 1372 3304 1372 3304 0 cap_shunt_n
rlabel metal2 2492 3668 2492 3668 0 cap_shunt_p
rlabel metal2 14420 1687 14420 1687 0 tune_series_gy[0]
rlabel metal2 15652 931 15652 931 0 tune_series_gy[1]
rlabel metal2 4060 2576 4060 2576 0 tune_series_gy[2]
rlabel metal2 24388 2352 24388 2352 0 tune_series_gy[3]
rlabel metal2 26404 1736 26404 1736 0 tune_series_gy[4]
rlabel metal2 11396 1792 11396 1792 0 tune_series_gy[5]
rlabel metal2 13076 1988 13076 1988 0 tune_series_gy[6]
rlabel metal3 13104 4116 13104 4116 0 tune_series_gy[7]
rlabel metal3 25228 3388 25228 3388 0 tune_series_gygy[0]
rlabel metal2 30716 2940 30716 2940 0 tune_series_gygy[1]
rlabel metal2 36148 2408 36148 2408 0 tune_series_gygy[2]
rlabel metal2 32844 9184 32844 9184 0 tune_series_gygy[3]
rlabel metal2 34412 8036 34412 8036 0 tune_series_gygy[4]
rlabel metal2 34188 9324 34188 9324 0 tune_series_gygy[5]
rlabel metal3 30996 3360 30996 3360 0 tune_series_gygy[6]
rlabel metal3 32816 7588 32816 7588 0 tune_series_gygy[7]
rlabel metal2 1204 2212 1204 2212 0 tune_shunt[0]
rlabel metal2 3724 11172 3724 11172 0 tune_shunt[10]
rlabel metal2 2100 1127 2100 1127 0 tune_shunt[1]
rlabel metal2 3332 1127 3332 1127 0 tune_shunt[2]
rlabel metal2 10556 5040 10556 5040 0 tune_shunt[3]
rlabel metal2 25088 13916 25088 13916 0 tune_shunt[4]
rlabel metal2 3724 14700 3724 14700 0 tune_shunt[5]
rlabel metal2 2492 3080 2492 3080 0 tune_shunt[6]
rlabel metal2 4116 2884 4116 2884 0 tune_shunt[7]
rlabel metal2 10724 1071 10724 1071 0 tune_shunt[8]
rlabel metal2 12236 2296 12236 2296 0 tune_shunt[9]
rlabel metal2 28364 2128 28364 2128 0 tune_shunt_gy[0]
rlabel metal2 35700 6300 35700 6300 0 tune_shunt_gy[1]
rlabel metal2 33936 7980 33936 7980 0 tune_shunt_gy[2]
rlabel metal3 29176 4844 29176 4844 0 tune_shunt_gy[3]
rlabel metal2 30100 2912 30100 2912 0 tune_shunt_gy[4]
<< properties >>
string FIXED_BBOX 0 0 40000 20000
<< end >>
