// This is the unpowered netlist.
module dlc (clk,
    clko,
    latch,
    on,
    op,
    rst,
    sdi,
    sig);
 input clk;
 output clko;
 input latch;
 output on;
 output op;
 input rst;
 input sdi;
 input sig;

 wire \trim_n[0] ;
 wire \trim_n[1] ;
 wire \trim_n[2] ;
 wire \trim_n[3] ;
 wire \trim_p[0] ;
 wire \trim_p[1] ;
 wire \trim_p[2] ;
 wire \trim_p[3] ;
 wire \u_trans0p.outn ;
 wire \u_trans0p.outp ;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0_ (.I(clk),
    .ZN(clko));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1_ (.ZN(\trim_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2_ (.ZN(\trim_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3_ (.ZN(\trim_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _4_ (.ZN(\trim_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _5_ (.ZN(\trim_p[0] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _6_ (.ZN(\trim_p[1] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _7_ (.ZN(\trim_p[2] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8_ (.ZN(\trim_p[3] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[0].fbn  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[0].fbp  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[1].fbn  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[1].fbp  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[2].fbn  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[2].fbp  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[3].fbn  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_FB[3].fbp  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[0].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[0].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[1].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[1].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[2].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[2].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[3].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[3].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[4].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[4].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[5].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[5].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[6].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[6].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[7].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[7].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[8].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[8].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[9].thrun  (.I(sdi),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_T[9].thrup  (.I(sig),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[0].crossn  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[0].crossp  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[1].crossn  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[1].crossp  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[2].crossn  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[2].crossp  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[3].crossn  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[3].crossp  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[4].crossn  (.I(\u_trans0p.outp ),
    .ZN(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans0p.gen_X[4].crossp  (.I(\u_trans0p.outn ),
    .ZN(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[0].fbn  (.I(on),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[0].fbp  (.I(op),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[1].fbn  (.I(on),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[1].fbp  (.I(op),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[2].fbn  (.I(on),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[2].fbp  (.I(op),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[3].fbn  (.I(on),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_FB[3].fbp  (.I(op),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[0].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[0].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[1].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[1].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[2].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[2].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[3].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[3].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[4].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[4].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[5].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[5].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[6].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[6].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[7].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[7].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[8].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[8].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[9].thrun  (.I(\u_trans0p.outp ),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_T[9].thrup  (.I(\u_trans0p.outn ),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[0].crossn  (.I(op),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[0].crossp  (.I(on),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[1].crossn  (.I(op),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[1].crossp  (.I(on),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[2].crossn  (.I(op),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[2].crossp  (.I(on),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[3].crossn  (.I(op),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[3].crossp  (.I(on),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[4].crossn  (.I(op),
    .ZN(on));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_trans1p.gen_X[4].crossp  (.I(on),
    .ZN(op));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0__I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[4].crossp_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[3].crossp_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[2].crossp_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[1].crossp_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[0].crossp_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[3].fbn_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[2].fbn_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[1].fbn_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[0].fbn_I  (.I(on));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[4].crossn_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[3].crossn_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[2].crossn_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[1].crossn_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_X[0].crossn_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[3].fbp_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[2].fbp_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[1].fbp_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_FB[0].fbp_I  (.I(op));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[9].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[8].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[7].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[6].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[5].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[4].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[3].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[2].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[1].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[0].thrun_I  (.I(sdi));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[9].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[8].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[7].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[6].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[5].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[4].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[3].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[2].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[1].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_T[0].thrup_I  (.I(sig));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[9].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[8].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[7].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[6].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[5].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[4].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[3].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[2].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[1].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[0].thrup_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[4].crossp_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[3].crossp_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[2].crossp_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[1].crossp_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[0].crossp_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[3].fbn_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[2].fbn_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[1].fbn_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[0].fbn_I  (.I(\u_trans0p.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[9].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[8].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[7].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[6].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[5].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[4].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[3].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[2].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[1].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans1p.gen_T[0].thrun_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[4].crossn_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[3].crossn_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[2].crossn_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[1].crossn_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_X[0].crossn_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[3].fbp_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[2].fbp_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[1].fbp_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_trans0p.gen_FB[0].fbp_I  (.I(\u_trans0p.outp ));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_329 ();
endmodule

