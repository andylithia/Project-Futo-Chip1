magic
tech gf180mcuC
magscale 1 10
timestamp 1669676130
<< metal1 >>
rect 1344 16490 178640 16524
rect 1344 16438 23376 16490
rect 23428 16438 23480 16490
rect 23532 16438 23584 16490
rect 23636 16438 67700 16490
rect 67752 16438 67804 16490
rect 67856 16438 67908 16490
rect 67960 16438 112024 16490
rect 112076 16438 112128 16490
rect 112180 16438 112232 16490
rect 112284 16438 156348 16490
rect 156400 16438 156452 16490
rect 156504 16438 156556 16490
rect 156608 16438 178640 16490
rect 1344 16404 178640 16438
rect 3166 15986 3218 15998
rect 3166 15922 3218 15934
rect 4734 15986 4786 15998
rect 4734 15922 4786 15934
rect 7870 15986 7922 15998
rect 7870 15922 7922 15934
rect 9662 15986 9714 15998
rect 9662 15922 9714 15934
rect 12574 15986 12626 15998
rect 12574 15922 12626 15934
rect 14142 15986 14194 15998
rect 14142 15922 14194 15934
rect 17502 15986 17554 15998
rect 17502 15922 17554 15934
rect 18846 15986 18898 15998
rect 18846 15922 18898 15934
rect 21982 15986 22034 15998
rect 21982 15922 22034 15934
rect 23550 15986 23602 15998
rect 23550 15922 23602 15934
rect 26686 15986 26738 15998
rect 26686 15922 26738 15934
rect 28254 15986 28306 15998
rect 28254 15922 28306 15934
rect 31390 15986 31442 15998
rect 31390 15922 31442 15934
rect 33182 15986 33234 15998
rect 33182 15922 33234 15934
rect 36094 15986 36146 15998
rect 36094 15922 36146 15934
rect 37662 15986 37714 15998
rect 37662 15922 37714 15934
rect 41022 15986 41074 15998
rect 41022 15922 41074 15934
rect 42366 15986 42418 15998
rect 42366 15922 42418 15934
rect 45502 15986 45554 15998
rect 45502 15922 45554 15934
rect 47070 15986 47122 15998
rect 47070 15922 47122 15934
rect 50206 15986 50258 15998
rect 50206 15922 50258 15934
rect 51774 15986 51826 15998
rect 51774 15922 51826 15934
rect 54910 15986 54962 15998
rect 54910 15922 54962 15934
rect 56702 15986 56754 15998
rect 56702 15922 56754 15934
rect 59614 15986 59666 15998
rect 59614 15922 59666 15934
rect 61182 15986 61234 15998
rect 61182 15922 61234 15934
rect 64542 15986 64594 15998
rect 64542 15922 64594 15934
rect 65886 15986 65938 15998
rect 65886 15922 65938 15934
rect 69022 15986 69074 15998
rect 69022 15922 69074 15934
rect 70590 15986 70642 15998
rect 70590 15922 70642 15934
rect 73726 15986 73778 15998
rect 73726 15922 73778 15934
rect 75294 15986 75346 15998
rect 75294 15922 75346 15934
rect 78430 15986 78482 15998
rect 78430 15922 78482 15934
rect 80222 15986 80274 15998
rect 80222 15922 80274 15934
rect 83134 15986 83186 15998
rect 83134 15922 83186 15934
rect 84702 15986 84754 15998
rect 84702 15922 84754 15934
rect 88062 15986 88114 15998
rect 88062 15922 88114 15934
rect 89406 15986 89458 15998
rect 89406 15922 89458 15934
rect 92542 15986 92594 15998
rect 92542 15922 92594 15934
rect 94110 15986 94162 15998
rect 94110 15922 94162 15934
rect 97246 15986 97298 15998
rect 97246 15922 97298 15934
rect 98814 15986 98866 15998
rect 98814 15922 98866 15934
rect 101950 15986 102002 15998
rect 101950 15922 102002 15934
rect 103742 15986 103794 15998
rect 103742 15922 103794 15934
rect 106654 15986 106706 15998
rect 106654 15922 106706 15934
rect 108222 15986 108274 15998
rect 108222 15922 108274 15934
rect 111582 15986 111634 15998
rect 111582 15922 111634 15934
rect 112926 15986 112978 15998
rect 112926 15922 112978 15934
rect 116062 15986 116114 15998
rect 116062 15922 116114 15934
rect 117630 15986 117682 15998
rect 117630 15922 117682 15934
rect 120766 15986 120818 15998
rect 120766 15922 120818 15934
rect 122334 15986 122386 15998
rect 122334 15922 122386 15934
rect 125470 15986 125522 15998
rect 125470 15922 125522 15934
rect 127262 15986 127314 15998
rect 127262 15922 127314 15934
rect 130174 15986 130226 15998
rect 130174 15922 130226 15934
rect 131742 15986 131794 15998
rect 131742 15922 131794 15934
rect 135102 15986 135154 15998
rect 135102 15922 135154 15934
rect 136446 15986 136498 15998
rect 136446 15922 136498 15934
rect 139582 15986 139634 15998
rect 139582 15922 139634 15934
rect 141150 15986 141202 15998
rect 141150 15922 141202 15934
rect 144286 15986 144338 15998
rect 144286 15922 144338 15934
rect 145854 15986 145906 15998
rect 145854 15922 145906 15934
rect 148990 15986 149042 15998
rect 148990 15922 149042 15934
rect 150782 15986 150834 15998
rect 150782 15922 150834 15934
rect 153694 15986 153746 15998
rect 153694 15922 153746 15934
rect 155262 15986 155314 15998
rect 155262 15922 155314 15934
rect 158622 15986 158674 15998
rect 158622 15922 158674 15934
rect 159966 15986 160018 15998
rect 159966 15922 160018 15934
rect 163102 15986 163154 15998
rect 163102 15922 163154 15934
rect 164670 15986 164722 15998
rect 164670 15922 164722 15934
rect 167806 15986 167858 15998
rect 167806 15922 167858 15934
rect 169374 15986 169426 15998
rect 169374 15922 169426 15934
rect 172510 15986 172562 15998
rect 172510 15922 172562 15934
rect 174302 15986 174354 15998
rect 174302 15922 174354 15934
rect 177214 15986 177266 15998
rect 177214 15922 177266 15934
rect 1344 15706 178800 15740
rect 1344 15654 45538 15706
rect 45590 15654 45642 15706
rect 45694 15654 45746 15706
rect 45798 15654 89862 15706
rect 89914 15654 89966 15706
rect 90018 15654 90070 15706
rect 90122 15654 134186 15706
rect 134238 15654 134290 15706
rect 134342 15654 134394 15706
rect 134446 15654 178510 15706
rect 178562 15654 178614 15706
rect 178666 15654 178718 15706
rect 178770 15654 178800 15706
rect 1344 15620 178800 15654
rect 178110 15538 178162 15550
rect 178110 15474 178162 15486
rect 1344 14922 178640 14956
rect 1344 14870 23376 14922
rect 23428 14870 23480 14922
rect 23532 14870 23584 14922
rect 23636 14870 67700 14922
rect 67752 14870 67804 14922
rect 67856 14870 67908 14922
rect 67960 14870 112024 14922
rect 112076 14870 112128 14922
rect 112180 14870 112232 14922
rect 112284 14870 156348 14922
rect 156400 14870 156452 14922
rect 156504 14870 156556 14922
rect 156608 14870 178640 14922
rect 1344 14836 178640 14870
rect 1344 14138 178800 14172
rect 1344 14086 45538 14138
rect 45590 14086 45642 14138
rect 45694 14086 45746 14138
rect 45798 14086 89862 14138
rect 89914 14086 89966 14138
rect 90018 14086 90070 14138
rect 90122 14086 134186 14138
rect 134238 14086 134290 14138
rect 134342 14086 134394 14138
rect 134446 14086 178510 14138
rect 178562 14086 178614 14138
rect 178666 14086 178718 14138
rect 178770 14086 178800 14138
rect 1344 14052 178800 14086
rect 1344 13354 178640 13388
rect 1344 13302 23376 13354
rect 23428 13302 23480 13354
rect 23532 13302 23584 13354
rect 23636 13302 67700 13354
rect 67752 13302 67804 13354
rect 67856 13302 67908 13354
rect 67960 13302 112024 13354
rect 112076 13302 112128 13354
rect 112180 13302 112232 13354
rect 112284 13302 156348 13354
rect 156400 13302 156452 13354
rect 156504 13302 156556 13354
rect 156608 13302 178640 13354
rect 1344 13268 178640 13302
rect 1344 12570 178800 12604
rect 1344 12518 45538 12570
rect 45590 12518 45642 12570
rect 45694 12518 45746 12570
rect 45798 12518 89862 12570
rect 89914 12518 89966 12570
rect 90018 12518 90070 12570
rect 90122 12518 134186 12570
rect 134238 12518 134290 12570
rect 134342 12518 134394 12570
rect 134446 12518 178510 12570
rect 178562 12518 178614 12570
rect 178666 12518 178718 12570
rect 178770 12518 178800 12570
rect 1344 12484 178800 12518
rect 1344 11786 178640 11820
rect 1344 11734 23376 11786
rect 23428 11734 23480 11786
rect 23532 11734 23584 11786
rect 23636 11734 67700 11786
rect 67752 11734 67804 11786
rect 67856 11734 67908 11786
rect 67960 11734 112024 11786
rect 112076 11734 112128 11786
rect 112180 11734 112232 11786
rect 112284 11734 156348 11786
rect 156400 11734 156452 11786
rect 156504 11734 156556 11786
rect 156608 11734 178640 11786
rect 1344 11700 178640 11734
rect 1344 11002 178800 11036
rect 1344 10950 45538 11002
rect 45590 10950 45642 11002
rect 45694 10950 45746 11002
rect 45798 10950 89862 11002
rect 89914 10950 89966 11002
rect 90018 10950 90070 11002
rect 90122 10950 134186 11002
rect 134238 10950 134290 11002
rect 134342 10950 134394 11002
rect 134446 10950 178510 11002
rect 178562 10950 178614 11002
rect 178666 10950 178718 11002
rect 178770 10950 178800 11002
rect 1344 10916 178800 10950
rect 1344 10218 178640 10252
rect 1344 10166 23376 10218
rect 23428 10166 23480 10218
rect 23532 10166 23584 10218
rect 23636 10166 67700 10218
rect 67752 10166 67804 10218
rect 67856 10166 67908 10218
rect 67960 10166 112024 10218
rect 112076 10166 112128 10218
rect 112180 10166 112232 10218
rect 112284 10166 156348 10218
rect 156400 10166 156452 10218
rect 156504 10166 156556 10218
rect 156608 10166 178640 10218
rect 1344 10132 178640 10166
rect 1344 9434 178800 9468
rect 1344 9382 45538 9434
rect 45590 9382 45642 9434
rect 45694 9382 45746 9434
rect 45798 9382 89862 9434
rect 89914 9382 89966 9434
rect 90018 9382 90070 9434
rect 90122 9382 134186 9434
rect 134238 9382 134290 9434
rect 134342 9382 134394 9434
rect 134446 9382 178510 9434
rect 178562 9382 178614 9434
rect 178666 9382 178718 9434
rect 178770 9382 178800 9434
rect 1344 9348 178800 9382
rect 1344 8650 178640 8684
rect 1344 8598 23376 8650
rect 23428 8598 23480 8650
rect 23532 8598 23584 8650
rect 23636 8598 67700 8650
rect 67752 8598 67804 8650
rect 67856 8598 67908 8650
rect 67960 8598 112024 8650
rect 112076 8598 112128 8650
rect 112180 8598 112232 8650
rect 112284 8598 156348 8650
rect 156400 8598 156452 8650
rect 156504 8598 156556 8650
rect 156608 8598 178640 8650
rect 1344 8564 178640 8598
rect 1344 7866 178800 7900
rect 1344 7814 45538 7866
rect 45590 7814 45642 7866
rect 45694 7814 45746 7866
rect 45798 7814 89862 7866
rect 89914 7814 89966 7866
rect 90018 7814 90070 7866
rect 90122 7814 134186 7866
rect 134238 7814 134290 7866
rect 134342 7814 134394 7866
rect 134446 7814 178510 7866
rect 178562 7814 178614 7866
rect 178666 7814 178718 7866
rect 178770 7814 178800 7866
rect 1344 7780 178800 7814
rect 58270 7362 58322 7374
rect 57922 7310 57934 7362
rect 57986 7310 57998 7362
rect 58270 7298 58322 7310
rect 65438 7362 65490 7374
rect 66334 7362 66386 7374
rect 66098 7310 66110 7362
rect 66162 7310 66174 7362
rect 65438 7298 65490 7310
rect 66334 7298 66386 7310
rect 66894 7362 66946 7374
rect 66894 7298 66946 7310
rect 67342 7362 67394 7374
rect 67342 7298 67394 7310
rect 67678 7362 67730 7374
rect 67678 7298 67730 7310
rect 1344 7082 178640 7116
rect 1344 7030 23376 7082
rect 23428 7030 23480 7082
rect 23532 7030 23584 7082
rect 23636 7030 67700 7082
rect 67752 7030 67804 7082
rect 67856 7030 67908 7082
rect 67960 7030 112024 7082
rect 112076 7030 112128 7082
rect 112180 7030 112232 7082
rect 112284 7030 156348 7082
rect 156400 7030 156452 7082
rect 156504 7030 156556 7082
rect 156608 7030 178640 7082
rect 1344 6996 178640 7030
rect 64094 6802 64146 6814
rect 64094 6738 64146 6750
rect 64542 6802 64594 6814
rect 64542 6738 64594 6750
rect 65102 6802 65154 6814
rect 65102 6738 65154 6750
rect 65998 6802 66050 6814
rect 65998 6738 66050 6750
rect 66894 6802 66946 6814
rect 66894 6738 66946 6750
rect 57486 6578 57538 6590
rect 58382 6578 58434 6590
rect 59614 6578 59666 6590
rect 96462 6578 96514 6590
rect 57810 6526 57822 6578
rect 57874 6526 57886 6578
rect 58706 6526 58718 6578
rect 58770 6526 58782 6578
rect 59266 6526 59278 6578
rect 59330 6526 59342 6578
rect 65426 6526 65438 6578
rect 65490 6526 65502 6578
rect 57486 6514 57538 6526
rect 58382 6514 58434 6526
rect 59614 6514 59666 6526
rect 96462 6514 96514 6526
rect 97134 6578 97186 6590
rect 97134 6514 97186 6526
rect 114830 6578 114882 6590
rect 114830 6514 114882 6526
rect 60062 6466 60114 6478
rect 60062 6402 60114 6414
rect 63758 6466 63810 6478
rect 63758 6402 63810 6414
rect 66110 6466 66162 6478
rect 66110 6402 66162 6414
rect 67006 6466 67058 6478
rect 67006 6402 67058 6414
rect 67678 6466 67730 6478
rect 67678 6402 67730 6414
rect 68126 6466 68178 6478
rect 68126 6402 68178 6414
rect 68574 6466 68626 6478
rect 68574 6402 68626 6414
rect 96350 6466 96402 6478
rect 96350 6402 96402 6414
rect 97022 6466 97074 6478
rect 97022 6402 97074 6414
rect 114718 6466 114770 6478
rect 114718 6402 114770 6414
rect 1344 6298 178800 6332
rect 1344 6246 45538 6298
rect 45590 6246 45642 6298
rect 45694 6246 45746 6298
rect 45798 6246 89862 6298
rect 89914 6246 89966 6298
rect 90018 6246 90070 6298
rect 90122 6246 134186 6298
rect 134238 6246 134290 6298
rect 134342 6246 134394 6298
rect 134446 6246 178510 6298
rect 178562 6246 178614 6298
rect 178666 6246 178718 6298
rect 178770 6246 178800 6298
rect 1344 6212 178800 6246
rect 61182 6130 61234 6142
rect 61182 6066 61234 6078
rect 68798 6130 68850 6142
rect 68798 6066 68850 6078
rect 69246 6130 69298 6142
rect 69246 6066 69298 6078
rect 96014 6130 96066 6142
rect 96014 6066 96066 6078
rect 114606 6130 114658 6142
rect 114606 6066 114658 6078
rect 59726 6018 59778 6030
rect 59726 5954 59778 5966
rect 107662 6018 107714 6030
rect 107662 5954 107714 5966
rect 60286 5906 60338 5918
rect 60286 5842 60338 5854
rect 60734 5906 60786 5918
rect 60734 5842 60786 5854
rect 63758 5906 63810 5918
rect 65662 5906 65714 5918
rect 64418 5854 64430 5906
rect 64482 5854 64494 5906
rect 63758 5842 63810 5854
rect 65662 5842 65714 5854
rect 66222 5906 66274 5918
rect 96126 5906 96178 5918
rect 67218 5854 67230 5906
rect 67282 5854 67294 5906
rect 68114 5854 68126 5906
rect 68178 5854 68190 5906
rect 66222 5842 66274 5854
rect 96126 5842 96178 5854
rect 97358 5906 97410 5918
rect 97358 5842 97410 5854
rect 98030 5906 98082 5918
rect 98030 5842 98082 5854
rect 113262 5906 113314 5918
rect 113262 5842 113314 5854
rect 113934 5906 113986 5918
rect 113934 5842 113986 5854
rect 115278 5906 115330 5918
rect 115278 5842 115330 5854
rect 56366 5794 56418 5806
rect 57598 5794 57650 5806
rect 58494 5794 58546 5806
rect 61966 5794 62018 5806
rect 56690 5742 56702 5794
rect 56754 5742 56766 5794
rect 57922 5742 57934 5794
rect 57986 5742 57998 5794
rect 58706 5742 58718 5794
rect 58770 5742 58782 5794
rect 56366 5730 56418 5742
rect 57598 5730 57650 5742
rect 58494 5730 58546 5742
rect 61966 5730 62018 5742
rect 62862 5794 62914 5806
rect 62862 5730 62914 5742
rect 63310 5794 63362 5806
rect 79326 5794 79378 5806
rect 64642 5742 64654 5794
rect 64706 5742 64718 5794
rect 66434 5742 66446 5794
rect 66498 5742 66510 5794
rect 67442 5742 67454 5794
rect 67506 5742 67518 5794
rect 68338 5742 68350 5794
rect 68402 5742 68414 5794
rect 63310 5730 63362 5742
rect 79326 5730 79378 5742
rect 97246 5682 97298 5694
rect 97246 5618 97298 5630
rect 97918 5682 97970 5694
rect 97918 5618 97970 5630
rect 113150 5682 113202 5694
rect 113150 5618 113202 5630
rect 113822 5682 113874 5694
rect 113822 5618 113874 5630
rect 115166 5682 115218 5694
rect 115166 5618 115218 5630
rect 1344 5514 178640 5548
rect 1344 5462 23376 5514
rect 23428 5462 23480 5514
rect 23532 5462 23584 5514
rect 23636 5462 67700 5514
rect 67752 5462 67804 5514
rect 67856 5462 67908 5514
rect 67960 5462 112024 5514
rect 112076 5462 112128 5514
rect 112180 5462 112232 5514
rect 112284 5462 156348 5514
rect 156400 5462 156452 5514
rect 156504 5462 156556 5514
rect 156608 5462 178640 5514
rect 1344 5428 178640 5462
rect 86606 5346 86658 5358
rect 86606 5282 86658 5294
rect 92318 5346 92370 5358
rect 92318 5282 92370 5294
rect 94782 5346 94834 5358
rect 94782 5282 94834 5294
rect 113710 5346 113762 5358
rect 113710 5282 113762 5294
rect 49198 5234 49250 5246
rect 60622 5234 60674 5246
rect 55458 5182 55470 5234
rect 55522 5182 55534 5234
rect 56578 5182 56590 5234
rect 56642 5182 56654 5234
rect 57474 5182 57486 5234
rect 57538 5182 57550 5234
rect 58370 5182 58382 5234
rect 58434 5182 58446 5234
rect 59266 5182 59278 5234
rect 59330 5182 59342 5234
rect 60162 5182 60174 5234
rect 60226 5182 60238 5234
rect 49198 5170 49250 5182
rect 60622 5170 60674 5182
rect 61406 5234 61458 5246
rect 62638 5234 62690 5246
rect 61730 5182 61742 5234
rect 61794 5182 61806 5234
rect 61406 5170 61458 5182
rect 62638 5170 62690 5182
rect 62974 5234 63026 5246
rect 62974 5170 63026 5182
rect 64430 5234 64482 5246
rect 65326 5234 65378 5246
rect 79886 5234 79938 5246
rect 64642 5182 64654 5234
rect 64706 5182 64718 5234
rect 78978 5182 78990 5234
rect 79042 5182 79054 5234
rect 64430 5170 64482 5182
rect 65326 5170 65378 5182
rect 79886 5170 79938 5182
rect 93214 5234 93266 5246
rect 93214 5170 93266 5182
rect 34302 5122 34354 5134
rect 33618 5070 33630 5122
rect 33682 5070 33694 5122
rect 34302 5058 34354 5070
rect 35198 5122 35250 5134
rect 35198 5058 35250 5070
rect 35534 5122 35586 5134
rect 50430 5122 50482 5134
rect 48514 5070 48526 5122
rect 48578 5070 48590 5122
rect 49746 5070 49758 5122
rect 49810 5070 49822 5122
rect 35534 5058 35586 5070
rect 50430 5058 50482 5070
rect 55694 5122 55746 5134
rect 69246 5122 69298 5134
rect 56354 5070 56366 5122
rect 56418 5070 56430 5122
rect 57250 5070 57262 5122
rect 57314 5070 57326 5122
rect 58146 5070 58158 5122
rect 58210 5070 58222 5122
rect 59042 5070 59054 5122
rect 59106 5070 59118 5122
rect 66322 5070 66334 5122
rect 66386 5070 66398 5122
rect 68226 5070 68238 5122
rect 68290 5070 68302 5122
rect 68450 5070 68462 5122
rect 68514 5070 68526 5122
rect 55694 5058 55746 5070
rect 69246 5058 69298 5070
rect 70366 5122 70418 5134
rect 70366 5058 70418 5070
rect 70702 5122 70754 5134
rect 70702 5058 70754 5070
rect 75854 5122 75906 5134
rect 79662 5122 79714 5134
rect 79090 5070 79102 5122
rect 79154 5070 79166 5122
rect 75854 5058 75906 5070
rect 79662 5058 79714 5070
rect 85934 5122 85986 5134
rect 85934 5058 85986 5070
rect 86494 5122 86546 5134
rect 86494 5058 86546 5070
rect 92430 5122 92482 5134
rect 98254 5122 98306 5134
rect 106766 5122 106818 5134
rect 96338 5070 96350 5122
rect 96402 5119 96414 5122
rect 96562 5119 96574 5122
rect 96402 5073 96574 5119
rect 96402 5070 96414 5073
rect 96562 5070 96574 5073
rect 96626 5070 96638 5122
rect 105970 5070 105982 5122
rect 106034 5070 106046 5122
rect 92430 5058 92482 5070
rect 98254 5058 98306 5070
rect 106766 5058 106818 5070
rect 107662 5122 107714 5134
rect 107662 5058 107714 5070
rect 112254 5122 112306 5134
rect 112254 5058 112306 5070
rect 115614 5122 115666 5134
rect 120542 5122 120594 5134
rect 118850 5070 118862 5122
rect 118914 5070 118926 5122
rect 115614 5058 115666 5070
rect 120542 5058 120594 5070
rect 59838 5010 59890 5022
rect 59838 4946 59890 4958
rect 63534 5010 63586 5022
rect 63534 4946 63586 4958
rect 67566 5010 67618 5022
rect 94894 5010 94946 5022
rect 83346 4958 83358 5010
rect 83410 4958 83422 5010
rect 67566 4946 67618 4958
rect 94894 4946 94946 4958
rect 95566 5010 95618 5022
rect 95566 4946 95618 4958
rect 96798 5010 96850 5022
rect 96798 4946 96850 4958
rect 97470 5010 97522 5022
rect 97470 4946 97522 4958
rect 98142 5010 98194 5022
rect 98142 4946 98194 4958
rect 112366 5010 112418 5022
rect 112366 4946 112418 4958
rect 113038 5010 113090 5022
rect 113038 4946 113090 4958
rect 113598 5010 113650 5022
rect 113598 4946 113650 4958
rect 114270 5010 114322 5022
rect 114270 4946 114322 4958
rect 119646 5010 119698 5022
rect 119646 4946 119698 4958
rect 120990 5010 121042 5022
rect 120990 4946 121042 4958
rect 63646 4898 63698 4910
rect 63646 4834 63698 4846
rect 65438 4898 65490 4910
rect 65438 4834 65490 4846
rect 66334 4898 66386 4910
rect 66334 4834 66386 4846
rect 67230 4898 67282 4910
rect 67230 4834 67282 4846
rect 69806 4898 69858 4910
rect 83022 4898 83074 4910
rect 80210 4846 80222 4898
rect 80274 4846 80286 4898
rect 69806 4834 69858 4846
rect 83022 4834 83074 4846
rect 84366 4898 84418 4910
rect 84366 4834 84418 4846
rect 85822 4898 85874 4910
rect 85822 4834 85874 4846
rect 96126 4898 96178 4910
rect 96126 4834 96178 4846
rect 98814 4898 98866 4910
rect 98814 4834 98866 4846
rect 105422 4898 105474 4910
rect 105422 4834 105474 4846
rect 108110 4898 108162 4910
rect 108110 4834 108162 4846
rect 114942 4898 114994 4910
rect 114942 4834 114994 4846
rect 115726 4898 115778 4910
rect 115726 4834 115778 4846
rect 118302 4898 118354 4910
rect 118302 4834 118354 4846
rect 141374 4898 141426 4910
rect 141374 4834 141426 4846
rect 1344 4730 178800 4764
rect 1344 4678 45538 4730
rect 45590 4678 45642 4730
rect 45694 4678 45746 4730
rect 45798 4678 89862 4730
rect 89914 4678 89966 4730
rect 90018 4678 90070 4730
rect 90122 4678 134186 4730
rect 134238 4678 134290 4730
rect 134342 4678 134394 4730
rect 134446 4678 178510 4730
rect 178562 4678 178614 4730
rect 178666 4678 178718 4730
rect 178770 4678 178800 4730
rect 1344 4644 178800 4678
rect 36430 4562 36482 4574
rect 36430 4498 36482 4510
rect 36878 4562 36930 4574
rect 36878 4498 36930 4510
rect 51550 4562 51602 4574
rect 51550 4498 51602 4510
rect 58382 4562 58434 4574
rect 58382 4498 58434 4510
rect 62190 4562 62242 4574
rect 62190 4498 62242 4510
rect 63534 4562 63586 4574
rect 63534 4498 63586 4510
rect 78990 4562 79042 4574
rect 78990 4498 79042 4510
rect 95902 4562 95954 4574
rect 95902 4498 95954 4510
rect 97246 4562 97298 4574
rect 97246 4498 97298 4510
rect 98030 4562 98082 4574
rect 98030 4498 98082 4510
rect 113150 4562 113202 4574
rect 113150 4498 113202 4510
rect 113934 4562 113986 4574
rect 113934 4498 113986 4510
rect 114494 4562 114546 4574
rect 114494 4498 114546 4510
rect 115278 4562 115330 4574
rect 115278 4498 115330 4510
rect 115838 4562 115890 4574
rect 115838 4498 115890 4510
rect 10670 4450 10722 4462
rect 10670 4386 10722 4398
rect 26350 4450 26402 4462
rect 26350 4386 26402 4398
rect 28030 4450 28082 4462
rect 28030 4386 28082 4398
rect 33518 4450 33570 4462
rect 33518 4386 33570 4398
rect 53230 4450 53282 4462
rect 53230 4386 53282 4398
rect 54910 4450 54962 4462
rect 57710 4450 57762 4462
rect 56690 4398 56702 4450
rect 56754 4398 56766 4450
rect 54910 4386 54962 4398
rect 57710 4386 57762 4398
rect 58270 4450 58322 4462
rect 58270 4386 58322 4398
rect 62862 4450 62914 4462
rect 62862 4386 62914 4398
rect 63422 4450 63474 4462
rect 63422 4386 63474 4398
rect 65550 4450 65602 4462
rect 65550 4386 65602 4398
rect 71150 4450 71202 4462
rect 71150 4386 71202 4398
rect 72606 4450 72658 4462
rect 72606 4386 72658 4398
rect 74286 4450 74338 4462
rect 74286 4386 74338 4398
rect 74846 4450 74898 4462
rect 74846 4386 74898 4398
rect 76190 4450 76242 4462
rect 76190 4386 76242 4398
rect 79662 4450 79714 4462
rect 79662 4386 79714 4398
rect 85822 4450 85874 4462
rect 85822 4386 85874 4398
rect 93662 4450 93714 4462
rect 93662 4386 93714 4398
rect 94670 4450 94722 4462
rect 94670 4386 94722 4398
rect 96014 4450 96066 4462
rect 96014 4386 96066 4398
rect 108110 4450 108162 4462
rect 108110 4386 108162 4398
rect 109790 4450 109842 4462
rect 109790 4386 109842 4398
rect 114606 4450 114658 4462
rect 114606 4386 114658 4398
rect 121102 4450 121154 4462
rect 121102 4386 121154 4398
rect 129054 4450 129106 4462
rect 129054 4386 129106 4398
rect 129950 4450 130002 4462
rect 129950 4386 130002 4398
rect 132750 4450 132802 4462
rect 132750 4386 132802 4398
rect 133422 4450 133474 4462
rect 133422 4386 133474 4398
rect 141262 4450 141314 4462
rect 141262 4386 141314 4398
rect 141934 4450 141986 4462
rect 141934 4386 141986 4398
rect 151790 4450 151842 4462
rect 151790 4386 151842 4398
rect 153470 4450 153522 4462
rect 153470 4386 153522 4398
rect 32958 4338 33010 4350
rect 35198 4338 35250 4350
rect 31266 4286 31278 4338
rect 31330 4286 31342 4338
rect 34402 4286 34414 4338
rect 34466 4286 34478 4338
rect 32958 4274 33010 4286
rect 35198 4274 35250 4286
rect 36094 4338 36146 4350
rect 51214 4338 51266 4350
rect 70142 4338 70194 4350
rect 49746 4286 49758 4338
rect 49810 4286 49822 4338
rect 56466 4286 56478 4338
rect 56530 4286 56542 4338
rect 61170 4286 61182 4338
rect 61234 4286 61246 4338
rect 64418 4286 64430 4338
rect 64482 4286 64494 4338
rect 64642 4286 64654 4338
rect 64706 4286 64718 4338
rect 66098 4286 66110 4338
rect 66162 4286 66174 4338
rect 69346 4286 69358 4338
rect 69410 4286 69422 4338
rect 36094 4274 36146 4286
rect 51214 4274 51266 4286
rect 70142 4274 70194 4286
rect 72270 4338 72322 4350
rect 72270 4274 72322 4286
rect 73950 4338 74002 4350
rect 73950 4274 74002 4286
rect 84030 4338 84082 4350
rect 92990 4338 93042 4350
rect 107438 4338 107490 4350
rect 120430 4338 120482 4350
rect 132302 4338 132354 4350
rect 140814 4338 140866 4350
rect 85026 4286 85038 4338
rect 85090 4286 85102 4338
rect 86482 4286 86494 4338
rect 86546 4286 86558 4338
rect 105746 4286 105758 4338
rect 105810 4286 105822 4338
rect 118738 4286 118750 4338
rect 118802 4286 118814 4338
rect 130722 4286 130734 4338
rect 130786 4286 130798 4338
rect 139346 4286 139358 4338
rect 139410 4286 139422 4338
rect 84030 4274 84082 4286
rect 92990 4274 93042 4286
rect 107438 4274 107490 4286
rect 120430 4274 120482 4286
rect 132302 4274 132354 4286
rect 140814 4274 140866 4286
rect 13022 4226 13074 4238
rect 13022 4162 13074 4174
rect 28702 4226 28754 4238
rect 28702 4162 28754 4174
rect 30830 4226 30882 4238
rect 30830 4162 30882 4174
rect 32062 4226 32114 4238
rect 32062 4162 32114 4174
rect 50318 4226 50370 4238
rect 50318 4162 50370 4174
rect 54350 4226 54402 4238
rect 54350 4162 54402 4174
rect 55806 4226 55858 4238
rect 71822 4226 71874 4238
rect 59826 4174 59838 4226
rect 59890 4174 59902 4226
rect 65762 4174 65774 4226
rect 65826 4223 65838 4226
rect 66098 4223 66110 4226
rect 65826 4177 66110 4223
rect 65826 4174 65838 4177
rect 66098 4174 66110 4177
rect 66162 4174 66174 4226
rect 68450 4174 68462 4226
rect 68514 4174 68526 4226
rect 69570 4174 69582 4226
rect 69634 4174 69646 4226
rect 70466 4174 70478 4226
rect 70530 4174 70542 4226
rect 55806 4162 55858 4174
rect 71822 4162 71874 4174
rect 73502 4226 73554 4238
rect 73502 4162 73554 4174
rect 75742 4226 75794 4238
rect 75742 4162 75794 4174
rect 77086 4226 77138 4238
rect 77086 4162 77138 4174
rect 78542 4226 78594 4238
rect 78542 4162 78594 4174
rect 83694 4226 83746 4238
rect 83694 4162 83746 4174
rect 84590 4226 84642 4238
rect 84590 4162 84642 4174
rect 91422 4226 91474 4238
rect 91422 4162 91474 4174
rect 92430 4226 92482 4238
rect 92430 4162 92482 4174
rect 105198 4226 105250 4238
rect 105198 4162 105250 4174
rect 106542 4226 106594 4238
rect 106542 4162 106594 4174
rect 118190 4226 118242 4238
rect 118190 4162 118242 4174
rect 119534 4226 119586 4238
rect 119534 4162 119586 4174
rect 126926 4226 126978 4238
rect 126926 4162 126978 4174
rect 127486 4226 127538 4238
rect 127486 4162 127538 4174
rect 131406 4226 131458 4238
rect 131406 4162 131458 4174
rect 139918 4226 139970 4238
rect 139918 4162 139970 4174
rect 142606 4226 142658 4238
rect 142606 4162 142658 4174
rect 150446 4226 150498 4238
rect 150446 4162 150498 4174
rect 151006 4226 151058 4238
rect 151006 4162 151058 4174
rect 93102 4114 93154 4126
rect 93102 4050 93154 4062
rect 1344 3946 178640 3980
rect 1344 3894 23376 3946
rect 23428 3894 23480 3946
rect 23532 3894 23584 3946
rect 23636 3894 67700 3946
rect 67752 3894 67804 3946
rect 67856 3894 67908 3946
rect 67960 3894 112024 3946
rect 112076 3894 112128 3946
rect 112180 3894 112232 3946
rect 112284 3894 156348 3946
rect 156400 3894 156452 3946
rect 156504 3894 156556 3946
rect 156608 3894 178640 3946
rect 1344 3860 178640 3894
rect 32510 3666 32562 3678
rect 9650 3614 9662 3666
rect 9714 3614 9726 3666
rect 28242 3614 28254 3666
rect 28306 3614 28318 3666
rect 32510 3602 32562 3614
rect 34862 3666 34914 3678
rect 57822 3666 57874 3678
rect 58718 3666 58770 3678
rect 59614 3666 59666 3678
rect 52770 3614 52782 3666
rect 52834 3614 52846 3666
rect 54898 3614 54910 3666
rect 54962 3614 54974 3666
rect 57474 3614 57486 3666
rect 57538 3614 57550 3666
rect 58370 3614 58382 3666
rect 58434 3614 58446 3666
rect 59266 3614 59278 3666
rect 59330 3614 59342 3666
rect 34862 3602 34914 3614
rect 57822 3602 57874 3614
rect 58718 3602 58770 3614
rect 59614 3602 59666 3614
rect 64654 3666 64706 3678
rect 68462 3666 68514 3678
rect 85710 3666 85762 3678
rect 64866 3614 64878 3666
rect 64930 3614 64942 3666
rect 66882 3614 66894 3666
rect 66946 3614 66958 3666
rect 73378 3614 73390 3666
rect 73442 3614 73454 3666
rect 75506 3614 75518 3666
rect 75570 3614 75582 3666
rect 64654 3602 64706 3614
rect 68462 3602 68514 3614
rect 85710 3602 85762 3614
rect 90638 3666 90690 3678
rect 121102 3666 121154 3678
rect 92754 3614 92766 3666
rect 92818 3614 92830 3666
rect 94882 3614 94894 3666
rect 94946 3614 94958 3666
rect 110562 3614 110574 3666
rect 110626 3614 110638 3666
rect 90638 3602 90690 3614
rect 121102 3602 121154 3614
rect 121550 3666 121602 3678
rect 131966 3666 132018 3678
rect 130386 3614 130398 3666
rect 130450 3614 130462 3666
rect 121550 3602 121602 3614
rect 131966 3602 132018 3614
rect 140366 3666 140418 3678
rect 153906 3614 153918 3666
rect 153970 3614 153982 3666
rect 140366 3602 140418 3614
rect 29262 3554 29314 3566
rect 62190 3554 62242 3566
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 25330 3502 25342 3554
rect 25394 3502 25406 3554
rect 34066 3502 34078 3554
rect 34130 3502 34142 3554
rect 35522 3502 35534 3554
rect 35586 3502 35598 3554
rect 55682 3502 55694 3554
rect 55746 3502 55758 3554
rect 57922 3502 57934 3554
rect 57986 3551 57998 3554
rect 58146 3551 58158 3554
rect 57986 3505 58158 3551
rect 57986 3502 57998 3505
rect 58146 3502 58158 3505
rect 58210 3502 58222 3554
rect 29262 3490 29314 3502
rect 62190 3490 62242 3502
rect 63758 3554 63810 3566
rect 81230 3554 81282 3566
rect 105982 3554 106034 3566
rect 132862 3554 132914 3566
rect 141262 3554 141314 3566
rect 65650 3502 65662 3554
rect 65714 3502 65726 3554
rect 69122 3502 69134 3554
rect 69186 3502 69198 3554
rect 70802 3502 70814 3554
rect 70866 3502 70878 3554
rect 72594 3502 72606 3554
rect 72658 3502 72670 3554
rect 84914 3502 84926 3554
rect 84978 3502 84990 3554
rect 86482 3502 86494 3554
rect 86546 3502 86558 3554
rect 92082 3502 92094 3554
rect 92146 3502 92158 3554
rect 107762 3502 107774 3554
rect 107826 3502 107838 3554
rect 119522 3502 119534 3554
rect 119586 3502 119598 3554
rect 120530 3502 120542 3554
rect 120594 3502 120606 3554
rect 127586 3502 127598 3554
rect 127650 3502 127662 3554
rect 128258 3502 128270 3554
rect 128322 3502 128334 3554
rect 131170 3502 131182 3554
rect 131234 3502 131246 3554
rect 139682 3502 139694 3554
rect 139746 3502 139758 3554
rect 151106 3502 151118 3554
rect 151170 3502 151182 3554
rect 151778 3502 151790 3554
rect 151842 3502 151854 3554
rect 63758 3490 63810 3502
rect 81230 3490 81282 3502
rect 105982 3490 106034 3502
rect 132862 3490 132914 3502
rect 141262 3490 141314 3502
rect 14254 3442 14306 3454
rect 62078 3442 62130 3454
rect 11778 3390 11790 3442
rect 11842 3390 11854 3442
rect 26114 3390 26126 3442
rect 26178 3390 26190 3442
rect 14254 3378 14306 3390
rect 62078 3378 62130 3390
rect 62862 3442 62914 3454
rect 62862 3378 62914 3390
rect 71598 3442 71650 3454
rect 71598 3378 71650 3390
rect 76302 3442 76354 3454
rect 76302 3378 76354 3390
rect 77310 3442 77362 3454
rect 77310 3378 77362 3390
rect 78990 3442 79042 3454
rect 78990 3378 79042 3390
rect 80222 3442 80274 3454
rect 80222 3378 80274 3390
rect 80670 3442 80722 3454
rect 80670 3378 80722 3390
rect 105534 3442 105586 3454
rect 142942 3442 142994 3454
rect 108434 3390 108446 3442
rect 108498 3390 108510 3442
rect 119746 3390 119758 3442
rect 119810 3390 119822 3442
rect 105534 3378 105586 3390
rect 142942 3378 142994 3390
rect 7310 3330 7362 3342
rect 7310 3266 7362 3278
rect 13582 3330 13634 3342
rect 13582 3266 13634 3278
rect 15150 3330 15202 3342
rect 15150 3266 15202 3278
rect 17502 3330 17554 3342
rect 17502 3266 17554 3278
rect 19630 3330 19682 3342
rect 19630 3266 19682 3278
rect 21422 3330 21474 3342
rect 21422 3266 21474 3278
rect 22990 3330 23042 3342
rect 22990 3266 23042 3278
rect 24446 3330 24498 3342
rect 24446 3266 24498 3278
rect 29710 3330 29762 3342
rect 29710 3266 29762 3278
rect 31390 3330 31442 3342
rect 31390 3266 31442 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 36206 3330 36258 3342
rect 36206 3266 36258 3278
rect 37102 3330 37154 3342
rect 37102 3266 37154 3278
rect 38110 3330 38162 3342
rect 38110 3266 38162 3278
rect 39790 3330 39842 3342
rect 39790 3266 39842 3278
rect 41470 3330 41522 3342
rect 41470 3266 41522 3278
rect 43150 3330 43202 3342
rect 43150 3266 43202 3278
rect 44942 3330 44994 3342
rect 44942 3266 44994 3278
rect 46510 3330 46562 3342
rect 46510 3266 46562 3278
rect 48862 3330 48914 3342
rect 48862 3266 48914 3278
rect 49870 3330 49922 3342
rect 49870 3266 49922 3278
rect 51550 3330 51602 3342
rect 51550 3266 51602 3278
rect 56702 3330 56754 3342
rect 56702 3266 56754 3278
rect 60622 3330 60674 3342
rect 60622 3266 60674 3278
rect 61406 3330 61458 3342
rect 61406 3266 61458 3278
rect 63422 3330 63474 3342
rect 63422 3266 63474 3278
rect 65662 3330 65714 3342
rect 65662 3266 65714 3278
rect 66446 3330 66498 3342
rect 66446 3266 66498 3278
rect 67566 3330 67618 3342
rect 67566 3266 67618 3278
rect 68910 3330 68962 3342
rect 68910 3266 68962 3278
rect 69806 3330 69858 3342
rect 69806 3266 69858 3278
rect 70590 3330 70642 3342
rect 70590 3266 70642 3278
rect 76638 3330 76690 3342
rect 76638 3266 76690 3278
rect 77646 3330 77698 3342
rect 77646 3266 77698 3278
rect 78206 3330 78258 3342
rect 78206 3266 78258 3278
rect 79326 3330 79378 3342
rect 79326 3266 79378 3278
rect 81790 3330 81842 3342
rect 81790 3266 81842 3278
rect 82910 3330 82962 3342
rect 82910 3266 82962 3278
rect 84366 3330 84418 3342
rect 84366 3266 84418 3278
rect 87054 3330 87106 3342
rect 87054 3266 87106 3278
rect 88062 3330 88114 3342
rect 88062 3266 88114 3278
rect 89630 3330 89682 3342
rect 89630 3266 89682 3278
rect 91086 3330 91138 3342
rect 91086 3266 91138 3278
rect 96574 3330 96626 3342
rect 96574 3266 96626 3278
rect 97246 3330 97298 3342
rect 97246 3266 97298 3278
rect 98030 3330 98082 3342
rect 98030 3266 98082 3278
rect 99822 3330 99874 3342
rect 99822 3266 99874 3278
rect 101390 3330 101442 3342
rect 101390 3266 101442 3278
rect 103742 3330 103794 3342
rect 103742 3266 103794 3278
rect 104750 3330 104802 3342
rect 104750 3266 104802 3278
rect 106430 3330 106482 3342
rect 106430 3266 106482 3278
rect 111582 3330 111634 3342
rect 111582 3266 111634 3278
rect 113150 3330 113202 3342
rect 113150 3266 113202 3278
rect 115502 3330 115554 3342
rect 115502 3266 115554 3278
rect 116510 3330 116562 3342
rect 116510 3266 116562 3278
rect 118190 3330 118242 3342
rect 123342 3330 123394 3342
rect 120306 3278 120318 3330
rect 120370 3278 120382 3330
rect 118190 3266 118242 3278
rect 123342 3266 123394 3278
rect 124910 3330 124962 3342
rect 124910 3266 124962 3278
rect 126366 3330 126418 3342
rect 126366 3266 126418 3278
rect 133310 3330 133362 3342
rect 133310 3266 133362 3278
rect 133982 3330 134034 3342
rect 133982 3266 134034 3278
rect 135102 3330 135154 3342
rect 135102 3266 135154 3278
rect 136670 3330 136722 3342
rect 136670 3266 136722 3278
rect 138126 3330 138178 3342
rect 138126 3266 138178 3278
rect 141710 3330 141762 3342
rect 141710 3266 141762 3278
rect 143390 3330 143442 3342
rect 143390 3266 143442 3278
rect 145070 3330 145122 3342
rect 145070 3266 145122 3278
rect 146862 3330 146914 3342
rect 146862 3266 146914 3278
rect 148430 3330 148482 3342
rect 148430 3266 148482 3278
rect 149886 3330 149938 3342
rect 149886 3266 149938 3278
rect 155150 3330 155202 3342
rect 155150 3266 155202 3278
rect 156830 3330 156882 3342
rect 156830 3266 156882 3278
rect 158622 3330 158674 3342
rect 158622 3266 158674 3278
rect 160190 3330 160242 3342
rect 160190 3266 160242 3278
rect 162542 3330 162594 3342
rect 162542 3266 162594 3278
rect 163550 3330 163602 3342
rect 163550 3266 163602 3278
rect 165230 3330 165282 3342
rect 165230 3266 165282 3278
rect 166910 3330 166962 3342
rect 166910 3266 166962 3278
rect 168590 3330 168642 3342
rect 168590 3266 168642 3278
rect 170382 3330 170434 3342
rect 170382 3266 170434 3278
rect 171950 3330 172002 3342
rect 171950 3266 172002 3278
rect 173070 3330 173122 3342
rect 173070 3266 173122 3278
rect 174302 3330 174354 3342
rect 174302 3266 174354 3278
rect 174974 3330 175026 3342
rect 174974 3266 175026 3278
rect 1344 3162 178800 3196
rect 1344 3110 45538 3162
rect 45590 3110 45642 3162
rect 45694 3110 45746 3162
rect 45798 3110 89862 3162
rect 89914 3110 89966 3162
rect 90018 3110 90070 3162
rect 90122 3110 134186 3162
rect 134238 3110 134290 3162
rect 134342 3110 134394 3162
rect 134446 3110 178510 3162
rect 178562 3110 178614 3162
rect 178666 3110 178718 3162
rect 178770 3110 178800 3162
rect 1344 3076 178800 3110
rect 69234 1710 69246 1762
rect 69298 1759 69310 1762
rect 69794 1759 69806 1762
rect 69298 1713 69806 1759
rect 69298 1710 69310 1713
rect 69794 1710 69806 1713
rect 69858 1710 69870 1762
rect 77634 1710 77646 1762
rect 77698 1759 77710 1762
rect 78194 1759 78206 1762
rect 77698 1713 78206 1759
rect 77698 1710 77710 1713
rect 78194 1710 78206 1713
rect 78258 1710 78270 1762
rect 80994 1710 81006 1762
rect 81058 1759 81070 1762
rect 81778 1759 81790 1762
rect 81058 1713 81790 1759
rect 81058 1710 81070 1713
rect 81778 1710 81790 1713
rect 81842 1710 81854 1762
rect 86034 1710 86046 1762
rect 86098 1759 86110 1762
rect 87042 1759 87054 1762
rect 86098 1713 87054 1759
rect 86098 1710 86110 1713
rect 87042 1710 87054 1713
rect 87106 1710 87118 1762
rect 96114 1710 96126 1762
rect 96178 1759 96190 1762
rect 97234 1759 97246 1762
rect 96178 1713 97246 1759
rect 96178 1710 96190 1713
rect 97234 1710 97246 1713
rect 97298 1710 97310 1762
rect 102834 1710 102846 1762
rect 102898 1759 102910 1762
rect 103730 1759 103742 1762
rect 102898 1713 103742 1759
rect 102898 1710 102910 1713
rect 103730 1710 103742 1713
rect 103794 1710 103806 1762
rect 114594 1710 114606 1762
rect 114658 1759 114670 1762
rect 115490 1759 115502 1762
rect 114658 1713 115502 1759
rect 114658 1710 114670 1713
rect 115490 1710 115502 1713
rect 115554 1710 115566 1762
rect 119634 1710 119646 1762
rect 119698 1759 119710 1762
rect 120306 1759 120318 1762
rect 119698 1713 120318 1759
rect 119698 1710 119710 1713
rect 120306 1710 120318 1713
rect 120370 1710 120382 1762
rect 133074 1710 133086 1762
rect 133138 1759 133150 1762
rect 133970 1759 133982 1762
rect 133138 1713 133982 1759
rect 133138 1710 133150 1713
rect 133970 1710 133982 1713
rect 134034 1710 134046 1762
rect 161634 1710 161646 1762
rect 161698 1759 161710 1762
rect 162530 1759 162542 1762
rect 161698 1713 162542 1759
rect 161698 1710 161710 1713
rect 162530 1710 162542 1713
rect 162594 1710 162606 1762
rect 173394 1710 173406 1762
rect 173458 1759 173470 1762
rect 174290 1759 174302 1762
rect 173458 1713 174302 1759
rect 173458 1710 173470 1713
rect 174290 1710 174302 1713
rect 174354 1710 174366 1762
<< via1 >>
rect 23376 16438 23428 16490
rect 23480 16438 23532 16490
rect 23584 16438 23636 16490
rect 67700 16438 67752 16490
rect 67804 16438 67856 16490
rect 67908 16438 67960 16490
rect 112024 16438 112076 16490
rect 112128 16438 112180 16490
rect 112232 16438 112284 16490
rect 156348 16438 156400 16490
rect 156452 16438 156504 16490
rect 156556 16438 156608 16490
rect 3166 15934 3218 15986
rect 4734 15934 4786 15986
rect 7870 15934 7922 15986
rect 9662 15934 9714 15986
rect 12574 15934 12626 15986
rect 14142 15934 14194 15986
rect 17502 15934 17554 15986
rect 18846 15934 18898 15986
rect 21982 15934 22034 15986
rect 23550 15934 23602 15986
rect 26686 15934 26738 15986
rect 28254 15934 28306 15986
rect 31390 15934 31442 15986
rect 33182 15934 33234 15986
rect 36094 15934 36146 15986
rect 37662 15934 37714 15986
rect 41022 15934 41074 15986
rect 42366 15934 42418 15986
rect 45502 15934 45554 15986
rect 47070 15934 47122 15986
rect 50206 15934 50258 15986
rect 51774 15934 51826 15986
rect 54910 15934 54962 15986
rect 56702 15934 56754 15986
rect 59614 15934 59666 15986
rect 61182 15934 61234 15986
rect 64542 15934 64594 15986
rect 65886 15934 65938 15986
rect 69022 15934 69074 15986
rect 70590 15934 70642 15986
rect 73726 15934 73778 15986
rect 75294 15934 75346 15986
rect 78430 15934 78482 15986
rect 80222 15934 80274 15986
rect 83134 15934 83186 15986
rect 84702 15934 84754 15986
rect 88062 15934 88114 15986
rect 89406 15934 89458 15986
rect 92542 15934 92594 15986
rect 94110 15934 94162 15986
rect 97246 15934 97298 15986
rect 98814 15934 98866 15986
rect 101950 15934 102002 15986
rect 103742 15934 103794 15986
rect 106654 15934 106706 15986
rect 108222 15934 108274 15986
rect 111582 15934 111634 15986
rect 112926 15934 112978 15986
rect 116062 15934 116114 15986
rect 117630 15934 117682 15986
rect 120766 15934 120818 15986
rect 122334 15934 122386 15986
rect 125470 15934 125522 15986
rect 127262 15934 127314 15986
rect 130174 15934 130226 15986
rect 131742 15934 131794 15986
rect 135102 15934 135154 15986
rect 136446 15934 136498 15986
rect 139582 15934 139634 15986
rect 141150 15934 141202 15986
rect 144286 15934 144338 15986
rect 145854 15934 145906 15986
rect 148990 15934 149042 15986
rect 150782 15934 150834 15986
rect 153694 15934 153746 15986
rect 155262 15934 155314 15986
rect 158622 15934 158674 15986
rect 159966 15934 160018 15986
rect 163102 15934 163154 15986
rect 164670 15934 164722 15986
rect 167806 15934 167858 15986
rect 169374 15934 169426 15986
rect 172510 15934 172562 15986
rect 174302 15934 174354 15986
rect 177214 15934 177266 15986
rect 45538 15654 45590 15706
rect 45642 15654 45694 15706
rect 45746 15654 45798 15706
rect 89862 15654 89914 15706
rect 89966 15654 90018 15706
rect 90070 15654 90122 15706
rect 134186 15654 134238 15706
rect 134290 15654 134342 15706
rect 134394 15654 134446 15706
rect 178510 15654 178562 15706
rect 178614 15654 178666 15706
rect 178718 15654 178770 15706
rect 178110 15486 178162 15538
rect 23376 14870 23428 14922
rect 23480 14870 23532 14922
rect 23584 14870 23636 14922
rect 67700 14870 67752 14922
rect 67804 14870 67856 14922
rect 67908 14870 67960 14922
rect 112024 14870 112076 14922
rect 112128 14870 112180 14922
rect 112232 14870 112284 14922
rect 156348 14870 156400 14922
rect 156452 14870 156504 14922
rect 156556 14870 156608 14922
rect 45538 14086 45590 14138
rect 45642 14086 45694 14138
rect 45746 14086 45798 14138
rect 89862 14086 89914 14138
rect 89966 14086 90018 14138
rect 90070 14086 90122 14138
rect 134186 14086 134238 14138
rect 134290 14086 134342 14138
rect 134394 14086 134446 14138
rect 178510 14086 178562 14138
rect 178614 14086 178666 14138
rect 178718 14086 178770 14138
rect 23376 13302 23428 13354
rect 23480 13302 23532 13354
rect 23584 13302 23636 13354
rect 67700 13302 67752 13354
rect 67804 13302 67856 13354
rect 67908 13302 67960 13354
rect 112024 13302 112076 13354
rect 112128 13302 112180 13354
rect 112232 13302 112284 13354
rect 156348 13302 156400 13354
rect 156452 13302 156504 13354
rect 156556 13302 156608 13354
rect 45538 12518 45590 12570
rect 45642 12518 45694 12570
rect 45746 12518 45798 12570
rect 89862 12518 89914 12570
rect 89966 12518 90018 12570
rect 90070 12518 90122 12570
rect 134186 12518 134238 12570
rect 134290 12518 134342 12570
rect 134394 12518 134446 12570
rect 178510 12518 178562 12570
rect 178614 12518 178666 12570
rect 178718 12518 178770 12570
rect 23376 11734 23428 11786
rect 23480 11734 23532 11786
rect 23584 11734 23636 11786
rect 67700 11734 67752 11786
rect 67804 11734 67856 11786
rect 67908 11734 67960 11786
rect 112024 11734 112076 11786
rect 112128 11734 112180 11786
rect 112232 11734 112284 11786
rect 156348 11734 156400 11786
rect 156452 11734 156504 11786
rect 156556 11734 156608 11786
rect 45538 10950 45590 11002
rect 45642 10950 45694 11002
rect 45746 10950 45798 11002
rect 89862 10950 89914 11002
rect 89966 10950 90018 11002
rect 90070 10950 90122 11002
rect 134186 10950 134238 11002
rect 134290 10950 134342 11002
rect 134394 10950 134446 11002
rect 178510 10950 178562 11002
rect 178614 10950 178666 11002
rect 178718 10950 178770 11002
rect 23376 10166 23428 10218
rect 23480 10166 23532 10218
rect 23584 10166 23636 10218
rect 67700 10166 67752 10218
rect 67804 10166 67856 10218
rect 67908 10166 67960 10218
rect 112024 10166 112076 10218
rect 112128 10166 112180 10218
rect 112232 10166 112284 10218
rect 156348 10166 156400 10218
rect 156452 10166 156504 10218
rect 156556 10166 156608 10218
rect 45538 9382 45590 9434
rect 45642 9382 45694 9434
rect 45746 9382 45798 9434
rect 89862 9382 89914 9434
rect 89966 9382 90018 9434
rect 90070 9382 90122 9434
rect 134186 9382 134238 9434
rect 134290 9382 134342 9434
rect 134394 9382 134446 9434
rect 178510 9382 178562 9434
rect 178614 9382 178666 9434
rect 178718 9382 178770 9434
rect 23376 8598 23428 8650
rect 23480 8598 23532 8650
rect 23584 8598 23636 8650
rect 67700 8598 67752 8650
rect 67804 8598 67856 8650
rect 67908 8598 67960 8650
rect 112024 8598 112076 8650
rect 112128 8598 112180 8650
rect 112232 8598 112284 8650
rect 156348 8598 156400 8650
rect 156452 8598 156504 8650
rect 156556 8598 156608 8650
rect 45538 7814 45590 7866
rect 45642 7814 45694 7866
rect 45746 7814 45798 7866
rect 89862 7814 89914 7866
rect 89966 7814 90018 7866
rect 90070 7814 90122 7866
rect 134186 7814 134238 7866
rect 134290 7814 134342 7866
rect 134394 7814 134446 7866
rect 178510 7814 178562 7866
rect 178614 7814 178666 7866
rect 178718 7814 178770 7866
rect 57934 7310 57986 7362
rect 58270 7310 58322 7362
rect 65438 7310 65490 7362
rect 66110 7310 66162 7362
rect 66334 7310 66386 7362
rect 66894 7310 66946 7362
rect 67342 7310 67394 7362
rect 67678 7310 67730 7362
rect 23376 7030 23428 7082
rect 23480 7030 23532 7082
rect 23584 7030 23636 7082
rect 67700 7030 67752 7082
rect 67804 7030 67856 7082
rect 67908 7030 67960 7082
rect 112024 7030 112076 7082
rect 112128 7030 112180 7082
rect 112232 7030 112284 7082
rect 156348 7030 156400 7082
rect 156452 7030 156504 7082
rect 156556 7030 156608 7082
rect 64094 6750 64146 6802
rect 64542 6750 64594 6802
rect 65102 6750 65154 6802
rect 65998 6750 66050 6802
rect 66894 6750 66946 6802
rect 57486 6526 57538 6578
rect 57822 6526 57874 6578
rect 58382 6526 58434 6578
rect 58718 6526 58770 6578
rect 59278 6526 59330 6578
rect 59614 6526 59666 6578
rect 65438 6526 65490 6578
rect 96462 6526 96514 6578
rect 97134 6526 97186 6578
rect 114830 6526 114882 6578
rect 60062 6414 60114 6466
rect 63758 6414 63810 6466
rect 66110 6414 66162 6466
rect 67006 6414 67058 6466
rect 67678 6414 67730 6466
rect 68126 6414 68178 6466
rect 68574 6414 68626 6466
rect 96350 6414 96402 6466
rect 97022 6414 97074 6466
rect 114718 6414 114770 6466
rect 45538 6246 45590 6298
rect 45642 6246 45694 6298
rect 45746 6246 45798 6298
rect 89862 6246 89914 6298
rect 89966 6246 90018 6298
rect 90070 6246 90122 6298
rect 134186 6246 134238 6298
rect 134290 6246 134342 6298
rect 134394 6246 134446 6298
rect 178510 6246 178562 6298
rect 178614 6246 178666 6298
rect 178718 6246 178770 6298
rect 61182 6078 61234 6130
rect 68798 6078 68850 6130
rect 69246 6078 69298 6130
rect 96014 6078 96066 6130
rect 114606 6078 114658 6130
rect 59726 5966 59778 6018
rect 107662 5966 107714 6018
rect 60286 5854 60338 5906
rect 60734 5854 60786 5906
rect 63758 5854 63810 5906
rect 64430 5854 64482 5906
rect 65662 5854 65714 5906
rect 66222 5854 66274 5906
rect 67230 5854 67282 5906
rect 68126 5854 68178 5906
rect 96126 5854 96178 5906
rect 97358 5854 97410 5906
rect 98030 5854 98082 5906
rect 113262 5854 113314 5906
rect 113934 5854 113986 5906
rect 115278 5854 115330 5906
rect 56366 5742 56418 5794
rect 56702 5742 56754 5794
rect 57598 5742 57650 5794
rect 57934 5742 57986 5794
rect 58494 5742 58546 5794
rect 58718 5742 58770 5794
rect 61966 5742 62018 5794
rect 62862 5742 62914 5794
rect 63310 5742 63362 5794
rect 64654 5742 64706 5794
rect 66446 5742 66498 5794
rect 67454 5742 67506 5794
rect 68350 5742 68402 5794
rect 79326 5742 79378 5794
rect 97246 5630 97298 5682
rect 97918 5630 97970 5682
rect 113150 5630 113202 5682
rect 113822 5630 113874 5682
rect 115166 5630 115218 5682
rect 23376 5462 23428 5514
rect 23480 5462 23532 5514
rect 23584 5462 23636 5514
rect 67700 5462 67752 5514
rect 67804 5462 67856 5514
rect 67908 5462 67960 5514
rect 112024 5462 112076 5514
rect 112128 5462 112180 5514
rect 112232 5462 112284 5514
rect 156348 5462 156400 5514
rect 156452 5462 156504 5514
rect 156556 5462 156608 5514
rect 86606 5294 86658 5346
rect 92318 5294 92370 5346
rect 94782 5294 94834 5346
rect 113710 5294 113762 5346
rect 49198 5182 49250 5234
rect 55470 5182 55522 5234
rect 56590 5182 56642 5234
rect 57486 5182 57538 5234
rect 58382 5182 58434 5234
rect 59278 5182 59330 5234
rect 60174 5182 60226 5234
rect 60622 5182 60674 5234
rect 61406 5182 61458 5234
rect 61742 5182 61794 5234
rect 62638 5182 62690 5234
rect 62974 5182 63026 5234
rect 64430 5182 64482 5234
rect 64654 5182 64706 5234
rect 65326 5182 65378 5234
rect 78990 5182 79042 5234
rect 79886 5182 79938 5234
rect 93214 5182 93266 5234
rect 33630 5070 33682 5122
rect 34302 5070 34354 5122
rect 35198 5070 35250 5122
rect 35534 5070 35586 5122
rect 48526 5070 48578 5122
rect 49758 5070 49810 5122
rect 50430 5070 50482 5122
rect 55694 5070 55746 5122
rect 56366 5070 56418 5122
rect 57262 5070 57314 5122
rect 58158 5070 58210 5122
rect 59054 5070 59106 5122
rect 66334 5070 66386 5122
rect 68238 5070 68290 5122
rect 68462 5070 68514 5122
rect 69246 5070 69298 5122
rect 70366 5070 70418 5122
rect 70702 5070 70754 5122
rect 75854 5070 75906 5122
rect 79102 5070 79154 5122
rect 79662 5070 79714 5122
rect 85934 5070 85986 5122
rect 86494 5070 86546 5122
rect 92430 5070 92482 5122
rect 96350 5070 96402 5122
rect 96574 5070 96626 5122
rect 98254 5070 98306 5122
rect 105982 5070 106034 5122
rect 106766 5070 106818 5122
rect 107662 5070 107714 5122
rect 112254 5070 112306 5122
rect 115614 5070 115666 5122
rect 118862 5070 118914 5122
rect 120542 5070 120594 5122
rect 59838 4958 59890 5010
rect 63534 4958 63586 5010
rect 67566 4958 67618 5010
rect 83358 4958 83410 5010
rect 94894 4958 94946 5010
rect 95566 4958 95618 5010
rect 96798 4958 96850 5010
rect 97470 4958 97522 5010
rect 98142 4958 98194 5010
rect 112366 4958 112418 5010
rect 113038 4958 113090 5010
rect 113598 4958 113650 5010
rect 114270 4958 114322 5010
rect 119646 4958 119698 5010
rect 120990 4958 121042 5010
rect 63646 4846 63698 4898
rect 65438 4846 65490 4898
rect 66334 4846 66386 4898
rect 67230 4846 67282 4898
rect 69806 4846 69858 4898
rect 80222 4846 80274 4898
rect 83022 4846 83074 4898
rect 84366 4846 84418 4898
rect 85822 4846 85874 4898
rect 96126 4846 96178 4898
rect 98814 4846 98866 4898
rect 105422 4846 105474 4898
rect 108110 4846 108162 4898
rect 114942 4846 114994 4898
rect 115726 4846 115778 4898
rect 118302 4846 118354 4898
rect 141374 4846 141426 4898
rect 45538 4678 45590 4730
rect 45642 4678 45694 4730
rect 45746 4678 45798 4730
rect 89862 4678 89914 4730
rect 89966 4678 90018 4730
rect 90070 4678 90122 4730
rect 134186 4678 134238 4730
rect 134290 4678 134342 4730
rect 134394 4678 134446 4730
rect 178510 4678 178562 4730
rect 178614 4678 178666 4730
rect 178718 4678 178770 4730
rect 36430 4510 36482 4562
rect 36878 4510 36930 4562
rect 51550 4510 51602 4562
rect 58382 4510 58434 4562
rect 62190 4510 62242 4562
rect 63534 4510 63586 4562
rect 78990 4510 79042 4562
rect 95902 4510 95954 4562
rect 97246 4510 97298 4562
rect 98030 4510 98082 4562
rect 113150 4510 113202 4562
rect 113934 4510 113986 4562
rect 114494 4510 114546 4562
rect 115278 4510 115330 4562
rect 115838 4510 115890 4562
rect 10670 4398 10722 4450
rect 26350 4398 26402 4450
rect 28030 4398 28082 4450
rect 33518 4398 33570 4450
rect 53230 4398 53282 4450
rect 54910 4398 54962 4450
rect 56702 4398 56754 4450
rect 57710 4398 57762 4450
rect 58270 4398 58322 4450
rect 62862 4398 62914 4450
rect 63422 4398 63474 4450
rect 65550 4398 65602 4450
rect 71150 4398 71202 4450
rect 72606 4398 72658 4450
rect 74286 4398 74338 4450
rect 74846 4398 74898 4450
rect 76190 4398 76242 4450
rect 79662 4398 79714 4450
rect 85822 4398 85874 4450
rect 93662 4398 93714 4450
rect 94670 4398 94722 4450
rect 96014 4398 96066 4450
rect 108110 4398 108162 4450
rect 109790 4398 109842 4450
rect 114606 4398 114658 4450
rect 121102 4398 121154 4450
rect 129054 4398 129106 4450
rect 129950 4398 130002 4450
rect 132750 4398 132802 4450
rect 133422 4398 133474 4450
rect 141262 4398 141314 4450
rect 141934 4398 141986 4450
rect 151790 4398 151842 4450
rect 153470 4398 153522 4450
rect 31278 4286 31330 4338
rect 32958 4286 33010 4338
rect 34414 4286 34466 4338
rect 35198 4286 35250 4338
rect 36094 4286 36146 4338
rect 49758 4286 49810 4338
rect 51214 4286 51266 4338
rect 56478 4286 56530 4338
rect 61182 4286 61234 4338
rect 64430 4286 64482 4338
rect 64654 4286 64706 4338
rect 66110 4286 66162 4338
rect 69358 4286 69410 4338
rect 70142 4286 70194 4338
rect 72270 4286 72322 4338
rect 73950 4286 74002 4338
rect 84030 4286 84082 4338
rect 85038 4286 85090 4338
rect 86494 4286 86546 4338
rect 92990 4286 93042 4338
rect 105758 4286 105810 4338
rect 107438 4286 107490 4338
rect 118750 4286 118802 4338
rect 120430 4286 120482 4338
rect 130734 4286 130786 4338
rect 132302 4286 132354 4338
rect 139358 4286 139410 4338
rect 140814 4286 140866 4338
rect 13022 4174 13074 4226
rect 28702 4174 28754 4226
rect 30830 4174 30882 4226
rect 32062 4174 32114 4226
rect 50318 4174 50370 4226
rect 54350 4174 54402 4226
rect 55806 4174 55858 4226
rect 59838 4174 59890 4226
rect 65774 4174 65826 4226
rect 66110 4174 66162 4226
rect 68462 4174 68514 4226
rect 69582 4174 69634 4226
rect 70478 4174 70530 4226
rect 71822 4174 71874 4226
rect 73502 4174 73554 4226
rect 75742 4174 75794 4226
rect 77086 4174 77138 4226
rect 78542 4174 78594 4226
rect 83694 4174 83746 4226
rect 84590 4174 84642 4226
rect 91422 4174 91474 4226
rect 92430 4174 92482 4226
rect 105198 4174 105250 4226
rect 106542 4174 106594 4226
rect 118190 4174 118242 4226
rect 119534 4174 119586 4226
rect 126926 4174 126978 4226
rect 127486 4174 127538 4226
rect 131406 4174 131458 4226
rect 139918 4174 139970 4226
rect 142606 4174 142658 4226
rect 150446 4174 150498 4226
rect 151006 4174 151058 4226
rect 93102 4062 93154 4114
rect 23376 3894 23428 3946
rect 23480 3894 23532 3946
rect 23584 3894 23636 3946
rect 67700 3894 67752 3946
rect 67804 3894 67856 3946
rect 67908 3894 67960 3946
rect 112024 3894 112076 3946
rect 112128 3894 112180 3946
rect 112232 3894 112284 3946
rect 156348 3894 156400 3946
rect 156452 3894 156504 3946
rect 156556 3894 156608 3946
rect 9662 3614 9714 3666
rect 28254 3614 28306 3666
rect 32510 3614 32562 3666
rect 34862 3614 34914 3666
rect 52782 3614 52834 3666
rect 54910 3614 54962 3666
rect 57486 3614 57538 3666
rect 57822 3614 57874 3666
rect 58382 3614 58434 3666
rect 58718 3614 58770 3666
rect 59278 3614 59330 3666
rect 59614 3614 59666 3666
rect 64654 3614 64706 3666
rect 64878 3614 64930 3666
rect 66894 3614 66946 3666
rect 68462 3614 68514 3666
rect 73390 3614 73442 3666
rect 75518 3614 75570 3666
rect 85710 3614 85762 3666
rect 90638 3614 90690 3666
rect 92766 3614 92818 3666
rect 94894 3614 94946 3666
rect 110574 3614 110626 3666
rect 121102 3614 121154 3666
rect 121550 3614 121602 3666
rect 130398 3614 130450 3666
rect 131966 3614 132018 3666
rect 140366 3614 140418 3666
rect 153918 3614 153970 3666
rect 12574 3502 12626 3554
rect 25342 3502 25394 3554
rect 29262 3502 29314 3554
rect 34078 3502 34130 3554
rect 35534 3502 35586 3554
rect 55694 3502 55746 3554
rect 57934 3502 57986 3554
rect 58158 3502 58210 3554
rect 62190 3502 62242 3554
rect 63758 3502 63810 3554
rect 65662 3502 65714 3554
rect 69134 3502 69186 3554
rect 70814 3502 70866 3554
rect 72606 3502 72658 3554
rect 81230 3502 81282 3554
rect 84926 3502 84978 3554
rect 86494 3502 86546 3554
rect 92094 3502 92146 3554
rect 105982 3502 106034 3554
rect 107774 3502 107826 3554
rect 119534 3502 119586 3554
rect 120542 3502 120594 3554
rect 127598 3502 127650 3554
rect 128270 3502 128322 3554
rect 131182 3502 131234 3554
rect 132862 3502 132914 3554
rect 139694 3502 139746 3554
rect 141262 3502 141314 3554
rect 151118 3502 151170 3554
rect 151790 3502 151842 3554
rect 11790 3390 11842 3442
rect 14254 3390 14306 3442
rect 26126 3390 26178 3442
rect 62078 3390 62130 3442
rect 62862 3390 62914 3442
rect 71598 3390 71650 3442
rect 76302 3390 76354 3442
rect 77310 3390 77362 3442
rect 78990 3390 79042 3442
rect 80222 3390 80274 3442
rect 80670 3390 80722 3442
rect 105534 3390 105586 3442
rect 108446 3390 108498 3442
rect 119758 3390 119810 3442
rect 142942 3390 142994 3442
rect 7310 3278 7362 3330
rect 13582 3278 13634 3330
rect 15150 3278 15202 3330
rect 17502 3278 17554 3330
rect 19630 3278 19682 3330
rect 21422 3278 21474 3330
rect 22990 3278 23042 3330
rect 24446 3278 24498 3330
rect 29710 3278 29762 3330
rect 31390 3278 31442 3330
rect 33182 3278 33234 3330
rect 36206 3278 36258 3330
rect 37102 3278 37154 3330
rect 38110 3278 38162 3330
rect 39790 3278 39842 3330
rect 41470 3278 41522 3330
rect 43150 3278 43202 3330
rect 44942 3278 44994 3330
rect 46510 3278 46562 3330
rect 48862 3278 48914 3330
rect 49870 3278 49922 3330
rect 51550 3278 51602 3330
rect 56702 3278 56754 3330
rect 60622 3278 60674 3330
rect 61406 3278 61458 3330
rect 63422 3278 63474 3330
rect 65662 3278 65714 3330
rect 66446 3278 66498 3330
rect 67566 3278 67618 3330
rect 68910 3278 68962 3330
rect 69806 3278 69858 3330
rect 70590 3278 70642 3330
rect 76638 3278 76690 3330
rect 77646 3278 77698 3330
rect 78206 3278 78258 3330
rect 79326 3278 79378 3330
rect 81790 3278 81842 3330
rect 82910 3278 82962 3330
rect 84366 3278 84418 3330
rect 87054 3278 87106 3330
rect 88062 3278 88114 3330
rect 89630 3278 89682 3330
rect 91086 3278 91138 3330
rect 96574 3278 96626 3330
rect 97246 3278 97298 3330
rect 98030 3278 98082 3330
rect 99822 3278 99874 3330
rect 101390 3278 101442 3330
rect 103742 3278 103794 3330
rect 104750 3278 104802 3330
rect 106430 3278 106482 3330
rect 111582 3278 111634 3330
rect 113150 3278 113202 3330
rect 115502 3278 115554 3330
rect 116510 3278 116562 3330
rect 118190 3278 118242 3330
rect 120318 3278 120370 3330
rect 123342 3278 123394 3330
rect 124910 3278 124962 3330
rect 126366 3278 126418 3330
rect 133310 3278 133362 3330
rect 133982 3278 134034 3330
rect 135102 3278 135154 3330
rect 136670 3278 136722 3330
rect 138126 3278 138178 3330
rect 141710 3278 141762 3330
rect 143390 3278 143442 3330
rect 145070 3278 145122 3330
rect 146862 3278 146914 3330
rect 148430 3278 148482 3330
rect 149886 3278 149938 3330
rect 155150 3278 155202 3330
rect 156830 3278 156882 3330
rect 158622 3278 158674 3330
rect 160190 3278 160242 3330
rect 162542 3278 162594 3330
rect 163550 3278 163602 3330
rect 165230 3278 165282 3330
rect 166910 3278 166962 3330
rect 168590 3278 168642 3330
rect 170382 3278 170434 3330
rect 171950 3278 172002 3330
rect 173070 3278 173122 3330
rect 174302 3278 174354 3330
rect 174974 3278 175026 3330
rect 45538 3110 45590 3162
rect 45642 3110 45694 3162
rect 45746 3110 45798 3162
rect 89862 3110 89914 3162
rect 89966 3110 90018 3162
rect 90070 3110 90122 3162
rect 134186 3110 134238 3162
rect 134290 3110 134342 3162
rect 134394 3110 134446 3162
rect 178510 3110 178562 3162
rect 178614 3110 178666 3162
rect 178718 3110 178770 3162
rect 69246 1710 69298 1762
rect 69806 1710 69858 1762
rect 77646 1710 77698 1762
rect 78206 1710 78258 1762
rect 81006 1710 81058 1762
rect 81790 1710 81842 1762
rect 86046 1710 86098 1762
rect 87054 1710 87106 1762
rect 96126 1710 96178 1762
rect 97246 1710 97298 1762
rect 102846 1710 102898 1762
rect 103742 1710 103794 1762
rect 114606 1710 114658 1762
rect 115502 1710 115554 1762
rect 119646 1710 119698 1762
rect 120318 1710 120370 1762
rect 133086 1710 133138 1762
rect 133982 1710 134034 1762
rect 161646 1710 161698 1762
rect 162542 1710 162594 1762
rect 173406 1710 173458 1762
rect 174302 1710 174354 1762
<< metal2 >>
rect 1344 19200 1456 20000
rect 2912 19200 3024 20000
rect 4480 19200 4592 20000
rect 6048 19200 6160 20000
rect 7616 19200 7728 20000
rect 9184 19200 9296 20000
rect 10752 19200 10864 20000
rect 12320 19200 12432 20000
rect 13888 19200 14000 20000
rect 15456 19200 15568 20000
rect 17024 19200 17136 20000
rect 18592 19200 18704 20000
rect 20160 19200 20272 20000
rect 21728 19200 21840 20000
rect 23296 19200 23408 20000
rect 24864 19200 24976 20000
rect 26432 19200 26544 20000
rect 28000 19200 28112 20000
rect 29568 19200 29680 20000
rect 31136 19200 31248 20000
rect 32704 19200 32816 20000
rect 34272 19200 34384 20000
rect 35840 19200 35952 20000
rect 37408 19200 37520 20000
rect 38976 19200 39088 20000
rect 40544 19200 40656 20000
rect 42112 19200 42224 20000
rect 43680 19200 43792 20000
rect 45248 19200 45360 20000
rect 46816 19200 46928 20000
rect 48384 19200 48496 20000
rect 49952 19200 50064 20000
rect 51520 19200 51632 20000
rect 53088 19200 53200 20000
rect 54656 19200 54768 20000
rect 56224 19200 56336 20000
rect 57792 19200 57904 20000
rect 59360 19200 59472 20000
rect 60928 19200 61040 20000
rect 62496 19200 62608 20000
rect 64064 19200 64176 20000
rect 65632 19200 65744 20000
rect 67200 19200 67312 20000
rect 68768 19200 68880 20000
rect 70336 19200 70448 20000
rect 71904 19200 72016 20000
rect 73472 19200 73584 20000
rect 75040 19200 75152 20000
rect 76608 19200 76720 20000
rect 78176 19200 78288 20000
rect 79744 19200 79856 20000
rect 81312 19200 81424 20000
rect 82880 19200 82992 20000
rect 84448 19200 84560 20000
rect 86016 19200 86128 20000
rect 87584 19200 87696 20000
rect 89152 19200 89264 20000
rect 90720 19200 90832 20000
rect 92288 19200 92400 20000
rect 93856 19200 93968 20000
rect 95424 19200 95536 20000
rect 96992 19200 97104 20000
rect 98560 19200 98672 20000
rect 100128 19200 100240 20000
rect 101696 19200 101808 20000
rect 103264 19200 103376 20000
rect 104832 19200 104944 20000
rect 106400 19200 106512 20000
rect 107968 19200 108080 20000
rect 109536 19200 109648 20000
rect 111104 19200 111216 20000
rect 112672 19200 112784 20000
rect 114240 19200 114352 20000
rect 115808 19200 115920 20000
rect 117376 19200 117488 20000
rect 118944 19200 119056 20000
rect 120512 19200 120624 20000
rect 122080 19200 122192 20000
rect 123648 19200 123760 20000
rect 125216 19200 125328 20000
rect 126784 19200 126896 20000
rect 128352 19200 128464 20000
rect 129920 19200 130032 20000
rect 131488 19200 131600 20000
rect 133056 19200 133168 20000
rect 134624 19200 134736 20000
rect 136192 19200 136304 20000
rect 137760 19200 137872 20000
rect 139328 19200 139440 20000
rect 140896 19200 141008 20000
rect 142464 19200 142576 20000
rect 144032 19200 144144 20000
rect 145600 19200 145712 20000
rect 147168 19200 147280 20000
rect 148736 19200 148848 20000
rect 150304 19200 150416 20000
rect 151872 19200 151984 20000
rect 153440 19200 153552 20000
rect 155008 19200 155120 20000
rect 156576 19200 156688 20000
rect 158144 19200 158256 20000
rect 159712 19200 159824 20000
rect 161280 19200 161392 20000
rect 162848 19200 162960 20000
rect 164416 19200 164528 20000
rect 165984 19200 166096 20000
rect 167552 19200 167664 20000
rect 169120 19200 169232 20000
rect 170688 19200 170800 20000
rect 172256 19200 172368 20000
rect 173824 19200 173936 20000
rect 175392 19200 175504 20000
rect 176960 19200 177072 20000
rect 178528 19200 178640 20000
rect 2940 15988 2996 19200
rect 3164 15988 3220 15998
rect 2940 15986 3220 15988
rect 2940 15934 3166 15986
rect 3218 15934 3220 15986
rect 2940 15932 3220 15934
rect 4508 15988 4564 19200
rect 4732 15988 4788 15998
rect 4508 15986 4788 15988
rect 4508 15934 4734 15986
rect 4786 15934 4788 15986
rect 4508 15932 4788 15934
rect 7644 15988 7700 19200
rect 9212 17668 9268 19200
rect 9212 17612 9716 17668
rect 7868 15988 7924 15998
rect 7644 15986 7924 15988
rect 7644 15934 7870 15986
rect 7922 15934 7924 15986
rect 7644 15932 7924 15934
rect 3164 15922 3220 15932
rect 4732 15922 4788 15932
rect 7868 15922 7924 15932
rect 9660 15986 9716 17612
rect 9660 15934 9662 15986
rect 9714 15934 9716 15986
rect 9660 15922 9716 15934
rect 12348 15988 12404 19200
rect 12572 15988 12628 15998
rect 12348 15986 12628 15988
rect 12348 15934 12574 15986
rect 12626 15934 12628 15986
rect 12348 15932 12628 15934
rect 13916 15988 13972 19200
rect 17052 17668 17108 19200
rect 17052 17612 17556 17668
rect 14140 15988 14196 15998
rect 13916 15986 14196 15988
rect 13916 15934 14142 15986
rect 14194 15934 14196 15986
rect 13916 15932 14196 15934
rect 12572 15922 12628 15932
rect 14140 15922 14196 15932
rect 17500 15986 17556 17612
rect 17500 15934 17502 15986
rect 17554 15934 17556 15986
rect 17500 15922 17556 15934
rect 18620 15988 18676 19200
rect 21756 16660 21812 19200
rect 23324 17444 23380 19200
rect 23212 17388 23380 17444
rect 21756 16604 22036 16660
rect 18844 15988 18900 15998
rect 18620 15986 18900 15988
rect 18620 15934 18846 15986
rect 18898 15934 18900 15986
rect 18620 15932 18900 15934
rect 18844 15922 18900 15932
rect 21980 15986 22036 16604
rect 21980 15934 21982 15986
rect 22034 15934 22036 15986
rect 21980 15922 22036 15934
rect 23212 15988 23268 17388
rect 23374 16492 23638 16502
rect 23430 16436 23478 16492
rect 23534 16436 23582 16492
rect 23374 16426 23638 16436
rect 23548 15988 23604 15998
rect 23212 15986 23604 15988
rect 23212 15934 23550 15986
rect 23602 15934 23604 15986
rect 23212 15932 23604 15934
rect 26460 15988 26516 19200
rect 26684 15988 26740 15998
rect 26460 15986 26740 15988
rect 26460 15934 26686 15986
rect 26738 15934 26740 15986
rect 26460 15932 26740 15934
rect 28028 15988 28084 19200
rect 28252 15988 28308 15998
rect 28028 15986 28308 15988
rect 28028 15934 28254 15986
rect 28306 15934 28308 15986
rect 28028 15932 28308 15934
rect 31164 15988 31220 19200
rect 32732 17668 32788 19200
rect 32732 17612 33236 17668
rect 31388 15988 31444 15998
rect 31164 15986 31444 15988
rect 31164 15934 31390 15986
rect 31442 15934 31444 15986
rect 31164 15932 31444 15934
rect 23548 15922 23604 15932
rect 26684 15922 26740 15932
rect 28252 15922 28308 15932
rect 31388 15922 31444 15932
rect 33180 15986 33236 17612
rect 33180 15934 33182 15986
rect 33234 15934 33236 15986
rect 33180 15922 33236 15934
rect 35868 15988 35924 19200
rect 36092 15988 36148 15998
rect 35868 15986 36148 15988
rect 35868 15934 36094 15986
rect 36146 15934 36148 15986
rect 35868 15932 36148 15934
rect 37436 15988 37492 19200
rect 40572 17668 40628 19200
rect 40572 17612 41076 17668
rect 37660 15988 37716 15998
rect 37436 15986 37716 15988
rect 37436 15934 37662 15986
rect 37714 15934 37716 15986
rect 37436 15932 37716 15934
rect 36092 15922 36148 15932
rect 37660 15922 37716 15932
rect 41020 15986 41076 17612
rect 41020 15934 41022 15986
rect 41074 15934 41076 15986
rect 41020 15922 41076 15934
rect 42140 15988 42196 19200
rect 45276 16660 45332 19200
rect 45276 16604 45556 16660
rect 42364 15988 42420 15998
rect 42140 15986 42420 15988
rect 42140 15934 42366 15986
rect 42418 15934 42420 15986
rect 42140 15932 42420 15934
rect 42364 15922 42420 15932
rect 45500 15986 45556 16604
rect 45500 15934 45502 15986
rect 45554 15934 45556 15986
rect 45500 15922 45556 15934
rect 46844 15988 46900 19200
rect 47068 15988 47124 15998
rect 46844 15986 47124 15988
rect 46844 15934 47070 15986
rect 47122 15934 47124 15986
rect 46844 15932 47124 15934
rect 49980 15988 50036 19200
rect 50204 15988 50260 15998
rect 49980 15986 50260 15988
rect 49980 15934 50206 15986
rect 50258 15934 50260 15986
rect 49980 15932 50260 15934
rect 51548 15988 51604 19200
rect 51772 15988 51828 15998
rect 51548 15986 51828 15988
rect 51548 15934 51774 15986
rect 51826 15934 51828 15986
rect 51548 15932 51828 15934
rect 54684 15988 54740 19200
rect 56252 17668 56308 19200
rect 56252 17612 56756 17668
rect 54908 15988 54964 15998
rect 54684 15986 54964 15988
rect 54684 15934 54910 15986
rect 54962 15934 54964 15986
rect 54684 15932 54964 15934
rect 47068 15922 47124 15932
rect 50204 15922 50260 15932
rect 51772 15922 51828 15932
rect 54908 15922 54964 15932
rect 56700 15986 56756 17612
rect 56700 15934 56702 15986
rect 56754 15934 56756 15986
rect 56700 15922 56756 15934
rect 59388 15988 59444 19200
rect 59612 15988 59668 15998
rect 59388 15986 59668 15988
rect 59388 15934 59614 15986
rect 59666 15934 59668 15986
rect 59388 15932 59668 15934
rect 60956 15988 61012 19200
rect 64092 17668 64148 19200
rect 64092 17612 64596 17668
rect 61180 15988 61236 15998
rect 60956 15986 61236 15988
rect 60956 15934 61182 15986
rect 61234 15934 61236 15986
rect 60956 15932 61236 15934
rect 59612 15922 59668 15932
rect 61180 15922 61236 15932
rect 64540 15986 64596 17612
rect 64540 15934 64542 15986
rect 64594 15934 64596 15986
rect 64540 15922 64596 15934
rect 65660 15988 65716 19200
rect 68796 16660 68852 19200
rect 68796 16604 69076 16660
rect 67698 16492 67962 16502
rect 67754 16436 67802 16492
rect 67858 16436 67906 16492
rect 67698 16426 67962 16436
rect 65884 15988 65940 15998
rect 65660 15986 65940 15988
rect 65660 15934 65886 15986
rect 65938 15934 65940 15986
rect 65660 15932 65940 15934
rect 65884 15922 65940 15932
rect 69020 15986 69076 16604
rect 69020 15934 69022 15986
rect 69074 15934 69076 15986
rect 69020 15922 69076 15934
rect 70364 15988 70420 19200
rect 70588 15988 70644 15998
rect 70364 15986 70644 15988
rect 70364 15934 70590 15986
rect 70642 15934 70644 15986
rect 70364 15932 70644 15934
rect 73500 15988 73556 19200
rect 73724 15988 73780 15998
rect 73500 15986 73780 15988
rect 73500 15934 73726 15986
rect 73778 15934 73780 15986
rect 73500 15932 73780 15934
rect 75068 15988 75124 19200
rect 75292 15988 75348 15998
rect 75068 15986 75348 15988
rect 75068 15934 75294 15986
rect 75346 15934 75348 15986
rect 75068 15932 75348 15934
rect 78204 15988 78260 19200
rect 79772 17668 79828 19200
rect 79772 17612 80276 17668
rect 78428 15988 78484 15998
rect 78204 15986 78484 15988
rect 78204 15934 78430 15986
rect 78482 15934 78484 15986
rect 78204 15932 78484 15934
rect 70588 15922 70644 15932
rect 73724 15922 73780 15932
rect 75292 15922 75348 15932
rect 78428 15922 78484 15932
rect 80220 15986 80276 17612
rect 80220 15934 80222 15986
rect 80274 15934 80276 15986
rect 80220 15922 80276 15934
rect 82908 15988 82964 19200
rect 83132 15988 83188 15998
rect 82908 15986 83188 15988
rect 82908 15934 83134 15986
rect 83186 15934 83188 15986
rect 82908 15932 83188 15934
rect 84476 15988 84532 19200
rect 87612 17668 87668 19200
rect 87612 17612 88116 17668
rect 84700 15988 84756 15998
rect 84476 15986 84756 15988
rect 84476 15934 84702 15986
rect 84754 15934 84756 15986
rect 84476 15932 84756 15934
rect 83132 15922 83188 15932
rect 84700 15922 84756 15932
rect 88060 15986 88116 17612
rect 88060 15934 88062 15986
rect 88114 15934 88116 15986
rect 88060 15922 88116 15934
rect 89180 15988 89236 19200
rect 92316 16660 92372 19200
rect 92316 16604 92596 16660
rect 89404 15988 89460 15998
rect 89180 15986 89460 15988
rect 89180 15934 89406 15986
rect 89458 15934 89460 15986
rect 89180 15932 89460 15934
rect 89404 15922 89460 15932
rect 92540 15986 92596 16604
rect 92540 15934 92542 15986
rect 92594 15934 92596 15986
rect 92540 15922 92596 15934
rect 93884 15988 93940 19200
rect 94108 15988 94164 15998
rect 93884 15986 94164 15988
rect 93884 15934 94110 15986
rect 94162 15934 94164 15986
rect 93884 15932 94164 15934
rect 97020 15988 97076 19200
rect 97244 15988 97300 15998
rect 97020 15986 97300 15988
rect 97020 15934 97246 15986
rect 97298 15934 97300 15986
rect 97020 15932 97300 15934
rect 98588 15988 98644 19200
rect 98812 15988 98868 15998
rect 98588 15986 98868 15988
rect 98588 15934 98814 15986
rect 98866 15934 98868 15986
rect 98588 15932 98868 15934
rect 101724 15988 101780 19200
rect 103292 17668 103348 19200
rect 103292 17612 103796 17668
rect 101948 15988 102004 15998
rect 101724 15986 102004 15988
rect 101724 15934 101950 15986
rect 102002 15934 102004 15986
rect 101724 15932 102004 15934
rect 94108 15922 94164 15932
rect 97244 15922 97300 15932
rect 98812 15922 98868 15932
rect 101948 15922 102004 15932
rect 103740 15986 103796 17612
rect 103740 15934 103742 15986
rect 103794 15934 103796 15986
rect 103740 15922 103796 15934
rect 106428 15988 106484 19200
rect 106652 15988 106708 15998
rect 106428 15986 106708 15988
rect 106428 15934 106654 15986
rect 106706 15934 106708 15986
rect 106428 15932 106708 15934
rect 107996 15988 108052 19200
rect 111132 17668 111188 19200
rect 111132 17612 111636 17668
rect 108220 15988 108276 15998
rect 107996 15986 108276 15988
rect 107996 15934 108222 15986
rect 108274 15934 108276 15986
rect 107996 15932 108276 15934
rect 106652 15922 106708 15932
rect 108220 15922 108276 15932
rect 111580 15986 111636 17612
rect 112022 16492 112286 16502
rect 112078 16436 112126 16492
rect 112182 16436 112230 16492
rect 112022 16426 112286 16436
rect 111580 15934 111582 15986
rect 111634 15934 111636 15986
rect 111580 15922 111636 15934
rect 112700 15988 112756 19200
rect 115836 16660 115892 19200
rect 115836 16604 116116 16660
rect 112924 15988 112980 15998
rect 112700 15986 112980 15988
rect 112700 15934 112926 15986
rect 112978 15934 112980 15986
rect 112700 15932 112980 15934
rect 112924 15922 112980 15932
rect 116060 15986 116116 16604
rect 116060 15934 116062 15986
rect 116114 15934 116116 15986
rect 116060 15922 116116 15934
rect 117404 15988 117460 19200
rect 117628 15988 117684 15998
rect 117404 15986 117684 15988
rect 117404 15934 117630 15986
rect 117682 15934 117684 15986
rect 117404 15932 117684 15934
rect 120540 15988 120596 19200
rect 120764 15988 120820 15998
rect 120540 15986 120820 15988
rect 120540 15934 120766 15986
rect 120818 15934 120820 15986
rect 120540 15932 120820 15934
rect 122108 15988 122164 19200
rect 122332 15988 122388 15998
rect 122108 15986 122388 15988
rect 122108 15934 122334 15986
rect 122386 15934 122388 15986
rect 122108 15932 122388 15934
rect 125244 15988 125300 19200
rect 126812 17668 126868 19200
rect 126812 17612 127316 17668
rect 125468 15988 125524 15998
rect 125244 15986 125524 15988
rect 125244 15934 125470 15986
rect 125522 15934 125524 15986
rect 125244 15932 125524 15934
rect 117628 15922 117684 15932
rect 120764 15922 120820 15932
rect 122332 15922 122388 15932
rect 125468 15922 125524 15932
rect 127260 15986 127316 17612
rect 127260 15934 127262 15986
rect 127314 15934 127316 15986
rect 127260 15922 127316 15934
rect 129948 15988 130004 19200
rect 130172 15988 130228 15998
rect 129948 15986 130228 15988
rect 129948 15934 130174 15986
rect 130226 15934 130228 15986
rect 129948 15932 130228 15934
rect 131516 15988 131572 19200
rect 134652 17668 134708 19200
rect 134652 17612 135156 17668
rect 131740 15988 131796 15998
rect 131516 15986 131796 15988
rect 131516 15934 131742 15986
rect 131794 15934 131796 15986
rect 131516 15932 131796 15934
rect 130172 15922 130228 15932
rect 131740 15922 131796 15932
rect 135100 15986 135156 17612
rect 135100 15934 135102 15986
rect 135154 15934 135156 15986
rect 135100 15922 135156 15934
rect 136220 15988 136276 19200
rect 139356 16660 139412 19200
rect 139356 16604 139636 16660
rect 136444 15988 136500 15998
rect 136220 15986 136500 15988
rect 136220 15934 136446 15986
rect 136498 15934 136500 15986
rect 136220 15932 136500 15934
rect 136444 15922 136500 15932
rect 139580 15986 139636 16604
rect 139580 15934 139582 15986
rect 139634 15934 139636 15986
rect 139580 15922 139636 15934
rect 140924 15988 140980 19200
rect 141148 15988 141204 15998
rect 140924 15986 141204 15988
rect 140924 15934 141150 15986
rect 141202 15934 141204 15986
rect 140924 15932 141204 15934
rect 144060 15988 144116 19200
rect 144284 15988 144340 15998
rect 144060 15986 144340 15988
rect 144060 15934 144286 15986
rect 144338 15934 144340 15986
rect 144060 15932 144340 15934
rect 145628 15988 145684 19200
rect 145852 15988 145908 15998
rect 145628 15986 145908 15988
rect 145628 15934 145854 15986
rect 145906 15934 145908 15986
rect 145628 15932 145908 15934
rect 148764 15988 148820 19200
rect 150332 17668 150388 19200
rect 150332 17612 150836 17668
rect 148988 15988 149044 15998
rect 148764 15986 149044 15988
rect 148764 15934 148990 15986
rect 149042 15934 149044 15986
rect 148764 15932 149044 15934
rect 141148 15922 141204 15932
rect 144284 15922 144340 15932
rect 145852 15922 145908 15932
rect 148988 15922 149044 15932
rect 150780 15986 150836 17612
rect 150780 15934 150782 15986
rect 150834 15934 150836 15986
rect 150780 15922 150836 15934
rect 153468 15988 153524 19200
rect 153692 15988 153748 15998
rect 153468 15986 153748 15988
rect 153468 15934 153694 15986
rect 153746 15934 153748 15986
rect 153468 15932 153748 15934
rect 155036 15988 155092 19200
rect 158172 17668 158228 19200
rect 158172 17612 158676 17668
rect 156346 16492 156610 16502
rect 156402 16436 156450 16492
rect 156506 16436 156554 16492
rect 156346 16426 156610 16436
rect 155260 15988 155316 15998
rect 155036 15986 155316 15988
rect 155036 15934 155262 15986
rect 155314 15934 155316 15986
rect 155036 15932 155316 15934
rect 153692 15922 153748 15932
rect 155260 15922 155316 15932
rect 158620 15986 158676 17612
rect 158620 15934 158622 15986
rect 158674 15934 158676 15986
rect 158620 15922 158676 15934
rect 159740 15988 159796 19200
rect 162876 16660 162932 19200
rect 162876 16604 163156 16660
rect 159964 15988 160020 15998
rect 159740 15986 160020 15988
rect 159740 15934 159966 15986
rect 160018 15934 160020 15986
rect 159740 15932 160020 15934
rect 159964 15922 160020 15932
rect 163100 15986 163156 16604
rect 163100 15934 163102 15986
rect 163154 15934 163156 15986
rect 163100 15922 163156 15934
rect 164444 15988 164500 19200
rect 164668 15988 164724 15998
rect 164444 15986 164724 15988
rect 164444 15934 164670 15986
rect 164722 15934 164724 15986
rect 164444 15932 164724 15934
rect 167580 15988 167636 19200
rect 167804 15988 167860 15998
rect 167580 15986 167860 15988
rect 167580 15934 167806 15986
rect 167858 15934 167860 15986
rect 167580 15932 167860 15934
rect 169148 15988 169204 19200
rect 169372 15988 169428 15998
rect 169148 15986 169428 15988
rect 169148 15934 169374 15986
rect 169426 15934 169428 15986
rect 169148 15932 169428 15934
rect 172284 15988 172340 19200
rect 173852 17668 173908 19200
rect 173852 17612 174356 17668
rect 172508 15988 172564 15998
rect 172284 15986 172564 15988
rect 172284 15934 172510 15986
rect 172562 15934 172564 15986
rect 172284 15932 172564 15934
rect 164668 15922 164724 15932
rect 167804 15922 167860 15932
rect 169372 15922 169428 15932
rect 172508 15922 172564 15932
rect 174300 15986 174356 17612
rect 174300 15934 174302 15986
rect 174354 15934 174356 15986
rect 174300 15922 174356 15934
rect 176988 15988 177044 19200
rect 178556 17444 178612 19200
rect 178108 17388 178612 17444
rect 177212 15988 177268 15998
rect 176988 15986 177268 15988
rect 176988 15934 177214 15986
rect 177266 15934 177268 15986
rect 176988 15932 177268 15934
rect 177212 15922 177268 15932
rect 45536 15708 45800 15718
rect 45592 15652 45640 15708
rect 45696 15652 45744 15708
rect 45536 15642 45800 15652
rect 89860 15708 90124 15718
rect 89916 15652 89964 15708
rect 90020 15652 90068 15708
rect 89860 15642 90124 15652
rect 134184 15708 134448 15718
rect 134240 15652 134288 15708
rect 134344 15652 134392 15708
rect 134184 15642 134448 15652
rect 178108 15538 178164 17388
rect 178508 15708 178772 15718
rect 178564 15652 178612 15708
rect 178668 15652 178716 15708
rect 178508 15642 178772 15652
rect 178108 15486 178110 15538
rect 178162 15486 178164 15538
rect 178108 15474 178164 15486
rect 23374 14924 23638 14934
rect 23430 14868 23478 14924
rect 23534 14868 23582 14924
rect 23374 14858 23638 14868
rect 67698 14924 67962 14934
rect 67754 14868 67802 14924
rect 67858 14868 67906 14924
rect 67698 14858 67962 14868
rect 112022 14924 112286 14934
rect 112078 14868 112126 14924
rect 112182 14868 112230 14924
rect 112022 14858 112286 14868
rect 156346 14924 156610 14934
rect 156402 14868 156450 14924
rect 156506 14868 156554 14924
rect 156346 14858 156610 14868
rect 45536 14140 45800 14150
rect 45592 14084 45640 14140
rect 45696 14084 45744 14140
rect 45536 14074 45800 14084
rect 89860 14140 90124 14150
rect 89916 14084 89964 14140
rect 90020 14084 90068 14140
rect 89860 14074 90124 14084
rect 134184 14140 134448 14150
rect 134240 14084 134288 14140
rect 134344 14084 134392 14140
rect 134184 14074 134448 14084
rect 178508 14140 178772 14150
rect 178564 14084 178612 14140
rect 178668 14084 178716 14140
rect 178508 14074 178772 14084
rect 23374 13356 23638 13366
rect 23430 13300 23478 13356
rect 23534 13300 23582 13356
rect 23374 13290 23638 13300
rect 67698 13356 67962 13366
rect 67754 13300 67802 13356
rect 67858 13300 67906 13356
rect 67698 13290 67962 13300
rect 112022 13356 112286 13366
rect 112078 13300 112126 13356
rect 112182 13300 112230 13356
rect 112022 13290 112286 13300
rect 156346 13356 156610 13366
rect 156402 13300 156450 13356
rect 156506 13300 156554 13356
rect 156346 13290 156610 13300
rect 45536 12572 45800 12582
rect 45592 12516 45640 12572
rect 45696 12516 45744 12572
rect 45536 12506 45800 12516
rect 89860 12572 90124 12582
rect 89916 12516 89964 12572
rect 90020 12516 90068 12572
rect 89860 12506 90124 12516
rect 134184 12572 134448 12582
rect 134240 12516 134288 12572
rect 134344 12516 134392 12572
rect 134184 12506 134448 12516
rect 178508 12572 178772 12582
rect 178564 12516 178612 12572
rect 178668 12516 178716 12572
rect 178508 12506 178772 12516
rect 23374 11788 23638 11798
rect 23430 11732 23478 11788
rect 23534 11732 23582 11788
rect 23374 11722 23638 11732
rect 67698 11788 67962 11798
rect 67754 11732 67802 11788
rect 67858 11732 67906 11788
rect 67698 11722 67962 11732
rect 112022 11788 112286 11798
rect 112078 11732 112126 11788
rect 112182 11732 112230 11788
rect 112022 11722 112286 11732
rect 156346 11788 156610 11798
rect 156402 11732 156450 11788
rect 156506 11732 156554 11788
rect 156346 11722 156610 11732
rect 45536 11004 45800 11014
rect 45592 10948 45640 11004
rect 45696 10948 45744 11004
rect 45536 10938 45800 10948
rect 89860 11004 90124 11014
rect 89916 10948 89964 11004
rect 90020 10948 90068 11004
rect 89860 10938 90124 10948
rect 134184 11004 134448 11014
rect 134240 10948 134288 11004
rect 134344 10948 134392 11004
rect 134184 10938 134448 10948
rect 178508 11004 178772 11014
rect 178564 10948 178612 11004
rect 178668 10948 178716 11004
rect 178508 10938 178772 10948
rect 23374 10220 23638 10230
rect 23430 10164 23478 10220
rect 23534 10164 23582 10220
rect 23374 10154 23638 10164
rect 67698 10220 67962 10230
rect 67754 10164 67802 10220
rect 67858 10164 67906 10220
rect 67698 10154 67962 10164
rect 112022 10220 112286 10230
rect 112078 10164 112126 10220
rect 112182 10164 112230 10220
rect 112022 10154 112286 10164
rect 156346 10220 156610 10230
rect 156402 10164 156450 10220
rect 156506 10164 156554 10220
rect 156346 10154 156610 10164
rect 45536 9436 45800 9446
rect 45592 9380 45640 9436
rect 45696 9380 45744 9436
rect 45536 9370 45800 9380
rect 89860 9436 90124 9446
rect 89916 9380 89964 9436
rect 90020 9380 90068 9436
rect 89860 9370 90124 9380
rect 134184 9436 134448 9446
rect 134240 9380 134288 9436
rect 134344 9380 134392 9436
rect 134184 9370 134448 9380
rect 178508 9436 178772 9446
rect 178564 9380 178612 9436
rect 178668 9380 178716 9436
rect 178508 9370 178772 9380
rect 23374 8652 23638 8662
rect 23430 8596 23478 8652
rect 23534 8596 23582 8652
rect 23374 8586 23638 8596
rect 67698 8652 67962 8662
rect 67754 8596 67802 8652
rect 67858 8596 67906 8652
rect 67698 8586 67962 8596
rect 112022 8652 112286 8662
rect 112078 8596 112126 8652
rect 112182 8596 112230 8652
rect 112022 8586 112286 8596
rect 156346 8652 156610 8662
rect 156402 8596 156450 8652
rect 156506 8596 156554 8652
rect 156346 8586 156610 8596
rect 45536 7868 45800 7878
rect 45592 7812 45640 7868
rect 45696 7812 45744 7868
rect 45536 7802 45800 7812
rect 89860 7868 90124 7878
rect 89916 7812 89964 7868
rect 90020 7812 90068 7868
rect 89860 7802 90124 7812
rect 134184 7868 134448 7878
rect 134240 7812 134288 7868
rect 134344 7812 134392 7868
rect 134184 7802 134448 7812
rect 178508 7868 178772 7878
rect 178564 7812 178612 7868
rect 178668 7812 178716 7868
rect 178508 7802 178772 7812
rect 57932 7362 57988 7374
rect 57932 7310 57934 7362
rect 57986 7310 57988 7362
rect 23374 7084 23638 7094
rect 23430 7028 23478 7084
rect 23534 7028 23582 7084
rect 23374 7018 23638 7028
rect 57484 6578 57540 6590
rect 57484 6526 57486 6578
rect 57538 6526 57540 6578
rect 51548 6468 51604 6478
rect 45536 6300 45800 6310
rect 45592 6244 45640 6300
rect 45696 6244 45744 6300
rect 45536 6234 45800 6244
rect 23374 5516 23638 5526
rect 23430 5460 23478 5516
rect 23534 5460 23582 5516
rect 23374 5450 23638 5460
rect 49196 5236 49252 5246
rect 33628 5122 33684 5134
rect 33628 5070 33630 5122
rect 33682 5070 33684 5122
rect 10668 4452 10724 4462
rect 10444 4450 10724 4452
rect 10444 4398 10670 4450
rect 10722 4398 10724 4450
rect 10444 4396 10724 4398
rect 9660 3780 9716 3790
rect 9660 3666 9716 3724
rect 9660 3614 9662 3666
rect 9714 3614 9716 3666
rect 9660 3602 9716 3614
rect 7308 3332 7364 3342
rect 7084 3330 7364 3332
rect 7084 3278 7310 3330
rect 7362 3278 7364 3330
rect 7084 3276 7364 3278
rect 7084 800 7140 3276
rect 7308 3266 7364 3276
rect 10444 800 10500 4396
rect 10668 4386 10724 4396
rect 26348 4450 26404 4462
rect 28028 4452 28084 4462
rect 26348 4398 26350 4450
rect 26402 4398 26404 4450
rect 13020 4226 13076 4238
rect 13020 4174 13022 4226
rect 13074 4174 13076 4226
rect 12572 3556 12628 3566
rect 12572 3462 12628 3500
rect 13020 3556 13076 4174
rect 23374 3948 23638 3958
rect 23430 3892 23478 3948
rect 23534 3892 23582 3948
rect 23374 3882 23638 3892
rect 13020 3490 13076 3500
rect 25340 3556 25396 3566
rect 25340 3462 25396 3500
rect 11788 3444 11844 3454
rect 11788 3350 11844 3388
rect 14252 3444 14308 3454
rect 12684 3332 12740 3342
rect 12684 800 12740 3276
rect 13580 3332 13636 3342
rect 13580 3238 13636 3276
rect 14252 2996 14308 3388
rect 26124 3444 26180 3454
rect 26124 3350 26180 3388
rect 15148 3332 15204 3342
rect 17500 3332 17556 3342
rect 19628 3332 19684 3342
rect 21420 3332 21476 3342
rect 22988 3332 23044 3342
rect 14252 2930 14308 2940
rect 14924 3330 15204 3332
rect 14924 3278 15150 3330
rect 15202 3278 15204 3330
rect 14924 3276 15204 3278
rect 14924 800 14980 3276
rect 15148 3266 15204 3276
rect 17164 3330 17556 3332
rect 17164 3278 17502 3330
rect 17554 3278 17556 3330
rect 17164 3276 17556 3278
rect 17164 800 17220 3276
rect 17500 3266 17556 3276
rect 19404 3330 19684 3332
rect 19404 3278 19630 3330
rect 19682 3278 19684 3330
rect 19404 3276 19684 3278
rect 19404 800 19460 3276
rect 19628 3266 19684 3276
rect 21084 3330 21476 3332
rect 21084 3278 21422 3330
rect 21474 3278 21476 3330
rect 21084 3276 21476 3278
rect 21084 800 21140 3276
rect 21420 3266 21476 3276
rect 22764 3330 23044 3332
rect 22764 3278 22990 3330
rect 23042 3278 23044 3330
rect 22764 3276 23044 3278
rect 22764 800 22820 3276
rect 22988 3266 23044 3276
rect 24444 3330 24500 3342
rect 24444 3278 24446 3330
rect 24498 3278 24500 3330
rect 24444 800 24500 3278
rect 26348 980 26404 4398
rect 26124 924 26404 980
rect 27804 4450 28084 4452
rect 27804 4398 28030 4450
rect 28082 4398 28084 4450
rect 27804 4396 28084 4398
rect 26124 800 26180 924
rect 27804 800 27860 4396
rect 28028 4386 28084 4396
rect 32956 4452 33012 4462
rect 31276 4338 31332 4350
rect 31276 4286 31278 4338
rect 31330 4286 31332 4338
rect 28700 4226 28756 4238
rect 28700 4174 28702 4226
rect 28754 4174 28756 4226
rect 28252 3668 28308 3678
rect 28252 3574 28308 3612
rect 28700 3444 28756 4174
rect 30828 4226 30884 4238
rect 30828 4174 30830 4226
rect 30882 4174 30884 4226
rect 30828 3780 30884 4174
rect 30828 3714 30884 3724
rect 31276 3780 31332 4286
rect 32956 4338 33012 4396
rect 33516 4452 33572 4462
rect 33516 4358 33572 4396
rect 32956 4286 32958 4338
rect 33010 4286 33012 4338
rect 32956 4274 33012 4286
rect 32060 4228 32116 4238
rect 32060 4134 32116 4172
rect 33628 4004 33684 5070
rect 34300 5122 34356 5134
rect 34300 5070 34302 5122
rect 34354 5070 34356 5122
rect 34300 4228 34356 5070
rect 35196 5124 35252 5134
rect 35196 5030 35252 5068
rect 35532 5124 35588 5134
rect 35532 4452 35588 5068
rect 36876 5124 36932 5134
rect 36428 4564 36484 4574
rect 36876 4564 36932 5068
rect 48524 5124 48580 5134
rect 48524 5030 48580 5068
rect 45536 4732 45800 4742
rect 45592 4676 45640 4732
rect 45696 4676 45744 4732
rect 45536 4666 45800 4676
rect 34300 4162 34356 4172
rect 34412 4338 34468 4350
rect 34412 4286 34414 4338
rect 34466 4286 34468 4338
rect 33628 3938 33684 3948
rect 34412 4004 34468 4286
rect 34412 3938 34468 3948
rect 34860 4340 34916 4350
rect 31276 3714 31332 3724
rect 31948 3780 32004 3790
rect 32004 3724 32564 3780
rect 31948 3714 32004 3724
rect 32508 3668 32564 3724
rect 32508 3574 32564 3612
rect 34076 3668 34132 3678
rect 29260 3556 29316 3566
rect 29260 3462 29316 3500
rect 34076 3554 34132 3612
rect 34860 3666 34916 4284
rect 35196 4340 35252 4350
rect 35196 4246 35252 4284
rect 34860 3614 34862 3666
rect 34914 3614 34916 3666
rect 34860 3602 34916 3614
rect 34076 3502 34078 3554
rect 34130 3502 34132 3554
rect 34076 3490 34132 3502
rect 35532 3554 35588 4396
rect 36092 4562 36932 4564
rect 36092 4510 36430 4562
rect 36482 4510 36878 4562
rect 36930 4510 36932 4562
rect 36092 4508 36932 4510
rect 36092 4338 36148 4508
rect 36428 4498 36484 4508
rect 36876 4498 36932 4508
rect 36092 4286 36094 4338
rect 36146 4286 36148 4338
rect 36092 4274 36148 4286
rect 49196 4340 49252 5180
rect 49196 4274 49252 4284
rect 49756 5122 49812 5134
rect 49756 5070 49758 5122
rect 49810 5070 49812 5122
rect 49756 4338 49812 5070
rect 50428 5124 50484 5134
rect 50428 5030 50484 5068
rect 51548 5124 51604 6412
rect 56364 5794 56420 5806
rect 56364 5742 56366 5794
rect 56418 5742 56420 5794
rect 55468 5348 55524 5358
rect 55468 5234 55524 5292
rect 55468 5182 55470 5234
rect 55522 5182 55524 5234
rect 55468 5170 55524 5182
rect 51548 4562 51604 5068
rect 55692 5124 55748 5134
rect 55692 5030 55748 5068
rect 56364 5124 56420 5742
rect 56700 5794 56756 5806
rect 56700 5742 56702 5794
rect 56754 5742 56756 5794
rect 56700 5348 56756 5742
rect 57484 5796 57540 6526
rect 57820 6580 57876 6590
rect 57932 6580 57988 7310
rect 57820 6578 57988 6580
rect 57820 6526 57822 6578
rect 57874 6526 57988 6578
rect 57820 6524 57988 6526
rect 58268 7362 58324 7374
rect 58268 7310 58270 7362
rect 58322 7310 58324 7362
rect 58268 6580 58324 7310
rect 65436 7362 65492 7374
rect 65436 7310 65438 7362
rect 65490 7310 65492 7362
rect 64092 6804 64148 6814
rect 64540 6804 64596 6814
rect 64092 6710 64148 6748
rect 64428 6748 64540 6804
rect 58380 6580 58436 6590
rect 58268 6578 58436 6580
rect 58268 6526 58382 6578
rect 58434 6526 58436 6578
rect 58268 6524 58436 6526
rect 57820 6514 57876 6524
rect 57596 5796 57652 5806
rect 57484 5794 57652 5796
rect 57484 5742 57598 5794
rect 57650 5742 57652 5794
rect 57484 5740 57652 5742
rect 56588 5236 56644 5246
rect 56700 5236 56756 5292
rect 56588 5234 56756 5236
rect 56588 5182 56590 5234
rect 56642 5182 56756 5234
rect 56588 5180 56756 5182
rect 56588 5170 56644 5180
rect 56420 5068 56532 5124
rect 56364 5058 56420 5068
rect 51548 4510 51550 4562
rect 51602 4510 51604 4562
rect 49756 4286 49758 4338
rect 49810 4286 49812 4338
rect 49756 3668 49812 4286
rect 51212 4340 51268 4350
rect 51548 4340 51604 4510
rect 53228 4452 53284 4462
rect 54908 4452 54964 4462
rect 51212 4338 51604 4340
rect 51212 4286 51214 4338
rect 51266 4286 51604 4338
rect 51212 4284 51604 4286
rect 53004 4450 53284 4452
rect 53004 4398 53230 4450
rect 53282 4398 53284 4450
rect 53004 4396 53284 4398
rect 51212 4274 51268 4284
rect 50316 4228 50372 4238
rect 50316 4134 50372 4172
rect 49756 3602 49812 3612
rect 52780 3668 52836 3678
rect 52780 3574 52836 3612
rect 35532 3502 35534 3554
rect 35586 3502 35588 3554
rect 35532 3490 35588 3502
rect 28700 2884 28756 3388
rect 29708 3332 29764 3342
rect 31388 3332 31444 3342
rect 33180 3332 33236 3342
rect 28700 2818 28756 2828
rect 29484 3330 29764 3332
rect 29484 3278 29710 3330
rect 29762 3278 29764 3330
rect 29484 3276 29764 3278
rect 29484 800 29540 3276
rect 29708 3266 29764 3276
rect 31164 3330 31444 3332
rect 31164 3278 31390 3330
rect 31442 3278 31444 3330
rect 31164 3276 31444 3278
rect 31164 800 31220 3276
rect 31388 3266 31444 3276
rect 32844 3330 33236 3332
rect 32844 3278 33182 3330
rect 33234 3278 33236 3330
rect 32844 3276 33236 3278
rect 32844 800 32900 3276
rect 33180 3266 33236 3276
rect 34524 3332 34580 3342
rect 34524 800 34580 3276
rect 36204 3332 36260 3342
rect 36204 3238 36260 3276
rect 37100 3330 37156 3342
rect 38108 3332 38164 3342
rect 39788 3332 39844 3342
rect 41468 3332 41524 3342
rect 43148 3332 43204 3342
rect 44940 3332 44996 3342
rect 46508 3332 46564 3342
rect 37100 3278 37102 3330
rect 37154 3278 37156 3330
rect 36204 1764 36260 1774
rect 36204 800 36260 1708
rect 37100 1764 37156 3278
rect 37100 1698 37156 1708
rect 37884 3330 38164 3332
rect 37884 3278 38110 3330
rect 38162 3278 38164 3330
rect 37884 3276 38164 3278
rect 37884 800 37940 3276
rect 38108 3266 38164 3276
rect 39564 3330 39844 3332
rect 39564 3278 39790 3330
rect 39842 3278 39844 3330
rect 39564 3276 39844 3278
rect 39564 800 39620 3276
rect 39788 3266 39844 3276
rect 41244 3330 41524 3332
rect 41244 3278 41470 3330
rect 41522 3278 41524 3330
rect 41244 3276 41524 3278
rect 41244 800 41300 3276
rect 41468 3266 41524 3276
rect 42924 3330 43204 3332
rect 42924 3278 43150 3330
rect 43202 3278 43204 3330
rect 42924 3276 43204 3278
rect 42924 800 42980 3276
rect 43148 3266 43204 3276
rect 44604 3330 44996 3332
rect 44604 3278 44942 3330
rect 44994 3278 44996 3330
rect 44604 3276 44996 3278
rect 44604 800 44660 3276
rect 44940 3266 44996 3276
rect 46284 3330 46564 3332
rect 46284 3278 46510 3330
rect 46562 3278 46564 3330
rect 46284 3276 46564 3278
rect 45536 3164 45800 3174
rect 45592 3108 45640 3164
rect 45696 3108 45744 3164
rect 45536 3098 45800 3108
rect 46284 800 46340 3276
rect 46508 3266 46564 3276
rect 47964 3332 48020 3342
rect 47964 800 48020 3276
rect 48860 3332 48916 3342
rect 49868 3332 49924 3342
rect 51548 3332 51604 3342
rect 48860 3238 48916 3276
rect 49644 3330 49924 3332
rect 49644 3278 49870 3330
rect 49922 3278 49924 3330
rect 49644 3276 49924 3278
rect 49644 800 49700 3276
rect 49868 3266 49924 3276
rect 51324 3330 51604 3332
rect 51324 3278 51550 3330
rect 51602 3278 51604 3330
rect 51324 3276 51604 3278
rect 51324 800 51380 3276
rect 51548 3266 51604 3276
rect 53004 800 53060 4396
rect 53228 4386 53284 4396
rect 54684 4450 54964 4452
rect 54684 4398 54910 4450
rect 54962 4398 54964 4450
rect 54684 4396 54964 4398
rect 54348 4226 54404 4238
rect 54348 4174 54350 4226
rect 54402 4174 54404 4226
rect 54348 3668 54404 4174
rect 54348 3602 54404 3612
rect 54684 800 54740 4396
rect 54908 4386 54964 4396
rect 56476 4338 56532 5068
rect 56700 4450 56756 5180
rect 57484 5348 57540 5358
rect 57484 5234 57540 5292
rect 57484 5182 57486 5234
rect 57538 5182 57540 5234
rect 57260 5124 57316 5162
rect 57260 5058 57316 5068
rect 56700 4398 56702 4450
rect 56754 4398 56756 4450
rect 56700 4386 56756 4398
rect 56476 4286 56478 4338
rect 56530 4286 56532 4338
rect 56476 4274 56532 4286
rect 55804 4228 55860 4238
rect 55692 4172 55804 4228
rect 54908 4116 54964 4126
rect 54908 3668 54964 4060
rect 54908 3574 54964 3612
rect 55692 3556 55748 4172
rect 55804 4134 55860 4172
rect 57484 3666 57540 5182
rect 57596 5124 57652 5740
rect 57932 5794 57988 6524
rect 57932 5742 57934 5794
rect 57986 5742 57988 5794
rect 57932 5348 57988 5742
rect 58380 5796 58436 6524
rect 58716 6578 58772 6590
rect 58716 6526 58718 6578
rect 58770 6526 58772 6578
rect 58492 5796 58548 5806
rect 58380 5794 58548 5796
rect 58380 5742 58494 5794
rect 58546 5742 58548 5794
rect 58380 5740 58548 5742
rect 57932 5282 57988 5292
rect 58380 5348 58436 5358
rect 58380 5234 58436 5292
rect 58380 5182 58382 5234
rect 58434 5182 58436 5234
rect 57596 5058 57652 5068
rect 58156 5124 58212 5134
rect 58268 5124 58324 5134
rect 58156 5122 58268 5124
rect 58156 5070 58158 5122
rect 58210 5070 58268 5122
rect 58156 5068 58268 5070
rect 58156 5058 58212 5068
rect 57708 4452 57764 4462
rect 58268 4452 58324 5068
rect 57708 4450 58100 4452
rect 57708 4398 57710 4450
rect 57762 4398 58100 4450
rect 57708 4396 58100 4398
rect 57708 4386 57764 4396
rect 57484 3614 57486 3666
rect 57538 3614 57540 3666
rect 57484 3602 57540 3614
rect 57820 3666 57876 3678
rect 57820 3614 57822 3666
rect 57874 3614 57876 3666
rect 57820 3556 57876 3614
rect 57932 3556 57988 3566
rect 57820 3554 57988 3556
rect 57820 3502 57934 3554
rect 57986 3502 57988 3554
rect 57820 3500 57988 3502
rect 55692 3424 55748 3500
rect 57932 3490 57988 3500
rect 56700 3332 56756 3342
rect 56364 3330 56756 3332
rect 56364 3278 56702 3330
rect 56754 3278 56756 3330
rect 56364 3276 56756 3278
rect 56364 800 56420 3276
rect 56700 3266 56756 3276
rect 58044 800 58100 4396
rect 58156 4450 58324 4452
rect 58156 4398 58270 4450
rect 58322 4398 58324 4450
rect 58156 4396 58324 4398
rect 58156 3554 58212 4396
rect 58268 4386 58324 4396
rect 58380 4562 58436 5182
rect 58492 5124 58548 5740
rect 58716 5794 58772 6526
rect 58716 5742 58718 5794
rect 58770 5742 58772 5794
rect 58716 5348 58772 5742
rect 58716 5282 58772 5292
rect 59276 6578 59332 6590
rect 59276 6526 59278 6578
rect 59330 6526 59332 6578
rect 59276 5348 59332 6526
rect 59276 5234 59332 5292
rect 59276 5182 59278 5234
rect 59330 5182 59332 5234
rect 58492 5058 58548 5068
rect 58716 5124 58772 5134
rect 58380 4510 58382 4562
rect 58434 4510 58436 4562
rect 58380 3666 58436 4510
rect 58380 3614 58382 3666
rect 58434 3614 58436 3666
rect 58380 3602 58436 3614
rect 58716 3666 58772 5068
rect 59052 5124 59108 5162
rect 59052 5058 59108 5068
rect 58716 3614 58718 3666
rect 58770 3614 58772 3666
rect 58716 3602 58772 3614
rect 59276 3666 59332 5182
rect 59276 3614 59278 3666
rect 59330 3614 59332 3666
rect 59276 3602 59332 3614
rect 59612 6578 59668 6590
rect 59612 6526 59614 6578
rect 59666 6526 59668 6578
rect 59612 6468 59668 6526
rect 59612 6020 59668 6412
rect 60060 6468 60116 6478
rect 60060 6374 60116 6412
rect 61180 6468 61236 6478
rect 63756 6468 63812 6478
rect 61180 6130 61236 6412
rect 61180 6078 61182 6130
rect 61234 6078 61236 6130
rect 59724 6020 59780 6030
rect 59612 6018 59780 6020
rect 59612 5966 59726 6018
rect 59778 5966 59780 6018
rect 59612 5964 59780 5966
rect 59612 3666 59668 5964
rect 59724 5954 59780 5964
rect 60284 5908 60340 5918
rect 60732 5908 60788 5918
rect 60284 5906 60732 5908
rect 60284 5854 60286 5906
rect 60338 5854 60732 5906
rect 60284 5852 60732 5854
rect 60284 5842 60340 5852
rect 60732 5776 60788 5852
rect 60172 5348 60228 5358
rect 60172 5234 60228 5292
rect 60172 5182 60174 5234
rect 60226 5182 60228 5234
rect 60172 5170 60228 5182
rect 60620 5236 60676 5246
rect 60620 5142 60676 5180
rect 61180 5236 61236 6078
rect 63644 6466 63812 6468
rect 63644 6414 63758 6466
rect 63810 6414 63812 6466
rect 63644 6412 63812 6414
rect 62188 5908 62244 5918
rect 61964 5794 62020 5806
rect 61964 5742 61966 5794
rect 62018 5742 62020 5794
rect 61740 5348 61796 5358
rect 59836 5124 59892 5134
rect 59836 5010 59892 5068
rect 59836 4958 59838 5010
rect 59890 4958 59892 5010
rect 59836 4226 59892 4958
rect 61180 4338 61236 5180
rect 61404 5236 61460 5246
rect 61404 5142 61460 5180
rect 61740 5234 61796 5292
rect 61740 5182 61742 5234
rect 61794 5182 61796 5234
rect 61740 5170 61796 5182
rect 61964 5236 62020 5742
rect 61964 5170 62020 5180
rect 62188 4562 62244 5852
rect 62860 5796 62916 5806
rect 62860 5794 63028 5796
rect 62860 5742 62862 5794
rect 62914 5742 63028 5794
rect 62860 5740 63028 5742
rect 62860 5730 62916 5740
rect 62636 5236 62692 5246
rect 62972 5236 63028 5740
rect 63308 5794 63364 5806
rect 63308 5742 63310 5794
rect 63362 5742 63364 5794
rect 63308 5236 63364 5742
rect 63644 5572 63700 6412
rect 63756 6402 63812 6412
rect 63756 5908 63812 5918
rect 63756 5814 63812 5852
rect 64428 5906 64484 6748
rect 64540 6710 64596 6748
rect 65100 6804 65156 6814
rect 65100 6710 65156 6748
rect 65436 6804 65492 7310
rect 66108 7362 66164 7374
rect 66108 7310 66110 7362
rect 66162 7310 66164 7362
rect 65436 6738 65492 6748
rect 65996 6804 66052 6814
rect 65996 6710 66052 6748
rect 65436 6578 65492 6590
rect 65436 6526 65438 6578
rect 65490 6526 65492 6578
rect 65436 6468 65492 6526
rect 64428 5854 64430 5906
rect 64482 5854 64484 5906
rect 63644 5516 63812 5572
rect 62636 5234 63364 5236
rect 62636 5182 62638 5234
rect 62690 5182 62974 5234
rect 63026 5182 63364 5234
rect 62636 5180 63364 5182
rect 62636 5170 62692 5180
rect 62972 5170 63028 5180
rect 63308 5012 63364 5180
rect 63532 5012 63588 5022
rect 63308 4956 63532 5012
rect 62188 4510 62190 4562
rect 62242 4510 62244 4562
rect 62188 4498 62244 4510
rect 62860 4452 62916 4462
rect 62860 4450 63140 4452
rect 62860 4398 62862 4450
rect 62914 4398 63140 4450
rect 62860 4396 63140 4398
rect 62860 4386 62916 4396
rect 61180 4286 61182 4338
rect 61234 4286 61236 4338
rect 61180 4274 61236 4286
rect 59836 4174 59838 4226
rect 59890 4174 59892 4226
rect 59836 4162 59892 4174
rect 59612 3614 59614 3666
rect 59666 3614 59668 3666
rect 59612 3602 59668 3614
rect 58156 3502 58158 3554
rect 58210 3502 58212 3554
rect 58156 3490 58212 3502
rect 62188 3556 62244 3566
rect 62188 3462 62244 3500
rect 62076 3442 62132 3454
rect 62076 3390 62078 3442
rect 62130 3390 62132 3442
rect 59724 3332 59780 3342
rect 59724 800 59780 3276
rect 60620 3332 60676 3342
rect 60620 3238 60676 3276
rect 61404 3330 61460 3342
rect 61404 3278 61406 3330
rect 61458 3278 61460 3330
rect 61404 800 61460 3278
rect 62076 3332 62132 3390
rect 62860 3444 62916 3454
rect 62860 3350 62916 3388
rect 62076 3266 62132 3276
rect 63084 800 63140 4396
rect 63420 4450 63476 4956
rect 63532 4918 63588 4956
rect 63644 4898 63700 4910
rect 63644 4846 63646 4898
rect 63698 4846 63700 4898
rect 63420 4398 63422 4450
rect 63474 4398 63476 4450
rect 63420 4386 63476 4398
rect 63532 4564 63588 4574
rect 63644 4564 63700 4846
rect 63532 4562 63700 4564
rect 63532 4510 63534 4562
rect 63586 4510 63700 4562
rect 63532 4508 63700 4510
rect 63532 4340 63588 4508
rect 63756 4452 63812 5516
rect 63532 4274 63588 4284
rect 63644 4396 63812 4452
rect 64428 5234 64484 5854
rect 65324 5908 65380 5918
rect 64428 5182 64430 5234
rect 64482 5182 64484 5234
rect 64428 5012 64484 5182
rect 63644 3668 63700 4396
rect 64428 4340 64484 4956
rect 64652 5794 64708 5806
rect 64652 5742 64654 5794
rect 64706 5742 64708 5794
rect 64652 5234 64708 5742
rect 64652 5182 64654 5234
rect 64706 5182 64708 5234
rect 64652 4340 64708 5182
rect 65324 5234 65380 5852
rect 65324 5182 65326 5234
rect 65378 5182 65380 5234
rect 65324 5170 65380 5182
rect 65436 4900 65492 6412
rect 66108 6468 66164 7310
rect 66108 6374 66164 6412
rect 66332 7362 66388 7374
rect 66332 7310 66334 7362
rect 66386 7310 66388 7362
rect 66332 6804 66388 7310
rect 65660 5908 65716 5918
rect 66220 5908 66276 5918
rect 65660 5814 65716 5852
rect 66108 5852 66220 5908
rect 64428 4338 64596 4340
rect 64428 4286 64430 4338
rect 64482 4286 64596 4338
rect 64428 4284 64596 4286
rect 64428 4274 64484 4284
rect 63756 3668 63812 3678
rect 63644 3612 63756 3668
rect 64540 3668 64596 4284
rect 64652 4246 64708 4284
rect 64876 4340 64932 4350
rect 64652 3668 64708 3678
rect 64540 3666 64708 3668
rect 64540 3614 64654 3666
rect 64706 3614 64708 3666
rect 64540 3612 64708 3614
rect 63756 3554 63812 3612
rect 64652 3602 64708 3612
rect 64876 3666 64932 4284
rect 65436 4340 65492 4844
rect 66108 5124 66164 5852
rect 66220 5814 66276 5852
rect 65548 4452 65604 4462
rect 65548 4450 65940 4452
rect 65548 4398 65550 4450
rect 65602 4398 65940 4450
rect 65548 4396 65940 4398
rect 65548 4386 65604 4396
rect 64876 3614 64878 3666
rect 64930 3614 64932 3666
rect 64876 3602 64932 3614
rect 65324 3668 65380 3678
rect 63756 3502 63758 3554
rect 63810 3502 63812 3554
rect 63756 3490 63812 3502
rect 64876 3444 64932 3454
rect 63420 3332 63476 3342
rect 63420 3238 63476 3276
rect 64876 1652 64932 3388
rect 64764 1596 64932 1652
rect 64764 800 64820 1596
rect 65324 800 65380 3612
rect 65436 3556 65492 4284
rect 65772 4226 65828 4238
rect 65772 4174 65774 4226
rect 65826 4174 65828 4226
rect 65660 3556 65716 3566
rect 65772 3556 65828 4174
rect 65436 3500 65604 3556
rect 65548 3332 65604 3500
rect 65660 3554 65828 3556
rect 65660 3502 65662 3554
rect 65714 3502 65828 3554
rect 65660 3500 65828 3502
rect 65660 3490 65716 3500
rect 65660 3332 65716 3342
rect 65548 3330 65716 3332
rect 65548 3278 65662 3330
rect 65714 3278 65716 3330
rect 65548 3276 65716 3278
rect 65660 3266 65716 3276
rect 65884 800 65940 4396
rect 66108 4338 66164 5068
rect 66332 5122 66388 6748
rect 66892 7362 66948 7374
rect 67340 7364 67396 7374
rect 67676 7364 67732 7374
rect 66892 7310 66894 7362
rect 66946 7310 66948 7362
rect 66892 6802 66948 7310
rect 66892 6750 66894 6802
rect 66946 6750 66948 6802
rect 66892 6692 66948 6750
rect 67228 7362 67396 7364
rect 67228 7310 67342 7362
rect 67394 7310 67396 7362
rect 67228 7308 67396 7310
rect 67228 6804 67284 7308
rect 67340 7298 67396 7308
rect 67564 7362 67732 7364
rect 67564 7310 67678 7362
rect 67730 7310 67732 7362
rect 67564 7308 67732 7310
rect 67228 6692 67284 6748
rect 66892 6636 67284 6692
rect 67004 6468 67060 6478
rect 67004 6374 67060 6412
rect 67228 5906 67284 6636
rect 67228 5854 67230 5906
rect 67282 5854 67284 5906
rect 67228 5842 67284 5854
rect 67452 6468 67508 6478
rect 66332 5070 66334 5122
rect 66386 5070 66388 5122
rect 66332 5058 66388 5070
rect 66444 5794 66500 5806
rect 66444 5742 66446 5794
rect 66498 5742 66500 5794
rect 66332 4900 66388 4910
rect 66444 4900 66500 5742
rect 67452 5796 67508 6412
rect 67452 5702 67508 5740
rect 66388 4844 66500 4900
rect 67116 5012 67172 5022
rect 66332 4806 66388 4844
rect 66108 4286 66110 4338
rect 66162 4286 66164 4338
rect 66108 4228 66164 4286
rect 66108 4226 66948 4228
rect 66108 4174 66110 4226
rect 66162 4174 66948 4226
rect 66108 4172 66948 4174
rect 66108 4162 66164 4172
rect 66892 3666 66948 4172
rect 66892 3614 66894 3666
rect 66946 3614 66948 3666
rect 66892 3602 66948 3614
rect 66444 3556 66500 3566
rect 66444 3330 66500 3500
rect 66444 3278 66446 3330
rect 66498 3278 66500 3330
rect 66444 3266 66500 3278
rect 67116 2548 67172 4956
rect 67564 5012 67620 7308
rect 67676 7298 67732 7308
rect 67698 7084 67962 7094
rect 67754 7028 67802 7084
rect 67858 7028 67906 7084
rect 67698 7018 67962 7028
rect 112022 7084 112286 7094
rect 112078 7028 112126 7084
rect 112182 7028 112230 7084
rect 112022 7018 112286 7028
rect 156346 7084 156610 7094
rect 156402 7028 156450 7084
rect 156506 7028 156554 7084
rect 156346 7018 156610 7028
rect 67676 6804 67732 6814
rect 67676 6468 67732 6748
rect 96460 6578 96516 6590
rect 96460 6526 96462 6578
rect 96514 6526 96516 6578
rect 68124 6468 68180 6478
rect 68572 6468 68628 6478
rect 67676 6466 68628 6468
rect 67676 6414 67678 6466
rect 67730 6414 68126 6466
rect 68178 6414 68574 6466
rect 68626 6414 68628 6466
rect 67676 6412 68628 6414
rect 67676 6402 67732 6412
rect 68124 5908 68180 6412
rect 68572 6132 68628 6412
rect 96012 6468 96068 6478
rect 89860 6300 90124 6310
rect 89916 6244 89964 6300
rect 90020 6244 90068 6300
rect 89860 6234 90124 6244
rect 68796 6132 68852 6142
rect 69244 6132 69300 6142
rect 96012 6132 96068 6412
rect 96348 6468 96404 6478
rect 96348 6374 96404 6412
rect 68572 6130 69300 6132
rect 68572 6078 68798 6130
rect 68850 6078 69246 6130
rect 69298 6078 69300 6130
rect 68572 6076 69300 6078
rect 68796 6066 68852 6076
rect 69244 6066 69300 6076
rect 95900 6130 96068 6132
rect 95900 6078 96014 6130
rect 96066 6078 96068 6130
rect 95900 6076 96068 6078
rect 68124 5906 68292 5908
rect 68124 5854 68126 5906
rect 68178 5854 68292 5906
rect 68124 5852 68292 5854
rect 68124 5842 68180 5852
rect 67698 5516 67962 5526
rect 67754 5460 67802 5516
rect 67858 5460 67906 5516
rect 67698 5450 67962 5460
rect 68236 5124 68292 5852
rect 68348 5796 68404 5806
rect 68404 5740 68516 5796
rect 68348 5664 68404 5740
rect 68236 5122 68404 5124
rect 68236 5070 68238 5122
rect 68290 5070 68404 5122
rect 68236 5068 68404 5070
rect 68236 5058 68292 5068
rect 67228 4898 67284 4910
rect 67228 4846 67230 4898
rect 67282 4846 67284 4898
rect 67564 4880 67620 4956
rect 67228 4116 67284 4846
rect 68348 4340 68404 5068
rect 68460 5122 68516 5740
rect 79324 5794 79380 5806
rect 79324 5742 79326 5794
rect 79378 5742 79380 5794
rect 75852 5460 75908 5470
rect 68460 5070 68462 5122
rect 68514 5070 68516 5122
rect 68460 5012 68516 5070
rect 69244 5124 69300 5134
rect 69244 5030 69300 5068
rect 70364 5122 70420 5134
rect 70364 5070 70366 5122
rect 70418 5070 70420 5122
rect 68460 4946 68516 4956
rect 69580 5012 69636 5022
rect 68460 4340 68516 4350
rect 68348 4284 68460 4340
rect 67228 4050 67284 4060
rect 68460 4226 68516 4284
rect 69356 4340 69412 4350
rect 69356 4246 69412 4284
rect 68460 4174 68462 4226
rect 68514 4174 68516 4226
rect 67698 3948 67962 3958
rect 67754 3892 67802 3948
rect 67858 3892 67906 3948
rect 67698 3882 67962 3892
rect 68460 3666 68516 4174
rect 69580 4226 69636 4956
rect 69804 4898 69860 4910
rect 69804 4846 69806 4898
rect 69858 4846 69860 4898
rect 69804 4340 69860 4846
rect 69804 4274 69860 4284
rect 70140 4340 70196 4350
rect 70140 4246 70196 4284
rect 69580 4174 69582 4226
rect 69634 4174 69636 4226
rect 69580 4116 69636 4174
rect 69580 4050 69636 4060
rect 68460 3614 68462 3666
rect 68514 3614 68516 3666
rect 68460 3602 68516 3614
rect 69132 3780 69188 3790
rect 69132 3556 69188 3724
rect 68684 3554 69188 3556
rect 68684 3502 69134 3554
rect 69186 3502 69188 3554
rect 68684 3500 69188 3502
rect 67004 2492 67172 2548
rect 67564 3330 67620 3342
rect 67564 3278 67566 3330
rect 67618 3278 67620 3330
rect 67004 800 67060 2492
rect 67564 800 67620 3278
rect 68684 800 68740 3500
rect 69132 3490 69188 3500
rect 70364 3556 70420 5070
rect 70700 5122 70756 5134
rect 70700 5070 70702 5122
rect 70754 5070 70756 5122
rect 70476 4226 70532 4238
rect 70476 4174 70478 4226
rect 70530 4174 70532 4226
rect 70476 4116 70532 4174
rect 70476 4050 70532 4060
rect 70700 3780 70756 5070
rect 75852 5122 75908 5404
rect 78988 5236 79044 5246
rect 78988 5142 79044 5180
rect 75852 5070 75854 5122
rect 75906 5070 75908 5122
rect 71148 4452 71204 4462
rect 70700 3714 70756 3724
rect 70924 4450 71204 4452
rect 70924 4398 71150 4450
rect 71202 4398 71204 4450
rect 70924 4396 71204 4398
rect 70812 3556 70868 3566
rect 70364 3554 70868 3556
rect 70364 3502 70814 3554
rect 70866 3502 70868 3554
rect 70364 3500 70868 3502
rect 68908 3330 68964 3342
rect 68908 3278 68910 3330
rect 68962 3278 68964 3330
rect 68908 2884 68964 3278
rect 68908 2818 68964 2828
rect 69804 3330 69860 3342
rect 69804 3278 69806 3330
rect 69858 3278 69860 3330
rect 69244 1762 69300 1774
rect 69244 1710 69246 1762
rect 69298 1710 69300 1762
rect 69244 800 69300 1710
rect 69804 1762 69860 3278
rect 69804 1710 69806 1762
rect 69858 1710 69860 1762
rect 69804 1698 69860 1710
rect 70364 800 70420 3500
rect 70812 3490 70868 3500
rect 70588 3330 70644 3342
rect 70588 3278 70590 3330
rect 70642 3278 70644 3330
rect 70588 2996 70644 3278
rect 70588 2930 70644 2940
rect 70924 800 70980 4396
rect 71148 4386 71204 4396
rect 72604 4452 72660 4462
rect 74284 4452 74340 4462
rect 72604 4450 73444 4452
rect 72604 4398 72606 4450
rect 72658 4398 73444 4450
rect 72604 4396 73444 4398
rect 72604 4386 72660 4396
rect 72268 4338 72324 4350
rect 72268 4286 72270 4338
rect 72322 4286 72324 4338
rect 71820 4228 71876 4238
rect 72268 4228 72324 4286
rect 71820 4226 72324 4228
rect 71820 4174 71822 4226
rect 71874 4174 72324 4226
rect 71820 4172 72324 4174
rect 72604 4228 72660 4238
rect 71820 4162 71876 4172
rect 71596 3444 71652 3454
rect 71596 3350 71652 3388
rect 72044 800 72100 4172
rect 72604 3554 72660 4172
rect 73388 3666 73444 4396
rect 74284 4358 74340 4396
rect 74844 4450 74900 4462
rect 74844 4398 74846 4450
rect 74898 4398 74900 4450
rect 73948 4338 74004 4350
rect 73948 4286 73950 4338
rect 74002 4286 74004 4338
rect 73500 4228 73556 4238
rect 73948 4228 74004 4286
rect 73500 4226 74004 4228
rect 73500 4174 73502 4226
rect 73554 4174 74004 4226
rect 73500 4172 74004 4174
rect 73500 4162 73556 4172
rect 73388 3614 73390 3666
rect 73442 3614 73444 3666
rect 73388 3602 73444 3614
rect 72604 3502 72606 3554
rect 72658 3502 72660 3554
rect 72604 3490 72660 3502
rect 72492 3444 72548 3454
rect 72492 1652 72548 3388
rect 72492 1596 72660 1652
rect 72604 800 72660 1596
rect 73724 800 73780 4172
rect 74284 3444 74340 3454
rect 74284 800 74340 3388
rect 74844 3444 74900 4398
rect 75740 4226 75796 4238
rect 75740 4174 75742 4226
rect 75794 4174 75796 4226
rect 75516 3668 75572 3678
rect 75516 3574 75572 3612
rect 74844 3378 74900 3388
rect 75404 3444 75460 3454
rect 75404 800 75460 3388
rect 75740 3444 75796 4174
rect 75852 4228 75908 5070
rect 79100 5122 79156 5134
rect 79100 5070 79102 5122
rect 79154 5070 79156 5122
rect 78988 4564 79044 4574
rect 79100 4564 79156 5070
rect 79324 5124 79380 5742
rect 81228 5460 81284 5470
rect 79884 5236 79940 5246
rect 79884 5142 79940 5180
rect 79324 5058 79380 5068
rect 79660 5124 79716 5134
rect 79660 5030 79716 5068
rect 80220 4900 80276 4910
rect 80220 4806 80276 4844
rect 78988 4562 79156 4564
rect 78988 4510 78990 4562
rect 79042 4510 79156 4562
rect 78988 4508 79156 4510
rect 78988 4498 79044 4508
rect 76188 4452 76244 4462
rect 79660 4452 79716 4462
rect 75852 4162 75908 4172
rect 75964 4450 76244 4452
rect 75964 4398 76190 4450
rect 76242 4398 76244 4450
rect 75964 4396 76244 4398
rect 75740 3378 75796 3388
rect 75964 800 76020 4396
rect 76188 4386 76244 4396
rect 79436 4450 79716 4452
rect 79436 4398 79662 4450
rect 79714 4398 79716 4450
rect 79436 4396 79716 4398
rect 77084 4228 77140 4238
rect 78540 4228 78596 4238
rect 77084 4226 77252 4228
rect 77084 4174 77086 4226
rect 77138 4174 77252 4226
rect 77084 4172 77252 4174
rect 77084 4162 77140 4172
rect 76300 3444 76356 3454
rect 76300 3350 76356 3388
rect 77196 3444 77252 4172
rect 78540 4226 78820 4228
rect 78540 4174 78542 4226
rect 78594 4174 78820 4226
rect 78540 4172 78820 4174
rect 78540 4162 78596 4172
rect 77308 3444 77364 3454
rect 77196 3442 77364 3444
rect 77196 3390 77310 3442
rect 77362 3390 77364 3442
rect 77196 3388 77364 3390
rect 76636 3332 76692 3342
rect 76636 3238 76692 3276
rect 77196 2548 77252 3388
rect 77308 3378 77364 3388
rect 78764 3444 78820 4172
rect 78988 3444 79044 3454
rect 78764 3442 79044 3444
rect 78764 3390 78990 3442
rect 79042 3390 79044 3442
rect 78764 3388 79044 3390
rect 77644 3330 77700 3342
rect 77644 3278 77646 3330
rect 77698 3278 77700 3330
rect 77644 2884 77700 3278
rect 77644 2818 77700 2828
rect 78204 3330 78260 3342
rect 78204 3278 78206 3330
rect 78258 3278 78260 3330
rect 77084 2492 77252 2548
rect 77084 800 77140 2492
rect 77644 1762 77700 1774
rect 77644 1710 77646 1762
rect 77698 1710 77700 1762
rect 77644 800 77700 1710
rect 78204 1762 78260 3278
rect 78204 1710 78206 1762
rect 78258 1710 78260 1762
rect 78204 1698 78260 1710
rect 78764 800 78820 3388
rect 78988 3378 79044 3388
rect 79324 3330 79380 3342
rect 79324 3278 79326 3330
rect 79378 3278 79380 3330
rect 79324 2996 79380 3278
rect 79324 2930 79380 2940
rect 79436 2212 79492 4396
rect 79660 4386 79716 4396
rect 81228 3556 81284 5404
rect 85708 5348 85764 5358
rect 84364 5124 84420 5134
rect 83356 5012 83412 5022
rect 83356 4918 83412 4956
rect 83020 4900 83076 4910
rect 83020 4806 83076 4844
rect 84364 4898 84420 5068
rect 84364 4846 84366 4898
rect 84418 4846 84420 4898
rect 84028 4340 84084 4350
rect 84028 4246 84084 4284
rect 84364 4340 84420 4846
rect 85708 4452 85764 5292
rect 86604 5348 86660 5358
rect 86604 5254 86660 5292
rect 92316 5348 92372 5358
rect 92316 5254 92372 5292
rect 94780 5348 94836 5358
rect 94780 5254 94836 5292
rect 95900 5348 95956 6076
rect 96012 6066 96068 6076
rect 96124 5908 96180 5918
rect 96124 5906 96404 5908
rect 96124 5854 96126 5906
rect 96178 5854 96404 5906
rect 96124 5852 96404 5854
rect 96124 5842 96180 5852
rect 93212 5236 93268 5246
rect 92428 5234 93268 5236
rect 92428 5182 93214 5234
rect 93266 5182 93268 5234
rect 92428 5180 93268 5182
rect 85932 5122 85988 5134
rect 85932 5070 85934 5122
rect 85986 5070 85988 5122
rect 85932 5012 85988 5070
rect 85932 4946 85988 4956
rect 86492 5122 86548 5134
rect 86492 5070 86494 5122
rect 86546 5070 86548 5122
rect 86492 5012 86548 5070
rect 92428 5122 92484 5180
rect 93212 5170 93268 5180
rect 92428 5070 92430 5122
rect 92482 5070 92484 5122
rect 92428 5058 92484 5070
rect 86492 4946 86548 4956
rect 94892 5010 94948 5022
rect 94892 4958 94894 5010
rect 94946 4958 94948 5010
rect 85820 4898 85876 4910
rect 85820 4846 85822 4898
rect 85874 4846 85876 4898
rect 85820 4676 85876 4846
rect 89860 4732 90124 4742
rect 89916 4676 89964 4732
rect 90020 4676 90068 4732
rect 85820 4620 85988 4676
rect 89860 4666 90124 4676
rect 85820 4452 85876 4462
rect 85708 4450 85876 4452
rect 85708 4398 85822 4450
rect 85874 4398 85876 4450
rect 85708 4396 85876 4398
rect 85820 4386 85876 4396
rect 85036 4340 85092 4350
rect 84364 4274 84420 4284
rect 84924 4338 85092 4340
rect 84924 4286 85038 4338
rect 85090 4286 85092 4338
rect 84924 4284 85092 4286
rect 83692 4228 83748 4238
rect 83692 3668 83748 4172
rect 84588 4228 84644 4238
rect 84588 4134 84644 4172
rect 84924 4228 84980 4284
rect 85036 4274 85092 4284
rect 83692 3602 83748 3612
rect 81228 3462 81284 3500
rect 84924 3554 84980 4172
rect 85708 4116 85764 4126
rect 85932 4116 85988 4620
rect 94892 4564 94948 4958
rect 95564 5012 95620 5022
rect 95564 4918 95620 4956
rect 94892 4498 94948 4508
rect 95900 4562 95956 5292
rect 96348 5122 96404 5852
rect 96348 5070 96350 5122
rect 96402 5070 96404 5122
rect 96348 5058 96404 5070
rect 95900 4510 95902 4562
rect 95954 4510 95956 4562
rect 95900 4498 95956 4510
rect 96124 4898 96180 4910
rect 96124 4846 96126 4898
rect 96178 4846 96180 4898
rect 89068 4452 89124 4462
rect 85764 4060 85988 4116
rect 86492 4340 86548 4350
rect 85708 3666 85764 4060
rect 85708 3614 85710 3666
rect 85762 3614 85764 3666
rect 85708 3602 85764 3614
rect 84924 3502 84926 3554
rect 84978 3502 84980 3554
rect 84924 3490 84980 3502
rect 86492 3554 86548 4284
rect 89068 3668 89124 4396
rect 93660 4450 93716 4462
rect 94668 4452 94724 4462
rect 93660 4398 93662 4450
rect 93714 4398 93716 4450
rect 92988 4340 93044 4350
rect 92428 4338 93044 4340
rect 92428 4286 92990 4338
rect 93042 4286 93044 4338
rect 92428 4284 93044 4286
rect 91420 4228 91476 4238
rect 91420 4134 91476 4172
rect 92092 4228 92148 4238
rect 89068 3602 89124 3612
rect 90636 3668 90692 3678
rect 90636 3574 90692 3612
rect 86492 3502 86494 3554
rect 86546 3502 86548 3554
rect 86492 3490 86548 3502
rect 92092 3556 92148 4172
rect 92428 4226 92484 4284
rect 92988 4274 93044 4284
rect 92428 4174 92430 4226
rect 92482 4174 92484 4226
rect 92428 4162 92484 4174
rect 93100 4116 93156 4126
rect 93100 4022 93156 4060
rect 92764 3668 92820 3678
rect 92764 3574 92820 3612
rect 80220 3444 80276 3454
rect 80668 3444 80724 3454
rect 80220 3442 80724 3444
rect 80220 3390 80222 3442
rect 80274 3390 80670 3442
rect 80722 3390 80724 3442
rect 92092 3424 92148 3500
rect 92764 3444 92820 3454
rect 80220 3388 80724 3390
rect 80220 3378 80276 3388
rect 79324 2156 79492 2212
rect 79324 800 79380 2156
rect 80444 800 80500 3388
rect 80668 3378 80724 3388
rect 81788 3330 81844 3342
rect 82908 3332 82964 3342
rect 81788 3278 81790 3330
rect 81842 3278 81844 3330
rect 81004 1762 81060 1774
rect 81004 1710 81006 1762
rect 81058 1710 81060 1762
rect 81004 800 81060 1710
rect 81788 1762 81844 3278
rect 81788 1710 81790 1762
rect 81842 1710 81844 1762
rect 81788 1698 81844 1710
rect 82684 3330 82964 3332
rect 82684 3278 82910 3330
rect 82962 3278 82964 3330
rect 82684 3276 82964 3278
rect 82684 800 82740 3276
rect 82908 3266 82964 3276
rect 84364 3330 84420 3342
rect 84364 3278 84366 3330
rect 84418 3278 84420 3330
rect 84364 800 84420 3278
rect 87052 3330 87108 3342
rect 88060 3332 88116 3342
rect 89628 3332 89684 3342
rect 87052 3278 87054 3330
rect 87106 3278 87108 3330
rect 86044 1762 86100 1774
rect 86044 1710 86046 1762
rect 86098 1710 86100 1762
rect 86044 800 86100 1710
rect 87052 1762 87108 3278
rect 87052 1710 87054 1762
rect 87106 1710 87108 1762
rect 87052 1698 87108 1710
rect 87724 3330 88116 3332
rect 87724 3278 88062 3330
rect 88114 3278 88116 3330
rect 87724 3276 88116 3278
rect 87724 800 87780 3276
rect 88060 3266 88116 3276
rect 89404 3330 89684 3332
rect 89404 3278 89630 3330
rect 89682 3278 89684 3330
rect 89404 3276 89684 3278
rect 89404 800 89460 3276
rect 89628 3266 89684 3276
rect 91084 3330 91140 3342
rect 91084 3278 91086 3330
rect 91138 3278 91140 3330
rect 89860 3164 90124 3174
rect 89916 3108 89964 3164
rect 90020 3108 90068 3164
rect 89860 3098 90124 3108
rect 91084 800 91140 3278
rect 92764 800 92820 3388
rect 93660 3444 93716 4398
rect 93660 3378 93716 3388
rect 94444 4450 94724 4452
rect 94444 4398 94670 4450
rect 94722 4398 94724 4450
rect 94444 4396 94724 4398
rect 94444 800 94500 4396
rect 94668 4386 94724 4396
rect 96012 4452 96068 4462
rect 96124 4452 96180 4846
rect 96012 4450 96180 4452
rect 96012 4398 96014 4450
rect 96066 4398 96180 4450
rect 96012 4396 96180 4398
rect 96012 4386 96068 4396
rect 94892 3668 94948 3678
rect 94892 3574 94948 3612
rect 96460 3332 96516 6526
rect 97132 6578 97188 6590
rect 97132 6526 97134 6578
rect 97186 6526 97188 6578
rect 97020 6468 97076 6478
rect 97020 5684 97076 6412
rect 97020 5618 97076 5628
rect 96572 5124 96628 5134
rect 96572 5122 96852 5124
rect 96572 5070 96574 5122
rect 96626 5070 96852 5122
rect 96572 5068 96852 5070
rect 96572 5058 96628 5068
rect 96796 5010 96852 5068
rect 96796 4958 96798 5010
rect 96850 4958 96852 5010
rect 96796 4946 96852 4958
rect 97132 4900 97188 6526
rect 114828 6580 114884 6590
rect 114828 6578 115892 6580
rect 114828 6526 114830 6578
rect 114882 6526 115892 6578
rect 114828 6524 115892 6526
rect 114828 6514 114884 6524
rect 114716 6466 114772 6478
rect 114716 6414 114718 6466
rect 114770 6414 114772 6466
rect 114716 6356 114772 6414
rect 114492 6300 114772 6356
rect 107660 6018 107716 6030
rect 107660 5966 107662 6018
rect 107714 5966 107716 6018
rect 97356 5906 97412 5918
rect 97356 5854 97358 5906
rect 97410 5854 97412 5906
rect 97244 5684 97300 5694
rect 97244 5590 97300 5628
rect 97356 5012 97412 5854
rect 98028 5906 98084 5918
rect 98028 5854 98030 5906
rect 98082 5854 98084 5906
rect 97916 5684 97972 5694
rect 97916 5124 97972 5628
rect 97916 5058 97972 5068
rect 97468 5012 97524 5022
rect 97356 5010 97524 5012
rect 97356 4958 97470 5010
rect 97522 4958 97524 5010
rect 97356 4956 97524 4958
rect 97468 4946 97524 4956
rect 97132 4834 97188 4844
rect 97244 4564 97300 4574
rect 97244 4470 97300 4508
rect 98028 4562 98084 5854
rect 98252 5124 98308 5134
rect 105980 5124 106036 5134
rect 98252 5030 98308 5068
rect 105756 5122 106036 5124
rect 105756 5070 105982 5122
rect 106034 5070 106036 5122
rect 105756 5068 106036 5070
rect 98140 5012 98196 5022
rect 98140 4918 98196 4956
rect 98812 4900 98868 4910
rect 98812 4806 98868 4844
rect 105420 4898 105476 4910
rect 105420 4846 105422 4898
rect 105474 4846 105476 4898
rect 98028 4510 98030 4562
rect 98082 4510 98084 4562
rect 98028 4498 98084 4510
rect 105196 4340 105252 4350
rect 105196 4226 105252 4284
rect 105420 4340 105476 4846
rect 105420 4274 105476 4284
rect 105756 4340 105812 5068
rect 105980 5058 106036 5068
rect 106540 5124 106596 5134
rect 105756 4246 105812 4284
rect 105196 4174 105198 4226
rect 105250 4174 105252 4226
rect 105196 3668 105252 4174
rect 105196 3602 105252 3612
rect 105980 4228 106036 4238
rect 105980 3556 106036 4172
rect 106540 4228 106596 5068
rect 106540 4134 106596 4172
rect 106764 5124 106820 5134
rect 106764 4116 106820 5068
rect 107660 5122 107716 5966
rect 113260 5906 113316 5918
rect 113260 5854 113262 5906
rect 113314 5854 113316 5906
rect 113148 5682 113204 5694
rect 113148 5630 113150 5682
rect 113202 5630 113204 5682
rect 112022 5516 112286 5526
rect 112078 5460 112126 5516
rect 112182 5460 112230 5516
rect 112022 5450 112286 5460
rect 113148 5348 113204 5630
rect 113148 5282 113204 5292
rect 113260 5236 113316 5854
rect 113932 5906 113988 5918
rect 113932 5854 113934 5906
rect 113986 5854 113988 5906
rect 113820 5684 113876 5694
rect 113708 5682 113876 5684
rect 113708 5630 113822 5682
rect 113874 5630 113876 5682
rect 113708 5628 113876 5630
rect 113708 5348 113764 5628
rect 113820 5618 113876 5628
rect 113708 5254 113764 5292
rect 113260 5170 113316 5180
rect 107660 5070 107662 5122
rect 107714 5070 107716 5122
rect 107660 5058 107716 5070
rect 112252 5124 112308 5134
rect 112252 5030 112308 5068
rect 112364 5010 112420 5022
rect 112364 4958 112366 5010
rect 112418 4958 112420 5010
rect 107436 4900 107492 4910
rect 107436 4338 107492 4844
rect 108108 4900 108164 4910
rect 108108 4806 108164 4844
rect 112364 4564 112420 4958
rect 113036 5012 113092 5022
rect 113596 5012 113652 5022
rect 113036 5010 113652 5012
rect 113036 4958 113038 5010
rect 113090 4958 113598 5010
rect 113650 4958 113652 5010
rect 113036 4956 113652 4958
rect 113036 4946 113092 4956
rect 113596 4946 113652 4956
rect 112364 4498 112420 4508
rect 113148 4564 113204 4574
rect 113148 4470 113204 4508
rect 113932 4562 113988 5854
rect 114492 5348 114548 6300
rect 114604 6132 114660 6142
rect 114604 6130 115668 6132
rect 114604 6078 114606 6130
rect 114658 6078 115668 6130
rect 114604 6076 115668 6078
rect 114604 6066 114660 6076
rect 115276 5906 115332 5918
rect 115276 5854 115278 5906
rect 115330 5854 115332 5906
rect 114268 5012 114324 5022
rect 114268 4918 114324 4956
rect 113932 4510 113934 4562
rect 113986 4510 113988 4562
rect 113932 4498 113988 4510
rect 114492 4900 114548 5292
rect 115164 5682 115220 5694
rect 115164 5630 115166 5682
rect 115218 5630 115220 5682
rect 114940 4900 114996 4910
rect 114492 4562 114548 4844
rect 114492 4510 114494 4562
rect 114546 4510 114548 4562
rect 114492 4498 114548 4510
rect 114604 4898 114996 4900
rect 114604 4846 114942 4898
rect 114994 4846 114996 4898
rect 114604 4844 114996 4846
rect 108108 4452 108164 4462
rect 109788 4452 109844 4462
rect 107436 4286 107438 4338
rect 107490 4286 107492 4338
rect 107436 4274 107492 4286
rect 107884 4450 108164 4452
rect 107884 4398 108110 4450
rect 108162 4398 108164 4450
rect 107884 4396 108164 4398
rect 106764 4050 106820 4060
rect 105980 3462 106036 3500
rect 107772 3556 107828 3566
rect 107772 3462 107828 3500
rect 105532 3442 105588 3454
rect 105532 3390 105534 3442
rect 105586 3390 105588 3442
rect 96572 3332 96628 3342
rect 96460 3330 96628 3332
rect 96460 3278 96574 3330
rect 96626 3278 96628 3330
rect 96460 3276 96628 3278
rect 96572 3266 96628 3276
rect 97244 3330 97300 3342
rect 98028 3332 98084 3342
rect 99820 3332 99876 3342
rect 101388 3332 101444 3342
rect 97244 3278 97246 3330
rect 97298 3278 97300 3330
rect 96124 1762 96180 1774
rect 96124 1710 96126 1762
rect 96178 1710 96180 1762
rect 96124 800 96180 1710
rect 97244 1762 97300 3278
rect 97244 1710 97246 1762
rect 97298 1710 97300 1762
rect 97244 1698 97300 1710
rect 97804 3330 98084 3332
rect 97804 3278 98030 3330
rect 98082 3278 98084 3330
rect 97804 3276 98084 3278
rect 97804 800 97860 3276
rect 98028 3266 98084 3276
rect 99484 3330 99876 3332
rect 99484 3278 99822 3330
rect 99874 3278 99876 3330
rect 99484 3276 99876 3278
rect 99484 800 99540 3276
rect 99820 3266 99876 3276
rect 101164 3330 101444 3332
rect 101164 3278 101390 3330
rect 101442 3278 101444 3330
rect 101164 3276 101444 3278
rect 101164 800 101220 3276
rect 101388 3266 101444 3276
rect 103740 3330 103796 3342
rect 104748 3332 104804 3342
rect 103740 3278 103742 3330
rect 103794 3278 103796 3330
rect 102844 1762 102900 1774
rect 102844 1710 102846 1762
rect 102898 1710 102900 1762
rect 102844 800 102900 1710
rect 103740 1762 103796 3278
rect 103740 1710 103742 1762
rect 103794 1710 103796 1762
rect 103740 1698 103796 1710
rect 104524 3330 104804 3332
rect 104524 3278 104750 3330
rect 104802 3278 104804 3330
rect 104524 3276 104804 3278
rect 104524 800 104580 3276
rect 104748 3266 104804 3276
rect 105532 3332 105588 3390
rect 106428 3332 106484 3342
rect 105532 3266 105588 3276
rect 106204 3330 106484 3332
rect 106204 3278 106430 3330
rect 106482 3278 106484 3330
rect 106204 3276 106484 3278
rect 106204 800 106260 3276
rect 106428 3266 106484 3276
rect 107884 800 107940 4396
rect 108108 4386 108164 4396
rect 109564 4450 109844 4452
rect 109564 4398 109790 4450
rect 109842 4398 109844 4450
rect 109564 4396 109844 4398
rect 108444 3444 108500 3454
rect 108444 3350 108500 3388
rect 109564 800 109620 4396
rect 109788 4386 109844 4396
rect 114604 4450 114660 4844
rect 114940 4834 114996 4844
rect 115164 4900 115220 5630
rect 115164 4834 115220 4844
rect 115276 4562 115332 5854
rect 115612 5122 115668 6076
rect 115612 5070 115614 5122
rect 115666 5070 115668 5122
rect 115612 5058 115668 5070
rect 115724 4900 115780 4910
rect 115724 4806 115780 4844
rect 115276 4510 115278 4562
rect 115330 4510 115332 4562
rect 115276 4498 115332 4510
rect 115836 4562 115892 6524
rect 134184 6300 134448 6310
rect 134240 6244 134288 6300
rect 134344 6244 134392 6300
rect 134184 6234 134448 6244
rect 178508 6300 178772 6310
rect 178564 6244 178612 6300
rect 178668 6244 178716 6300
rect 178508 6234 178772 6244
rect 156346 5516 156610 5526
rect 156402 5460 156450 5516
rect 156506 5460 156554 5516
rect 156346 5450 156610 5460
rect 118860 5124 118916 5134
rect 118748 5122 118916 5124
rect 118748 5070 118862 5122
rect 118914 5070 118916 5122
rect 118748 5068 118916 5070
rect 118300 4900 118356 4910
rect 115836 4510 115838 4562
rect 115890 4510 115892 4562
rect 115836 4498 115892 4510
rect 118188 4898 118356 4900
rect 118188 4846 118302 4898
rect 118354 4846 118356 4898
rect 118188 4844 118356 4846
rect 114604 4398 114606 4450
rect 114658 4398 114660 4450
rect 114604 4386 114660 4398
rect 118188 4340 118244 4844
rect 118300 4834 118356 4844
rect 118188 4226 118244 4284
rect 118748 4340 118804 5068
rect 118860 5058 118916 5068
rect 120540 5122 120596 5134
rect 120540 5070 120542 5122
rect 120594 5070 120596 5122
rect 118748 4246 118804 4284
rect 119644 5010 119700 5022
rect 119644 4958 119646 5010
rect 119698 4958 119700 5010
rect 119644 4900 119700 4958
rect 120540 5012 120596 5070
rect 120540 4946 120596 4956
rect 120988 5012 121044 5022
rect 120988 4918 121044 4956
rect 118188 4174 118190 4226
rect 118242 4174 118244 4226
rect 112022 3948 112286 3958
rect 112078 3892 112126 3948
rect 112182 3892 112230 3948
rect 112022 3882 112286 3892
rect 110572 3668 110628 3678
rect 110572 3574 110628 3612
rect 118188 3668 118244 4174
rect 119532 4228 119588 4238
rect 119532 4134 119588 4172
rect 118188 3602 118244 3612
rect 119532 3780 119588 3790
rect 119644 3780 119700 4844
rect 141372 4898 141428 4910
rect 141372 4846 141374 4898
rect 141426 4846 141428 4898
rect 134184 4732 134448 4742
rect 134240 4676 134288 4732
rect 134344 4676 134392 4732
rect 134184 4666 134448 4676
rect 120428 4452 120484 4462
rect 120428 4338 120484 4396
rect 121100 4452 121156 4462
rect 121100 4358 121156 4396
rect 128044 4452 128100 4462
rect 120428 4286 120430 4338
rect 120482 4286 120484 4338
rect 120428 4274 120484 4286
rect 119588 3724 119700 3780
rect 120540 4228 120596 4238
rect 119532 3554 119588 3724
rect 119532 3502 119534 3554
rect 119586 3502 119588 3554
rect 119532 3490 119588 3502
rect 120540 3668 120596 4172
rect 126924 4226 126980 4238
rect 127484 4228 127540 4238
rect 126924 4174 126926 4226
rect 126978 4174 126980 4226
rect 126924 4116 126980 4174
rect 120540 3554 120596 3612
rect 121100 3780 121156 3790
rect 121100 3666 121156 3724
rect 121100 3614 121102 3666
rect 121154 3614 121156 3666
rect 121100 3602 121156 3614
rect 121548 3668 121604 3678
rect 121548 3574 121604 3612
rect 120540 3502 120542 3554
rect 120594 3502 120596 3554
rect 120540 3490 120596 3502
rect 126924 3556 126980 4060
rect 126924 3490 126980 3500
rect 127372 4226 127540 4228
rect 127372 4174 127486 4226
rect 127538 4174 127540 4226
rect 127372 4172 127540 4174
rect 127372 3556 127428 4172
rect 127484 4162 127540 4172
rect 119756 3444 119812 3454
rect 119756 3350 119812 3388
rect 121324 3444 121380 3454
rect 111580 3332 111636 3342
rect 113148 3332 113204 3342
rect 111244 3330 111636 3332
rect 111244 3278 111582 3330
rect 111634 3278 111636 3330
rect 111244 3276 111636 3278
rect 111244 800 111300 3276
rect 111580 3266 111636 3276
rect 112924 3330 113204 3332
rect 112924 3278 113150 3330
rect 113202 3278 113204 3330
rect 112924 3276 113204 3278
rect 112924 800 112980 3276
rect 113148 3266 113204 3276
rect 115500 3330 115556 3342
rect 116508 3332 116564 3342
rect 118188 3332 118244 3342
rect 115500 3278 115502 3330
rect 115554 3278 115556 3330
rect 114604 1762 114660 1774
rect 114604 1710 114606 1762
rect 114658 1710 114660 1762
rect 114604 800 114660 1710
rect 115500 1762 115556 3278
rect 115500 1710 115502 1762
rect 115554 1710 115556 1762
rect 115500 1698 115556 1710
rect 116284 3330 116564 3332
rect 116284 3278 116510 3330
rect 116562 3278 116564 3330
rect 116284 3276 116564 3278
rect 116284 800 116340 3276
rect 116508 3266 116564 3276
rect 117964 3330 118244 3332
rect 117964 3278 118190 3330
rect 118242 3278 118244 3330
rect 117964 3276 118244 3278
rect 117964 800 118020 3276
rect 118188 3266 118244 3276
rect 120316 3330 120372 3342
rect 120316 3278 120318 3330
rect 120370 3278 120372 3330
rect 119644 1762 119700 1774
rect 119644 1710 119646 1762
rect 119698 1710 119700 1762
rect 119644 800 119700 1710
rect 120316 1762 120372 3278
rect 120316 1710 120318 1762
rect 120370 1710 120372 1762
rect 120316 1698 120372 1710
rect 121324 800 121380 3388
rect 123340 3332 123396 3342
rect 124908 3332 124964 3342
rect 123004 3330 123396 3332
rect 123004 3278 123342 3330
rect 123394 3278 123396 3330
rect 123004 3276 123396 3278
rect 123004 800 123060 3276
rect 123340 3266 123396 3276
rect 124684 3330 124964 3332
rect 124684 3278 124910 3330
rect 124962 3278 124964 3330
rect 124684 3276 124964 3278
rect 124684 800 124740 3276
rect 124908 3266 124964 3276
rect 126364 3330 126420 3342
rect 126364 3278 126366 3330
rect 126418 3278 126420 3330
rect 126364 800 126420 3278
rect 127372 2884 127428 3500
rect 127596 4116 127652 4126
rect 127596 3554 127652 4060
rect 127596 3502 127598 3554
rect 127650 3502 127652 3554
rect 127596 3490 127652 3502
rect 127372 2818 127428 2828
rect 128044 800 128100 4396
rect 129052 4452 129108 4462
rect 129948 4452 130004 4462
rect 129052 4358 129108 4396
rect 129724 4450 130004 4452
rect 129724 4398 129950 4450
rect 130002 4398 130004 4450
rect 129724 4396 130004 4398
rect 128268 3556 128324 3566
rect 128268 3462 128324 3500
rect 129724 800 129780 4396
rect 129948 4386 130004 4396
rect 132748 4450 132804 4462
rect 133420 4452 133476 4462
rect 132748 4398 132750 4450
rect 132802 4398 132804 4450
rect 130732 4338 130788 4350
rect 130732 4286 130734 4338
rect 130786 4286 130788 4338
rect 130396 3668 130452 3678
rect 130396 3574 130452 3612
rect 130732 3668 130788 4286
rect 132300 4340 132356 4350
rect 132748 4340 132804 4398
rect 132300 4338 132804 4340
rect 132300 4286 132302 4338
rect 132354 4286 132804 4338
rect 132300 4284 132804 4286
rect 132860 4450 133476 4452
rect 132860 4398 133422 4450
rect 133474 4398 133476 4450
rect 132860 4396 133476 4398
rect 132300 4274 132356 4284
rect 131404 4226 131460 4238
rect 131404 4174 131406 4226
rect 131458 4174 131460 4226
rect 130732 3602 130788 3612
rect 131180 3668 131236 3678
rect 131180 3554 131236 3612
rect 131404 3668 131460 4174
rect 131404 3602 131460 3612
rect 131964 4228 132020 4238
rect 131964 3780 132020 4172
rect 131964 3666 132020 3724
rect 131964 3614 131966 3666
rect 132018 3614 132020 3666
rect 131964 3602 132020 3614
rect 131180 3502 131182 3554
rect 131234 3502 131236 3554
rect 131180 3490 131236 3502
rect 132860 3554 132916 4396
rect 133420 4386 133476 4396
rect 141260 4450 141316 4462
rect 141260 4398 141262 4450
rect 141314 4398 141316 4450
rect 132860 3502 132862 3554
rect 132914 3502 132916 3554
rect 132860 3490 132916 3502
rect 139356 4338 139412 4350
rect 139356 4286 139358 4338
rect 139410 4286 139412 4338
rect 139356 3444 139412 4286
rect 140812 4340 140868 4350
rect 141260 4340 141316 4398
rect 140812 4338 141316 4340
rect 140812 4286 140814 4338
rect 140866 4286 141316 4338
rect 140812 4284 141316 4286
rect 140812 4274 140868 4284
rect 139916 4228 139972 4238
rect 139916 4134 139972 4172
rect 140364 3668 140420 3678
rect 140364 3574 140420 3612
rect 139356 3378 139412 3388
rect 139692 3554 139748 3566
rect 139692 3502 139694 3554
rect 139746 3502 139748 3554
rect 139692 3444 139748 3502
rect 141260 3556 141316 3566
rect 141372 3556 141428 4846
rect 178508 4732 178772 4742
rect 178564 4676 178612 4732
rect 178668 4676 178716 4732
rect 178508 4666 178772 4676
rect 141932 4452 141988 4462
rect 151788 4452 151844 4462
rect 153468 4452 153524 4462
rect 141260 3554 141428 3556
rect 141260 3502 141262 3554
rect 141314 3502 141428 3554
rect 141260 3500 141428 3502
rect 141820 4450 141988 4452
rect 141820 4398 141934 4450
rect 141986 4398 141988 4450
rect 141820 4396 141988 4398
rect 141260 3490 141316 3500
rect 139692 3378 139748 3388
rect 131404 3332 131460 3342
rect 131404 800 131460 3276
rect 133308 3332 133364 3342
rect 133308 3238 133364 3276
rect 133980 3330 134036 3342
rect 135100 3332 135156 3342
rect 136668 3332 136724 3342
rect 133980 3278 133982 3330
rect 134034 3278 134036 3330
rect 133084 1762 133140 1774
rect 133084 1710 133086 1762
rect 133138 1710 133140 1762
rect 133084 800 133140 1710
rect 133980 1762 134036 3278
rect 134764 3330 135156 3332
rect 134764 3278 135102 3330
rect 135154 3278 135156 3330
rect 134764 3276 135156 3278
rect 134184 3164 134448 3174
rect 134240 3108 134288 3164
rect 134344 3108 134392 3164
rect 134184 3098 134448 3108
rect 133980 1710 133982 1762
rect 134034 1710 134036 1762
rect 133980 1698 134036 1710
rect 134764 800 134820 3276
rect 135100 3266 135156 3276
rect 136444 3330 136724 3332
rect 136444 3278 136670 3330
rect 136722 3278 136724 3330
rect 136444 3276 136724 3278
rect 136444 800 136500 3276
rect 136668 3266 136724 3276
rect 138124 3330 138180 3342
rect 138124 3278 138126 3330
rect 138178 3278 138180 3330
rect 138124 800 138180 3278
rect 139804 3332 139860 3342
rect 139804 800 139860 3276
rect 141708 3332 141764 3342
rect 141708 3238 141764 3276
rect 141820 980 141876 4396
rect 141932 4386 141988 4396
rect 151564 4450 151844 4452
rect 151564 4398 151790 4450
rect 151842 4398 151844 4450
rect 151564 4396 151844 4398
rect 142604 4226 142660 4238
rect 142604 4174 142606 4226
rect 142658 4174 142660 4226
rect 142604 3444 142660 4174
rect 150444 4226 150500 4238
rect 150444 4174 150446 4226
rect 150498 4174 150500 4226
rect 150444 4116 150500 4174
rect 150444 4050 150500 4060
rect 151004 4226 151060 4238
rect 151004 4174 151006 4226
rect 151058 4174 151060 4226
rect 151004 3556 151060 4174
rect 142604 3378 142660 3388
rect 142940 3444 142996 3454
rect 142940 3350 142996 3388
rect 143388 3332 143444 3342
rect 145068 3332 145124 3342
rect 146860 3332 146916 3342
rect 148428 3332 148484 3342
rect 141484 924 141876 980
rect 143164 3330 143444 3332
rect 143164 3278 143390 3330
rect 143442 3278 143444 3330
rect 143164 3276 143444 3278
rect 141484 800 141540 924
rect 143164 800 143220 3276
rect 143388 3266 143444 3276
rect 144844 3330 145124 3332
rect 144844 3278 145070 3330
rect 145122 3278 145124 3330
rect 144844 3276 145124 3278
rect 144844 800 144900 3276
rect 145068 3266 145124 3276
rect 146524 3330 146916 3332
rect 146524 3278 146862 3330
rect 146914 3278 146916 3330
rect 146524 3276 146916 3278
rect 146524 800 146580 3276
rect 146860 3266 146916 3276
rect 148204 3330 148484 3332
rect 148204 3278 148430 3330
rect 148482 3278 148484 3330
rect 148204 3276 148484 3278
rect 148204 800 148260 3276
rect 148428 3266 148484 3276
rect 149884 3330 149940 3342
rect 149884 3278 149886 3330
rect 149938 3278 149940 3330
rect 149884 800 149940 3278
rect 151004 2996 151060 3500
rect 151116 4116 151172 4126
rect 151116 3554 151172 4060
rect 151116 3502 151118 3554
rect 151170 3502 151172 3554
rect 151116 3490 151172 3502
rect 151004 2930 151060 2940
rect 151564 800 151620 4396
rect 151788 4386 151844 4396
rect 153244 4450 153524 4452
rect 153244 4398 153470 4450
rect 153522 4398 153524 4450
rect 153244 4396 153524 4398
rect 151788 3556 151844 3566
rect 151788 3462 151844 3500
rect 153244 800 153300 4396
rect 153468 4386 153524 4396
rect 156346 3948 156610 3958
rect 156402 3892 156450 3948
rect 156506 3892 156554 3948
rect 156346 3882 156610 3892
rect 153916 3666 153972 3678
rect 153916 3614 153918 3666
rect 153970 3614 153972 3666
rect 153916 3444 153972 3614
rect 153916 3378 153972 3388
rect 155148 3332 155204 3342
rect 156828 3332 156884 3342
rect 158620 3332 158676 3342
rect 160188 3332 160244 3342
rect 154924 3330 155204 3332
rect 154924 3278 155150 3330
rect 155202 3278 155204 3330
rect 154924 3276 155204 3278
rect 154924 800 154980 3276
rect 155148 3266 155204 3276
rect 156604 3330 156884 3332
rect 156604 3278 156830 3330
rect 156882 3278 156884 3330
rect 156604 3276 156884 3278
rect 156604 800 156660 3276
rect 156828 3266 156884 3276
rect 158284 3330 158676 3332
rect 158284 3278 158622 3330
rect 158674 3278 158676 3330
rect 158284 3276 158676 3278
rect 158284 800 158340 3276
rect 158620 3266 158676 3276
rect 159964 3330 160244 3332
rect 159964 3278 160190 3330
rect 160242 3278 160244 3330
rect 159964 3276 160244 3278
rect 159964 800 160020 3276
rect 160188 3266 160244 3276
rect 162540 3330 162596 3342
rect 163548 3332 163604 3342
rect 165228 3332 165284 3342
rect 166908 3332 166964 3342
rect 168588 3332 168644 3342
rect 170380 3332 170436 3342
rect 171948 3332 172004 3342
rect 173068 3332 173124 3342
rect 162540 3278 162542 3330
rect 162594 3278 162596 3330
rect 161644 1762 161700 1774
rect 161644 1710 161646 1762
rect 161698 1710 161700 1762
rect 161644 800 161700 1710
rect 162540 1762 162596 3278
rect 162540 1710 162542 1762
rect 162594 1710 162596 1762
rect 162540 1698 162596 1710
rect 163324 3330 163604 3332
rect 163324 3278 163550 3330
rect 163602 3278 163604 3330
rect 163324 3276 163604 3278
rect 163324 800 163380 3276
rect 163548 3266 163604 3276
rect 165004 3330 165284 3332
rect 165004 3278 165230 3330
rect 165282 3278 165284 3330
rect 165004 3276 165284 3278
rect 165004 800 165060 3276
rect 165228 3266 165284 3276
rect 166684 3330 166964 3332
rect 166684 3278 166910 3330
rect 166962 3278 166964 3330
rect 166684 3276 166964 3278
rect 166684 800 166740 3276
rect 166908 3266 166964 3276
rect 168364 3330 168644 3332
rect 168364 3278 168590 3330
rect 168642 3278 168644 3330
rect 168364 3276 168644 3278
rect 168364 800 168420 3276
rect 168588 3266 168644 3276
rect 170044 3330 170436 3332
rect 170044 3278 170382 3330
rect 170434 3278 170436 3330
rect 170044 3276 170436 3278
rect 170044 800 170100 3276
rect 170380 3266 170436 3276
rect 171724 3330 172004 3332
rect 171724 3278 171950 3330
rect 172002 3278 172004 3330
rect 171724 3276 172004 3278
rect 171724 800 171780 3276
rect 171948 3266 172004 3276
rect 172844 3330 173124 3332
rect 172844 3278 173070 3330
rect 173122 3278 173124 3330
rect 172844 3276 173124 3278
rect 172844 800 172900 3276
rect 173068 3266 173124 3276
rect 173964 3332 174020 3342
rect 173404 1762 173460 1774
rect 173404 1710 173406 1762
rect 173458 1710 173460 1762
rect 173404 800 173460 1710
rect 173964 800 174020 3276
rect 174300 3330 174356 3342
rect 174300 3278 174302 3330
rect 174354 3278 174356 3330
rect 174300 1762 174356 3278
rect 174972 3332 175028 3342
rect 174972 3238 175028 3276
rect 178508 3164 178772 3174
rect 178564 3108 178612 3164
rect 178668 3108 178716 3164
rect 178508 3098 178772 3108
rect 174300 1710 174302 1762
rect 174354 1710 174356 1762
rect 174300 1698 174356 1710
rect 5936 0 6048 800
rect 6496 0 6608 800
rect 7056 0 7168 800
rect 7616 0 7728 800
rect 8176 0 8288 800
rect 8736 0 8848 800
rect 9296 0 9408 800
rect 9856 0 9968 800
rect 10416 0 10528 800
rect 10976 0 11088 800
rect 11536 0 11648 800
rect 12096 0 12208 800
rect 12656 0 12768 800
rect 13216 0 13328 800
rect 13776 0 13888 800
rect 14336 0 14448 800
rect 14896 0 15008 800
rect 15456 0 15568 800
rect 16016 0 16128 800
rect 16576 0 16688 800
rect 17136 0 17248 800
rect 17696 0 17808 800
rect 18256 0 18368 800
rect 18816 0 18928 800
rect 19376 0 19488 800
rect 19936 0 20048 800
rect 20496 0 20608 800
rect 21056 0 21168 800
rect 21616 0 21728 800
rect 22176 0 22288 800
rect 22736 0 22848 800
rect 23296 0 23408 800
rect 23856 0 23968 800
rect 24416 0 24528 800
rect 24976 0 25088 800
rect 25536 0 25648 800
rect 26096 0 26208 800
rect 26656 0 26768 800
rect 27216 0 27328 800
rect 27776 0 27888 800
rect 28336 0 28448 800
rect 28896 0 29008 800
rect 29456 0 29568 800
rect 30016 0 30128 800
rect 30576 0 30688 800
rect 31136 0 31248 800
rect 31696 0 31808 800
rect 32256 0 32368 800
rect 32816 0 32928 800
rect 33376 0 33488 800
rect 33936 0 34048 800
rect 34496 0 34608 800
rect 35056 0 35168 800
rect 35616 0 35728 800
rect 36176 0 36288 800
rect 36736 0 36848 800
rect 37296 0 37408 800
rect 37856 0 37968 800
rect 38416 0 38528 800
rect 38976 0 39088 800
rect 39536 0 39648 800
rect 40096 0 40208 800
rect 40656 0 40768 800
rect 41216 0 41328 800
rect 41776 0 41888 800
rect 42336 0 42448 800
rect 42896 0 43008 800
rect 43456 0 43568 800
rect 44016 0 44128 800
rect 44576 0 44688 800
rect 45136 0 45248 800
rect 45696 0 45808 800
rect 46256 0 46368 800
rect 46816 0 46928 800
rect 47376 0 47488 800
rect 47936 0 48048 800
rect 48496 0 48608 800
rect 49056 0 49168 800
rect 49616 0 49728 800
rect 50176 0 50288 800
rect 50736 0 50848 800
rect 51296 0 51408 800
rect 51856 0 51968 800
rect 52416 0 52528 800
rect 52976 0 53088 800
rect 53536 0 53648 800
rect 54096 0 54208 800
rect 54656 0 54768 800
rect 55216 0 55328 800
rect 55776 0 55888 800
rect 56336 0 56448 800
rect 56896 0 57008 800
rect 57456 0 57568 800
rect 58016 0 58128 800
rect 58576 0 58688 800
rect 59136 0 59248 800
rect 59696 0 59808 800
rect 60256 0 60368 800
rect 60816 0 60928 800
rect 61376 0 61488 800
rect 61936 0 62048 800
rect 62496 0 62608 800
rect 63056 0 63168 800
rect 63616 0 63728 800
rect 64176 0 64288 800
rect 64736 0 64848 800
rect 65296 0 65408 800
rect 65856 0 65968 800
rect 66416 0 66528 800
rect 66976 0 67088 800
rect 67536 0 67648 800
rect 68096 0 68208 800
rect 68656 0 68768 800
rect 69216 0 69328 800
rect 69776 0 69888 800
rect 70336 0 70448 800
rect 70896 0 71008 800
rect 71456 0 71568 800
rect 72016 0 72128 800
rect 72576 0 72688 800
rect 73136 0 73248 800
rect 73696 0 73808 800
rect 74256 0 74368 800
rect 74816 0 74928 800
rect 75376 0 75488 800
rect 75936 0 76048 800
rect 76496 0 76608 800
rect 77056 0 77168 800
rect 77616 0 77728 800
rect 78176 0 78288 800
rect 78736 0 78848 800
rect 79296 0 79408 800
rect 79856 0 79968 800
rect 80416 0 80528 800
rect 80976 0 81088 800
rect 81536 0 81648 800
rect 82096 0 82208 800
rect 82656 0 82768 800
rect 83216 0 83328 800
rect 83776 0 83888 800
rect 84336 0 84448 800
rect 84896 0 85008 800
rect 85456 0 85568 800
rect 86016 0 86128 800
rect 86576 0 86688 800
rect 87136 0 87248 800
rect 87696 0 87808 800
rect 88256 0 88368 800
rect 88816 0 88928 800
rect 89376 0 89488 800
rect 89936 0 90048 800
rect 90496 0 90608 800
rect 91056 0 91168 800
rect 91616 0 91728 800
rect 92176 0 92288 800
rect 92736 0 92848 800
rect 93296 0 93408 800
rect 93856 0 93968 800
rect 94416 0 94528 800
rect 94976 0 95088 800
rect 95536 0 95648 800
rect 96096 0 96208 800
rect 96656 0 96768 800
rect 97216 0 97328 800
rect 97776 0 97888 800
rect 98336 0 98448 800
rect 98896 0 99008 800
rect 99456 0 99568 800
rect 100016 0 100128 800
rect 100576 0 100688 800
rect 101136 0 101248 800
rect 101696 0 101808 800
rect 102256 0 102368 800
rect 102816 0 102928 800
rect 103376 0 103488 800
rect 103936 0 104048 800
rect 104496 0 104608 800
rect 105056 0 105168 800
rect 105616 0 105728 800
rect 106176 0 106288 800
rect 106736 0 106848 800
rect 107296 0 107408 800
rect 107856 0 107968 800
rect 108416 0 108528 800
rect 108976 0 109088 800
rect 109536 0 109648 800
rect 110096 0 110208 800
rect 110656 0 110768 800
rect 111216 0 111328 800
rect 111776 0 111888 800
rect 112336 0 112448 800
rect 112896 0 113008 800
rect 113456 0 113568 800
rect 114016 0 114128 800
rect 114576 0 114688 800
rect 115136 0 115248 800
rect 115696 0 115808 800
rect 116256 0 116368 800
rect 116816 0 116928 800
rect 117376 0 117488 800
rect 117936 0 118048 800
rect 118496 0 118608 800
rect 119056 0 119168 800
rect 119616 0 119728 800
rect 120176 0 120288 800
rect 120736 0 120848 800
rect 121296 0 121408 800
rect 121856 0 121968 800
rect 122416 0 122528 800
rect 122976 0 123088 800
rect 123536 0 123648 800
rect 124096 0 124208 800
rect 124656 0 124768 800
rect 125216 0 125328 800
rect 125776 0 125888 800
rect 126336 0 126448 800
rect 126896 0 127008 800
rect 127456 0 127568 800
rect 128016 0 128128 800
rect 128576 0 128688 800
rect 129136 0 129248 800
rect 129696 0 129808 800
rect 130256 0 130368 800
rect 130816 0 130928 800
rect 131376 0 131488 800
rect 131936 0 132048 800
rect 132496 0 132608 800
rect 133056 0 133168 800
rect 133616 0 133728 800
rect 134176 0 134288 800
rect 134736 0 134848 800
rect 135296 0 135408 800
rect 135856 0 135968 800
rect 136416 0 136528 800
rect 136976 0 137088 800
rect 137536 0 137648 800
rect 138096 0 138208 800
rect 138656 0 138768 800
rect 139216 0 139328 800
rect 139776 0 139888 800
rect 140336 0 140448 800
rect 140896 0 141008 800
rect 141456 0 141568 800
rect 142016 0 142128 800
rect 142576 0 142688 800
rect 143136 0 143248 800
rect 143696 0 143808 800
rect 144256 0 144368 800
rect 144816 0 144928 800
rect 145376 0 145488 800
rect 145936 0 146048 800
rect 146496 0 146608 800
rect 147056 0 147168 800
rect 147616 0 147728 800
rect 148176 0 148288 800
rect 148736 0 148848 800
rect 149296 0 149408 800
rect 149856 0 149968 800
rect 150416 0 150528 800
rect 150976 0 151088 800
rect 151536 0 151648 800
rect 152096 0 152208 800
rect 152656 0 152768 800
rect 153216 0 153328 800
rect 153776 0 153888 800
rect 154336 0 154448 800
rect 154896 0 155008 800
rect 155456 0 155568 800
rect 156016 0 156128 800
rect 156576 0 156688 800
rect 157136 0 157248 800
rect 157696 0 157808 800
rect 158256 0 158368 800
rect 158816 0 158928 800
rect 159376 0 159488 800
rect 159936 0 160048 800
rect 160496 0 160608 800
rect 161056 0 161168 800
rect 161616 0 161728 800
rect 162176 0 162288 800
rect 162736 0 162848 800
rect 163296 0 163408 800
rect 163856 0 163968 800
rect 164416 0 164528 800
rect 164976 0 165088 800
rect 165536 0 165648 800
rect 166096 0 166208 800
rect 166656 0 166768 800
rect 167216 0 167328 800
rect 167776 0 167888 800
rect 168336 0 168448 800
rect 168896 0 169008 800
rect 169456 0 169568 800
rect 170016 0 170128 800
rect 170576 0 170688 800
rect 171136 0 171248 800
rect 171696 0 171808 800
rect 172256 0 172368 800
rect 172816 0 172928 800
rect 173376 0 173488 800
rect 173936 0 174048 800
<< via2 >>
rect 23374 16490 23430 16492
rect 23374 16438 23376 16490
rect 23376 16438 23428 16490
rect 23428 16438 23430 16490
rect 23374 16436 23430 16438
rect 23478 16490 23534 16492
rect 23478 16438 23480 16490
rect 23480 16438 23532 16490
rect 23532 16438 23534 16490
rect 23478 16436 23534 16438
rect 23582 16490 23638 16492
rect 23582 16438 23584 16490
rect 23584 16438 23636 16490
rect 23636 16438 23638 16490
rect 23582 16436 23638 16438
rect 67698 16490 67754 16492
rect 67698 16438 67700 16490
rect 67700 16438 67752 16490
rect 67752 16438 67754 16490
rect 67698 16436 67754 16438
rect 67802 16490 67858 16492
rect 67802 16438 67804 16490
rect 67804 16438 67856 16490
rect 67856 16438 67858 16490
rect 67802 16436 67858 16438
rect 67906 16490 67962 16492
rect 67906 16438 67908 16490
rect 67908 16438 67960 16490
rect 67960 16438 67962 16490
rect 67906 16436 67962 16438
rect 112022 16490 112078 16492
rect 112022 16438 112024 16490
rect 112024 16438 112076 16490
rect 112076 16438 112078 16490
rect 112022 16436 112078 16438
rect 112126 16490 112182 16492
rect 112126 16438 112128 16490
rect 112128 16438 112180 16490
rect 112180 16438 112182 16490
rect 112126 16436 112182 16438
rect 112230 16490 112286 16492
rect 112230 16438 112232 16490
rect 112232 16438 112284 16490
rect 112284 16438 112286 16490
rect 112230 16436 112286 16438
rect 156346 16490 156402 16492
rect 156346 16438 156348 16490
rect 156348 16438 156400 16490
rect 156400 16438 156402 16490
rect 156346 16436 156402 16438
rect 156450 16490 156506 16492
rect 156450 16438 156452 16490
rect 156452 16438 156504 16490
rect 156504 16438 156506 16490
rect 156450 16436 156506 16438
rect 156554 16490 156610 16492
rect 156554 16438 156556 16490
rect 156556 16438 156608 16490
rect 156608 16438 156610 16490
rect 156554 16436 156610 16438
rect 45536 15706 45592 15708
rect 45536 15654 45538 15706
rect 45538 15654 45590 15706
rect 45590 15654 45592 15706
rect 45536 15652 45592 15654
rect 45640 15706 45696 15708
rect 45640 15654 45642 15706
rect 45642 15654 45694 15706
rect 45694 15654 45696 15706
rect 45640 15652 45696 15654
rect 45744 15706 45800 15708
rect 45744 15654 45746 15706
rect 45746 15654 45798 15706
rect 45798 15654 45800 15706
rect 45744 15652 45800 15654
rect 89860 15706 89916 15708
rect 89860 15654 89862 15706
rect 89862 15654 89914 15706
rect 89914 15654 89916 15706
rect 89860 15652 89916 15654
rect 89964 15706 90020 15708
rect 89964 15654 89966 15706
rect 89966 15654 90018 15706
rect 90018 15654 90020 15706
rect 89964 15652 90020 15654
rect 90068 15706 90124 15708
rect 90068 15654 90070 15706
rect 90070 15654 90122 15706
rect 90122 15654 90124 15706
rect 90068 15652 90124 15654
rect 134184 15706 134240 15708
rect 134184 15654 134186 15706
rect 134186 15654 134238 15706
rect 134238 15654 134240 15706
rect 134184 15652 134240 15654
rect 134288 15706 134344 15708
rect 134288 15654 134290 15706
rect 134290 15654 134342 15706
rect 134342 15654 134344 15706
rect 134288 15652 134344 15654
rect 134392 15706 134448 15708
rect 134392 15654 134394 15706
rect 134394 15654 134446 15706
rect 134446 15654 134448 15706
rect 134392 15652 134448 15654
rect 178508 15706 178564 15708
rect 178508 15654 178510 15706
rect 178510 15654 178562 15706
rect 178562 15654 178564 15706
rect 178508 15652 178564 15654
rect 178612 15706 178668 15708
rect 178612 15654 178614 15706
rect 178614 15654 178666 15706
rect 178666 15654 178668 15706
rect 178612 15652 178668 15654
rect 178716 15706 178772 15708
rect 178716 15654 178718 15706
rect 178718 15654 178770 15706
rect 178770 15654 178772 15706
rect 178716 15652 178772 15654
rect 23374 14922 23430 14924
rect 23374 14870 23376 14922
rect 23376 14870 23428 14922
rect 23428 14870 23430 14922
rect 23374 14868 23430 14870
rect 23478 14922 23534 14924
rect 23478 14870 23480 14922
rect 23480 14870 23532 14922
rect 23532 14870 23534 14922
rect 23478 14868 23534 14870
rect 23582 14922 23638 14924
rect 23582 14870 23584 14922
rect 23584 14870 23636 14922
rect 23636 14870 23638 14922
rect 23582 14868 23638 14870
rect 67698 14922 67754 14924
rect 67698 14870 67700 14922
rect 67700 14870 67752 14922
rect 67752 14870 67754 14922
rect 67698 14868 67754 14870
rect 67802 14922 67858 14924
rect 67802 14870 67804 14922
rect 67804 14870 67856 14922
rect 67856 14870 67858 14922
rect 67802 14868 67858 14870
rect 67906 14922 67962 14924
rect 67906 14870 67908 14922
rect 67908 14870 67960 14922
rect 67960 14870 67962 14922
rect 67906 14868 67962 14870
rect 112022 14922 112078 14924
rect 112022 14870 112024 14922
rect 112024 14870 112076 14922
rect 112076 14870 112078 14922
rect 112022 14868 112078 14870
rect 112126 14922 112182 14924
rect 112126 14870 112128 14922
rect 112128 14870 112180 14922
rect 112180 14870 112182 14922
rect 112126 14868 112182 14870
rect 112230 14922 112286 14924
rect 112230 14870 112232 14922
rect 112232 14870 112284 14922
rect 112284 14870 112286 14922
rect 112230 14868 112286 14870
rect 156346 14922 156402 14924
rect 156346 14870 156348 14922
rect 156348 14870 156400 14922
rect 156400 14870 156402 14922
rect 156346 14868 156402 14870
rect 156450 14922 156506 14924
rect 156450 14870 156452 14922
rect 156452 14870 156504 14922
rect 156504 14870 156506 14922
rect 156450 14868 156506 14870
rect 156554 14922 156610 14924
rect 156554 14870 156556 14922
rect 156556 14870 156608 14922
rect 156608 14870 156610 14922
rect 156554 14868 156610 14870
rect 45536 14138 45592 14140
rect 45536 14086 45538 14138
rect 45538 14086 45590 14138
rect 45590 14086 45592 14138
rect 45536 14084 45592 14086
rect 45640 14138 45696 14140
rect 45640 14086 45642 14138
rect 45642 14086 45694 14138
rect 45694 14086 45696 14138
rect 45640 14084 45696 14086
rect 45744 14138 45800 14140
rect 45744 14086 45746 14138
rect 45746 14086 45798 14138
rect 45798 14086 45800 14138
rect 45744 14084 45800 14086
rect 89860 14138 89916 14140
rect 89860 14086 89862 14138
rect 89862 14086 89914 14138
rect 89914 14086 89916 14138
rect 89860 14084 89916 14086
rect 89964 14138 90020 14140
rect 89964 14086 89966 14138
rect 89966 14086 90018 14138
rect 90018 14086 90020 14138
rect 89964 14084 90020 14086
rect 90068 14138 90124 14140
rect 90068 14086 90070 14138
rect 90070 14086 90122 14138
rect 90122 14086 90124 14138
rect 90068 14084 90124 14086
rect 134184 14138 134240 14140
rect 134184 14086 134186 14138
rect 134186 14086 134238 14138
rect 134238 14086 134240 14138
rect 134184 14084 134240 14086
rect 134288 14138 134344 14140
rect 134288 14086 134290 14138
rect 134290 14086 134342 14138
rect 134342 14086 134344 14138
rect 134288 14084 134344 14086
rect 134392 14138 134448 14140
rect 134392 14086 134394 14138
rect 134394 14086 134446 14138
rect 134446 14086 134448 14138
rect 134392 14084 134448 14086
rect 178508 14138 178564 14140
rect 178508 14086 178510 14138
rect 178510 14086 178562 14138
rect 178562 14086 178564 14138
rect 178508 14084 178564 14086
rect 178612 14138 178668 14140
rect 178612 14086 178614 14138
rect 178614 14086 178666 14138
rect 178666 14086 178668 14138
rect 178612 14084 178668 14086
rect 178716 14138 178772 14140
rect 178716 14086 178718 14138
rect 178718 14086 178770 14138
rect 178770 14086 178772 14138
rect 178716 14084 178772 14086
rect 23374 13354 23430 13356
rect 23374 13302 23376 13354
rect 23376 13302 23428 13354
rect 23428 13302 23430 13354
rect 23374 13300 23430 13302
rect 23478 13354 23534 13356
rect 23478 13302 23480 13354
rect 23480 13302 23532 13354
rect 23532 13302 23534 13354
rect 23478 13300 23534 13302
rect 23582 13354 23638 13356
rect 23582 13302 23584 13354
rect 23584 13302 23636 13354
rect 23636 13302 23638 13354
rect 23582 13300 23638 13302
rect 67698 13354 67754 13356
rect 67698 13302 67700 13354
rect 67700 13302 67752 13354
rect 67752 13302 67754 13354
rect 67698 13300 67754 13302
rect 67802 13354 67858 13356
rect 67802 13302 67804 13354
rect 67804 13302 67856 13354
rect 67856 13302 67858 13354
rect 67802 13300 67858 13302
rect 67906 13354 67962 13356
rect 67906 13302 67908 13354
rect 67908 13302 67960 13354
rect 67960 13302 67962 13354
rect 67906 13300 67962 13302
rect 112022 13354 112078 13356
rect 112022 13302 112024 13354
rect 112024 13302 112076 13354
rect 112076 13302 112078 13354
rect 112022 13300 112078 13302
rect 112126 13354 112182 13356
rect 112126 13302 112128 13354
rect 112128 13302 112180 13354
rect 112180 13302 112182 13354
rect 112126 13300 112182 13302
rect 112230 13354 112286 13356
rect 112230 13302 112232 13354
rect 112232 13302 112284 13354
rect 112284 13302 112286 13354
rect 112230 13300 112286 13302
rect 156346 13354 156402 13356
rect 156346 13302 156348 13354
rect 156348 13302 156400 13354
rect 156400 13302 156402 13354
rect 156346 13300 156402 13302
rect 156450 13354 156506 13356
rect 156450 13302 156452 13354
rect 156452 13302 156504 13354
rect 156504 13302 156506 13354
rect 156450 13300 156506 13302
rect 156554 13354 156610 13356
rect 156554 13302 156556 13354
rect 156556 13302 156608 13354
rect 156608 13302 156610 13354
rect 156554 13300 156610 13302
rect 45536 12570 45592 12572
rect 45536 12518 45538 12570
rect 45538 12518 45590 12570
rect 45590 12518 45592 12570
rect 45536 12516 45592 12518
rect 45640 12570 45696 12572
rect 45640 12518 45642 12570
rect 45642 12518 45694 12570
rect 45694 12518 45696 12570
rect 45640 12516 45696 12518
rect 45744 12570 45800 12572
rect 45744 12518 45746 12570
rect 45746 12518 45798 12570
rect 45798 12518 45800 12570
rect 45744 12516 45800 12518
rect 89860 12570 89916 12572
rect 89860 12518 89862 12570
rect 89862 12518 89914 12570
rect 89914 12518 89916 12570
rect 89860 12516 89916 12518
rect 89964 12570 90020 12572
rect 89964 12518 89966 12570
rect 89966 12518 90018 12570
rect 90018 12518 90020 12570
rect 89964 12516 90020 12518
rect 90068 12570 90124 12572
rect 90068 12518 90070 12570
rect 90070 12518 90122 12570
rect 90122 12518 90124 12570
rect 90068 12516 90124 12518
rect 134184 12570 134240 12572
rect 134184 12518 134186 12570
rect 134186 12518 134238 12570
rect 134238 12518 134240 12570
rect 134184 12516 134240 12518
rect 134288 12570 134344 12572
rect 134288 12518 134290 12570
rect 134290 12518 134342 12570
rect 134342 12518 134344 12570
rect 134288 12516 134344 12518
rect 134392 12570 134448 12572
rect 134392 12518 134394 12570
rect 134394 12518 134446 12570
rect 134446 12518 134448 12570
rect 134392 12516 134448 12518
rect 178508 12570 178564 12572
rect 178508 12518 178510 12570
rect 178510 12518 178562 12570
rect 178562 12518 178564 12570
rect 178508 12516 178564 12518
rect 178612 12570 178668 12572
rect 178612 12518 178614 12570
rect 178614 12518 178666 12570
rect 178666 12518 178668 12570
rect 178612 12516 178668 12518
rect 178716 12570 178772 12572
rect 178716 12518 178718 12570
rect 178718 12518 178770 12570
rect 178770 12518 178772 12570
rect 178716 12516 178772 12518
rect 23374 11786 23430 11788
rect 23374 11734 23376 11786
rect 23376 11734 23428 11786
rect 23428 11734 23430 11786
rect 23374 11732 23430 11734
rect 23478 11786 23534 11788
rect 23478 11734 23480 11786
rect 23480 11734 23532 11786
rect 23532 11734 23534 11786
rect 23478 11732 23534 11734
rect 23582 11786 23638 11788
rect 23582 11734 23584 11786
rect 23584 11734 23636 11786
rect 23636 11734 23638 11786
rect 23582 11732 23638 11734
rect 67698 11786 67754 11788
rect 67698 11734 67700 11786
rect 67700 11734 67752 11786
rect 67752 11734 67754 11786
rect 67698 11732 67754 11734
rect 67802 11786 67858 11788
rect 67802 11734 67804 11786
rect 67804 11734 67856 11786
rect 67856 11734 67858 11786
rect 67802 11732 67858 11734
rect 67906 11786 67962 11788
rect 67906 11734 67908 11786
rect 67908 11734 67960 11786
rect 67960 11734 67962 11786
rect 67906 11732 67962 11734
rect 112022 11786 112078 11788
rect 112022 11734 112024 11786
rect 112024 11734 112076 11786
rect 112076 11734 112078 11786
rect 112022 11732 112078 11734
rect 112126 11786 112182 11788
rect 112126 11734 112128 11786
rect 112128 11734 112180 11786
rect 112180 11734 112182 11786
rect 112126 11732 112182 11734
rect 112230 11786 112286 11788
rect 112230 11734 112232 11786
rect 112232 11734 112284 11786
rect 112284 11734 112286 11786
rect 112230 11732 112286 11734
rect 156346 11786 156402 11788
rect 156346 11734 156348 11786
rect 156348 11734 156400 11786
rect 156400 11734 156402 11786
rect 156346 11732 156402 11734
rect 156450 11786 156506 11788
rect 156450 11734 156452 11786
rect 156452 11734 156504 11786
rect 156504 11734 156506 11786
rect 156450 11732 156506 11734
rect 156554 11786 156610 11788
rect 156554 11734 156556 11786
rect 156556 11734 156608 11786
rect 156608 11734 156610 11786
rect 156554 11732 156610 11734
rect 45536 11002 45592 11004
rect 45536 10950 45538 11002
rect 45538 10950 45590 11002
rect 45590 10950 45592 11002
rect 45536 10948 45592 10950
rect 45640 11002 45696 11004
rect 45640 10950 45642 11002
rect 45642 10950 45694 11002
rect 45694 10950 45696 11002
rect 45640 10948 45696 10950
rect 45744 11002 45800 11004
rect 45744 10950 45746 11002
rect 45746 10950 45798 11002
rect 45798 10950 45800 11002
rect 45744 10948 45800 10950
rect 89860 11002 89916 11004
rect 89860 10950 89862 11002
rect 89862 10950 89914 11002
rect 89914 10950 89916 11002
rect 89860 10948 89916 10950
rect 89964 11002 90020 11004
rect 89964 10950 89966 11002
rect 89966 10950 90018 11002
rect 90018 10950 90020 11002
rect 89964 10948 90020 10950
rect 90068 11002 90124 11004
rect 90068 10950 90070 11002
rect 90070 10950 90122 11002
rect 90122 10950 90124 11002
rect 90068 10948 90124 10950
rect 134184 11002 134240 11004
rect 134184 10950 134186 11002
rect 134186 10950 134238 11002
rect 134238 10950 134240 11002
rect 134184 10948 134240 10950
rect 134288 11002 134344 11004
rect 134288 10950 134290 11002
rect 134290 10950 134342 11002
rect 134342 10950 134344 11002
rect 134288 10948 134344 10950
rect 134392 11002 134448 11004
rect 134392 10950 134394 11002
rect 134394 10950 134446 11002
rect 134446 10950 134448 11002
rect 134392 10948 134448 10950
rect 178508 11002 178564 11004
rect 178508 10950 178510 11002
rect 178510 10950 178562 11002
rect 178562 10950 178564 11002
rect 178508 10948 178564 10950
rect 178612 11002 178668 11004
rect 178612 10950 178614 11002
rect 178614 10950 178666 11002
rect 178666 10950 178668 11002
rect 178612 10948 178668 10950
rect 178716 11002 178772 11004
rect 178716 10950 178718 11002
rect 178718 10950 178770 11002
rect 178770 10950 178772 11002
rect 178716 10948 178772 10950
rect 23374 10218 23430 10220
rect 23374 10166 23376 10218
rect 23376 10166 23428 10218
rect 23428 10166 23430 10218
rect 23374 10164 23430 10166
rect 23478 10218 23534 10220
rect 23478 10166 23480 10218
rect 23480 10166 23532 10218
rect 23532 10166 23534 10218
rect 23478 10164 23534 10166
rect 23582 10218 23638 10220
rect 23582 10166 23584 10218
rect 23584 10166 23636 10218
rect 23636 10166 23638 10218
rect 23582 10164 23638 10166
rect 67698 10218 67754 10220
rect 67698 10166 67700 10218
rect 67700 10166 67752 10218
rect 67752 10166 67754 10218
rect 67698 10164 67754 10166
rect 67802 10218 67858 10220
rect 67802 10166 67804 10218
rect 67804 10166 67856 10218
rect 67856 10166 67858 10218
rect 67802 10164 67858 10166
rect 67906 10218 67962 10220
rect 67906 10166 67908 10218
rect 67908 10166 67960 10218
rect 67960 10166 67962 10218
rect 67906 10164 67962 10166
rect 112022 10218 112078 10220
rect 112022 10166 112024 10218
rect 112024 10166 112076 10218
rect 112076 10166 112078 10218
rect 112022 10164 112078 10166
rect 112126 10218 112182 10220
rect 112126 10166 112128 10218
rect 112128 10166 112180 10218
rect 112180 10166 112182 10218
rect 112126 10164 112182 10166
rect 112230 10218 112286 10220
rect 112230 10166 112232 10218
rect 112232 10166 112284 10218
rect 112284 10166 112286 10218
rect 112230 10164 112286 10166
rect 156346 10218 156402 10220
rect 156346 10166 156348 10218
rect 156348 10166 156400 10218
rect 156400 10166 156402 10218
rect 156346 10164 156402 10166
rect 156450 10218 156506 10220
rect 156450 10166 156452 10218
rect 156452 10166 156504 10218
rect 156504 10166 156506 10218
rect 156450 10164 156506 10166
rect 156554 10218 156610 10220
rect 156554 10166 156556 10218
rect 156556 10166 156608 10218
rect 156608 10166 156610 10218
rect 156554 10164 156610 10166
rect 45536 9434 45592 9436
rect 45536 9382 45538 9434
rect 45538 9382 45590 9434
rect 45590 9382 45592 9434
rect 45536 9380 45592 9382
rect 45640 9434 45696 9436
rect 45640 9382 45642 9434
rect 45642 9382 45694 9434
rect 45694 9382 45696 9434
rect 45640 9380 45696 9382
rect 45744 9434 45800 9436
rect 45744 9382 45746 9434
rect 45746 9382 45798 9434
rect 45798 9382 45800 9434
rect 45744 9380 45800 9382
rect 89860 9434 89916 9436
rect 89860 9382 89862 9434
rect 89862 9382 89914 9434
rect 89914 9382 89916 9434
rect 89860 9380 89916 9382
rect 89964 9434 90020 9436
rect 89964 9382 89966 9434
rect 89966 9382 90018 9434
rect 90018 9382 90020 9434
rect 89964 9380 90020 9382
rect 90068 9434 90124 9436
rect 90068 9382 90070 9434
rect 90070 9382 90122 9434
rect 90122 9382 90124 9434
rect 90068 9380 90124 9382
rect 134184 9434 134240 9436
rect 134184 9382 134186 9434
rect 134186 9382 134238 9434
rect 134238 9382 134240 9434
rect 134184 9380 134240 9382
rect 134288 9434 134344 9436
rect 134288 9382 134290 9434
rect 134290 9382 134342 9434
rect 134342 9382 134344 9434
rect 134288 9380 134344 9382
rect 134392 9434 134448 9436
rect 134392 9382 134394 9434
rect 134394 9382 134446 9434
rect 134446 9382 134448 9434
rect 134392 9380 134448 9382
rect 178508 9434 178564 9436
rect 178508 9382 178510 9434
rect 178510 9382 178562 9434
rect 178562 9382 178564 9434
rect 178508 9380 178564 9382
rect 178612 9434 178668 9436
rect 178612 9382 178614 9434
rect 178614 9382 178666 9434
rect 178666 9382 178668 9434
rect 178612 9380 178668 9382
rect 178716 9434 178772 9436
rect 178716 9382 178718 9434
rect 178718 9382 178770 9434
rect 178770 9382 178772 9434
rect 178716 9380 178772 9382
rect 23374 8650 23430 8652
rect 23374 8598 23376 8650
rect 23376 8598 23428 8650
rect 23428 8598 23430 8650
rect 23374 8596 23430 8598
rect 23478 8650 23534 8652
rect 23478 8598 23480 8650
rect 23480 8598 23532 8650
rect 23532 8598 23534 8650
rect 23478 8596 23534 8598
rect 23582 8650 23638 8652
rect 23582 8598 23584 8650
rect 23584 8598 23636 8650
rect 23636 8598 23638 8650
rect 23582 8596 23638 8598
rect 67698 8650 67754 8652
rect 67698 8598 67700 8650
rect 67700 8598 67752 8650
rect 67752 8598 67754 8650
rect 67698 8596 67754 8598
rect 67802 8650 67858 8652
rect 67802 8598 67804 8650
rect 67804 8598 67856 8650
rect 67856 8598 67858 8650
rect 67802 8596 67858 8598
rect 67906 8650 67962 8652
rect 67906 8598 67908 8650
rect 67908 8598 67960 8650
rect 67960 8598 67962 8650
rect 67906 8596 67962 8598
rect 112022 8650 112078 8652
rect 112022 8598 112024 8650
rect 112024 8598 112076 8650
rect 112076 8598 112078 8650
rect 112022 8596 112078 8598
rect 112126 8650 112182 8652
rect 112126 8598 112128 8650
rect 112128 8598 112180 8650
rect 112180 8598 112182 8650
rect 112126 8596 112182 8598
rect 112230 8650 112286 8652
rect 112230 8598 112232 8650
rect 112232 8598 112284 8650
rect 112284 8598 112286 8650
rect 112230 8596 112286 8598
rect 156346 8650 156402 8652
rect 156346 8598 156348 8650
rect 156348 8598 156400 8650
rect 156400 8598 156402 8650
rect 156346 8596 156402 8598
rect 156450 8650 156506 8652
rect 156450 8598 156452 8650
rect 156452 8598 156504 8650
rect 156504 8598 156506 8650
rect 156450 8596 156506 8598
rect 156554 8650 156610 8652
rect 156554 8598 156556 8650
rect 156556 8598 156608 8650
rect 156608 8598 156610 8650
rect 156554 8596 156610 8598
rect 45536 7866 45592 7868
rect 45536 7814 45538 7866
rect 45538 7814 45590 7866
rect 45590 7814 45592 7866
rect 45536 7812 45592 7814
rect 45640 7866 45696 7868
rect 45640 7814 45642 7866
rect 45642 7814 45694 7866
rect 45694 7814 45696 7866
rect 45640 7812 45696 7814
rect 45744 7866 45800 7868
rect 45744 7814 45746 7866
rect 45746 7814 45798 7866
rect 45798 7814 45800 7866
rect 45744 7812 45800 7814
rect 89860 7866 89916 7868
rect 89860 7814 89862 7866
rect 89862 7814 89914 7866
rect 89914 7814 89916 7866
rect 89860 7812 89916 7814
rect 89964 7866 90020 7868
rect 89964 7814 89966 7866
rect 89966 7814 90018 7866
rect 90018 7814 90020 7866
rect 89964 7812 90020 7814
rect 90068 7866 90124 7868
rect 90068 7814 90070 7866
rect 90070 7814 90122 7866
rect 90122 7814 90124 7866
rect 90068 7812 90124 7814
rect 134184 7866 134240 7868
rect 134184 7814 134186 7866
rect 134186 7814 134238 7866
rect 134238 7814 134240 7866
rect 134184 7812 134240 7814
rect 134288 7866 134344 7868
rect 134288 7814 134290 7866
rect 134290 7814 134342 7866
rect 134342 7814 134344 7866
rect 134288 7812 134344 7814
rect 134392 7866 134448 7868
rect 134392 7814 134394 7866
rect 134394 7814 134446 7866
rect 134446 7814 134448 7866
rect 134392 7812 134448 7814
rect 178508 7866 178564 7868
rect 178508 7814 178510 7866
rect 178510 7814 178562 7866
rect 178562 7814 178564 7866
rect 178508 7812 178564 7814
rect 178612 7866 178668 7868
rect 178612 7814 178614 7866
rect 178614 7814 178666 7866
rect 178666 7814 178668 7866
rect 178612 7812 178668 7814
rect 178716 7866 178772 7868
rect 178716 7814 178718 7866
rect 178718 7814 178770 7866
rect 178770 7814 178772 7866
rect 178716 7812 178772 7814
rect 23374 7082 23430 7084
rect 23374 7030 23376 7082
rect 23376 7030 23428 7082
rect 23428 7030 23430 7082
rect 23374 7028 23430 7030
rect 23478 7082 23534 7084
rect 23478 7030 23480 7082
rect 23480 7030 23532 7082
rect 23532 7030 23534 7082
rect 23478 7028 23534 7030
rect 23582 7082 23638 7084
rect 23582 7030 23584 7082
rect 23584 7030 23636 7082
rect 23636 7030 23638 7082
rect 23582 7028 23638 7030
rect 51548 6412 51604 6468
rect 45536 6298 45592 6300
rect 45536 6246 45538 6298
rect 45538 6246 45590 6298
rect 45590 6246 45592 6298
rect 45536 6244 45592 6246
rect 45640 6298 45696 6300
rect 45640 6246 45642 6298
rect 45642 6246 45694 6298
rect 45694 6246 45696 6298
rect 45640 6244 45696 6246
rect 45744 6298 45800 6300
rect 45744 6246 45746 6298
rect 45746 6246 45798 6298
rect 45798 6246 45800 6298
rect 45744 6244 45800 6246
rect 23374 5514 23430 5516
rect 23374 5462 23376 5514
rect 23376 5462 23428 5514
rect 23428 5462 23430 5514
rect 23374 5460 23430 5462
rect 23478 5514 23534 5516
rect 23478 5462 23480 5514
rect 23480 5462 23532 5514
rect 23532 5462 23534 5514
rect 23478 5460 23534 5462
rect 23582 5514 23638 5516
rect 23582 5462 23584 5514
rect 23584 5462 23636 5514
rect 23636 5462 23638 5514
rect 23582 5460 23638 5462
rect 49196 5234 49252 5236
rect 49196 5182 49198 5234
rect 49198 5182 49250 5234
rect 49250 5182 49252 5234
rect 49196 5180 49252 5182
rect 9660 3724 9716 3780
rect 12572 3554 12628 3556
rect 12572 3502 12574 3554
rect 12574 3502 12626 3554
rect 12626 3502 12628 3554
rect 12572 3500 12628 3502
rect 23374 3946 23430 3948
rect 23374 3894 23376 3946
rect 23376 3894 23428 3946
rect 23428 3894 23430 3946
rect 23374 3892 23430 3894
rect 23478 3946 23534 3948
rect 23478 3894 23480 3946
rect 23480 3894 23532 3946
rect 23532 3894 23534 3946
rect 23478 3892 23534 3894
rect 23582 3946 23638 3948
rect 23582 3894 23584 3946
rect 23584 3894 23636 3946
rect 23636 3894 23638 3946
rect 23582 3892 23638 3894
rect 13020 3500 13076 3556
rect 25340 3554 25396 3556
rect 25340 3502 25342 3554
rect 25342 3502 25394 3554
rect 25394 3502 25396 3554
rect 25340 3500 25396 3502
rect 11788 3442 11844 3444
rect 11788 3390 11790 3442
rect 11790 3390 11842 3442
rect 11842 3390 11844 3442
rect 11788 3388 11844 3390
rect 14252 3442 14308 3444
rect 14252 3390 14254 3442
rect 14254 3390 14306 3442
rect 14306 3390 14308 3442
rect 14252 3388 14308 3390
rect 12684 3276 12740 3332
rect 13580 3330 13636 3332
rect 13580 3278 13582 3330
rect 13582 3278 13634 3330
rect 13634 3278 13636 3330
rect 13580 3276 13636 3278
rect 26124 3442 26180 3444
rect 26124 3390 26126 3442
rect 26126 3390 26178 3442
rect 26178 3390 26180 3442
rect 26124 3388 26180 3390
rect 14252 2940 14308 2996
rect 32956 4396 33012 4452
rect 28252 3666 28308 3668
rect 28252 3614 28254 3666
rect 28254 3614 28306 3666
rect 28306 3614 28308 3666
rect 28252 3612 28308 3614
rect 30828 3724 30884 3780
rect 33516 4450 33572 4452
rect 33516 4398 33518 4450
rect 33518 4398 33570 4450
rect 33570 4398 33572 4450
rect 33516 4396 33572 4398
rect 32060 4226 32116 4228
rect 32060 4174 32062 4226
rect 32062 4174 32114 4226
rect 32114 4174 32116 4226
rect 32060 4172 32116 4174
rect 35196 5122 35252 5124
rect 35196 5070 35198 5122
rect 35198 5070 35250 5122
rect 35250 5070 35252 5122
rect 35196 5068 35252 5070
rect 35532 5122 35588 5124
rect 35532 5070 35534 5122
rect 35534 5070 35586 5122
rect 35586 5070 35588 5122
rect 35532 5068 35588 5070
rect 36876 5068 36932 5124
rect 48524 5122 48580 5124
rect 48524 5070 48526 5122
rect 48526 5070 48578 5122
rect 48578 5070 48580 5122
rect 48524 5068 48580 5070
rect 45536 4730 45592 4732
rect 45536 4678 45538 4730
rect 45538 4678 45590 4730
rect 45590 4678 45592 4730
rect 45536 4676 45592 4678
rect 45640 4730 45696 4732
rect 45640 4678 45642 4730
rect 45642 4678 45694 4730
rect 45694 4678 45696 4730
rect 45640 4676 45696 4678
rect 45744 4730 45800 4732
rect 45744 4678 45746 4730
rect 45746 4678 45798 4730
rect 45798 4678 45800 4730
rect 45744 4676 45800 4678
rect 35532 4396 35588 4452
rect 34300 4172 34356 4228
rect 33628 3948 33684 4004
rect 34412 3948 34468 4004
rect 34860 4284 34916 4340
rect 31276 3724 31332 3780
rect 31948 3724 32004 3780
rect 32508 3666 32564 3668
rect 32508 3614 32510 3666
rect 32510 3614 32562 3666
rect 32562 3614 32564 3666
rect 32508 3612 32564 3614
rect 34076 3612 34132 3668
rect 29260 3554 29316 3556
rect 29260 3502 29262 3554
rect 29262 3502 29314 3554
rect 29314 3502 29316 3554
rect 29260 3500 29316 3502
rect 35196 4338 35252 4340
rect 35196 4286 35198 4338
rect 35198 4286 35250 4338
rect 35250 4286 35252 4338
rect 35196 4284 35252 4286
rect 49196 4284 49252 4340
rect 50428 5122 50484 5124
rect 50428 5070 50430 5122
rect 50430 5070 50482 5122
rect 50482 5070 50484 5122
rect 50428 5068 50484 5070
rect 55468 5292 55524 5348
rect 51548 5068 51604 5124
rect 55692 5122 55748 5124
rect 55692 5070 55694 5122
rect 55694 5070 55746 5122
rect 55746 5070 55748 5122
rect 55692 5068 55748 5070
rect 64092 6802 64148 6804
rect 64092 6750 64094 6802
rect 64094 6750 64146 6802
rect 64146 6750 64148 6802
rect 64092 6748 64148 6750
rect 64540 6802 64596 6804
rect 64540 6750 64542 6802
rect 64542 6750 64594 6802
rect 64594 6750 64596 6802
rect 64540 6748 64596 6750
rect 56700 5292 56756 5348
rect 56364 5122 56420 5124
rect 56364 5070 56366 5122
rect 56366 5070 56418 5122
rect 56418 5070 56420 5122
rect 56364 5068 56420 5070
rect 50316 4226 50372 4228
rect 50316 4174 50318 4226
rect 50318 4174 50370 4226
rect 50370 4174 50372 4226
rect 50316 4172 50372 4174
rect 49756 3612 49812 3668
rect 52780 3666 52836 3668
rect 52780 3614 52782 3666
rect 52782 3614 52834 3666
rect 52834 3614 52836 3666
rect 52780 3612 52836 3614
rect 28700 3388 28756 3444
rect 28700 2828 28756 2884
rect 34524 3276 34580 3332
rect 36204 3330 36260 3332
rect 36204 3278 36206 3330
rect 36206 3278 36258 3330
rect 36258 3278 36260 3330
rect 36204 3276 36260 3278
rect 36204 1708 36260 1764
rect 37100 1708 37156 1764
rect 45536 3162 45592 3164
rect 45536 3110 45538 3162
rect 45538 3110 45590 3162
rect 45590 3110 45592 3162
rect 45536 3108 45592 3110
rect 45640 3162 45696 3164
rect 45640 3110 45642 3162
rect 45642 3110 45694 3162
rect 45694 3110 45696 3162
rect 45640 3108 45696 3110
rect 45744 3162 45800 3164
rect 45744 3110 45746 3162
rect 45746 3110 45798 3162
rect 45798 3110 45800 3162
rect 45744 3108 45800 3110
rect 47964 3276 48020 3332
rect 48860 3330 48916 3332
rect 48860 3278 48862 3330
rect 48862 3278 48914 3330
rect 48914 3278 48916 3330
rect 48860 3276 48916 3278
rect 54348 3612 54404 3668
rect 57484 5292 57540 5348
rect 57260 5122 57316 5124
rect 57260 5070 57262 5122
rect 57262 5070 57314 5122
rect 57314 5070 57316 5122
rect 57260 5068 57316 5070
rect 55804 4226 55860 4228
rect 55804 4174 55806 4226
rect 55806 4174 55858 4226
rect 55858 4174 55860 4226
rect 55804 4172 55860 4174
rect 54908 4060 54964 4116
rect 54908 3666 54964 3668
rect 54908 3614 54910 3666
rect 54910 3614 54962 3666
rect 54962 3614 54964 3666
rect 54908 3612 54964 3614
rect 57932 5292 57988 5348
rect 58380 5292 58436 5348
rect 57596 5068 57652 5124
rect 58268 5068 58324 5124
rect 55692 3554 55748 3556
rect 55692 3502 55694 3554
rect 55694 3502 55746 3554
rect 55746 3502 55748 3554
rect 55692 3500 55748 3502
rect 58716 5292 58772 5348
rect 59276 5292 59332 5348
rect 58492 5068 58548 5124
rect 58716 5068 58772 5124
rect 59052 5122 59108 5124
rect 59052 5070 59054 5122
rect 59054 5070 59106 5122
rect 59106 5070 59108 5122
rect 59052 5068 59108 5070
rect 59612 6412 59668 6468
rect 60060 6466 60116 6468
rect 60060 6414 60062 6466
rect 60062 6414 60114 6466
rect 60114 6414 60116 6466
rect 60060 6412 60116 6414
rect 61180 6412 61236 6468
rect 60732 5906 60788 5908
rect 60732 5854 60734 5906
rect 60734 5854 60786 5906
rect 60786 5854 60788 5906
rect 60732 5852 60788 5854
rect 60172 5292 60228 5348
rect 60620 5234 60676 5236
rect 60620 5182 60622 5234
rect 60622 5182 60674 5234
rect 60674 5182 60676 5234
rect 60620 5180 60676 5182
rect 62188 5852 62244 5908
rect 61740 5292 61796 5348
rect 61180 5180 61236 5236
rect 59836 5068 59892 5124
rect 61404 5234 61460 5236
rect 61404 5182 61406 5234
rect 61406 5182 61458 5234
rect 61458 5182 61460 5234
rect 61404 5180 61460 5182
rect 61964 5180 62020 5236
rect 63756 5906 63812 5908
rect 63756 5854 63758 5906
rect 63758 5854 63810 5906
rect 63810 5854 63812 5906
rect 63756 5852 63812 5854
rect 65100 6802 65156 6804
rect 65100 6750 65102 6802
rect 65102 6750 65154 6802
rect 65154 6750 65156 6802
rect 65100 6748 65156 6750
rect 65436 6748 65492 6804
rect 65996 6802 66052 6804
rect 65996 6750 65998 6802
rect 65998 6750 66050 6802
rect 66050 6750 66052 6802
rect 65996 6748 66052 6750
rect 65436 6412 65492 6468
rect 63532 5010 63588 5012
rect 63532 4958 63534 5010
rect 63534 4958 63586 5010
rect 63586 4958 63588 5010
rect 63532 4956 63588 4958
rect 62188 3554 62244 3556
rect 62188 3502 62190 3554
rect 62190 3502 62242 3554
rect 62242 3502 62244 3554
rect 62188 3500 62244 3502
rect 59724 3276 59780 3332
rect 60620 3330 60676 3332
rect 60620 3278 60622 3330
rect 60622 3278 60674 3330
rect 60674 3278 60676 3330
rect 60620 3276 60676 3278
rect 62860 3442 62916 3444
rect 62860 3390 62862 3442
rect 62862 3390 62914 3442
rect 62914 3390 62916 3442
rect 62860 3388 62916 3390
rect 62076 3276 62132 3332
rect 63532 4284 63588 4340
rect 65324 5852 65380 5908
rect 64428 4956 64484 5012
rect 66108 6466 66164 6468
rect 66108 6414 66110 6466
rect 66110 6414 66162 6466
rect 66162 6414 66164 6466
rect 66108 6412 66164 6414
rect 66332 6748 66388 6804
rect 65660 5906 65716 5908
rect 65660 5854 65662 5906
rect 65662 5854 65714 5906
rect 65714 5854 65716 5906
rect 65660 5852 65716 5854
rect 66220 5906 66276 5908
rect 66220 5854 66222 5906
rect 66222 5854 66274 5906
rect 66274 5854 66276 5906
rect 66220 5852 66276 5854
rect 65436 4898 65492 4900
rect 65436 4846 65438 4898
rect 65438 4846 65490 4898
rect 65490 4846 65492 4898
rect 65436 4844 65492 4846
rect 63756 3612 63812 3668
rect 64652 4338 64708 4340
rect 64652 4286 64654 4338
rect 64654 4286 64706 4338
rect 64706 4286 64708 4338
rect 64652 4284 64708 4286
rect 64876 4284 64932 4340
rect 66108 5068 66164 5124
rect 65436 4284 65492 4340
rect 65324 3612 65380 3668
rect 64876 3388 64932 3444
rect 63420 3330 63476 3332
rect 63420 3278 63422 3330
rect 63422 3278 63474 3330
rect 63474 3278 63476 3330
rect 63420 3276 63476 3278
rect 67228 6748 67284 6804
rect 67004 6466 67060 6468
rect 67004 6414 67006 6466
rect 67006 6414 67058 6466
rect 67058 6414 67060 6466
rect 67004 6412 67060 6414
rect 67452 6412 67508 6468
rect 67452 5794 67508 5796
rect 67452 5742 67454 5794
rect 67454 5742 67506 5794
rect 67506 5742 67508 5794
rect 67452 5740 67508 5742
rect 66332 4898 66388 4900
rect 66332 4846 66334 4898
rect 66334 4846 66386 4898
rect 66386 4846 66388 4898
rect 66332 4844 66388 4846
rect 67116 4956 67172 5012
rect 66444 3500 66500 3556
rect 67698 7082 67754 7084
rect 67698 7030 67700 7082
rect 67700 7030 67752 7082
rect 67752 7030 67754 7082
rect 67698 7028 67754 7030
rect 67802 7082 67858 7084
rect 67802 7030 67804 7082
rect 67804 7030 67856 7082
rect 67856 7030 67858 7082
rect 67802 7028 67858 7030
rect 67906 7082 67962 7084
rect 67906 7030 67908 7082
rect 67908 7030 67960 7082
rect 67960 7030 67962 7082
rect 67906 7028 67962 7030
rect 112022 7082 112078 7084
rect 112022 7030 112024 7082
rect 112024 7030 112076 7082
rect 112076 7030 112078 7082
rect 112022 7028 112078 7030
rect 112126 7082 112182 7084
rect 112126 7030 112128 7082
rect 112128 7030 112180 7082
rect 112180 7030 112182 7082
rect 112126 7028 112182 7030
rect 112230 7082 112286 7084
rect 112230 7030 112232 7082
rect 112232 7030 112284 7082
rect 112284 7030 112286 7082
rect 112230 7028 112286 7030
rect 156346 7082 156402 7084
rect 156346 7030 156348 7082
rect 156348 7030 156400 7082
rect 156400 7030 156402 7082
rect 156346 7028 156402 7030
rect 156450 7082 156506 7084
rect 156450 7030 156452 7082
rect 156452 7030 156504 7082
rect 156504 7030 156506 7082
rect 156450 7028 156506 7030
rect 156554 7082 156610 7084
rect 156554 7030 156556 7082
rect 156556 7030 156608 7082
rect 156608 7030 156610 7082
rect 156554 7028 156610 7030
rect 67676 6748 67732 6804
rect 96012 6412 96068 6468
rect 89860 6298 89916 6300
rect 89860 6246 89862 6298
rect 89862 6246 89914 6298
rect 89914 6246 89916 6298
rect 89860 6244 89916 6246
rect 89964 6298 90020 6300
rect 89964 6246 89966 6298
rect 89966 6246 90018 6298
rect 90018 6246 90020 6298
rect 89964 6244 90020 6246
rect 90068 6298 90124 6300
rect 90068 6246 90070 6298
rect 90070 6246 90122 6298
rect 90122 6246 90124 6298
rect 90068 6244 90124 6246
rect 96348 6466 96404 6468
rect 96348 6414 96350 6466
rect 96350 6414 96402 6466
rect 96402 6414 96404 6466
rect 96348 6412 96404 6414
rect 67698 5514 67754 5516
rect 67698 5462 67700 5514
rect 67700 5462 67752 5514
rect 67752 5462 67754 5514
rect 67698 5460 67754 5462
rect 67802 5514 67858 5516
rect 67802 5462 67804 5514
rect 67804 5462 67856 5514
rect 67856 5462 67858 5514
rect 67802 5460 67858 5462
rect 67906 5514 67962 5516
rect 67906 5462 67908 5514
rect 67908 5462 67960 5514
rect 67960 5462 67962 5514
rect 67906 5460 67962 5462
rect 68348 5794 68404 5796
rect 68348 5742 68350 5794
rect 68350 5742 68402 5794
rect 68402 5742 68404 5794
rect 68348 5740 68404 5742
rect 67564 5010 67620 5012
rect 67564 4958 67566 5010
rect 67566 4958 67618 5010
rect 67618 4958 67620 5010
rect 67564 4956 67620 4958
rect 75852 5404 75908 5460
rect 69244 5122 69300 5124
rect 69244 5070 69246 5122
rect 69246 5070 69298 5122
rect 69298 5070 69300 5122
rect 69244 5068 69300 5070
rect 68460 4956 68516 5012
rect 69580 4956 69636 5012
rect 68460 4284 68516 4340
rect 67228 4060 67284 4116
rect 69356 4338 69412 4340
rect 69356 4286 69358 4338
rect 69358 4286 69410 4338
rect 69410 4286 69412 4338
rect 69356 4284 69412 4286
rect 67698 3946 67754 3948
rect 67698 3894 67700 3946
rect 67700 3894 67752 3946
rect 67752 3894 67754 3946
rect 67698 3892 67754 3894
rect 67802 3946 67858 3948
rect 67802 3894 67804 3946
rect 67804 3894 67856 3946
rect 67856 3894 67858 3946
rect 67802 3892 67858 3894
rect 67906 3946 67962 3948
rect 67906 3894 67908 3946
rect 67908 3894 67960 3946
rect 67960 3894 67962 3946
rect 67906 3892 67962 3894
rect 69804 4284 69860 4340
rect 70140 4338 70196 4340
rect 70140 4286 70142 4338
rect 70142 4286 70194 4338
rect 70194 4286 70196 4338
rect 70140 4284 70196 4286
rect 69580 4060 69636 4116
rect 69132 3724 69188 3780
rect 70476 4060 70532 4116
rect 78988 5234 79044 5236
rect 78988 5182 78990 5234
rect 78990 5182 79042 5234
rect 79042 5182 79044 5234
rect 78988 5180 79044 5182
rect 70700 3724 70756 3780
rect 68908 2828 68964 2884
rect 70588 2940 70644 2996
rect 72604 4172 72660 4228
rect 71596 3442 71652 3444
rect 71596 3390 71598 3442
rect 71598 3390 71650 3442
rect 71650 3390 71652 3442
rect 71596 3388 71652 3390
rect 74284 4450 74340 4452
rect 74284 4398 74286 4450
rect 74286 4398 74338 4450
rect 74338 4398 74340 4450
rect 74284 4396 74340 4398
rect 72492 3388 72548 3444
rect 74284 3388 74340 3444
rect 75516 3666 75572 3668
rect 75516 3614 75518 3666
rect 75518 3614 75570 3666
rect 75570 3614 75572 3666
rect 75516 3612 75572 3614
rect 74844 3388 74900 3444
rect 75404 3388 75460 3444
rect 81228 5404 81284 5460
rect 79884 5234 79940 5236
rect 79884 5182 79886 5234
rect 79886 5182 79938 5234
rect 79938 5182 79940 5234
rect 79884 5180 79940 5182
rect 79324 5068 79380 5124
rect 79660 5122 79716 5124
rect 79660 5070 79662 5122
rect 79662 5070 79714 5122
rect 79714 5070 79716 5122
rect 79660 5068 79716 5070
rect 80220 4898 80276 4900
rect 80220 4846 80222 4898
rect 80222 4846 80274 4898
rect 80274 4846 80276 4898
rect 80220 4844 80276 4846
rect 75852 4172 75908 4228
rect 75740 3388 75796 3444
rect 76300 3442 76356 3444
rect 76300 3390 76302 3442
rect 76302 3390 76354 3442
rect 76354 3390 76356 3442
rect 76300 3388 76356 3390
rect 76636 3330 76692 3332
rect 76636 3278 76638 3330
rect 76638 3278 76690 3330
rect 76690 3278 76692 3330
rect 76636 3276 76692 3278
rect 77644 2828 77700 2884
rect 79324 2940 79380 2996
rect 85708 5292 85764 5348
rect 84364 5068 84420 5124
rect 83356 5010 83412 5012
rect 83356 4958 83358 5010
rect 83358 4958 83410 5010
rect 83410 4958 83412 5010
rect 83356 4956 83412 4958
rect 83020 4898 83076 4900
rect 83020 4846 83022 4898
rect 83022 4846 83074 4898
rect 83074 4846 83076 4898
rect 83020 4844 83076 4846
rect 84028 4338 84084 4340
rect 84028 4286 84030 4338
rect 84030 4286 84082 4338
rect 84082 4286 84084 4338
rect 84028 4284 84084 4286
rect 86604 5346 86660 5348
rect 86604 5294 86606 5346
rect 86606 5294 86658 5346
rect 86658 5294 86660 5346
rect 86604 5292 86660 5294
rect 92316 5346 92372 5348
rect 92316 5294 92318 5346
rect 92318 5294 92370 5346
rect 92370 5294 92372 5346
rect 92316 5292 92372 5294
rect 94780 5346 94836 5348
rect 94780 5294 94782 5346
rect 94782 5294 94834 5346
rect 94834 5294 94836 5346
rect 94780 5292 94836 5294
rect 95900 5292 95956 5348
rect 85932 4956 85988 5012
rect 86492 4956 86548 5012
rect 89860 4730 89916 4732
rect 89860 4678 89862 4730
rect 89862 4678 89914 4730
rect 89914 4678 89916 4730
rect 89860 4676 89916 4678
rect 89964 4730 90020 4732
rect 89964 4678 89966 4730
rect 89966 4678 90018 4730
rect 90018 4678 90020 4730
rect 89964 4676 90020 4678
rect 90068 4730 90124 4732
rect 90068 4678 90070 4730
rect 90070 4678 90122 4730
rect 90122 4678 90124 4730
rect 90068 4676 90124 4678
rect 84364 4284 84420 4340
rect 83692 4226 83748 4228
rect 83692 4174 83694 4226
rect 83694 4174 83746 4226
rect 83746 4174 83748 4226
rect 83692 4172 83748 4174
rect 84588 4226 84644 4228
rect 84588 4174 84590 4226
rect 84590 4174 84642 4226
rect 84642 4174 84644 4226
rect 84588 4172 84644 4174
rect 84924 4172 84980 4228
rect 83692 3612 83748 3668
rect 81228 3554 81284 3556
rect 81228 3502 81230 3554
rect 81230 3502 81282 3554
rect 81282 3502 81284 3554
rect 81228 3500 81284 3502
rect 95564 5010 95620 5012
rect 95564 4958 95566 5010
rect 95566 4958 95618 5010
rect 95618 4958 95620 5010
rect 95564 4956 95620 4958
rect 94892 4508 94948 4564
rect 89068 4396 89124 4452
rect 85708 4060 85764 4116
rect 86492 4338 86548 4340
rect 86492 4286 86494 4338
rect 86494 4286 86546 4338
rect 86546 4286 86548 4338
rect 86492 4284 86548 4286
rect 91420 4226 91476 4228
rect 91420 4174 91422 4226
rect 91422 4174 91474 4226
rect 91474 4174 91476 4226
rect 91420 4172 91476 4174
rect 92092 4172 92148 4228
rect 89068 3612 89124 3668
rect 90636 3666 90692 3668
rect 90636 3614 90638 3666
rect 90638 3614 90690 3666
rect 90690 3614 90692 3666
rect 90636 3612 90692 3614
rect 93100 4114 93156 4116
rect 93100 4062 93102 4114
rect 93102 4062 93154 4114
rect 93154 4062 93156 4114
rect 93100 4060 93156 4062
rect 92764 3666 92820 3668
rect 92764 3614 92766 3666
rect 92766 3614 92818 3666
rect 92818 3614 92820 3666
rect 92764 3612 92820 3614
rect 92092 3554 92148 3556
rect 92092 3502 92094 3554
rect 92094 3502 92146 3554
rect 92146 3502 92148 3554
rect 92092 3500 92148 3502
rect 92764 3388 92820 3444
rect 89860 3162 89916 3164
rect 89860 3110 89862 3162
rect 89862 3110 89914 3162
rect 89914 3110 89916 3162
rect 89860 3108 89916 3110
rect 89964 3162 90020 3164
rect 89964 3110 89966 3162
rect 89966 3110 90018 3162
rect 90018 3110 90020 3162
rect 89964 3108 90020 3110
rect 90068 3162 90124 3164
rect 90068 3110 90070 3162
rect 90070 3110 90122 3162
rect 90122 3110 90124 3162
rect 90068 3108 90124 3110
rect 93660 3388 93716 3444
rect 94892 3666 94948 3668
rect 94892 3614 94894 3666
rect 94894 3614 94946 3666
rect 94946 3614 94948 3666
rect 94892 3612 94948 3614
rect 97020 6466 97076 6468
rect 97020 6414 97022 6466
rect 97022 6414 97074 6466
rect 97074 6414 97076 6466
rect 97020 6412 97076 6414
rect 97020 5628 97076 5684
rect 97244 5682 97300 5684
rect 97244 5630 97246 5682
rect 97246 5630 97298 5682
rect 97298 5630 97300 5682
rect 97244 5628 97300 5630
rect 97916 5682 97972 5684
rect 97916 5630 97918 5682
rect 97918 5630 97970 5682
rect 97970 5630 97972 5682
rect 97916 5628 97972 5630
rect 97916 5068 97972 5124
rect 97132 4844 97188 4900
rect 97244 4562 97300 4564
rect 97244 4510 97246 4562
rect 97246 4510 97298 4562
rect 97298 4510 97300 4562
rect 97244 4508 97300 4510
rect 98252 5122 98308 5124
rect 98252 5070 98254 5122
rect 98254 5070 98306 5122
rect 98306 5070 98308 5122
rect 98252 5068 98308 5070
rect 98140 5010 98196 5012
rect 98140 4958 98142 5010
rect 98142 4958 98194 5010
rect 98194 4958 98196 5010
rect 98140 4956 98196 4958
rect 98812 4898 98868 4900
rect 98812 4846 98814 4898
rect 98814 4846 98866 4898
rect 98866 4846 98868 4898
rect 98812 4844 98868 4846
rect 105196 4284 105252 4340
rect 105420 4284 105476 4340
rect 106540 5068 106596 5124
rect 105756 4338 105812 4340
rect 105756 4286 105758 4338
rect 105758 4286 105810 4338
rect 105810 4286 105812 4338
rect 105756 4284 105812 4286
rect 105196 3612 105252 3668
rect 105980 4172 106036 4228
rect 106540 4226 106596 4228
rect 106540 4174 106542 4226
rect 106542 4174 106594 4226
rect 106594 4174 106596 4226
rect 106540 4172 106596 4174
rect 106764 5122 106820 5124
rect 106764 5070 106766 5122
rect 106766 5070 106818 5122
rect 106818 5070 106820 5122
rect 106764 5068 106820 5070
rect 112022 5514 112078 5516
rect 112022 5462 112024 5514
rect 112024 5462 112076 5514
rect 112076 5462 112078 5514
rect 112022 5460 112078 5462
rect 112126 5514 112182 5516
rect 112126 5462 112128 5514
rect 112128 5462 112180 5514
rect 112180 5462 112182 5514
rect 112126 5460 112182 5462
rect 112230 5514 112286 5516
rect 112230 5462 112232 5514
rect 112232 5462 112284 5514
rect 112284 5462 112286 5514
rect 112230 5460 112286 5462
rect 113148 5292 113204 5348
rect 113708 5346 113764 5348
rect 113708 5294 113710 5346
rect 113710 5294 113762 5346
rect 113762 5294 113764 5346
rect 113708 5292 113764 5294
rect 113260 5180 113316 5236
rect 112252 5122 112308 5124
rect 112252 5070 112254 5122
rect 112254 5070 112306 5122
rect 112306 5070 112308 5122
rect 112252 5068 112308 5070
rect 107436 4844 107492 4900
rect 108108 4898 108164 4900
rect 108108 4846 108110 4898
rect 108110 4846 108162 4898
rect 108162 4846 108164 4898
rect 108108 4844 108164 4846
rect 112364 4508 112420 4564
rect 113148 4562 113204 4564
rect 113148 4510 113150 4562
rect 113150 4510 113202 4562
rect 113202 4510 113204 4562
rect 113148 4508 113204 4510
rect 114492 5292 114548 5348
rect 114268 5010 114324 5012
rect 114268 4958 114270 5010
rect 114270 4958 114322 5010
rect 114322 4958 114324 5010
rect 114268 4956 114324 4958
rect 114492 4844 114548 4900
rect 106764 4060 106820 4116
rect 105980 3554 106036 3556
rect 105980 3502 105982 3554
rect 105982 3502 106034 3554
rect 106034 3502 106036 3554
rect 105980 3500 106036 3502
rect 107772 3554 107828 3556
rect 107772 3502 107774 3554
rect 107774 3502 107826 3554
rect 107826 3502 107828 3554
rect 107772 3500 107828 3502
rect 105532 3276 105588 3332
rect 108444 3442 108500 3444
rect 108444 3390 108446 3442
rect 108446 3390 108498 3442
rect 108498 3390 108500 3442
rect 108444 3388 108500 3390
rect 115164 4844 115220 4900
rect 115724 4898 115780 4900
rect 115724 4846 115726 4898
rect 115726 4846 115778 4898
rect 115778 4846 115780 4898
rect 115724 4844 115780 4846
rect 134184 6298 134240 6300
rect 134184 6246 134186 6298
rect 134186 6246 134238 6298
rect 134238 6246 134240 6298
rect 134184 6244 134240 6246
rect 134288 6298 134344 6300
rect 134288 6246 134290 6298
rect 134290 6246 134342 6298
rect 134342 6246 134344 6298
rect 134288 6244 134344 6246
rect 134392 6298 134448 6300
rect 134392 6246 134394 6298
rect 134394 6246 134446 6298
rect 134446 6246 134448 6298
rect 134392 6244 134448 6246
rect 178508 6298 178564 6300
rect 178508 6246 178510 6298
rect 178510 6246 178562 6298
rect 178562 6246 178564 6298
rect 178508 6244 178564 6246
rect 178612 6298 178668 6300
rect 178612 6246 178614 6298
rect 178614 6246 178666 6298
rect 178666 6246 178668 6298
rect 178612 6244 178668 6246
rect 178716 6298 178772 6300
rect 178716 6246 178718 6298
rect 178718 6246 178770 6298
rect 178770 6246 178772 6298
rect 178716 6244 178772 6246
rect 156346 5514 156402 5516
rect 156346 5462 156348 5514
rect 156348 5462 156400 5514
rect 156400 5462 156402 5514
rect 156346 5460 156402 5462
rect 156450 5514 156506 5516
rect 156450 5462 156452 5514
rect 156452 5462 156504 5514
rect 156504 5462 156506 5514
rect 156450 5460 156506 5462
rect 156554 5514 156610 5516
rect 156554 5462 156556 5514
rect 156556 5462 156608 5514
rect 156608 5462 156610 5514
rect 156554 5460 156610 5462
rect 118188 4284 118244 4340
rect 118748 4338 118804 4340
rect 118748 4286 118750 4338
rect 118750 4286 118802 4338
rect 118802 4286 118804 4338
rect 118748 4284 118804 4286
rect 120540 4956 120596 5012
rect 120988 5010 121044 5012
rect 120988 4958 120990 5010
rect 120990 4958 121042 5010
rect 121042 4958 121044 5010
rect 120988 4956 121044 4958
rect 119644 4844 119700 4900
rect 112022 3946 112078 3948
rect 112022 3894 112024 3946
rect 112024 3894 112076 3946
rect 112076 3894 112078 3946
rect 112022 3892 112078 3894
rect 112126 3946 112182 3948
rect 112126 3894 112128 3946
rect 112128 3894 112180 3946
rect 112180 3894 112182 3946
rect 112126 3892 112182 3894
rect 112230 3946 112286 3948
rect 112230 3894 112232 3946
rect 112232 3894 112284 3946
rect 112284 3894 112286 3946
rect 112230 3892 112286 3894
rect 110572 3666 110628 3668
rect 110572 3614 110574 3666
rect 110574 3614 110626 3666
rect 110626 3614 110628 3666
rect 110572 3612 110628 3614
rect 119532 4226 119588 4228
rect 119532 4174 119534 4226
rect 119534 4174 119586 4226
rect 119586 4174 119588 4226
rect 119532 4172 119588 4174
rect 118188 3612 118244 3668
rect 134184 4730 134240 4732
rect 134184 4678 134186 4730
rect 134186 4678 134238 4730
rect 134238 4678 134240 4730
rect 134184 4676 134240 4678
rect 134288 4730 134344 4732
rect 134288 4678 134290 4730
rect 134290 4678 134342 4730
rect 134342 4678 134344 4730
rect 134288 4676 134344 4678
rect 134392 4730 134448 4732
rect 134392 4678 134394 4730
rect 134394 4678 134446 4730
rect 134446 4678 134448 4730
rect 134392 4676 134448 4678
rect 120428 4396 120484 4452
rect 121100 4450 121156 4452
rect 121100 4398 121102 4450
rect 121102 4398 121154 4450
rect 121154 4398 121156 4450
rect 121100 4396 121156 4398
rect 128044 4396 128100 4452
rect 119532 3724 119588 3780
rect 120540 4172 120596 4228
rect 126924 4060 126980 4116
rect 120540 3612 120596 3668
rect 121100 3724 121156 3780
rect 121548 3666 121604 3668
rect 121548 3614 121550 3666
rect 121550 3614 121602 3666
rect 121602 3614 121604 3666
rect 121548 3612 121604 3614
rect 126924 3500 126980 3556
rect 127372 3500 127428 3556
rect 119756 3442 119812 3444
rect 119756 3390 119758 3442
rect 119758 3390 119810 3442
rect 119810 3390 119812 3442
rect 119756 3388 119812 3390
rect 121324 3388 121380 3444
rect 127596 4060 127652 4116
rect 127372 2828 127428 2884
rect 129052 4450 129108 4452
rect 129052 4398 129054 4450
rect 129054 4398 129106 4450
rect 129106 4398 129108 4450
rect 129052 4396 129108 4398
rect 128268 3554 128324 3556
rect 128268 3502 128270 3554
rect 128270 3502 128322 3554
rect 128322 3502 128324 3554
rect 128268 3500 128324 3502
rect 130396 3666 130452 3668
rect 130396 3614 130398 3666
rect 130398 3614 130450 3666
rect 130450 3614 130452 3666
rect 130396 3612 130452 3614
rect 130732 3612 130788 3668
rect 131180 3612 131236 3668
rect 131404 3612 131460 3668
rect 131964 4172 132020 4228
rect 131964 3724 132020 3780
rect 139916 4226 139972 4228
rect 139916 4174 139918 4226
rect 139918 4174 139970 4226
rect 139970 4174 139972 4226
rect 139916 4172 139972 4174
rect 140364 3666 140420 3668
rect 140364 3614 140366 3666
rect 140366 3614 140418 3666
rect 140418 3614 140420 3666
rect 140364 3612 140420 3614
rect 139356 3388 139412 3444
rect 178508 4730 178564 4732
rect 178508 4678 178510 4730
rect 178510 4678 178562 4730
rect 178562 4678 178564 4730
rect 178508 4676 178564 4678
rect 178612 4730 178668 4732
rect 178612 4678 178614 4730
rect 178614 4678 178666 4730
rect 178666 4678 178668 4730
rect 178612 4676 178668 4678
rect 178716 4730 178772 4732
rect 178716 4678 178718 4730
rect 178718 4678 178770 4730
rect 178770 4678 178772 4730
rect 178716 4676 178772 4678
rect 139692 3388 139748 3444
rect 131404 3276 131460 3332
rect 133308 3330 133364 3332
rect 133308 3278 133310 3330
rect 133310 3278 133362 3330
rect 133362 3278 133364 3330
rect 133308 3276 133364 3278
rect 134184 3162 134240 3164
rect 134184 3110 134186 3162
rect 134186 3110 134238 3162
rect 134238 3110 134240 3162
rect 134184 3108 134240 3110
rect 134288 3162 134344 3164
rect 134288 3110 134290 3162
rect 134290 3110 134342 3162
rect 134342 3110 134344 3162
rect 134288 3108 134344 3110
rect 134392 3162 134448 3164
rect 134392 3110 134394 3162
rect 134394 3110 134446 3162
rect 134446 3110 134448 3162
rect 134392 3108 134448 3110
rect 139804 3276 139860 3332
rect 141708 3330 141764 3332
rect 141708 3278 141710 3330
rect 141710 3278 141762 3330
rect 141762 3278 141764 3330
rect 141708 3276 141764 3278
rect 150444 4060 150500 4116
rect 151004 3500 151060 3556
rect 142604 3388 142660 3444
rect 142940 3442 142996 3444
rect 142940 3390 142942 3442
rect 142942 3390 142994 3442
rect 142994 3390 142996 3442
rect 142940 3388 142996 3390
rect 151116 4060 151172 4116
rect 151004 2940 151060 2996
rect 151788 3554 151844 3556
rect 151788 3502 151790 3554
rect 151790 3502 151842 3554
rect 151842 3502 151844 3554
rect 151788 3500 151844 3502
rect 156346 3946 156402 3948
rect 156346 3894 156348 3946
rect 156348 3894 156400 3946
rect 156400 3894 156402 3946
rect 156346 3892 156402 3894
rect 156450 3946 156506 3948
rect 156450 3894 156452 3946
rect 156452 3894 156504 3946
rect 156504 3894 156506 3946
rect 156450 3892 156506 3894
rect 156554 3946 156610 3948
rect 156554 3894 156556 3946
rect 156556 3894 156608 3946
rect 156608 3894 156610 3946
rect 156554 3892 156610 3894
rect 153916 3388 153972 3444
rect 173964 3276 174020 3332
rect 174972 3330 175028 3332
rect 174972 3278 174974 3330
rect 174974 3278 175026 3330
rect 175026 3278 175028 3330
rect 174972 3276 175028 3278
rect 178508 3162 178564 3164
rect 178508 3110 178510 3162
rect 178510 3110 178562 3162
rect 178562 3110 178564 3162
rect 178508 3108 178564 3110
rect 178612 3162 178668 3164
rect 178612 3110 178614 3162
rect 178614 3110 178666 3162
rect 178666 3110 178668 3162
rect 178612 3108 178668 3110
rect 178716 3162 178772 3164
rect 178716 3110 178718 3162
rect 178718 3110 178770 3162
rect 178770 3110 178772 3162
rect 178716 3108 178772 3110
<< metal3 >>
rect 23364 16436 23374 16492
rect 23430 16436 23478 16492
rect 23534 16436 23582 16492
rect 23638 16436 23648 16492
rect 67688 16436 67698 16492
rect 67754 16436 67802 16492
rect 67858 16436 67906 16492
rect 67962 16436 67972 16492
rect 112012 16436 112022 16492
rect 112078 16436 112126 16492
rect 112182 16436 112230 16492
rect 112286 16436 112296 16492
rect 156336 16436 156346 16492
rect 156402 16436 156450 16492
rect 156506 16436 156554 16492
rect 156610 16436 156620 16492
rect 45526 15652 45536 15708
rect 45592 15652 45640 15708
rect 45696 15652 45744 15708
rect 45800 15652 45810 15708
rect 89850 15652 89860 15708
rect 89916 15652 89964 15708
rect 90020 15652 90068 15708
rect 90124 15652 90134 15708
rect 134174 15652 134184 15708
rect 134240 15652 134288 15708
rect 134344 15652 134392 15708
rect 134448 15652 134458 15708
rect 178498 15652 178508 15708
rect 178564 15652 178612 15708
rect 178668 15652 178716 15708
rect 178772 15652 178782 15708
rect 23364 14868 23374 14924
rect 23430 14868 23478 14924
rect 23534 14868 23582 14924
rect 23638 14868 23648 14924
rect 67688 14868 67698 14924
rect 67754 14868 67802 14924
rect 67858 14868 67906 14924
rect 67962 14868 67972 14924
rect 112012 14868 112022 14924
rect 112078 14868 112126 14924
rect 112182 14868 112230 14924
rect 112286 14868 112296 14924
rect 156336 14868 156346 14924
rect 156402 14868 156450 14924
rect 156506 14868 156554 14924
rect 156610 14868 156620 14924
rect 45526 14084 45536 14140
rect 45592 14084 45640 14140
rect 45696 14084 45744 14140
rect 45800 14084 45810 14140
rect 89850 14084 89860 14140
rect 89916 14084 89964 14140
rect 90020 14084 90068 14140
rect 90124 14084 90134 14140
rect 134174 14084 134184 14140
rect 134240 14084 134288 14140
rect 134344 14084 134392 14140
rect 134448 14084 134458 14140
rect 178498 14084 178508 14140
rect 178564 14084 178612 14140
rect 178668 14084 178716 14140
rect 178772 14084 178782 14140
rect 23364 13300 23374 13356
rect 23430 13300 23478 13356
rect 23534 13300 23582 13356
rect 23638 13300 23648 13356
rect 67688 13300 67698 13356
rect 67754 13300 67802 13356
rect 67858 13300 67906 13356
rect 67962 13300 67972 13356
rect 112012 13300 112022 13356
rect 112078 13300 112126 13356
rect 112182 13300 112230 13356
rect 112286 13300 112296 13356
rect 156336 13300 156346 13356
rect 156402 13300 156450 13356
rect 156506 13300 156554 13356
rect 156610 13300 156620 13356
rect 45526 12516 45536 12572
rect 45592 12516 45640 12572
rect 45696 12516 45744 12572
rect 45800 12516 45810 12572
rect 89850 12516 89860 12572
rect 89916 12516 89964 12572
rect 90020 12516 90068 12572
rect 90124 12516 90134 12572
rect 134174 12516 134184 12572
rect 134240 12516 134288 12572
rect 134344 12516 134392 12572
rect 134448 12516 134458 12572
rect 178498 12516 178508 12572
rect 178564 12516 178612 12572
rect 178668 12516 178716 12572
rect 178772 12516 178782 12572
rect 23364 11732 23374 11788
rect 23430 11732 23478 11788
rect 23534 11732 23582 11788
rect 23638 11732 23648 11788
rect 67688 11732 67698 11788
rect 67754 11732 67802 11788
rect 67858 11732 67906 11788
rect 67962 11732 67972 11788
rect 112012 11732 112022 11788
rect 112078 11732 112126 11788
rect 112182 11732 112230 11788
rect 112286 11732 112296 11788
rect 156336 11732 156346 11788
rect 156402 11732 156450 11788
rect 156506 11732 156554 11788
rect 156610 11732 156620 11788
rect 45526 10948 45536 11004
rect 45592 10948 45640 11004
rect 45696 10948 45744 11004
rect 45800 10948 45810 11004
rect 89850 10948 89860 11004
rect 89916 10948 89964 11004
rect 90020 10948 90068 11004
rect 90124 10948 90134 11004
rect 134174 10948 134184 11004
rect 134240 10948 134288 11004
rect 134344 10948 134392 11004
rect 134448 10948 134458 11004
rect 178498 10948 178508 11004
rect 178564 10948 178612 11004
rect 178668 10948 178716 11004
rect 178772 10948 178782 11004
rect 23364 10164 23374 10220
rect 23430 10164 23478 10220
rect 23534 10164 23582 10220
rect 23638 10164 23648 10220
rect 67688 10164 67698 10220
rect 67754 10164 67802 10220
rect 67858 10164 67906 10220
rect 67962 10164 67972 10220
rect 112012 10164 112022 10220
rect 112078 10164 112126 10220
rect 112182 10164 112230 10220
rect 112286 10164 112296 10220
rect 156336 10164 156346 10220
rect 156402 10164 156450 10220
rect 156506 10164 156554 10220
rect 156610 10164 156620 10220
rect 45526 9380 45536 9436
rect 45592 9380 45640 9436
rect 45696 9380 45744 9436
rect 45800 9380 45810 9436
rect 89850 9380 89860 9436
rect 89916 9380 89964 9436
rect 90020 9380 90068 9436
rect 90124 9380 90134 9436
rect 134174 9380 134184 9436
rect 134240 9380 134288 9436
rect 134344 9380 134392 9436
rect 134448 9380 134458 9436
rect 178498 9380 178508 9436
rect 178564 9380 178612 9436
rect 178668 9380 178716 9436
rect 178772 9380 178782 9436
rect 23364 8596 23374 8652
rect 23430 8596 23478 8652
rect 23534 8596 23582 8652
rect 23638 8596 23648 8652
rect 67688 8596 67698 8652
rect 67754 8596 67802 8652
rect 67858 8596 67906 8652
rect 67962 8596 67972 8652
rect 112012 8596 112022 8652
rect 112078 8596 112126 8652
rect 112182 8596 112230 8652
rect 112286 8596 112296 8652
rect 156336 8596 156346 8652
rect 156402 8596 156450 8652
rect 156506 8596 156554 8652
rect 156610 8596 156620 8652
rect 45526 7812 45536 7868
rect 45592 7812 45640 7868
rect 45696 7812 45744 7868
rect 45800 7812 45810 7868
rect 89850 7812 89860 7868
rect 89916 7812 89964 7868
rect 90020 7812 90068 7868
rect 90124 7812 90134 7868
rect 134174 7812 134184 7868
rect 134240 7812 134288 7868
rect 134344 7812 134392 7868
rect 134448 7812 134458 7868
rect 178498 7812 178508 7868
rect 178564 7812 178612 7868
rect 178668 7812 178716 7868
rect 178772 7812 178782 7868
rect 23364 7028 23374 7084
rect 23430 7028 23478 7084
rect 23534 7028 23582 7084
rect 23638 7028 23648 7084
rect 67688 7028 67698 7084
rect 67754 7028 67802 7084
rect 67858 7028 67906 7084
rect 67962 7028 67972 7084
rect 112012 7028 112022 7084
rect 112078 7028 112126 7084
rect 112182 7028 112230 7084
rect 112286 7028 112296 7084
rect 156336 7028 156346 7084
rect 156402 7028 156450 7084
rect 156506 7028 156554 7084
rect 156610 7028 156620 7084
rect 64082 6748 64092 6804
rect 64148 6748 64540 6804
rect 64596 6748 65100 6804
rect 65156 6748 65436 6804
rect 65492 6748 65996 6804
rect 66052 6748 66332 6804
rect 66388 6748 67228 6804
rect 67284 6748 67676 6804
rect 67732 6748 67742 6804
rect 51538 6412 51548 6468
rect 51604 6412 59612 6468
rect 59668 6412 60060 6468
rect 60116 6412 61180 6468
rect 61236 6412 61246 6468
rect 65426 6412 65436 6468
rect 65492 6412 66108 6468
rect 66164 6412 67004 6468
rect 67060 6412 67452 6468
rect 67508 6412 67518 6468
rect 96002 6412 96012 6468
rect 96068 6412 96348 6468
rect 96404 6412 97020 6468
rect 97076 6412 97086 6468
rect 45526 6244 45536 6300
rect 45592 6244 45640 6300
rect 45696 6244 45744 6300
rect 45800 6244 45810 6300
rect 89850 6244 89860 6300
rect 89916 6244 89964 6300
rect 90020 6244 90068 6300
rect 90124 6244 90134 6300
rect 134174 6244 134184 6300
rect 134240 6244 134288 6300
rect 134344 6244 134392 6300
rect 134448 6244 134458 6300
rect 178498 6244 178508 6300
rect 178564 6244 178612 6300
rect 178668 6244 178716 6300
rect 178772 6244 178782 6300
rect 60722 5852 60732 5908
rect 60788 5852 62188 5908
rect 62244 5852 63756 5908
rect 63812 5852 65324 5908
rect 65380 5852 65660 5908
rect 65716 5852 66220 5908
rect 66276 5852 66286 5908
rect 67442 5740 67452 5796
rect 67508 5740 68348 5796
rect 68404 5740 68414 5796
rect 97010 5628 97020 5684
rect 97076 5628 97244 5684
rect 97300 5628 97916 5684
rect 97972 5628 97982 5684
rect 23364 5460 23374 5516
rect 23430 5460 23478 5516
rect 23534 5460 23582 5516
rect 23638 5460 23648 5516
rect 67688 5460 67698 5516
rect 67754 5460 67802 5516
rect 67858 5460 67906 5516
rect 67962 5460 67972 5516
rect 112012 5460 112022 5516
rect 112078 5460 112126 5516
rect 112182 5460 112230 5516
rect 112286 5460 112296 5516
rect 156336 5460 156346 5516
rect 156402 5460 156450 5516
rect 156506 5460 156554 5516
rect 156610 5460 156620 5516
rect 75842 5404 75852 5460
rect 75908 5404 81228 5460
rect 81284 5404 81294 5460
rect 55412 5236 55468 5348
rect 55524 5292 56700 5348
rect 56756 5292 57484 5348
rect 57540 5292 57932 5348
rect 57988 5292 58380 5348
rect 58436 5292 58716 5348
rect 58772 5292 59276 5348
rect 59332 5292 60172 5348
rect 60228 5292 61740 5348
rect 61796 5292 85708 5348
rect 85764 5292 86604 5348
rect 86660 5292 92316 5348
rect 92372 5292 94780 5348
rect 94836 5292 95900 5348
rect 95956 5292 95966 5348
rect 112252 5292 113148 5348
rect 113204 5292 113708 5348
rect 113764 5292 114492 5348
rect 114548 5292 114558 5348
rect 49186 5180 49196 5236
rect 49252 5180 55468 5236
rect 60610 5180 60620 5236
rect 60676 5180 61180 5236
rect 61236 5180 61404 5236
rect 61460 5180 61964 5236
rect 62020 5180 62030 5236
rect 78978 5180 78988 5236
rect 79044 5180 79884 5236
rect 79940 5180 79950 5236
rect 112252 5124 112308 5292
rect 113250 5180 113260 5236
rect 113316 5180 113326 5236
rect 35186 5068 35196 5124
rect 35252 5068 35532 5124
rect 35588 5068 36876 5124
rect 36932 5068 48524 5124
rect 48580 5068 50428 5124
rect 50484 5068 51548 5124
rect 51604 5068 51614 5124
rect 55682 5068 55692 5124
rect 55748 5068 56364 5124
rect 56420 5068 57260 5124
rect 57316 5068 57596 5124
rect 57652 5068 58268 5124
rect 58324 5068 58492 5124
rect 58548 5068 58716 5124
rect 58772 5068 59052 5124
rect 59108 5068 59836 5124
rect 59892 5068 59902 5124
rect 66098 5068 66108 5124
rect 66164 5068 69244 5124
rect 69300 5068 79324 5124
rect 79380 5068 79660 5124
rect 79716 5068 84364 5124
rect 84420 5068 84430 5124
rect 97906 5068 97916 5124
rect 97972 5068 98252 5124
rect 98308 5068 106540 5124
rect 106596 5068 106606 5124
rect 106754 5068 106764 5124
rect 106820 5068 112252 5124
rect 112308 5068 112318 5124
rect 113260 5012 113316 5180
rect 63522 4956 63532 5012
rect 63588 4956 64428 5012
rect 64484 4956 64494 5012
rect 67106 4956 67116 5012
rect 67172 4956 67564 5012
rect 67620 4956 67630 5012
rect 68450 4956 68460 5012
rect 68516 4956 69580 5012
rect 69636 4956 69646 5012
rect 83346 4956 83356 5012
rect 83412 4956 85932 5012
rect 85988 4956 86492 5012
rect 86548 4956 86558 5012
rect 95554 4956 95564 5012
rect 95620 4956 98140 5012
rect 98196 4956 98206 5012
rect 113260 4956 114268 5012
rect 114324 4956 114334 5012
rect 120530 4956 120540 5012
rect 120596 4956 120988 5012
rect 121044 4956 121054 5012
rect 65426 4844 65436 4900
rect 65492 4844 66332 4900
rect 66388 4844 66398 4900
rect 80210 4844 80220 4900
rect 80276 4844 83020 4900
rect 83076 4844 83086 4900
rect 97122 4844 97132 4900
rect 97188 4844 98812 4900
rect 98868 4844 98878 4900
rect 107426 4844 107436 4900
rect 107492 4844 108108 4900
rect 108164 4844 108174 4900
rect 114482 4844 114492 4900
rect 114548 4844 115164 4900
rect 115220 4844 115724 4900
rect 115780 4844 119644 4900
rect 119700 4844 119710 4900
rect 45526 4676 45536 4732
rect 45592 4676 45640 4732
rect 45696 4676 45744 4732
rect 45800 4676 45810 4732
rect 89850 4676 89860 4732
rect 89916 4676 89964 4732
rect 90020 4676 90068 4732
rect 90124 4676 90134 4732
rect 134174 4676 134184 4732
rect 134240 4676 134288 4732
rect 134344 4676 134392 4732
rect 134448 4676 134458 4732
rect 178498 4676 178508 4732
rect 178564 4676 178612 4732
rect 178668 4676 178716 4732
rect 178772 4676 178782 4732
rect 94882 4508 94892 4564
rect 94948 4508 97244 4564
rect 97300 4508 97310 4564
rect 112354 4508 112364 4564
rect 112420 4508 113148 4564
rect 113204 4508 113214 4564
rect 32946 4396 32956 4452
rect 33012 4396 33516 4452
rect 33572 4396 35532 4452
rect 35588 4396 35598 4452
rect 74274 4396 74284 4452
rect 74340 4396 89068 4452
rect 89124 4396 89134 4452
rect 120418 4396 120428 4452
rect 120484 4396 121100 4452
rect 121156 4396 121166 4452
rect 128034 4396 128044 4452
rect 128100 4396 129052 4452
rect 129108 4396 129118 4452
rect 34850 4284 34860 4340
rect 34916 4284 35196 4340
rect 35252 4284 49196 4340
rect 49252 4284 49262 4340
rect 55412 4284 63532 4340
rect 63588 4284 64652 4340
rect 64708 4284 64876 4340
rect 64932 4284 65436 4340
rect 65492 4284 65502 4340
rect 68450 4284 68460 4340
rect 68516 4284 69356 4340
rect 69412 4284 69804 4340
rect 69860 4284 70140 4340
rect 70196 4284 70206 4340
rect 84018 4284 84028 4340
rect 84084 4284 84364 4340
rect 84420 4284 86492 4340
rect 86548 4284 86558 4340
rect 105186 4284 105196 4340
rect 105252 4284 105420 4340
rect 105476 4284 105756 4340
rect 105812 4284 105822 4340
rect 118178 4284 118188 4340
rect 118244 4284 118748 4340
rect 118804 4284 118814 4340
rect 55412 4228 55468 4284
rect 32050 4172 32060 4228
rect 32116 4172 34300 4228
rect 34356 4172 50316 4228
rect 50372 4172 55468 4228
rect 55794 4172 55804 4228
rect 55860 4172 72604 4228
rect 72660 4172 75852 4228
rect 75908 4172 75918 4228
rect 83682 4172 83692 4228
rect 83748 4172 84588 4228
rect 84644 4172 84924 4228
rect 84980 4172 84990 4228
rect 91410 4172 91420 4228
rect 91476 4172 92092 4228
rect 92148 4172 105980 4228
rect 106036 4172 106046 4228
rect 106530 4172 106540 4228
rect 106596 4172 119532 4228
rect 119588 4172 120540 4228
rect 120596 4172 120606 4228
rect 131954 4172 131964 4228
rect 132020 4172 139916 4228
rect 139972 4172 139982 4228
rect 54898 4060 54908 4116
rect 54964 4060 67228 4116
rect 67284 4060 67294 4116
rect 69570 4060 69580 4116
rect 69636 4060 70476 4116
rect 70532 4060 85708 4116
rect 85764 4060 93100 4116
rect 93156 4060 106764 4116
rect 106820 4060 106830 4116
rect 126914 4060 126924 4116
rect 126980 4060 127596 4116
rect 127652 4060 150444 4116
rect 150500 4060 151116 4116
rect 151172 4060 151182 4116
rect 32172 3948 33628 4004
rect 33684 3948 34412 4004
rect 34468 3948 34478 4004
rect 23364 3892 23374 3948
rect 23430 3892 23478 3948
rect 23534 3892 23582 3948
rect 23638 3892 23648 3948
rect 9650 3724 9660 3780
rect 9716 3724 30828 3780
rect 30884 3724 31276 3780
rect 31332 3724 31948 3780
rect 32004 3724 32014 3780
rect 32172 3668 32228 3948
rect 67688 3892 67698 3948
rect 67754 3892 67802 3948
rect 67858 3892 67906 3948
rect 67962 3892 67972 3948
rect 112012 3892 112022 3948
rect 112078 3892 112126 3948
rect 112182 3892 112230 3948
rect 112286 3892 112296 3948
rect 156336 3892 156346 3948
rect 156402 3892 156450 3948
rect 156506 3892 156554 3948
rect 156610 3892 156620 3948
rect 69122 3724 69132 3780
rect 69188 3724 70700 3780
rect 70756 3724 70766 3780
rect 119522 3724 119532 3780
rect 119588 3724 121100 3780
rect 121156 3724 131964 3780
rect 132020 3724 132030 3780
rect 28242 3612 28252 3668
rect 28308 3612 32228 3668
rect 32498 3612 32508 3668
rect 32564 3612 34076 3668
rect 34132 3612 34142 3668
rect 49746 3612 49756 3668
rect 49812 3612 52780 3668
rect 52836 3612 52846 3668
rect 54338 3612 54348 3668
rect 54404 3612 54908 3668
rect 54964 3612 54974 3668
rect 63746 3612 63756 3668
rect 63812 3612 65324 3668
rect 65380 3612 65390 3668
rect 75506 3612 75516 3668
rect 75572 3612 83692 3668
rect 83748 3612 83758 3668
rect 89058 3612 89068 3668
rect 89124 3612 90636 3668
rect 90692 3612 92764 3668
rect 92820 3612 92830 3668
rect 94882 3612 94892 3668
rect 94948 3612 105196 3668
rect 105252 3612 105262 3668
rect 110562 3612 110572 3668
rect 110628 3612 118188 3668
rect 118244 3612 118254 3668
rect 120530 3612 120540 3668
rect 120596 3612 121548 3668
rect 121604 3612 130228 3668
rect 130386 3612 130396 3668
rect 130452 3612 130732 3668
rect 130788 3612 131180 3668
rect 131236 3612 131246 3668
rect 131394 3612 131404 3668
rect 131460 3612 140364 3668
rect 140420 3612 140430 3668
rect 130172 3556 130228 3612
rect 131404 3556 131460 3612
rect 12562 3500 12572 3556
rect 12628 3500 13020 3556
rect 13076 3500 25340 3556
rect 25396 3500 29260 3556
rect 29316 3500 55692 3556
rect 55748 3500 55758 3556
rect 62178 3500 62188 3556
rect 62244 3500 66444 3556
rect 66500 3500 66510 3556
rect 81218 3500 81228 3556
rect 81284 3500 92092 3556
rect 92148 3500 92158 3556
rect 105970 3500 105980 3556
rect 106036 3500 107772 3556
rect 107828 3500 126924 3556
rect 126980 3500 126990 3556
rect 127362 3500 127372 3556
rect 127428 3500 128268 3556
rect 128324 3500 128334 3556
rect 130172 3500 131460 3556
rect 150994 3500 151004 3556
rect 151060 3500 151788 3556
rect 151844 3500 151854 3556
rect 11778 3388 11788 3444
rect 11844 3388 14252 3444
rect 14308 3388 14318 3444
rect 26114 3388 26124 3444
rect 26180 3388 28700 3444
rect 28756 3388 28766 3444
rect 62850 3388 62860 3444
rect 62916 3388 64876 3444
rect 64932 3388 64942 3444
rect 71586 3388 71596 3444
rect 71652 3388 72492 3444
rect 72548 3388 72558 3444
rect 74274 3388 74284 3444
rect 74340 3388 74844 3444
rect 74900 3388 74910 3444
rect 75394 3388 75404 3444
rect 75460 3388 75740 3444
rect 75796 3388 76300 3444
rect 76356 3388 76366 3444
rect 92754 3388 92764 3444
rect 92820 3388 93660 3444
rect 93716 3388 93726 3444
rect 105532 3388 108444 3444
rect 108500 3388 108510 3444
rect 119746 3388 119756 3444
rect 119812 3388 121324 3444
rect 121380 3388 121390 3444
rect 139346 3388 139356 3444
rect 139412 3388 139692 3444
rect 139748 3388 142604 3444
rect 142660 3388 142940 3444
rect 142996 3388 153916 3444
rect 153972 3388 153982 3444
rect 105532 3332 105588 3388
rect 12674 3276 12684 3332
rect 12740 3276 13580 3332
rect 13636 3276 13646 3332
rect 34514 3276 34524 3332
rect 34580 3276 36204 3332
rect 36260 3276 36270 3332
rect 47954 3276 47964 3332
rect 48020 3276 48860 3332
rect 48916 3276 48926 3332
rect 59714 3276 59724 3332
rect 59780 3276 60620 3332
rect 60676 3276 60686 3332
rect 62066 3276 62076 3332
rect 62132 3276 63420 3332
rect 63476 3276 63486 3332
rect 76626 3276 76636 3332
rect 76692 3276 105532 3332
rect 105588 3276 105598 3332
rect 131394 3276 131404 3332
rect 131460 3276 133308 3332
rect 133364 3276 133374 3332
rect 139794 3276 139804 3332
rect 139860 3276 141708 3332
rect 141764 3276 141774 3332
rect 173954 3276 173964 3332
rect 174020 3276 174972 3332
rect 175028 3276 175038 3332
rect 45526 3108 45536 3164
rect 45592 3108 45640 3164
rect 45696 3108 45744 3164
rect 45800 3108 45810 3164
rect 89850 3108 89860 3164
rect 89916 3108 89964 3164
rect 90020 3108 90068 3164
rect 90124 3108 90134 3164
rect 134174 3108 134184 3164
rect 134240 3108 134288 3164
rect 134344 3108 134392 3164
rect 134448 3108 134458 3164
rect 178498 3108 178508 3164
rect 178564 3108 178612 3164
rect 178668 3108 178716 3164
rect 178772 3108 178782 3164
rect 14242 2940 14252 2996
rect 14308 2940 70588 2996
rect 70644 2940 70654 2996
rect 79314 2940 79324 2996
rect 79380 2940 151004 2996
rect 151060 2940 151070 2996
rect 28690 2828 28700 2884
rect 28756 2828 68908 2884
rect 68964 2828 68974 2884
rect 77634 2828 77644 2884
rect 77700 2828 127372 2884
rect 127428 2828 127438 2884
rect 36194 1708 36204 1764
rect 36260 1708 37100 1764
rect 37156 1708 37166 1764
<< via3 >>
rect 23374 16436 23430 16492
rect 23478 16436 23534 16492
rect 23582 16436 23638 16492
rect 67698 16436 67754 16492
rect 67802 16436 67858 16492
rect 67906 16436 67962 16492
rect 112022 16436 112078 16492
rect 112126 16436 112182 16492
rect 112230 16436 112286 16492
rect 156346 16436 156402 16492
rect 156450 16436 156506 16492
rect 156554 16436 156610 16492
rect 45536 15652 45592 15708
rect 45640 15652 45696 15708
rect 45744 15652 45800 15708
rect 89860 15652 89916 15708
rect 89964 15652 90020 15708
rect 90068 15652 90124 15708
rect 134184 15652 134240 15708
rect 134288 15652 134344 15708
rect 134392 15652 134448 15708
rect 178508 15652 178564 15708
rect 178612 15652 178668 15708
rect 178716 15652 178772 15708
rect 23374 14868 23430 14924
rect 23478 14868 23534 14924
rect 23582 14868 23638 14924
rect 67698 14868 67754 14924
rect 67802 14868 67858 14924
rect 67906 14868 67962 14924
rect 112022 14868 112078 14924
rect 112126 14868 112182 14924
rect 112230 14868 112286 14924
rect 156346 14868 156402 14924
rect 156450 14868 156506 14924
rect 156554 14868 156610 14924
rect 45536 14084 45592 14140
rect 45640 14084 45696 14140
rect 45744 14084 45800 14140
rect 89860 14084 89916 14140
rect 89964 14084 90020 14140
rect 90068 14084 90124 14140
rect 134184 14084 134240 14140
rect 134288 14084 134344 14140
rect 134392 14084 134448 14140
rect 178508 14084 178564 14140
rect 178612 14084 178668 14140
rect 178716 14084 178772 14140
rect 23374 13300 23430 13356
rect 23478 13300 23534 13356
rect 23582 13300 23638 13356
rect 67698 13300 67754 13356
rect 67802 13300 67858 13356
rect 67906 13300 67962 13356
rect 112022 13300 112078 13356
rect 112126 13300 112182 13356
rect 112230 13300 112286 13356
rect 156346 13300 156402 13356
rect 156450 13300 156506 13356
rect 156554 13300 156610 13356
rect 45536 12516 45592 12572
rect 45640 12516 45696 12572
rect 45744 12516 45800 12572
rect 89860 12516 89916 12572
rect 89964 12516 90020 12572
rect 90068 12516 90124 12572
rect 134184 12516 134240 12572
rect 134288 12516 134344 12572
rect 134392 12516 134448 12572
rect 178508 12516 178564 12572
rect 178612 12516 178668 12572
rect 178716 12516 178772 12572
rect 23374 11732 23430 11788
rect 23478 11732 23534 11788
rect 23582 11732 23638 11788
rect 67698 11732 67754 11788
rect 67802 11732 67858 11788
rect 67906 11732 67962 11788
rect 112022 11732 112078 11788
rect 112126 11732 112182 11788
rect 112230 11732 112286 11788
rect 156346 11732 156402 11788
rect 156450 11732 156506 11788
rect 156554 11732 156610 11788
rect 45536 10948 45592 11004
rect 45640 10948 45696 11004
rect 45744 10948 45800 11004
rect 89860 10948 89916 11004
rect 89964 10948 90020 11004
rect 90068 10948 90124 11004
rect 134184 10948 134240 11004
rect 134288 10948 134344 11004
rect 134392 10948 134448 11004
rect 178508 10948 178564 11004
rect 178612 10948 178668 11004
rect 178716 10948 178772 11004
rect 23374 10164 23430 10220
rect 23478 10164 23534 10220
rect 23582 10164 23638 10220
rect 67698 10164 67754 10220
rect 67802 10164 67858 10220
rect 67906 10164 67962 10220
rect 112022 10164 112078 10220
rect 112126 10164 112182 10220
rect 112230 10164 112286 10220
rect 156346 10164 156402 10220
rect 156450 10164 156506 10220
rect 156554 10164 156610 10220
rect 45536 9380 45592 9436
rect 45640 9380 45696 9436
rect 45744 9380 45800 9436
rect 89860 9380 89916 9436
rect 89964 9380 90020 9436
rect 90068 9380 90124 9436
rect 134184 9380 134240 9436
rect 134288 9380 134344 9436
rect 134392 9380 134448 9436
rect 178508 9380 178564 9436
rect 178612 9380 178668 9436
rect 178716 9380 178772 9436
rect 23374 8596 23430 8652
rect 23478 8596 23534 8652
rect 23582 8596 23638 8652
rect 67698 8596 67754 8652
rect 67802 8596 67858 8652
rect 67906 8596 67962 8652
rect 112022 8596 112078 8652
rect 112126 8596 112182 8652
rect 112230 8596 112286 8652
rect 156346 8596 156402 8652
rect 156450 8596 156506 8652
rect 156554 8596 156610 8652
rect 45536 7812 45592 7868
rect 45640 7812 45696 7868
rect 45744 7812 45800 7868
rect 89860 7812 89916 7868
rect 89964 7812 90020 7868
rect 90068 7812 90124 7868
rect 134184 7812 134240 7868
rect 134288 7812 134344 7868
rect 134392 7812 134448 7868
rect 178508 7812 178564 7868
rect 178612 7812 178668 7868
rect 178716 7812 178772 7868
rect 23374 7028 23430 7084
rect 23478 7028 23534 7084
rect 23582 7028 23638 7084
rect 67698 7028 67754 7084
rect 67802 7028 67858 7084
rect 67906 7028 67962 7084
rect 112022 7028 112078 7084
rect 112126 7028 112182 7084
rect 112230 7028 112286 7084
rect 156346 7028 156402 7084
rect 156450 7028 156506 7084
rect 156554 7028 156610 7084
rect 45536 6244 45592 6300
rect 45640 6244 45696 6300
rect 45744 6244 45800 6300
rect 89860 6244 89916 6300
rect 89964 6244 90020 6300
rect 90068 6244 90124 6300
rect 134184 6244 134240 6300
rect 134288 6244 134344 6300
rect 134392 6244 134448 6300
rect 178508 6244 178564 6300
rect 178612 6244 178668 6300
rect 178716 6244 178772 6300
rect 23374 5460 23430 5516
rect 23478 5460 23534 5516
rect 23582 5460 23638 5516
rect 67698 5460 67754 5516
rect 67802 5460 67858 5516
rect 67906 5460 67962 5516
rect 112022 5460 112078 5516
rect 112126 5460 112182 5516
rect 112230 5460 112286 5516
rect 156346 5460 156402 5516
rect 156450 5460 156506 5516
rect 156554 5460 156610 5516
rect 45536 4676 45592 4732
rect 45640 4676 45696 4732
rect 45744 4676 45800 4732
rect 89860 4676 89916 4732
rect 89964 4676 90020 4732
rect 90068 4676 90124 4732
rect 134184 4676 134240 4732
rect 134288 4676 134344 4732
rect 134392 4676 134448 4732
rect 178508 4676 178564 4732
rect 178612 4676 178668 4732
rect 178716 4676 178772 4732
rect 23374 3892 23430 3948
rect 23478 3892 23534 3948
rect 23582 3892 23638 3948
rect 67698 3892 67754 3948
rect 67802 3892 67858 3948
rect 67906 3892 67962 3948
rect 112022 3892 112078 3948
rect 112126 3892 112182 3948
rect 112230 3892 112286 3948
rect 156346 3892 156402 3948
rect 156450 3892 156506 3948
rect 156554 3892 156610 3948
rect 45536 3108 45592 3164
rect 45640 3108 45696 3164
rect 45744 3108 45800 3164
rect 89860 3108 89916 3164
rect 89964 3108 90020 3164
rect 90068 3108 90124 3164
rect 134184 3108 134240 3164
rect 134288 3108 134344 3164
rect 134392 3108 134448 3164
rect 178508 3108 178564 3164
rect 178612 3108 178668 3164
rect 178716 3108 178772 3164
<< metal4 >>
rect 23346 16492 23666 16524
rect 23346 16436 23374 16492
rect 23430 16436 23478 16492
rect 23534 16436 23582 16492
rect 23638 16436 23666 16492
rect 23346 14924 23666 16436
rect 23346 14868 23374 14924
rect 23430 14868 23478 14924
rect 23534 14868 23582 14924
rect 23638 14868 23666 14924
rect 23346 13356 23666 14868
rect 23346 13300 23374 13356
rect 23430 13300 23478 13356
rect 23534 13300 23582 13356
rect 23638 13300 23666 13356
rect 23346 11788 23666 13300
rect 23346 11732 23374 11788
rect 23430 11732 23478 11788
rect 23534 11732 23582 11788
rect 23638 11732 23666 11788
rect 23346 10220 23666 11732
rect 23346 10164 23374 10220
rect 23430 10164 23478 10220
rect 23534 10164 23582 10220
rect 23638 10164 23666 10220
rect 23346 8652 23666 10164
rect 23346 8596 23374 8652
rect 23430 8596 23478 8652
rect 23534 8596 23582 8652
rect 23638 8596 23666 8652
rect 23346 7084 23666 8596
rect 23346 7028 23374 7084
rect 23430 7028 23478 7084
rect 23534 7028 23582 7084
rect 23638 7028 23666 7084
rect 23346 5516 23666 7028
rect 23346 5460 23374 5516
rect 23430 5460 23478 5516
rect 23534 5460 23582 5516
rect 23638 5460 23666 5516
rect 23346 3948 23666 5460
rect 23346 3892 23374 3948
rect 23430 3892 23478 3948
rect 23534 3892 23582 3948
rect 23638 3892 23666 3948
rect 23346 3076 23666 3892
rect 45508 15708 45828 16524
rect 45508 15652 45536 15708
rect 45592 15652 45640 15708
rect 45696 15652 45744 15708
rect 45800 15652 45828 15708
rect 45508 14140 45828 15652
rect 45508 14084 45536 14140
rect 45592 14084 45640 14140
rect 45696 14084 45744 14140
rect 45800 14084 45828 14140
rect 45508 12572 45828 14084
rect 45508 12516 45536 12572
rect 45592 12516 45640 12572
rect 45696 12516 45744 12572
rect 45800 12516 45828 12572
rect 45508 11004 45828 12516
rect 45508 10948 45536 11004
rect 45592 10948 45640 11004
rect 45696 10948 45744 11004
rect 45800 10948 45828 11004
rect 45508 9436 45828 10948
rect 45508 9380 45536 9436
rect 45592 9380 45640 9436
rect 45696 9380 45744 9436
rect 45800 9380 45828 9436
rect 45508 7868 45828 9380
rect 45508 7812 45536 7868
rect 45592 7812 45640 7868
rect 45696 7812 45744 7868
rect 45800 7812 45828 7868
rect 45508 6300 45828 7812
rect 45508 6244 45536 6300
rect 45592 6244 45640 6300
rect 45696 6244 45744 6300
rect 45800 6244 45828 6300
rect 45508 4732 45828 6244
rect 45508 4676 45536 4732
rect 45592 4676 45640 4732
rect 45696 4676 45744 4732
rect 45800 4676 45828 4732
rect 45508 3164 45828 4676
rect 45508 3108 45536 3164
rect 45592 3108 45640 3164
rect 45696 3108 45744 3164
rect 45800 3108 45828 3164
rect 45508 3076 45828 3108
rect 67670 16492 67990 16524
rect 67670 16436 67698 16492
rect 67754 16436 67802 16492
rect 67858 16436 67906 16492
rect 67962 16436 67990 16492
rect 67670 14924 67990 16436
rect 67670 14868 67698 14924
rect 67754 14868 67802 14924
rect 67858 14868 67906 14924
rect 67962 14868 67990 14924
rect 67670 13356 67990 14868
rect 67670 13300 67698 13356
rect 67754 13300 67802 13356
rect 67858 13300 67906 13356
rect 67962 13300 67990 13356
rect 67670 11788 67990 13300
rect 67670 11732 67698 11788
rect 67754 11732 67802 11788
rect 67858 11732 67906 11788
rect 67962 11732 67990 11788
rect 67670 10220 67990 11732
rect 67670 10164 67698 10220
rect 67754 10164 67802 10220
rect 67858 10164 67906 10220
rect 67962 10164 67990 10220
rect 67670 8652 67990 10164
rect 67670 8596 67698 8652
rect 67754 8596 67802 8652
rect 67858 8596 67906 8652
rect 67962 8596 67990 8652
rect 67670 7084 67990 8596
rect 67670 7028 67698 7084
rect 67754 7028 67802 7084
rect 67858 7028 67906 7084
rect 67962 7028 67990 7084
rect 67670 5516 67990 7028
rect 67670 5460 67698 5516
rect 67754 5460 67802 5516
rect 67858 5460 67906 5516
rect 67962 5460 67990 5516
rect 67670 3948 67990 5460
rect 67670 3892 67698 3948
rect 67754 3892 67802 3948
rect 67858 3892 67906 3948
rect 67962 3892 67990 3948
rect 67670 3076 67990 3892
rect 89832 15708 90152 16524
rect 89832 15652 89860 15708
rect 89916 15652 89964 15708
rect 90020 15652 90068 15708
rect 90124 15652 90152 15708
rect 89832 14140 90152 15652
rect 89832 14084 89860 14140
rect 89916 14084 89964 14140
rect 90020 14084 90068 14140
rect 90124 14084 90152 14140
rect 89832 12572 90152 14084
rect 89832 12516 89860 12572
rect 89916 12516 89964 12572
rect 90020 12516 90068 12572
rect 90124 12516 90152 12572
rect 89832 11004 90152 12516
rect 89832 10948 89860 11004
rect 89916 10948 89964 11004
rect 90020 10948 90068 11004
rect 90124 10948 90152 11004
rect 89832 9436 90152 10948
rect 89832 9380 89860 9436
rect 89916 9380 89964 9436
rect 90020 9380 90068 9436
rect 90124 9380 90152 9436
rect 89832 7868 90152 9380
rect 89832 7812 89860 7868
rect 89916 7812 89964 7868
rect 90020 7812 90068 7868
rect 90124 7812 90152 7868
rect 89832 6300 90152 7812
rect 89832 6244 89860 6300
rect 89916 6244 89964 6300
rect 90020 6244 90068 6300
rect 90124 6244 90152 6300
rect 89832 4732 90152 6244
rect 89832 4676 89860 4732
rect 89916 4676 89964 4732
rect 90020 4676 90068 4732
rect 90124 4676 90152 4732
rect 89832 3164 90152 4676
rect 89832 3108 89860 3164
rect 89916 3108 89964 3164
rect 90020 3108 90068 3164
rect 90124 3108 90152 3164
rect 89832 3076 90152 3108
rect 111994 16492 112314 16524
rect 111994 16436 112022 16492
rect 112078 16436 112126 16492
rect 112182 16436 112230 16492
rect 112286 16436 112314 16492
rect 111994 14924 112314 16436
rect 111994 14868 112022 14924
rect 112078 14868 112126 14924
rect 112182 14868 112230 14924
rect 112286 14868 112314 14924
rect 111994 13356 112314 14868
rect 111994 13300 112022 13356
rect 112078 13300 112126 13356
rect 112182 13300 112230 13356
rect 112286 13300 112314 13356
rect 111994 11788 112314 13300
rect 111994 11732 112022 11788
rect 112078 11732 112126 11788
rect 112182 11732 112230 11788
rect 112286 11732 112314 11788
rect 111994 10220 112314 11732
rect 111994 10164 112022 10220
rect 112078 10164 112126 10220
rect 112182 10164 112230 10220
rect 112286 10164 112314 10220
rect 111994 8652 112314 10164
rect 111994 8596 112022 8652
rect 112078 8596 112126 8652
rect 112182 8596 112230 8652
rect 112286 8596 112314 8652
rect 111994 7084 112314 8596
rect 111994 7028 112022 7084
rect 112078 7028 112126 7084
rect 112182 7028 112230 7084
rect 112286 7028 112314 7084
rect 111994 5516 112314 7028
rect 111994 5460 112022 5516
rect 112078 5460 112126 5516
rect 112182 5460 112230 5516
rect 112286 5460 112314 5516
rect 111994 3948 112314 5460
rect 111994 3892 112022 3948
rect 112078 3892 112126 3948
rect 112182 3892 112230 3948
rect 112286 3892 112314 3948
rect 111994 3076 112314 3892
rect 134156 15708 134476 16524
rect 134156 15652 134184 15708
rect 134240 15652 134288 15708
rect 134344 15652 134392 15708
rect 134448 15652 134476 15708
rect 134156 14140 134476 15652
rect 134156 14084 134184 14140
rect 134240 14084 134288 14140
rect 134344 14084 134392 14140
rect 134448 14084 134476 14140
rect 134156 12572 134476 14084
rect 134156 12516 134184 12572
rect 134240 12516 134288 12572
rect 134344 12516 134392 12572
rect 134448 12516 134476 12572
rect 134156 11004 134476 12516
rect 134156 10948 134184 11004
rect 134240 10948 134288 11004
rect 134344 10948 134392 11004
rect 134448 10948 134476 11004
rect 134156 9436 134476 10948
rect 134156 9380 134184 9436
rect 134240 9380 134288 9436
rect 134344 9380 134392 9436
rect 134448 9380 134476 9436
rect 134156 7868 134476 9380
rect 134156 7812 134184 7868
rect 134240 7812 134288 7868
rect 134344 7812 134392 7868
rect 134448 7812 134476 7868
rect 134156 6300 134476 7812
rect 134156 6244 134184 6300
rect 134240 6244 134288 6300
rect 134344 6244 134392 6300
rect 134448 6244 134476 6300
rect 134156 4732 134476 6244
rect 134156 4676 134184 4732
rect 134240 4676 134288 4732
rect 134344 4676 134392 4732
rect 134448 4676 134476 4732
rect 134156 3164 134476 4676
rect 134156 3108 134184 3164
rect 134240 3108 134288 3164
rect 134344 3108 134392 3164
rect 134448 3108 134476 3164
rect 134156 3076 134476 3108
rect 156318 16492 156638 16524
rect 156318 16436 156346 16492
rect 156402 16436 156450 16492
rect 156506 16436 156554 16492
rect 156610 16436 156638 16492
rect 156318 14924 156638 16436
rect 156318 14868 156346 14924
rect 156402 14868 156450 14924
rect 156506 14868 156554 14924
rect 156610 14868 156638 14924
rect 156318 13356 156638 14868
rect 156318 13300 156346 13356
rect 156402 13300 156450 13356
rect 156506 13300 156554 13356
rect 156610 13300 156638 13356
rect 156318 11788 156638 13300
rect 156318 11732 156346 11788
rect 156402 11732 156450 11788
rect 156506 11732 156554 11788
rect 156610 11732 156638 11788
rect 156318 10220 156638 11732
rect 156318 10164 156346 10220
rect 156402 10164 156450 10220
rect 156506 10164 156554 10220
rect 156610 10164 156638 10220
rect 156318 8652 156638 10164
rect 156318 8596 156346 8652
rect 156402 8596 156450 8652
rect 156506 8596 156554 8652
rect 156610 8596 156638 8652
rect 156318 7084 156638 8596
rect 156318 7028 156346 7084
rect 156402 7028 156450 7084
rect 156506 7028 156554 7084
rect 156610 7028 156638 7084
rect 156318 5516 156638 7028
rect 156318 5460 156346 5516
rect 156402 5460 156450 5516
rect 156506 5460 156554 5516
rect 156610 5460 156638 5516
rect 156318 3948 156638 5460
rect 156318 3892 156346 3948
rect 156402 3892 156450 3948
rect 156506 3892 156554 3948
rect 156610 3892 156638 3948
rect 156318 3076 156638 3892
rect 178480 15708 178800 16524
rect 178480 15652 178508 15708
rect 178564 15652 178612 15708
rect 178668 15652 178716 15708
rect 178772 15652 178800 15708
rect 178480 14140 178800 15652
rect 178480 14084 178508 14140
rect 178564 14084 178612 14140
rect 178668 14084 178716 14140
rect 178772 14084 178800 14140
rect 178480 12572 178800 14084
rect 178480 12516 178508 12572
rect 178564 12516 178612 12572
rect 178668 12516 178716 12572
rect 178772 12516 178800 12572
rect 178480 11004 178800 12516
rect 178480 10948 178508 11004
rect 178564 10948 178612 11004
rect 178668 10948 178716 11004
rect 178772 10948 178800 11004
rect 178480 9436 178800 10948
rect 178480 9380 178508 9436
rect 178564 9380 178612 9436
rect 178668 9380 178716 9436
rect 178772 9380 178800 9436
rect 178480 7868 178800 9380
rect 178480 7812 178508 7868
rect 178564 7812 178612 7868
rect 178668 7812 178716 7868
rect 178772 7812 178800 7868
rect 178480 6300 178800 7812
rect 178480 6244 178508 6300
rect 178564 6244 178612 6300
rect 178668 6244 178716 6300
rect 178772 6244 178800 6300
rect 178480 4732 178800 6244
rect 178480 4676 178508 4732
rect 178564 4676 178612 4732
rect 178668 4676 178716 4732
rect 178772 4676 178800 4732
rect 178480 3164 178800 4676
rect 178480 3108 178508 3164
rect 178564 3108 178612 3164
rect 178668 3108 178716 3164
rect 178772 3108 178800 3164
rect 178480 3076 178800 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__A1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 79296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__CLK
timestamp 1667941163
transform 1 0 55776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__D
timestamp 1667941163
transform 1 0 54320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__CLK
timestamp 1667941163
transform -1 0 29344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__D
timestamp 1667941163
transform -1 0 28784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__CLK
timestamp 1667941163
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__D
timestamp 1667941163
transform -1 0 14336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__CLK
timestamp 1667941163
transform -1 0 75936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__CLK
timestamp 1667941163
transform 1 0 91392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__D
timestamp 1667941163
transform -1 0 90720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__CLK
timestamp 1667941163
transform -1 0 106064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__D
timestamp 1667941163
transform -1 0 105616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__CLK
timestamp 1667941163
transform 1 0 126896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__D
timestamp 1667941163
transform -1 0 127568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__CLK
timestamp 1667941163
transform 1 0 150416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__D
timestamp 1667941163
transform -1 0 151088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__I
timestamp 1667941163
transform 1 0 121520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I
timestamp 1667941163
transform 1 0 121072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout11_I
timestamp 1667941163
transform 1 0 61936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout12_I
timestamp 1667941163
transform 1 0 60704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout13_I
timestamp 1667941163
transform 1 0 69216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1667941163
transform -1 0 63840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1667941163
transform 1 0 67648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1667941163
transform 1 0 70672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1667941163
transform -1 0 70448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1667941163
transform -1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1667941163
transform -1 0 73584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1667941163
transform -1 0 75824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1667941163
transform -1 0 77168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1667941163
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1667941163
transform -1 0 80304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[0\].pun_I
timestamp 1667941163
transform 1 0 69216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[1\].pun_I
timestamp 1667941163
transform 1 0 67648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[2\].pun_I
timestamp 1667941163
transform 1 0 68768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[3\].pun_I
timestamp 1667941163
transform 1 0 69776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[4\].pun_I
timestamp 1667941163
transform -1 0 66976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[5\].pun_I
timestamp 1667941163
transform 1 0 64512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[6\].pun_I
timestamp 1667941163
transform 1 0 64064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[6\].pup_I
timestamp 1667941163
transform 1 0 61152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[7\].pun_I
timestamp 1667941163
transform 1 0 65632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[7\].pup_I
timestamp 1667941163
transform 1 0 60032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[8\].pun_I
timestamp 1667941163
transform 1 0 63728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[9\].pun_I
timestamp 1667941163
transform -1 0 62720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[9\].pup_I
timestamp 1667941163
transform 1 0 60592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[10\].pun_I
timestamp 1667941163
transform -1 0 68544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[11\].pun_I
timestamp 1667941163
transform -1 0 65520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[12\].pun_I
timestamp 1667941163
transform 1 0 63280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[13\].pun_I
timestamp 1667941163
transform 1 0 62944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[14\].pun_I
timestamp 1667941163
transform -1 0 67424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[15\].pun_I
timestamp 1667941163
transform 1 0 62832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[16\].pun_I
timestamp 1667941163
transform 1 0 68096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[17\].pun_I
timestamp 1667941163
transform 1 0 68544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_PU\[18\].pun_I
timestamp 1667941163
transform 1 0 62160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[0\].ntrimn_EN
timestamp 1667941163
transform 1 0 105392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[0\].ntrimp_EN
timestamp 1667941163
transform 1 0 105168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[0\].ptrimn_I
timestamp 1667941163
transform 1 0 51520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[0\].ptrimp_I
timestamp 1667941163
transform 1 0 50400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[1\].ntrimn_EN
timestamp 1667941163
transform 1 0 118272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[1\].ntrimp_EN
timestamp 1667941163
transform 1 0 118160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[1\].ptrimn_I
timestamp 1667941163
transform 1 0 35504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[1\].ptrimp_I
timestamp 1667941163
transform 1 0 36400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[2\].ptrimn_EN
timestamp 1667941163
transform -1 0 30912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[2\].ptrimn_I
timestamp 1667941163
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[2\].ptrimp_EN
timestamp 1667941163
transform -1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[2\].ptrimp_I
timestamp 1667941163
transform 1 0 36848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ntrimn_EN
timestamp 1667941163
transform -1 0 142688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ntrimp_EN
timestamp 1667941163
transform -1 0 143024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ptrimn_EN
timestamp 1667941163
transform -1 0 83776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ptrimn_I
timestamp 1667941163
transform 1 0 84336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ptrimp_EN
timestamp 1667941163
transform -1 0 84672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_inj.gen_TRIM\[3\].ptrimp_I
timestamp 1667941163
transform 1 0 84000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 6384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 6832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51
timestamp 1667941163
transform 1 0 7056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56
timestamp 1667941163
transform 1 0 7616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64
timestamp 1667941163
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1667941163
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1667941163
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102
timestamp 1667941163
transform 1 0 12768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1667941163
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112
timestamp 1667941163
transform 1 0 13888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116
timestamp 1667941163
transform 1 0 14336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120
timestamp 1667941163
transform 1 0 14784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_126
timestamp 1667941163
transform 1 0 15456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134
timestamp 1667941163
transform 1 0 16352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 16800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1667941163
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_147
timestamp 1667941163
transform 1 0 17808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155
timestamp 1667941163
transform 1 0 18704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159
timestamp 1667941163
transform 1 0 19152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_161
timestamp 1667941163
transform 1 0 19376 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_166
timestamp 1667941163
transform 1 0 19936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_182
timestamp 1667941163
transform 1 0 21728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190
timestamp 1667941163
transform 1 0 22624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_196
timestamp 1667941163
transform 1 0 23296 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_204
timestamp 1667941163
transform 1 0 24192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1667941163
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1667941163
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_242
timestamp 1667941163
transform 1 0 28448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1667941163
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1667941163
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 29344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_256
timestamp 1667941163
transform 1 0 30016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_264
timestamp 1667941163
transform 1 0 30912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_266
timestamp 1667941163
transform 1 0 31136 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_271
timestamp 1667941163
transform 1 0 31696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_275
timestamp 1667941163
transform 1 0 32144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1667941163
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_287
timestamp 1667941163
transform 1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_308
timestamp 1667941163
transform 1 0 35840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1667941163
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1667941163
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_322
timestamp 1667941163
transform 1 0 37408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_326
timestamp 1667941163
transform 1 0 37856 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_331
timestamp 1667941163
transform 1 0 38416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_339
timestamp 1667941163
transform 1 0 39312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_341
timestamp 1667941163
transform 1 0 39536 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_346
timestamp 1667941163
transform 1 0 40096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1667941163
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_356
timestamp 1667941163
transform 1 0 41216 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_361
timestamp 1667941163
transform 1 0 41776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_369
timestamp 1667941163
transform 1 0 42672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_371
timestamp 1667941163
transform 1 0 42896 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_376
timestamp 1667941163
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1667941163
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1667941163
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_392
timestamp 1667941163
transform 1 0 45248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_400
timestamp 1667941163
transform 1 0 46144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_406
timestamp 1667941163
transform 1 0 46816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_414
timestamp 1667941163
transform 1 0 47712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1667941163
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1667941163
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_427
timestamp 1667941163
transform 1 0 49168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_431
timestamp 1667941163
transform 1 0 49616 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_436
timestamp 1667941163
transform 1 0 50176 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_444
timestamp 1667941163
transform 1 0 51072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_446
timestamp 1667941163
transform 1 0 51296 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_451
timestamp 1667941163
transform 1 0 51856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1667941163
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_487
timestamp 1667941163
transform 1 0 55888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1667941163
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1667941163
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_497
timestamp 1667941163
transform 1 0 57008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_499
timestamp 1667941163
transform 1 0 57232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_506
timestamp 1667941163
transform 1 0 58016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_514
timestamp 1667941163
transform 1 0 58912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_522
timestamp 1667941163
transform 1 0 59808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1667941163
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1667941163
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_532
timestamp 1667941163
transform 1 0 60928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_534
timestamp 1667941163
transform 1 0 61152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_539
timestamp 1667941163
transform 1 0 61712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_545
timestamp 1667941163
transform 1 0 62384 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_551
timestamp 1667941163
transform 1 0 63056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1667941163
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_562
timestamp 1667941163
transform 1 0 64288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_570
timestamp 1667941163
transform 1 0 65184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_578
timestamp 1667941163
transform 1 0 66080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_588
timestamp 1667941163
transform 1 0 67200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1667941163
transform 1 0 67872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1667941163
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_600
timestamp 1667941163
transform 1 0 68544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_608
timestamp 1667941163
transform 1 0 69440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_614
timestamp 1667941163
transform 1 0 70112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_616
timestamp 1667941163
transform 1 0 70336 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_623
timestamp 1667941163
transform 1 0 71120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1667941163
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_632
timestamp 1667941163
transform 1 0 72128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_634
timestamp 1667941163
transform 1 0 72352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1667941163
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1667941163
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_674
timestamp 1667941163
transform 1 0 76832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_676
timestamp 1667941163
transform 1 0 77056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_683
timestamp 1667941163
transform 1 0 77840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_689
timestamp 1667941163
transform 1 0 78512 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_691
timestamp 1667941163
transform 1 0 78736 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_698
timestamp 1667941163
transform 1 0 79520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1667941163
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_705
timestamp 1667941163
transform 1 0 80304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_715
timestamp 1667941163
transform 1 0 81424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_721
timestamp 1667941163
transform 1 0 82096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_725
timestamp 1667941163
transform 1 0 82544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_731
timestamp 1667941163
transform 1 0 83216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_737
timestamp 1667941163
transform 1 0 83888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_743
timestamp 1667941163
transform 1 0 84560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_762
timestamp 1667941163
transform 1 0 86688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_768
timestamp 1667941163
transform 1 0 87360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1667941163
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_777
timestamp 1667941163
transform 1 0 88368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_785
timestamp 1667941163
transform 1 0 89264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_791
timestamp 1667941163
transform 1 0 89936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_795
timestamp 1667941163
transform 1 0 90384 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_798
timestamp 1667941163
transform 1 0 90720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_804
timestamp 1667941163
transform 1 0 91392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1667941163
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_837
timestamp 1667941163
transform 1 0 95088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1667941163
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_842
timestamp 1667941163
transform 1 0 95648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_846
timestamp 1667941163
transform 1 0 96096 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_848
timestamp 1667941163
transform 1 0 96320 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_853
timestamp 1667941163
transform 1 0 96880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_859
timestamp 1667941163
transform 1 0 97552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_861
timestamp 1667941163
transform 1 0 97776 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_866
timestamp 1667941163
transform 1 0 98336 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1667941163
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1667941163
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_882
timestamp 1667941163
transform 1 0 100128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_890
timestamp 1667941163
transform 1 0 101024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_896
timestamp 1667941163
transform 1 0 101696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_904
timestamp 1667941163
transform 1 0 102592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_908
timestamp 1667941163
transform 1 0 103040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_912
timestamp 1667941163
transform 1 0 103488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_917
timestamp 1667941163
transform 1 0 104048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_921
timestamp 1667941163
transform 1 0 104496 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_926
timestamp 1667941163
transform 1 0 105056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_928
timestamp 1667941163
transform 1 0 105280 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_931
timestamp 1667941163
transform 1 0 105616 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_935
timestamp 1667941163
transform 1 0 106064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_941
timestamp 1667941163
transform 1 0 106736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_947
timestamp 1667941163
transform 1 0 107408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_977
timestamp 1667941163
transform 1 0 110768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1667941163
transform 1 0 110992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1667941163
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_987
timestamp 1667941163
transform 1 0 111888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_995
timestamp 1667941163
transform 1 0 112784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1001
timestamp 1667941163
transform 1 0 113456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1009
timestamp 1667941163
transform 1 0 114352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1013
timestamp 1667941163
transform 1 0 114800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1667941163
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1022
timestamp 1667941163
transform 1 0 115808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1026
timestamp 1667941163
transform 1 0 116256 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1031
timestamp 1667941163
transform 1 0 116816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1039
timestamp 1667941163
transform 1 0 117712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1041
timestamp 1667941163
transform 1 0 117936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1046
timestamp 1667941163
transform 1 0 118496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1052
timestamp 1667941163
transform 1 0 119168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1059
timestamp 1667941163
transform 1 0 119952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1067
timestamp 1667941163
transform 1 0 120848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1071
timestamp 1667941163
transform 1 0 121296 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1075
timestamp 1667941163
transform 1 0 121744 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1083
timestamp 1667941163
transform 1 0 122640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1667941163
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1092
timestamp 1667941163
transform 1 0 123648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1100
timestamp 1667941163
transform 1 0 124544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1106
timestamp 1667941163
transform 1 0 125216 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1114
timestamp 1667941163
transform 1 0 126112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1119
timestamp 1667941163
transform 1 0 126672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1122
timestamp 1667941163
transform 1 0 127008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1124
timestamp 1667941163
transform 1 0 127232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1667941163
transform 1 0 130592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1667941163
transform 1 0 130928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1175
timestamp 1667941163
transform 1 0 132944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1181
timestamp 1667941163
transform 1 0 133616 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1187
timestamp 1667941163
transform 1 0 134288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1189
timestamp 1667941163
transform 1 0 134512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1192
timestamp 1667941163
transform 1 0 134848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1197
timestamp 1667941163
transform 1 0 135408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1205
timestamp 1667941163
transform 1 0 136304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1211
timestamp 1667941163
transform 1 0 136976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1219
timestamp 1667941163
transform 1 0 137872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1224
timestamp 1667941163
transform 1 0 138432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1227
timestamp 1667941163
transform 1 0 138768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1231
timestamp 1667941163
transform 1 0 139216 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1250
timestamp 1667941163
transform 1 0 141344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1256
timestamp 1667941163
transform 1 0 142016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1262
timestamp 1667941163
transform 1 0 142688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1265
timestamp 1667941163
transform 1 0 143024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1271
timestamp 1667941163
transform 1 0 143696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1279
timestamp 1667941163
transform 1 0 144592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1281
timestamp 1667941163
transform 1 0 144816 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1286
timestamp 1667941163
transform 1 0 145376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1294
timestamp 1667941163
transform 1 0 146272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1297
timestamp 1667941163
transform 1 0 146608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1302
timestamp 1667941163
transform 1 0 147168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1310
timestamp 1667941163
transform 1 0 148064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1316
timestamp 1667941163
transform 1 0 148736 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1324
timestamp 1667941163
transform 1 0 149632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1329
timestamp 1667941163
transform 1 0 150192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1332
timestamp 1667941163
transform 1 0 150528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1334
timestamp 1667941163
transform 1 0 150752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1364
timestamp 1667941163
transform 1 0 154112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1367
timestamp 1667941163
transform 1 0 154448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1371
timestamp 1667941163
transform 1 0 154896 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1376
timestamp 1667941163
transform 1 0 155456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1384
timestamp 1667941163
transform 1 0 156352 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1386
timestamp 1667941163
transform 1 0 156576 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1391
timestamp 1667941163
transform 1 0 157136 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1399
timestamp 1667941163
transform 1 0 158032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1402
timestamp 1667941163
transform 1 0 158368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1407
timestamp 1667941163
transform 1 0 158928 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1415
timestamp 1667941163
transform 1 0 159824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1421
timestamp 1667941163
transform 1 0 160496 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1429
timestamp 1667941163
transform 1 0 161392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1433
timestamp 1667941163
transform 1 0 161840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1437
timestamp 1667941163
transform 1 0 162288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1442
timestamp 1667941163
transform 1 0 162848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1446
timestamp 1667941163
transform 1 0 163296 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1451
timestamp 1667941163
transform 1 0 163856 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1459
timestamp 1667941163
transform 1 0 164752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1461
timestamp 1667941163
transform 1 0 164976 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1466
timestamp 1667941163
transform 1 0 165536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1472
timestamp 1667941163
transform 1 0 166208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1476
timestamp 1667941163
transform 1 0 166656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1481
timestamp 1667941163
transform 1 0 167216 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1489
timestamp 1667941163
transform 1 0 168112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1491
timestamp 1667941163
transform 1 0 168336 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1496
timestamp 1667941163
transform 1 0 168896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1504
timestamp 1667941163
transform 1 0 169792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1507
timestamp 1667941163
transform 1 0 170128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1512
timestamp 1667941163
transform 1 0 170688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1520
timestamp 1667941163
transform 1 0 171584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1526
timestamp 1667941163
transform 1 0 172256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1530
timestamp 1667941163
transform 1 0 172704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1536
timestamp 1667941163
transform 1 0 173376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1542
timestamp 1667941163
transform 1 0 174048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1547
timestamp 1667941163
transform 1 0 174608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1553 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 175280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1569
timestamp 1667941163
transform 1 0 177072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1573
timestamp 1667941163
transform 1 0 177520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1577
timestamp 1667941163
transform 1 0 177968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_73
timestamp 1667941163
transform 1 0 9520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_81
timestamp 1667941163
transform 1 0 10416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_86
timestamp 1667941163
transform 1 0 10976 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_102
timestamp 1667941163
transform 1 0 12768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_106
timestamp 1667941163
transform 1 0 13216 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_138
timestamp 1667941163
transform 1 0 16800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1667941163
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1667941163
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_215
timestamp 1667941163
transform 1 0 25424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_219
timestamp 1667941163
transform 1 0 25872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_221
timestamp 1667941163
transform 1 0 26096 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_226
timestamp 1667941163
transform 1 0 26656 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_234
timestamp 1667941163
transform 1 0 27552 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_236
timestamp 1667941163
transform 1 0 27776 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_241
timestamp 1667941163
transform 1 0 28336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_245
timestamp 1667941163
transform 1 0 28784 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_261
timestamp 1667941163
transform 1 0 30576 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_264
timestamp 1667941163
transform 1 0 30912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1667941163
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1667941163
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_289
timestamp 1667941163
transform 1 0 33712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_293
timestamp 1667941163
transform 1 0 34160 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_311
timestamp 1667941163
transform 1 0 36176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_315
timestamp 1667941163
transform 1 0 36624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_319
timestamp 1667941163
transform 1 0 37072 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_351
timestamp 1667941163
transform 1 0 40656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1667941163
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1667941163
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1667941163
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1667941163
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_446
timestamp 1667941163
transform 1 0 51296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_450
timestamp 1667941163
transform 1 0 51744 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_458
timestamp 1667941163
transform 1 0 52640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_466
timestamp 1667941163
transform 1 0 53536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_470
timestamp 1667941163
transform 1 0 53984 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_472
timestamp 1667941163
transform 1 0 54208 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_475
timestamp 1667941163
transform 1 0 54544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_481
timestamp 1667941163
transform 1 0 55216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_485
timestamp 1667941163
transform 1 0 55664 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_488
timestamp 1667941163
transform 1 0 56000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1667941163
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_499
timestamp 1667941163
transform 1 0 57232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_505
timestamp 1667941163
transform 1 0 57904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_513
timestamp 1667941163
transform 1 0 58800 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_541
timestamp 1667941163
transform 1 0 61936 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_545
timestamp 1667941163
transform 1 0 62384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_551
timestamp 1667941163
transform 1 0 63056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_559
timestamp 1667941163
transform 1 0 63952 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1667941163
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1667941163
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_575
timestamp 1667941163
transform 1 0 65744 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_603
timestamp 1667941163
transform 1 0 68880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_611
timestamp 1667941163
transform 1 0 69776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_619
timestamp 1667941163
transform 1 0 70672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_621
timestamp 1667941163
transform 1 0 70896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_626
timestamp 1667941163
transform 1 0 71456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_630
timestamp 1667941163
transform 1 0 71904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1667941163
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_641
timestamp 1667941163
transform 1 0 73136 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_645
timestamp 1667941163
transform 1 0 73584 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_653
timestamp 1667941163
transform 1 0 74480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_659
timestamp 1667941163
transform 1 0 75152 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_665
timestamp 1667941163
transform 1 0 75824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_671
timestamp 1667941163
transform 1 0 76496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_677
timestamp 1667941163
transform 1 0 77168 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_685
timestamp 1667941163
transform 1 0 78064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_687
timestamp 1667941163
transform 1 0 78288 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_690
timestamp 1667941163
transform 1 0 78624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_696
timestamp 1667941163
transform 1 0 79296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_702
timestamp 1667941163
transform 1 0 79968 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_712
timestamp 1667941163
transform 1 0 81088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_728
timestamp 1667941163
transform 1 0 82880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_732
timestamp 1667941163
transform 1 0 83328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_736
timestamp 1667941163
transform 1 0 83776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_740
timestamp 1667941163
transform 1 0 84224 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_744
timestamp 1667941163
transform 1 0 84672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_763
timestamp 1667941163
transform 1 0 86800 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_779
timestamp 1667941163
transform 1 0 88592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_783
timestamp 1667941163
transform 1 0 89040 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_799
timestamp 1667941163
transform 1 0 90832 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_803
timestamp 1667941163
transform 1 0 91280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_806
timestamp 1667941163
transform 1 0 91616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_810
timestamp 1667941163
transform 1 0 92064 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_815
timestamp 1667941163
transform 1 0 92624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_821
timestamp 1667941163
transform 1 0 93296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_827
timestamp 1667941163
transform 1 0 93968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_831
timestamp 1667941163
transform 1 0 94416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_836
timestamp 1667941163
transform 1 0 94976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_840
timestamp 1667941163
transform 1 0 95424 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_842
timestamp 1667941163
transform 1 0 95648 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_847
timestamp 1667941163
transform 1 0 96208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1667941163
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_854
timestamp 1667941163
transform 1 0 96992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_859
timestamp 1667941163
transform 1 0 97552 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_865
timestamp 1667941163
transform 1 0 98224 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_897
timestamp 1667941163
transform 1 0 101808 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_913
timestamp 1667941163
transform 1 0 103600 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_921
timestamp 1667941163
transform 1 0 104496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_925
timestamp 1667941163
transform 1 0 104944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_929
timestamp 1667941163
transform 1 0 105392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_948
timestamp 1667941163
transform 1 0 107520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_956
timestamp 1667941163
transform 1 0 108416 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_964
timestamp 1667941163
transform 1 0 109312 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_966
timestamp 1667941163
transform 1 0 109536 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_971
timestamp 1667941163
transform 1 0 110096 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_987
timestamp 1667941163
transform 1 0 111888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_991
timestamp 1667941163
transform 1 0 112336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_993
timestamp 1667941163
transform 1 0 112560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1667941163
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1001
timestamp 1667941163
transform 1 0 113456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1007
timestamp 1667941163
transform 1 0 114128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1013
timestamp 1667941163
transform 1 0 114800 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1019
timestamp 1667941163
transform 1 0 115472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1025
timestamp 1667941163
transform 1 0 116144 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1041
timestamp 1667941163
transform 1 0 117936 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1045
timestamp 1667941163
transform 1 0 118384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1064
timestamp 1667941163
transform 1 0 120512 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1067
timestamp 1667941163
transform 1 0 120848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_1072
timestamp 1667941163
transform 1 0 121408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1104
timestamp 1667941163
transform 1 0 124992 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1120
timestamp 1667941163
transform 1 0 126784 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1123
timestamp 1667941163
transform 1 0 127120 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1127
timestamp 1667941163
transform 1 0 127568 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1135
timestamp 1667941163
transform 1 0 128464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1667941163
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1143
timestamp 1667941163
transform 1 0 129360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1151
timestamp 1667941163
transform 1 0 130256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1170
timestamp 1667941163
transform 1 0 132384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1176
timestamp 1667941163
transform 1 0 133056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1182
timestamp 1667941163
transform 1 0 133728 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1198
timestamp 1667941163
transform 1 0 135520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1667941163
transform 1 0 136416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1209
timestamp 1667941163
transform 1 0 136752 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1225
timestamp 1667941163
transform 1 0 138544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1246
timestamp 1667941163
transform 1 0 140896 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1252
timestamp 1667941163
transform 1 0 141568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1258
timestamp 1667941163
transform 1 0 142240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1262
timestamp 1667941163
transform 1 0 142688 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_1280
timestamp 1667941163
transform 1 0 144704 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1312
timestamp 1667941163
transform 1 0 148288 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1328
timestamp 1667941163
transform 1 0 150080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1330
timestamp 1667941163
transform 1 0 150304 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1333
timestamp 1667941163
transform 1 0 150640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1337
timestamp 1667941163
transform 1 0 151088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1341
timestamp 1667941163
transform 1 0 151536 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1346
timestamp 1667941163
transform 1 0 152096 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1348
timestamp 1667941163
transform 1 0 152320 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1351
timestamp 1667941163
transform 1 0 152656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1355
timestamp 1667941163
transform 1 0 153104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_1361
timestamp 1667941163
transform 1 0 153776 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1393
timestamp 1667941163
transform 1 0 157360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1409
timestamp 1667941163
transform 1 0 159152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1417
timestamp 1667941163
transform 1 0 160048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1419
timestamp 1667941163
transform 1 0 160272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1422
timestamp 1667941163
transform 1 0 160608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1486
timestamp 1667941163
transform 1 0 167776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1490
timestamp 1667941163
transform 1 0 168224 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_1493
timestamp 1667941163
transform 1 0 168560 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1557
timestamp 1667941163
transform 1 0 175728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1561
timestamp 1667941163
transform 1 0 176176 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1564
timestamp 1667941163
transform 1 0 176512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1580
timestamp 1667941163
transform 1 0 178304 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1667941163
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1667941163
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1667941163
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1667941163
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1667941163
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1667941163
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1667941163
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1667941163
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_250
timestamp 1667941163
transform 1 0 29344 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_282
timestamp 1667941163
transform 1 0 32928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_303
timestamp 1667941163
transform 1 0 35280 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_307
timestamp 1667941163
transform 1 0 35728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_315
timestamp 1667941163
transform 1 0 36624 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1667941163
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1667941163
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1667941163
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1667941163
transform 1 0 45248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_408
timestamp 1667941163
transform 1 0 47040 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_416
timestamp 1667941163
transform 1 0 47936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_418
timestamp 1667941163
transform 1 0 48160 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_436
timestamp 1667941163
transform 1 0 50176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_440
timestamp 1667941163
transform 1 0 50624 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1667941163
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1667941163
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_463
timestamp 1667941163
transform 1 0 53200 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_479
timestamp 1667941163
transform 1 0 54992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_487
timestamp 1667941163
transform 1 0 55888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_495
timestamp 1667941163
transform 1 0 56784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_503
timestamp 1667941163
transform 1 0 57680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_511
timestamp 1667941163
transform 1 0 58576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_519
timestamp 1667941163
transform 1 0 59472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_527
timestamp 1667941163
transform 1 0 60368 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1667941163
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1667941163
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_541
timestamp 1667941163
transform 1 0 61936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_545
timestamp 1667941163
transform 1 0 62384 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_548
timestamp 1667941163
transform 1 0 62720 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_552
timestamp 1667941163
transform 1 0 63168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_560
timestamp 1667941163
transform 1 0 64064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_568
timestamp 1667941163
transform 1 0 64960 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_576
timestamp 1667941163
transform 1 0 65856 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_584
timestamp 1667941163
transform 1 0 66752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_586
timestamp 1667941163
transform 1 0 66976 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_593
timestamp 1667941163
transform 1 0 67760 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_601
timestamp 1667941163
transform 1 0 68656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1667941163
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_608
timestamp 1667941163
transform 1 0 69440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_610
timestamp 1667941163
transform 1 0 69664 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_613
timestamp 1667941163
transform 1 0 70000 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_617
timestamp 1667941163
transform 1 0 70448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_621
timestamp 1667941163
transform 1 0 70896 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_653
timestamp 1667941163
transform 1 0 74480 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_661
timestamp 1667941163
transform 1 0 75376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_663
timestamp 1667941163
transform 1 0 75600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_666
timestamp 1667941163
transform 1 0 75936 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_676
timestamp 1667941163
transform 1 0 77056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_684
timestamp 1667941163
transform 1 0 77952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_688
timestamp 1667941163
transform 1 0 78400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_696
timestamp 1667941163
transform 1 0 79296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_706
timestamp 1667941163
transform 1 0 80416 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_722
timestamp 1667941163
transform 1 0 82208 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_726
timestamp 1667941163
transform 1 0 82656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_734
timestamp 1667941163
transform 1 0 83552 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_738
timestamp 1667941163
transform 1 0 84000 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_740
timestamp 1667941163
transform 1 0 84224 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_743
timestamp 1667941163
transform 1 0 84560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_747
timestamp 1667941163
transform 1 0 85008 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_751
timestamp 1667941163
transform 1 0 85456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_757
timestamp 1667941163
transform 1 0 86128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_763
timestamp 1667941163
transform 1 0 86800 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_795
timestamp 1667941163
transform 1 0 90384 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1667941163
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_818
timestamp 1667941163
transform 1 0 92960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_823
timestamp 1667941163
transform 1 0 93520 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_831
timestamp 1667941163
transform 1 0 94416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_837
timestamp 1667941163
transform 1 0 95088 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_843
timestamp 1667941163
transform 1 0 95760 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_849
timestamp 1667941163
transform 1 0 96432 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_855
timestamp 1667941163
transform 1 0 97104 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_861
timestamp 1667941163
transform 1 0 97776 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_867
timestamp 1667941163
transform 1 0 98448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_873
timestamp 1667941163
transform 1 0 99120 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_881
timestamp 1667941163
transform 1 0 100016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_885
timestamp 1667941163
transform 1 0 100464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_889
timestamp 1667941163
transform 1 0 100912 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_921
timestamp 1667941163
transform 1 0 104496 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_931
timestamp 1667941163
transform 1 0 105616 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_950
timestamp 1667941163
transform 1 0 107744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_956
timestamp 1667941163
transform 1 0 108416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_960
timestamp 1667941163
transform 1 0 108864 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_976
timestamp 1667941163
transform 1 0 110656 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_984
timestamp 1667941163
transform 1 0 111552 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_988
timestamp 1667941163
transform 1 0 112000 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_993
timestamp 1667941163
transform 1 0 112560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_999
timestamp 1667941163
transform 1 0 113232 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1005
timestamp 1667941163
transform 1 0 113904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1011
timestamp 1667941163
transform 1 0 114576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1017
timestamp 1667941163
transform 1 0 115248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1023
timestamp 1667941163
transform 1 0 115920 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1027
timestamp 1667941163
transform 1 0 116368 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1031
timestamp 1667941163
transform 1 0 116816 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1039
timestamp 1667941163
transform 1 0 117712 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1043
timestamp 1667941163
transform 1 0 118160 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1046
timestamp 1667941163
transform 1 0 118496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1065
timestamp 1667941163
transform 1 0 120624 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1071
timestamp 1667941163
transform 1 0 121296 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1087
timestamp 1667941163
transform 1 0 123088 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1095
timestamp 1667941163
transform 1 0 123984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1099
timestamp 1667941163
transform 1 0 124432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1102
timestamp 1667941163
transform 1 0 124768 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1166
timestamp 1667941163
transform 1 0 131936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1170
timestamp 1667941163
transform 1 0 132384 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1173
timestamp 1667941163
transform 1 0 132720 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1237
timestamp 1667941163
transform 1 0 139888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1241
timestamp 1667941163
transform 1 0 140336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1244
timestamp 1667941163
transform 1 0 140672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1248
timestamp 1667941163
transform 1 0 141120 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_1253
timestamp 1667941163
transform 1 0 141680 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1285
timestamp 1667941163
transform 1 0 145264 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1301
timestamp 1667941163
transform 1 0 147056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1309
timestamp 1667941163
transform 1 0 147952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1315
timestamp 1667941163
transform 1 0 148624 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1379
timestamp 1667941163
transform 1 0 155792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1383
timestamp 1667941163
transform 1 0 156240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1386
timestamp 1667941163
transform 1 0 156576 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1450
timestamp 1667941163
transform 1 0 163744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1454
timestamp 1667941163
transform 1 0 164192 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_1457
timestamp 1667941163
transform 1 0 164528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1521
timestamp 1667941163
transform 1 0 171696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1525
timestamp 1667941163
transform 1 0 172144 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_1528
timestamp 1667941163
transform 1 0 172480 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1560
timestamp 1667941163
transform 1 0 176064 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1576
timestamp 1667941163
transform 1 0 177856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1580
timestamp 1667941163
transform 1 0 178304 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1667941163
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1667941163
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1667941163
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1667941163
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1667941163
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1667941163
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1667941163
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1667941163
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1667941163
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1667941163
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1667941163
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1667941163
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1667941163
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_428
timestamp 1667941163
transform 1 0 49280 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_460
timestamp 1667941163
transform 1 0 52864 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_476
timestamp 1667941163
transform 1 0 54656 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_484
timestamp 1667941163
transform 1 0 55552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_488
timestamp 1667941163
transform 1 0 56000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1667941163
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_499
timestamp 1667941163
transform 1 0 57232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_507
timestamp 1667941163
transform 1 0 58128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_515
timestamp 1667941163
transform 1 0 59024 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_519
timestamp 1667941163
transform 1 0 59472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_528
timestamp 1667941163
transform 1 0 60480 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_532
timestamp 1667941163
transform 1 0 60928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_536
timestamp 1667941163
transform 1 0 61376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_540
timestamp 1667941163
transform 1 0 61824 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_543
timestamp 1667941163
transform 1 0 62160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_547
timestamp 1667941163
transform 1 0 62608 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_551
timestamp 1667941163
transform 1 0 63056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_555
timestamp 1667941163
transform 1 0 63504 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_559
timestamp 1667941163
transform 1 0 63952 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1667941163
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_570
timestamp 1667941163
transform 1 0 65184 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_576
timestamp 1667941163
transform 1 0 65856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_584
timestamp 1667941163
transform 1 0 66752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_592
timestamp 1667941163
transform 1 0 67648 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_600
timestamp 1667941163
transform 1 0 68544 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_604
timestamp 1667941163
transform 1 0 68992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_608
timestamp 1667941163
transform 1 0 69440 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_624
timestamp 1667941163
transform 1 0 71232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_632
timestamp 1667941163
transform 1 0 72128 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_636
timestamp 1667941163
transform 1 0 72576 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1667941163
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_641
timestamp 1667941163
transform 1 0 73136 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_673
timestamp 1667941163
transform 1 0 76720 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_689
timestamp 1667941163
transform 1 0 78512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_693
timestamp 1667941163
transform 1 0 78960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_695
timestamp 1667941163
transform 1 0 79184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_698
timestamp 1667941163
transform 1 0 79520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_706
timestamp 1667941163
transform 1 0 80416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_712
timestamp 1667941163
transform 1 0 81088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_776
timestamp 1667941163
transform 1 0 88256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1667941163
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_783
timestamp 1667941163
transform 1 0 89040 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_815
timestamp 1667941163
transform 1 0 92624 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_831
timestamp 1667941163
transform 1 0 94416 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_839
timestamp 1667941163
transform 1 0 95312 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_843
timestamp 1667941163
transform 1 0 95760 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_848
timestamp 1667941163
transform 1 0 96320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_854
timestamp 1667941163
transform 1 0 96992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_859
timestamp 1667941163
transform 1 0 97552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_865
timestamp 1667941163
transform 1 0 98224 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_897
timestamp 1667941163
transform 1 0 101808 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_913
timestamp 1667941163
transform 1 0 103600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_921
timestamp 1667941163
transform 1 0 104496 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_925
timestamp 1667941163
transform 1 0 104944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_941
timestamp 1667941163
transform 1 0 106736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_945
timestamp 1667941163
transform 1 0 107184 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_947
timestamp 1667941163
transform 1 0 107408 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_952
timestamp 1667941163
transform 1 0 107968 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_984
timestamp 1667941163
transform 1 0 111552 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_992
timestamp 1667941163
transform 1 0 112448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_996
timestamp 1667941163
transform 1 0 112896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1001
timestamp 1667941163
transform 1 0 113456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1007
timestamp 1667941163
transform 1 0 114128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1013
timestamp 1667941163
transform 1 0 114800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_1019
timestamp 1667941163
transform 1 0 115472 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1051
timestamp 1667941163
transform 1 0 119056 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1059
timestamp 1667941163
transform 1 0 119952 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1063
timestamp 1667941163
transform 1 0 120400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1067
timestamp 1667941163
transform 1 0 120848 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1131
timestamp 1667941163
transform 1 0 128016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1135
timestamp 1667941163
transform 1 0 128464 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1138
timestamp 1667941163
transform 1 0 128800 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1202
timestamp 1667941163
transform 1 0 135968 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1206
timestamp 1667941163
transform 1 0 136416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1209
timestamp 1667941163
transform 1 0 136752 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1273
timestamp 1667941163
transform 1 0 143920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1667941163
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1280
timestamp 1667941163
transform 1 0 144704 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1344
timestamp 1667941163
transform 1 0 151872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1348
timestamp 1667941163
transform 1 0 152320 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1351
timestamp 1667941163
transform 1 0 152656 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1415
timestamp 1667941163
transform 1 0 159824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1419
timestamp 1667941163
transform 1 0 160272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1422
timestamp 1667941163
transform 1 0 160608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1486
timestamp 1667941163
transform 1 0 167776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1490
timestamp 1667941163
transform 1 0 168224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1493
timestamp 1667941163
transform 1 0 168560 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1557
timestamp 1667941163
transform 1 0 175728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1561
timestamp 1667941163
transform 1 0 176176 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1564
timestamp 1667941163
transform 1 0 176512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1580
timestamp 1667941163
transform 1 0 178304 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1667941163
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1667941163
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1667941163
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1667941163
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1667941163
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1667941163
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1667941163
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1667941163
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1667941163
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1667941163
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1667941163
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1667941163
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1667941163
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1667941163
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1667941163
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1667941163
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_463
timestamp 1667941163
transform 1 0 53200 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_495
timestamp 1667941163
transform 1 0 56784 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_499
timestamp 1667941163
transform 1 0 57232 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_506
timestamp 1667941163
transform 1 0 58016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_514
timestamp 1667941163
transform 1 0 58912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_522
timestamp 1667941163
transform 1 0 59808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_526
timestamp 1667941163
transform 1 0 60256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_530
timestamp 1667941163
transform 1 0 60704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_534
timestamp 1667941163
transform 1 0 61152 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_550
timestamp 1667941163
transform 1 0 62944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_554
timestamp 1667941163
transform 1 0 63392 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_558
timestamp 1667941163
transform 1 0 63840 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_562
timestamp 1667941163
transform 1 0 64288 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_566
timestamp 1667941163
transform 1 0 64736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_574
timestamp 1667941163
transform 1 0 65632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_582
timestamp 1667941163
transform 1 0 66528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_590
timestamp 1667941163
transform 1 0 67424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_594
timestamp 1667941163
transform 1 0 67872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_598
timestamp 1667941163
transform 1 0 68320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1667941163
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1667941163
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1667941163
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1667941163
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1667941163
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1667941163
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1667941163
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1667941163
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1667941163
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1667941163
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_818
timestamp 1667941163
transform 1 0 92960 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_834
timestamp 1667941163
transform 1 0 94752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_842
timestamp 1667941163
transform 1 0 95648 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_846
timestamp 1667941163
transform 1 0 96096 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_851
timestamp 1667941163
transform 1 0 96656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_857
timestamp 1667941163
transform 1 0 97328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_873
timestamp 1667941163
transform 1 0 99120 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_881
timestamp 1667941163
transform 1 0 100016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_885
timestamp 1667941163
transform 1 0 100464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_889
timestamp 1667941163
transform 1 0 100912 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_953
timestamp 1667941163
transform 1 0 108080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1667941163
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_960
timestamp 1667941163
transform 1 0 108864 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_992
timestamp 1667941163
transform 1 0 112448 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1008
timestamp 1667941163
transform 1 0 114240 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1010
timestamp 1667941163
transform 1 0 114464 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1015
timestamp 1667941163
transform 1 0 115024 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1023
timestamp 1667941163
transform 1 0 115920 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1027
timestamp 1667941163
transform 1 0 116368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1031
timestamp 1667941163
transform 1 0 116816 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1095
timestamp 1667941163
transform 1 0 123984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1667941163
transform 1 0 124432 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1102
timestamp 1667941163
transform 1 0 124768 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1166
timestamp 1667941163
transform 1 0 131936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1170
timestamp 1667941163
transform 1 0 132384 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1173
timestamp 1667941163
transform 1 0 132720 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1237
timestamp 1667941163
transform 1 0 139888 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1241
timestamp 1667941163
transform 1 0 140336 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1244
timestamp 1667941163
transform 1 0 140672 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1308
timestamp 1667941163
transform 1 0 147840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1312
timestamp 1667941163
transform 1 0 148288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1315
timestamp 1667941163
transform 1 0 148624 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1379
timestamp 1667941163
transform 1 0 155792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1383
timestamp 1667941163
transform 1 0 156240 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1386
timestamp 1667941163
transform 1 0 156576 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1450
timestamp 1667941163
transform 1 0 163744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1454
timestamp 1667941163
transform 1 0 164192 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1457
timestamp 1667941163
transform 1 0 164528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1521
timestamp 1667941163
transform 1 0 171696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1525
timestamp 1667941163
transform 1 0 172144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1528
timestamp 1667941163
transform 1 0 172480 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1560
timestamp 1667941163
transform 1 0 176064 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1576
timestamp 1667941163
transform 1 0 177856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1580
timestamp 1667941163
transform 1 0 178304 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1667941163
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1667941163
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1667941163
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1667941163
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1667941163
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1667941163
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1667941163
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1667941163
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1667941163
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1667941163
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1667941163
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1667941163
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1667941163
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1667941163
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1667941163
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1667941163
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1667941163
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_499
timestamp 1667941163
transform 1 0 57232 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_503
timestamp 1667941163
transform 1 0 57680 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_510
timestamp 1667941163
transform 1 0 58464 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_542
timestamp 1667941163
transform 1 0 62048 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_558
timestamp 1667941163
transform 1 0 63840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_566
timestamp 1667941163
transform 1 0 64736 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1667941163
transform 1 0 65184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_573
timestamp 1667941163
transform 1 0 65520 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_575
timestamp 1667941163
transform 1 0 65744 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_582
timestamp 1667941163
transform 1 0 66528 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_586
timestamp 1667941163
transform 1 0 66976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_590
timestamp 1667941163
transform 1 0 67424 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_594
timestamp 1667941163
transform 1 0 67872 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_626
timestamp 1667941163
transform 1 0 71456 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1667941163
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1667941163
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1667941163
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1667941163
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1667941163
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1667941163
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1667941163
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1667941163
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1667941163
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1667941163
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1667941163
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_854
timestamp 1667941163
transform 1 0 96992 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_918
timestamp 1667941163
transform 1 0 104160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_922
timestamp 1667941163
transform 1 0 104608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_925
timestamp 1667941163
transform 1 0 104944 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1667941163
transform 1 0 112112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1667941163
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_996
timestamp 1667941163
transform 1 0 112896 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1060
timestamp 1667941163
transform 1 0 120064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1064
timestamp 1667941163
transform 1 0 120512 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1067
timestamp 1667941163
transform 1 0 120848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1131
timestamp 1667941163
transform 1 0 128016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1667941163
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1138
timestamp 1667941163
transform 1 0 128800 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1202
timestamp 1667941163
transform 1 0 135968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1667941163
transform 1 0 136416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1209
timestamp 1667941163
transform 1 0 136752 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1273
timestamp 1667941163
transform 1 0 143920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1277
timestamp 1667941163
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1280
timestamp 1667941163
transform 1 0 144704 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1344
timestamp 1667941163
transform 1 0 151872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1348
timestamp 1667941163
transform 1 0 152320 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1351
timestamp 1667941163
transform 1 0 152656 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1415
timestamp 1667941163
transform 1 0 159824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1419
timestamp 1667941163
transform 1 0 160272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1422
timestamp 1667941163
transform 1 0 160608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1486
timestamp 1667941163
transform 1 0 167776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1490
timestamp 1667941163
transform 1 0 168224 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1493
timestamp 1667941163
transform 1 0 168560 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1557
timestamp 1667941163
transform 1 0 175728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1561
timestamp 1667941163
transform 1 0 176176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1564
timestamp 1667941163
transform 1 0 176512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1580
timestamp 1667941163
transform 1 0 178304 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1667941163
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1667941163
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1667941163
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1667941163
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1667941163
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1667941163
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1667941163
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1667941163
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1667941163
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1667941163
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1667941163
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1667941163
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1667941163
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1667941163
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1667941163
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1667941163
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1667941163
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1667941163
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1667941163
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1667941163
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1667941163
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1667941163
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1667941163
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1667941163
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1667941163
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1667941163
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1667941163
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1667941163
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1667941163
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1667941163
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1667941163
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1667941163
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_818
timestamp 1667941163
transform 1 0 92960 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_882
timestamp 1667941163
transform 1 0 100128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1667941163
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1667941163
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1667941163
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1667941163
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1667941163
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1667941163
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1667941163
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1031
timestamp 1667941163
transform 1 0 116816 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1095
timestamp 1667941163
transform 1 0 123984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1099
timestamp 1667941163
transform 1 0 124432 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1102
timestamp 1667941163
transform 1 0 124768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1166
timestamp 1667941163
transform 1 0 131936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1170
timestamp 1667941163
transform 1 0 132384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1173
timestamp 1667941163
transform 1 0 132720 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1237
timestamp 1667941163
transform 1 0 139888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1241
timestamp 1667941163
transform 1 0 140336 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1244
timestamp 1667941163
transform 1 0 140672 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1308
timestamp 1667941163
transform 1 0 147840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1312
timestamp 1667941163
transform 1 0 148288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1315
timestamp 1667941163
transform 1 0 148624 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1379
timestamp 1667941163
transform 1 0 155792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1383
timestamp 1667941163
transform 1 0 156240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1386
timestamp 1667941163
transform 1 0 156576 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1450
timestamp 1667941163
transform 1 0 163744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1454
timestamp 1667941163
transform 1 0 164192 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1457
timestamp 1667941163
transform 1 0 164528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1521
timestamp 1667941163
transform 1 0 171696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1525
timestamp 1667941163
transform 1 0 172144 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1528
timestamp 1667941163
transform 1 0 172480 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1560
timestamp 1667941163
transform 1 0 176064 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1576
timestamp 1667941163
transform 1 0 177856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1580
timestamp 1667941163
transform 1 0 178304 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1667941163
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1667941163
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1667941163
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1667941163
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1667941163
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1667941163
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1667941163
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1667941163
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1667941163
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1667941163
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1667941163
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1667941163
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1667941163
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1667941163
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1667941163
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1667941163
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1667941163
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1667941163
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1667941163
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1667941163
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1667941163
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1667941163
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1667941163
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1667941163
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1667941163
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1667941163
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1667941163
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1667941163
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1667941163
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1667941163
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1667941163
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1667941163
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1667941163
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1667941163
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1667941163
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1667941163
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1667941163
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1667941163
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_996
timestamp 1667941163
transform 1 0 112896 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1060
timestamp 1667941163
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1667941163
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1067
timestamp 1667941163
transform 1 0 120848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1131
timestamp 1667941163
transform 1 0 128016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1135
timestamp 1667941163
transform 1 0 128464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1138
timestamp 1667941163
transform 1 0 128800 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1667941163
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1667941163
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1667941163
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1667941163
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1667941163
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1280
timestamp 1667941163
transform 1 0 144704 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1344
timestamp 1667941163
transform 1 0 151872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1348
timestamp 1667941163
transform 1 0 152320 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1351
timestamp 1667941163
transform 1 0 152656 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1415
timestamp 1667941163
transform 1 0 159824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1419
timestamp 1667941163
transform 1 0 160272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1422
timestamp 1667941163
transform 1 0 160608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1486
timestamp 1667941163
transform 1 0 167776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1490
timestamp 1667941163
transform 1 0 168224 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1493
timestamp 1667941163
transform 1 0 168560 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1557
timestamp 1667941163
transform 1 0 175728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1561
timestamp 1667941163
transform 1 0 176176 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1564
timestamp 1667941163
transform 1 0 176512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1580
timestamp 1667941163
transform 1 0 178304 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1667941163
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1667941163
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1667941163
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1667941163
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1667941163
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1667941163
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1667941163
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1667941163
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1667941163
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1667941163
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1667941163
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1667941163
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1667941163
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1667941163
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1667941163
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1667941163
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1667941163
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1667941163
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1667941163
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1667941163
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1667941163
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1667941163
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1667941163
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1667941163
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1667941163
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1667941163
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1667941163
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1667941163
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1667941163
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1667941163
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1667941163
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1667941163
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1667941163
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1667941163
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1667941163
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1667941163
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1667941163
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1667941163
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1667941163
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1667941163
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1031
timestamp 1667941163
transform 1 0 116816 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1095
timestamp 1667941163
transform 1 0 123984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1099
timestamp 1667941163
transform 1 0 124432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1102
timestamp 1667941163
transform 1 0 124768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1166
timestamp 1667941163
transform 1 0 131936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1170
timestamp 1667941163
transform 1 0 132384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1667941163
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1667941163
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1667941163
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1244
timestamp 1667941163
transform 1 0 140672 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1308
timestamp 1667941163
transform 1 0 147840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1312
timestamp 1667941163
transform 1 0 148288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1315
timestamp 1667941163
transform 1 0 148624 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1379
timestamp 1667941163
transform 1 0 155792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1383
timestamp 1667941163
transform 1 0 156240 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1386
timestamp 1667941163
transform 1 0 156576 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1450
timestamp 1667941163
transform 1 0 163744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1454
timestamp 1667941163
transform 1 0 164192 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1457
timestamp 1667941163
transform 1 0 164528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1521
timestamp 1667941163
transform 1 0 171696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1525
timestamp 1667941163
transform 1 0 172144 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1528
timestamp 1667941163
transform 1 0 172480 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_1560
timestamp 1667941163
transform 1 0 176064 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1576
timestamp 1667941163
transform 1 0 177856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1580
timestamp 1667941163
transform 1 0 178304 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1667941163
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1667941163
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1667941163
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1667941163
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1667941163
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1667941163
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1667941163
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1667941163
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1667941163
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1667941163
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1667941163
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1667941163
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1667941163
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1667941163
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1667941163
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1667941163
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1667941163
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1667941163
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1667941163
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1667941163
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1667941163
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1667941163
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1667941163
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1667941163
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1667941163
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1667941163
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1667941163
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1667941163
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1667941163
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1667941163
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1667941163
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1667941163
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1667941163
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1667941163
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1667941163
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1667941163
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1667941163
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1667941163
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_996
timestamp 1667941163
transform 1 0 112896 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1667941163
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1667941163
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1667941163
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1667941163
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1667941163
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1667941163
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1667941163
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1667941163
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1667941163
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1667941163
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1667941163
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1280
timestamp 1667941163
transform 1 0 144704 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1344
timestamp 1667941163
transform 1 0 151872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1348
timestamp 1667941163
transform 1 0 152320 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1351
timestamp 1667941163
transform 1 0 152656 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1415
timestamp 1667941163
transform 1 0 159824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1419
timestamp 1667941163
transform 1 0 160272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1422
timestamp 1667941163
transform 1 0 160608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1486
timestamp 1667941163
transform 1 0 167776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1490
timestamp 1667941163
transform 1 0 168224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1493
timestamp 1667941163
transform 1 0 168560 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1557
timestamp 1667941163
transform 1 0 175728 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1561
timestamp 1667941163
transform 1 0 176176 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_1564
timestamp 1667941163
transform 1 0 176512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1580
timestamp 1667941163
transform 1 0 178304 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1667941163
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1667941163
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1667941163
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1667941163
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1667941163
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1667941163
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1667941163
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1667941163
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1667941163
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1667941163
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1667941163
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1667941163
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1667941163
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1667941163
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1667941163
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1667941163
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1667941163
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1667941163
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1667941163
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1667941163
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1667941163
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1667941163
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1667941163
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1667941163
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1667941163
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1667941163
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1667941163
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1667941163
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1667941163
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1667941163
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1667941163
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_882
timestamp 1667941163
transform 1 0 100128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1667941163
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1667941163
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1667941163
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1667941163
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1667941163
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1667941163
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1667941163
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1667941163
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1667941163
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1667941163
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1667941163
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1667941163
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1667941163
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1667941163
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1667941163
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1667941163
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1244
timestamp 1667941163
transform 1 0 140672 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1308
timestamp 1667941163
transform 1 0 147840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1312
timestamp 1667941163
transform 1 0 148288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1315
timestamp 1667941163
transform 1 0 148624 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1379
timestamp 1667941163
transform 1 0 155792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1383
timestamp 1667941163
transform 1 0 156240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1386
timestamp 1667941163
transform 1 0 156576 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1450
timestamp 1667941163
transform 1 0 163744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1454
timestamp 1667941163
transform 1 0 164192 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1457
timestamp 1667941163
transform 1 0 164528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1521
timestamp 1667941163
transform 1 0 171696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1525
timestamp 1667941163
transform 1 0 172144 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_1528
timestamp 1667941163
transform 1 0 172480 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_1560
timestamp 1667941163
transform 1 0 176064 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1576
timestamp 1667941163
transform 1 0 177856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1580
timestamp 1667941163
transform 1 0 178304 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1667941163
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1667941163
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1667941163
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1667941163
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1667941163
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1667941163
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1667941163
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1667941163
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1667941163
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1667941163
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1667941163
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1667941163
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1667941163
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1667941163
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1667941163
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1667941163
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1667941163
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1667941163
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1667941163
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1667941163
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1667941163
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1667941163
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1667941163
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1667941163
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1667941163
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1667941163
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1667941163
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1667941163
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1667941163
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1667941163
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1667941163
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1667941163
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_854
timestamp 1667941163
transform 1 0 96992 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_918
timestamp 1667941163
transform 1 0 104160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1667941163
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1667941163
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1667941163
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1667941163
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1667941163
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1667941163
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1667941163
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1667941163
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1667941163
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1667941163
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1667941163
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1667941163
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1667941163
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1667941163
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1273
timestamp 1667941163
transform 1 0 143920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1667941163
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1280
timestamp 1667941163
transform 1 0 144704 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1344
timestamp 1667941163
transform 1 0 151872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1348
timestamp 1667941163
transform 1 0 152320 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1351
timestamp 1667941163
transform 1 0 152656 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1415
timestamp 1667941163
transform 1 0 159824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1419
timestamp 1667941163
transform 1 0 160272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1422
timestamp 1667941163
transform 1 0 160608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1486
timestamp 1667941163
transform 1 0 167776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1490
timestamp 1667941163
transform 1 0 168224 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1493
timestamp 1667941163
transform 1 0 168560 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1557
timestamp 1667941163
transform 1 0 175728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1561
timestamp 1667941163
transform 1 0 176176 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_1564
timestamp 1667941163
transform 1 0 176512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1580
timestamp 1667941163
transform 1 0 178304 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1667941163
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1667941163
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1667941163
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1667941163
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1667941163
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1667941163
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1667941163
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1667941163
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1667941163
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1667941163
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1667941163
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1667941163
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1667941163
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1667941163
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1667941163
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1667941163
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1667941163
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1667941163
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1667941163
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1667941163
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1667941163
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1667941163
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1667941163
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1667941163
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1667941163
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1667941163
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1667941163
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1667941163
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1667941163
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1667941163
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1667941163
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1667941163
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1667941163
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1667941163
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1667941163
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_889
timestamp 1667941163
transform 1 0 100912 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_953
timestamp 1667941163
transform 1 0 108080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1667941163
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1667941163
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1667941163
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1667941163
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1667941163
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1667941163
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1667941163
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1667941163
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1667941163
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1667941163
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1667941163
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1667941163
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1667941163
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1244
timestamp 1667941163
transform 1 0 140672 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1308
timestamp 1667941163
transform 1 0 147840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1312
timestamp 1667941163
transform 1 0 148288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1315
timestamp 1667941163
transform 1 0 148624 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1379
timestamp 1667941163
transform 1 0 155792 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1383
timestamp 1667941163
transform 1 0 156240 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1386
timestamp 1667941163
transform 1 0 156576 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1450
timestamp 1667941163
transform 1 0 163744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1454
timestamp 1667941163
transform 1 0 164192 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1457
timestamp 1667941163
transform 1 0 164528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1521
timestamp 1667941163
transform 1 0 171696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1525
timestamp 1667941163
transform 1 0 172144 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_1528
timestamp 1667941163
transform 1 0 172480 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_1560
timestamp 1667941163
transform 1 0 176064 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1576
timestamp 1667941163
transform 1 0 177856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1580
timestamp 1667941163
transform 1 0 178304 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1667941163
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1667941163
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1667941163
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1667941163
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1667941163
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1667941163
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1667941163
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1667941163
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1667941163
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1667941163
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1667941163
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1667941163
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1667941163
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1667941163
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1667941163
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1667941163
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1667941163
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1667941163
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1667941163
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1667941163
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1667941163
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1667941163
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1667941163
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1667941163
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1667941163
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1667941163
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1667941163
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1667941163
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1667941163
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1667941163
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1667941163
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1667941163
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1667941163
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1667941163
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1667941163
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1667941163
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1667941163
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1667941163
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1667941163
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1667941163
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1667941163
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1667941163
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1667941163
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1667941163
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1667941163
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1667941163
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1667941163
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1667941163
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1667941163
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1280
timestamp 1667941163
transform 1 0 144704 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1344
timestamp 1667941163
transform 1 0 151872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1348
timestamp 1667941163
transform 1 0 152320 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1351
timestamp 1667941163
transform 1 0 152656 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1415
timestamp 1667941163
transform 1 0 159824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1419
timestamp 1667941163
transform 1 0 160272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1422
timestamp 1667941163
transform 1 0 160608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1486
timestamp 1667941163
transform 1 0 167776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1490
timestamp 1667941163
transform 1 0 168224 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1493
timestamp 1667941163
transform 1 0 168560 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1557
timestamp 1667941163
transform 1 0 175728 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1561
timestamp 1667941163
transform 1 0 176176 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_1564
timestamp 1667941163
transform 1 0 176512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1580
timestamp 1667941163
transform 1 0 178304 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1667941163
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1667941163
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1667941163
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1667941163
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1667941163
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1667941163
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1667941163
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1667941163
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1667941163
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1667941163
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1667941163
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1667941163
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1667941163
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1667941163
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1667941163
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1667941163
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1667941163
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1667941163
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1667941163
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1667941163
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1667941163
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1667941163
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1667941163
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1667941163
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1667941163
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1667941163
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1667941163
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1667941163
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1667941163
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1667941163
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1667941163
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1667941163
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1667941163
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1667941163
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1667941163
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1667941163
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1667941163
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1667941163
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1667941163
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1667941163
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1667941163
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1667941163
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1667941163
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1667941163
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1667941163
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1667941163
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1667941163
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1667941163
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1667941163
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1667941163
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1667941163
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1244
timestamp 1667941163
transform 1 0 140672 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1308
timestamp 1667941163
transform 1 0 147840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1312
timestamp 1667941163
transform 1 0 148288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1315
timestamp 1667941163
transform 1 0 148624 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1379
timestamp 1667941163
transform 1 0 155792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1383
timestamp 1667941163
transform 1 0 156240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1386
timestamp 1667941163
transform 1 0 156576 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1450
timestamp 1667941163
transform 1 0 163744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1454
timestamp 1667941163
transform 1 0 164192 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1457
timestamp 1667941163
transform 1 0 164528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1521
timestamp 1667941163
transform 1 0 171696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1525
timestamp 1667941163
transform 1 0 172144 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_1528
timestamp 1667941163
transform 1 0 172480 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_1560
timestamp 1667941163
transform 1 0 176064 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1576
timestamp 1667941163
transform 1 0 177856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1580
timestamp 1667941163
transform 1 0 178304 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1667941163
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1667941163
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1667941163
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1667941163
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1667941163
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1667941163
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1667941163
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1667941163
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1667941163
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1667941163
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1667941163
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1667941163
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1667941163
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1667941163
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1667941163
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1667941163
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1667941163
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1667941163
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1667941163
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1667941163
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1667941163
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1667941163
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1667941163
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1667941163
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1667941163
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1667941163
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1667941163
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1667941163
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1667941163
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1667941163
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1667941163
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1667941163
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1667941163
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1667941163
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1667941163
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1667941163
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1667941163
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1667941163
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1667941163
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1667941163
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1667941163
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1667941163
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1667941163
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1667941163
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1667941163
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1667941163
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1667941163
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1667941163
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1273
timestamp 1667941163
transform 1 0 143920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1667941163
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1280
timestamp 1667941163
transform 1 0 144704 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1344
timestamp 1667941163
transform 1 0 151872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1348
timestamp 1667941163
transform 1 0 152320 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1351
timestamp 1667941163
transform 1 0 152656 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1415
timestamp 1667941163
transform 1 0 159824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1419
timestamp 1667941163
transform 1 0 160272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1422
timestamp 1667941163
transform 1 0 160608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1486
timestamp 1667941163
transform 1 0 167776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1490
timestamp 1667941163
transform 1 0 168224 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1493
timestamp 1667941163
transform 1 0 168560 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1557
timestamp 1667941163
transform 1 0 175728 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1561
timestamp 1667941163
transform 1 0 176176 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_1564
timestamp 1667941163
transform 1 0 176512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1572
timestamp 1667941163
transform 1 0 177408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1580
timestamp 1667941163
transform 1 0 178304 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_2
timestamp 1667941163
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_10
timestamp 1667941163
transform 1 0 2464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_14
timestamp 1667941163
transform 1 0 2912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_19
timestamp 1667941163
transform 1 0 3472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_27
timestamp 1667941163
transform 1 0 4368 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_33
timestamp 1667941163
transform 1 0 5040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_37
timestamp 1667941163
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_53
timestamp 1667941163
transform 1 0 7280 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_61
timestamp 1667941163
transform 1 0 8176 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_69
timestamp 1667941163
transform 1 0 9072 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_72
timestamp 1667941163
transform 1 0 9408 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_77
timestamp 1667941163
transform 1 0 9968 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_93
timestamp 1667941163
transform 1 0 11760 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_97
timestamp 1667941163
transform 1 0 12208 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_103
timestamp 1667941163
transform 1 0 12880 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_107
timestamp 1667941163
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_111
timestamp 1667941163
transform 1 0 13776 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_117
timestamp 1667941163
transform 1 0 14448 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_133
timestamp 1667941163
transform 1 0 16240 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_137
timestamp 1667941163
transform 1 0 16688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 16912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_142
timestamp 1667941163
transform 1 0 17248 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_147
timestamp 1667941163
transform 1 0 17808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_159
timestamp 1667941163
transform 1 0 19152 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_177
timestamp 1667941163
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_181
timestamp 1667941163
transform 1 0 21616 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_187
timestamp 1667941163
transform 1 0 22288 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_195
timestamp 1667941163
transform 1 0 23184 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_201
timestamp 1667941163
transform 1 0 23856 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_209
timestamp 1667941163
transform 1 0 24752 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_212
timestamp 1667941163
transform 1 0 25088 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_220
timestamp 1667941163
transform 1 0 25984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_224
timestamp 1667941163
transform 1 0 26432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_229
timestamp 1667941163
transform 1 0 26992 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_237
timestamp 1667941163
transform 1 0 27888 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_243
timestamp 1667941163
transform 1 0 28560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_247
timestamp 1667941163
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_263
timestamp 1667941163
transform 1 0 30800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_271
timestamp 1667941163
transform 1 0 31696 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_279
timestamp 1667941163
transform 1 0 32592 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_282
timestamp 1667941163
transform 1 0 32928 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_287
timestamp 1667941163
transform 1 0 33488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_303
timestamp 1667941163
transform 1 0 35280 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_307
timestamp 1667941163
transform 1 0 35728 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_313
timestamp 1667941163
transform 1 0 36400 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_317
timestamp 1667941163
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_321
timestamp 1667941163
transform 1 0 37296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_327
timestamp 1667941163
transform 1 0 37968 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_343
timestamp 1667941163
transform 1 0 39760 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_347
timestamp 1667941163
transform 1 0 40208 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_349
timestamp 1667941163
transform 1 0 40432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_352
timestamp 1667941163
transform 1 0 40768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_357
timestamp 1667941163
transform 1 0 41328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_369
timestamp 1667941163
transform 1 0 42672 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_387
timestamp 1667941163
transform 1 0 44688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_391
timestamp 1667941163
transform 1 0 45136 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_397
timestamp 1667941163
transform 1 0 45808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 46704 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_411
timestamp 1667941163
transform 1 0 47376 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_419
timestamp 1667941163
transform 1 0 48272 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_422
timestamp 1667941163
transform 1 0 48608 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_430
timestamp 1667941163
transform 1 0 49504 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_434
timestamp 1667941163
transform 1 0 49952 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_439
timestamp 1667941163
transform 1 0 50512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_447
timestamp 1667941163
transform 1 0 51408 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_453
timestamp 1667941163
transform 1 0 52080 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_457
timestamp 1667941163
transform 1 0 52528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_473
timestamp 1667941163
transform 1 0 54320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_481
timestamp 1667941163
transform 1 0 55216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_489
timestamp 1667941163
transform 1 0 56112 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_492
timestamp 1667941163
transform 1 0 56448 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_497
timestamp 1667941163
transform 1 0 57008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_513
timestamp 1667941163
transform 1 0 58800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_517
timestamp 1667941163
transform 1 0 59248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_523
timestamp 1667941163
transform 1 0 59920 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1667941163
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_531
timestamp 1667941163
transform 1 0 60816 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_537
timestamp 1667941163
transform 1 0 61488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_553
timestamp 1667941163
transform 1 0 63280 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_557
timestamp 1667941163
transform 1 0 63728 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_559
timestamp 1667941163
transform 1 0 63952 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_562
timestamp 1667941163
transform 1 0 64288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_567
timestamp 1667941163
transform 1 0 64848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_579
timestamp 1667941163
transform 1 0 66192 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_597
timestamp 1667941163
transform 1 0 68208 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_601
timestamp 1667941163
transform 1 0 68656 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_607
timestamp 1667941163
transform 1 0 69328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_615
timestamp 1667941163
transform 1 0 70224 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_621
timestamp 1667941163
transform 1 0 70896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_629
timestamp 1667941163
transform 1 0 71792 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_632
timestamp 1667941163
transform 1 0 72128 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_640
timestamp 1667941163
transform 1 0 73024 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_644
timestamp 1667941163
transform 1 0 73472 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_649
timestamp 1667941163
transform 1 0 74032 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_657
timestamp 1667941163
transform 1 0 74928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_663
timestamp 1667941163
transform 1 0 75600 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_667
timestamp 1667941163
transform 1 0 76048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_683
timestamp 1667941163
transform 1 0 77840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_691
timestamp 1667941163
transform 1 0 78736 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_699
timestamp 1667941163
transform 1 0 79632 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_702
timestamp 1667941163
transform 1 0 79968 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_707
timestamp 1667941163
transform 1 0 80528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_723
timestamp 1667941163
transform 1 0 82320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_727
timestamp 1667941163
transform 1 0 82768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_733
timestamp 1667941163
transform 1 0 83440 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_737
timestamp 1667941163
transform 1 0 83888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_741
timestamp 1667941163
transform 1 0 84336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_747
timestamp 1667941163
transform 1 0 85008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_763
timestamp 1667941163
transform 1 0 86800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_767
timestamp 1667941163
transform 1 0 87248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_769
timestamp 1667941163
transform 1 0 87472 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_772
timestamp 1667941163
transform 1 0 87808 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_777
timestamp 1667941163
transform 1 0 88368 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_789
timestamp 1667941163
transform 1 0 89712 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_807
timestamp 1667941163
transform 1 0 91728 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_811
timestamp 1667941163
transform 1 0 92176 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_817
timestamp 1667941163
transform 1 0 92848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_825
timestamp 1667941163
transform 1 0 93744 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_831
timestamp 1667941163
transform 1 0 94416 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_839
timestamp 1667941163
transform 1 0 95312 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_842
timestamp 1667941163
transform 1 0 95648 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_850
timestamp 1667941163
transform 1 0 96544 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_854
timestamp 1667941163
transform 1 0 96992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_859
timestamp 1667941163
transform 1 0 97552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_867
timestamp 1667941163
transform 1 0 98448 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_873
timestamp 1667941163
transform 1 0 99120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_877
timestamp 1667941163
transform 1 0 99568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_893
timestamp 1667941163
transform 1 0 101360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_901
timestamp 1667941163
transform 1 0 102256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_909
timestamp 1667941163
transform 1 0 103152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_912
timestamp 1667941163
transform 1 0 103488 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_917
timestamp 1667941163
transform 1 0 104048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_933
timestamp 1667941163
transform 1 0 105840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_937
timestamp 1667941163
transform 1 0 106288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_943
timestamp 1667941163
transform 1 0 106960 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_947
timestamp 1667941163
transform 1 0 107408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_951
timestamp 1667941163
transform 1 0 107856 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_957
timestamp 1667941163
transform 1 0 108528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_973
timestamp 1667941163
transform 1 0 110320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_977
timestamp 1667941163
transform 1 0 110768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_979
timestamp 1667941163
transform 1 0 110992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_982
timestamp 1667941163
transform 1 0 111328 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_987
timestamp 1667941163
transform 1 0 111888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_999
timestamp 1667941163
transform 1 0 113232 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1017
timestamp 1667941163
transform 1 0 115248 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1021
timestamp 1667941163
transform 1 0 115696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1027
timestamp 1667941163
transform 1 0 116368 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1035
timestamp 1667941163
transform 1 0 117264 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1041
timestamp 1667941163
transform 1 0 117936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1049
timestamp 1667941163
transform 1 0 118832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1052
timestamp 1667941163
transform 1 0 119168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1060
timestamp 1667941163
transform 1 0 120064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1064
timestamp 1667941163
transform 1 0 120512 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1069
timestamp 1667941163
transform 1 0 121072 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1077
timestamp 1667941163
transform 1 0 121968 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1083
timestamp 1667941163
transform 1 0 122640 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1087
timestamp 1667941163
transform 1 0 123088 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1103
timestamp 1667941163
transform 1 0 124880 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1111
timestamp 1667941163
transform 1 0 125776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1119
timestamp 1667941163
transform 1 0 126672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1122
timestamp 1667941163
transform 1 0 127008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1127
timestamp 1667941163
transform 1 0 127568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1143
timestamp 1667941163
transform 1 0 129360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1147
timestamp 1667941163
transform 1 0 129808 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1153
timestamp 1667941163
transform 1 0 130480 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1157
timestamp 1667941163
transform 1 0 130928 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1161
timestamp 1667941163
transform 1 0 131376 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1167
timestamp 1667941163
transform 1 0 132048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1183
timestamp 1667941163
transform 1 0 133840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1187
timestamp 1667941163
transform 1 0 134288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1189
timestamp 1667941163
transform 1 0 134512 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1192
timestamp 1667941163
transform 1 0 134848 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1197
timestamp 1667941163
transform 1 0 135408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1209
timestamp 1667941163
transform 1 0 136752 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1227
timestamp 1667941163
transform 1 0 138768 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1231
timestamp 1667941163
transform 1 0 139216 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1237
timestamp 1667941163
transform 1 0 139888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1245
timestamp 1667941163
transform 1 0 140784 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1251
timestamp 1667941163
transform 1 0 141456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1259
timestamp 1667941163
transform 1 0 142352 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1262
timestamp 1667941163
transform 1 0 142688 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1270
timestamp 1667941163
transform 1 0 143584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1274
timestamp 1667941163
transform 1 0 144032 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1279
timestamp 1667941163
transform 1 0 144592 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1287
timestamp 1667941163
transform 1 0 145488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1293
timestamp 1667941163
transform 1 0 146160 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1297
timestamp 1667941163
transform 1 0 146608 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1313
timestamp 1667941163
transform 1 0 148400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1321
timestamp 1667941163
transform 1 0 149296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1329
timestamp 1667941163
transform 1 0 150192 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1332
timestamp 1667941163
transform 1 0 150528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1337
timestamp 1667941163
transform 1 0 151088 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1353
timestamp 1667941163
transform 1 0 152880 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1357
timestamp 1667941163
transform 1 0 153328 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1363
timestamp 1667941163
transform 1 0 154000 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1367
timestamp 1667941163
transform 1 0 154448 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1371
timestamp 1667941163
transform 1 0 154896 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1377
timestamp 1667941163
transform 1 0 155568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1393
timestamp 1667941163
transform 1 0 157360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1397
timestamp 1667941163
transform 1 0 157808 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1399
timestamp 1667941163
transform 1 0 158032 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1402
timestamp 1667941163
transform 1 0 158368 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1407
timestamp 1667941163
transform 1 0 158928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1419
timestamp 1667941163
transform 1 0 160272 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1437
timestamp 1667941163
transform 1 0 162288 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1441
timestamp 1667941163
transform 1 0 162736 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1447
timestamp 1667941163
transform 1 0 163408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1455
timestamp 1667941163
transform 1 0 164304 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1461
timestamp 1667941163
transform 1 0 164976 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1469
timestamp 1667941163
transform 1 0 165872 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1472
timestamp 1667941163
transform 1 0 166208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1480
timestamp 1667941163
transform 1 0 167104 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1484
timestamp 1667941163
transform 1 0 167552 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1489
timestamp 1667941163
transform 1 0 168112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1497
timestamp 1667941163
transform 1 0 169008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1503
timestamp 1667941163
transform 1 0 169680 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1507
timestamp 1667941163
transform 1 0 170128 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1523
timestamp 1667941163
transform 1 0 171920 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1531
timestamp 1667941163
transform 1 0 172816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1539
timestamp 1667941163
transform 1 0 173712 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1542
timestamp 1667941163
transform 1 0 174048 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1547
timestamp 1667941163
transform 1 0 174608 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1563
timestamp 1667941163
transform 1 0 176400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1567
timestamp 1667941163
transform 1 0 176848 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1573
timestamp 1667941163
transform 1 0 177520 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1577
timestamp 1667941163
transform 1 0 177968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 178640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 178640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 178640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 178640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 178640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 178640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 178640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 178640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 178640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 178640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 178640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 178640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 178640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 178640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 178640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 178640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 178640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1667941163
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1667941163
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1667941163
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1667941163
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1667941163
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1667941163
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1667941163
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1667941163
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1667941163
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1667941163
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1667941163
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1667941163
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1667941163
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1667941163
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1667941163
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1667941163
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1667941163
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1667941163
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1667941163
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1667941163
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1667941163
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1667941163
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1667941163
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1667941163
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1667941163
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1667941163
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1667941163
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1667941163
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1667941163
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1667941163
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1667941163
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1667941163
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1667941163
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1667941163
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1667941163
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1667941163
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1667941163
transform 1 0 150304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1667941163
transform 1 0 154224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1667941163
transform 1 0 158144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1667941163
transform 1 0 162064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1667941163
transform 1 0 165984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1667941163
transform 1 0 169904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1667941163
transform 1 0 173824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1667941163
transform 1 0 177744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1667941163
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_81
timestamp 1667941163
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_82
timestamp 1667941163
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_83
timestamp 1667941163
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1667941163
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1667941163
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1667941163
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1667941163
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1667941163
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1667941163
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1667941163
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1667941163
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1667941163
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1667941163
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1667941163
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1667941163
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1667941163
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1667941163
transform 1 0 152432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1667941163
transform 1 0 160384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1667941163
transform 1 0 168336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1667941163
transform 1 0 176288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1667941163
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1667941163
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1667941163
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1667941163
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1667941163
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1667941163
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1667941163
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1667941163
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1667941163
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1667941163
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1667941163
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1667941163
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1667941163
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1667941163
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1667941163
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1667941163
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1667941163
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1667941163
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1667941163
transform 1 0 148400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1667941163
transform 1 0 156352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1667941163
transform 1 0 164304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1667941163
transform 1 0 172256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1667941163
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1667941163
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1667941163
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1667941163
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1667941163
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1667941163
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1667941163
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1667941163
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1667941163
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1667941163
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1667941163
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1667941163
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1667941163
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1667941163
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1667941163
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1667941163
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1667941163
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1667941163
transform 1 0 152432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1667941163
transform 1 0 160384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1667941163
transform 1 0 168336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1667941163
transform 1 0 176288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1667941163
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1667941163
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1667941163
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1667941163
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1667941163
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1667941163
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1667941163
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1667941163
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1667941163
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1667941163
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1667941163
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1667941163
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1667941163
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1667941163
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1667941163
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1667941163
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1667941163
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1667941163
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 148400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 156352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 164304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 172256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 152432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 160384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 168336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 176288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 148400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 156352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 164304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 172256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 152432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 160384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 168336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 176288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 148400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 156352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 164304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 172256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 152432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 160384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 168336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 176288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1667941163
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1667941163
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1667941163
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1667941163
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1667941163
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1667941163
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1667941163
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1667941163
transform 1 0 148400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1667941163
transform 1 0 156352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1667941163
transform 1 0 164304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1667941163
transform 1 0 172256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1667941163
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1667941163
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1667941163
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1667941163
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1667941163
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1667941163
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1667941163
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1667941163
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1667941163
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1667941163
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1667941163
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1667941163
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1667941163
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1667941163
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1667941163
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1667941163
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1667941163
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1667941163
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1667941163
transform 1 0 152432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1667941163
transform 1 0 160384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1667941163
transform 1 0 168336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1667941163
transform 1 0 176288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1667941163
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1667941163
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1667941163
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1667941163
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1667941163
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1667941163
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1667941163
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1667941163
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1667941163
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1667941163
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1667941163
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1667941163
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1667941163
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1667941163
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1667941163
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1667941163
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1667941163
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1667941163
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1667941163
transform 1 0 148400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1667941163
transform 1 0 156352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1667941163
transform 1 0 164304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1667941163
transform 1 0 172256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1667941163
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1667941163
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1667941163
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1667941163
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1667941163
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1667941163
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1667941163
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1667941163
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1667941163
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1667941163
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1667941163
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1667941163
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1667941163
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1667941163
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1667941163
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1667941163
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1667941163
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1667941163
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1667941163
transform 1 0 152432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1667941163
transform 1 0 160384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1667941163
transform 1 0 168336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1667941163
transform 1 0 176288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1667941163
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1667941163
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1667941163
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1667941163
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1667941163
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1667941163
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1667941163
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1667941163
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1667941163
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1667941163
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1667941163
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1667941163
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1667941163
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1667941163
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1667941163
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1667941163
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1667941163
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1667941163
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1667941163
transform 1 0 148400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1667941163
transform 1 0 156352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1667941163
transform 1 0 164304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1667941163
transform 1 0 172256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1667941163
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1667941163
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1667941163
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1667941163
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1667941163
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1667941163
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1667941163
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1667941163
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1667941163
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1667941163
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1667941163
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1667941163
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1667941163
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1667941163
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1667941163
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1667941163
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1667941163
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1667941163
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1667941163
transform 1 0 152432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1667941163
transform 1 0 160384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1667941163
transform 1 0 168336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1667941163
transform 1 0 176288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1667941163
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1667941163
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1667941163
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1667941163
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1667941163
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1667941163
transform 1 0 24864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1667941163
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1667941163
transform 1 0 32704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1667941163
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1667941163
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1667941163
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1667941163
transform 1 0 48384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1667941163
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1667941163
transform 1 0 56224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1667941163
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1667941163
transform 1 0 64064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1667941163
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1667941163
transform 1 0 71904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1667941163
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1667941163
transform 1 0 79744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1667941163
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1667941163
transform 1 0 87584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1667941163
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1667941163
transform 1 0 95424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1667941163
transform 1 0 99344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1667941163
transform 1 0 103264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1667941163
transform 1 0 107184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1667941163
transform 1 0 111104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1667941163
transform 1 0 115024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1667941163
transform 1 0 118944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1667941163
transform 1 0 122864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1667941163
transform 1 0 126784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1667941163
transform 1 0 130704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1667941163
transform 1 0 134624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1667941163
transform 1 0 138544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1667941163
transform 1 0 142464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1667941163
transform 1 0 146384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1667941163
transform 1 0 150304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1667941163
transform 1 0 154224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1667941163
transform 1 0 158144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1667941163
transform 1 0 162064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1667941163
transform 1 0 165984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1667941163
transform 1 0 169904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1667941163
transform 1 0 173824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1667941163
transform 1 0 177744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _030_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 61936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _031_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 79520 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _032_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 82880 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _033_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 55888 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _034_
timestamp 1667941163
transform 1 0 25200 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _035_
timestamp 1667941163
transform -1 0 12768 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _036_
timestamp 1667941163
transform 1 0 72464 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _037_
timestamp 1667941163
transform 1 0 91840 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _038_
timestamp 1667941163
transform 1 0 107520 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _039_
timestamp 1667941163
transform 1 0 127344 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _040_
timestamp 1667941163
transform 1 0 150864 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _242_
timestamp 1667941163
transform -1 0 120848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _243_
timestamp 1667941163
transform 1 0 119280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout11 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 61936 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout12 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 60480 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout13
timestamp 1667941163
transform 1 0 65968 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout14
timestamp 1667941163
transform 1 0 66304 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 63952 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1667941163
transform -1 0 67760 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1667941163
transform -1 0 69440 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1667941163
transform -1 0 71120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1667941163
transform 1 0 72128 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1667941163
transform 1 0 73808 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1667941163
transform 1 0 76160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1667941163
transform 1 0 77168 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1667941163
transform 1 0 78848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 80528 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[0\].pdn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 113456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[0\].pdn_15 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 114576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[0\].pdp
timestamp 1667941163
transform -1 0 96320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[0\].pdp_16
timestamp 1667941163
transform -1 0 97104 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[1\].pdn_17
timestamp 1667941163
transform -1 0 115248 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[1\].pdn
timestamp 1667941163
transform -1 0 114800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[1\].pdp
timestamp 1667941163
transform -1 0 97552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[1\].pdp_18
timestamp 1667941163
transform -1 0 97776 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[2\].pdn_19
timestamp 1667941163
transform 1 0 114352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[2\].pdn
timestamp 1667941163
transform 1 0 115472 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[2\].pdp
timestamp 1667941163
transform 1 0 98000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[2\].pdp_20
timestamp 1667941163
transform 1 0 95312 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[3\].pdn
timestamp 1667941163
transform -1 0 115024 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[3\].pdn_21
timestamp 1667941163
transform -1 0 116144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[3\].pdp
timestamp 1667941163
transform -1 0 98224 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[3\].pdp_22
timestamp 1667941163
transform 1 0 97776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[4\].pdn
timestamp 1667941163
transform -1 0 112560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[4\].pdn_23
timestamp 1667941163
transform -1 0 113456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[4\].pdp
timestamp 1667941163
transform -1 0 96656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[4\].pdp_24
timestamp 1667941163
transform -1 0 96880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[5\].pdn
timestamp 1667941163
transform -1 0 114128 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[5\].pdn_25
timestamp 1667941163
transform 1 0 113680 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[5\].pdp_26
timestamp 1667941163
transform -1 0 96432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[5\].pdp
timestamp 1667941163
transform -1 0 96208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[6\].pdn
timestamp 1667941163
transform 1 0 113456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[6\].pdn_27
timestamp 1667941163
transform 1 0 112784 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[6\].pdp
timestamp 1667941163
transform -1 0 97328 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[6\].pdp_28
timestamp 1667941163
transform -1 0 99120 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[7\].pdn
timestamp 1667941163
transform -1 0 115472 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[7\].pdn_29
timestamp 1667941163
transform 1 0 115024 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.gen_PD\[7\].pdp
timestamp 1667941163
transform -1 0 95088 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_PD\[7\].pdp_30
timestamp 1667941163
transform -1 0 97552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[0\].pun pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 67984 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[0\].pup
timestamp 1667941163
transform -1 0 58016 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[1\].pun
timestamp 1667941163
transform 1 0 66752 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[1\].pup
timestamp 1667941163
transform -1 0 55888 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[2\].pun
timestamp 1667941163
transform 1 0 67872 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[2\].pup
timestamp 1667941163
transform 1 0 56224 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[3\].pun
timestamp 1667941163
transform 1 0 70000 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[3\].pup
timestamp 1667941163
transform 1 0 56112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[4\].pun
timestamp 1667941163
transform -1 0 66528 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[4\].pup
timestamp 1667941163
transform 1 0 57904 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[5\].pun
timestamp 1667941163
transform 1 0 64960 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[5\].pup
timestamp 1667941163
transform 1 0 59696 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[6\].pun
timestamp 1667941163
transform 1 0 64176 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[6\].pup
timestamp 1667941163
transform -1 0 59808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[7\].pun
timestamp 1667941163
transform 1 0 66080 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[7\].pup
timestamp 1667941163
transform -1 0 59808 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[8\].pun
timestamp 1667941163
transform 1 0 65184 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[8\].pup
timestamp 1667941163
transform -1 0 58464 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[9\].pun
timestamp 1667941163
transform 1 0 63392 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[9\].pup
timestamp 1667941163
transform 1 0 61264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[10\].pun
timestamp 1667941163
transform 1 0 69104 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[10\].pup
timestamp 1667941163
transform 1 0 57008 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[11\].pun
timestamp 1667941163
transform 1 0 64512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[11\].pup
timestamp 1667941163
transform 1 0 57344 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[12\].pun
timestamp 1667941163
transform 1 0 64176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[12\].pup
timestamp 1667941163
transform 1 0 58800 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[13\].pun
timestamp 1667941163
transform 1 0 64288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[13\].pup
timestamp 1667941163
transform 1 0 56224 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[14\].pun
timestamp 1667941163
transform 1 0 65856 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[14\].pup
timestamp 1667941163
transform 1 0 57456 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[15\].pun
timestamp 1667941163
transform 1 0 63280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[15\].pup
timestamp 1667941163
transform 1 0 58352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[16\].pun
timestamp 1667941163
transform 1 0 66976 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[16\].pup
timestamp 1667941163
transform -1 0 58912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[17\].pun
timestamp 1667941163
transform 1 0 66080 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[17\].pup
timestamp 1667941163
transform 1 0 58128 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[18\].pun
timestamp 1667941163
transform 1 0 65408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_inj.gen_PU\[18\].pup
timestamp 1667941163
transform 1 0 58240 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[0\].ntrimn_31
timestamp 1667941163
transform -1 0 107968 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ntrimn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 105840 0 1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[0\].ntrimp_32
timestamp 1667941163
transform -1 0 108416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ntrimp
timestamp 1667941163
transform 1 0 105616 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ptrimn
timestamp 1667941163
transform 1 0 49392 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[0\].ptrimp
timestamp 1667941163
transform -1 0 50176 0 1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[1\].ntrimn_33
timestamp 1667941163
transform -1 0 121296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ntrimn
timestamp 1667941163
transform 1 0 118720 0 1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[1\].ntrimp_34
timestamp 1667941163
transform -1 0 121408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ntrimp
timestamp 1667941163
transform 1 0 118608 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ptrimn
timestamp 1667941163
transform 1 0 33376 0 1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[1\].ptrimp
timestamp 1667941163
transform 1 0 34272 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[2\].ntrimn_35
timestamp 1667941163
transform -1 0 133728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ntrimn
timestamp 1667941163
transform 1 0 131040 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ntrimp
timestamp 1667941163
transform 1 0 130480 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[2\].ntrimp_36
timestamp 1667941163
transform -1 0 133056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ptrimn
timestamp 1667941163
transform 1 0 31136 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[2\].ptrimp
timestamp 1667941163
transform 1 0 33936 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[3\].ntrimn_37
timestamp 1667941163
transform -1 0 141568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ntrimn
timestamp 1667941163
transform 1 0 138992 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.gen_TRIM\[3\].ntrimp_38
timestamp 1667941163
transform -1 0 141680 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ntrimp
timestamp 1667941163
transform 1 0 139440 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ptrimn
timestamp 1667941163
transform 1 0 84784 0 1 3136
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  u_inj.gen_TRIM\[3\].ptrimp
timestamp 1667941163
transform 1 0 84896 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.nsijn
timestamp 1667941163
transform -1 0 86128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.nsijp
timestamp 1667941163
transform -1 0 92624 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_inj.nsijp_214 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 93520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.psijn
timestamp 1667941163
transform 1 0 92848 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_inj.psijn_215
timestamp 1667941163
transform 1 0 92176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_inj.psijp
timestamp 1667941163
transform 1 0 86352 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  u_inj.siginv pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 79296 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_inj.siginv_39
timestamp 1667941163
transform -1 0 79296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_40
timestamp 1667941163
transform 1 0 65296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_41
timestamp 1667941163
transform -1 0 67872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_42
timestamp 1667941163
transform -1 0 70112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_43
timestamp 1667941163
transform -1 0 71456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_44
timestamp 1667941163
transform 1 0 71344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_45
timestamp 1667941163
transform -1 0 75152 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_46
timestamp 1667941163
transform -1 0 76496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_47
timestamp 1667941163
transform -1 0 78512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_48
timestamp 1667941163
transform -1 0 79968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_49
timestamp 1667941163
transform -1 0 82096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_50
timestamp 1667941163
transform -1 0 83216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_51
timestamp 1667941163
transform 1 0 84112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_52
timestamp 1667941163
transform -1 0 87360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_53
timestamp 1667941163
transform -1 0 88368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_54
timestamp 1667941163
transform -1 0 89936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_55
timestamp 1667941163
transform -1 0 91392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_56
timestamp 1667941163
transform -1 0 93968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_57
timestamp 1667941163
transform -1 0 94976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_58
timestamp 1667941163
transform -1 0 97552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_59
timestamp 1667941163
transform -1 0 98336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_60
timestamp 1667941163
transform -1 0 100128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_61
timestamp 1667941163
transform -1 0 101696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_62
timestamp 1667941163
transform -1 0 104048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_63
timestamp 1667941163
transform -1 0 105056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_64
timestamp 1667941163
transform -1 0 106736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_65
timestamp 1667941163
transform -1 0 108416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_66
timestamp 1667941163
transform -1 0 110096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_67
timestamp 1667941163
transform -1 0 111888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_68
timestamp 1667941163
transform -1 0 113456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_69
timestamp 1667941163
transform -1 0 115808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_70
timestamp 1667941163
transform -1 0 116816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_71
timestamp 1667941163
transform -1 0 118496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_72
timestamp 1667941163
transform -1 0 123648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_73
timestamp 1667941163
transform -1 0 125216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_74
timestamp 1667941163
transform -1 0 126672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_75
timestamp 1667941163
transform -1 0 129360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_76
timestamp 1667941163
transform -1 0 130256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_77
timestamp 1667941163
transform -1 0 133616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_78
timestamp 1667941163
transform -1 0 134288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_79
timestamp 1667941163
transform -1 0 135408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_80
timestamp 1667941163
transform -1 0 136976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_81
timestamp 1667941163
transform -1 0 138432 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_82
timestamp 1667941163
transform -1 0 142016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_83
timestamp 1667941163
transform -1 0 142240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_84
timestamp 1667941163
transform -1 0 143696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_85
timestamp 1667941163
transform -1 0 145376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_86
timestamp 1667941163
transform -1 0 147168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_87
timestamp 1667941163
transform -1 0 148736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_88
timestamp 1667941163
transform -1 0 150192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_89
timestamp 1667941163
transform -1 0 152096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_90
timestamp 1667941163
transform -1 0 153776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_91
timestamp 1667941163
transform -1 0 155456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_92
timestamp 1667941163
transform -1 0 157136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_93
timestamp 1667941163
transform -1 0 158928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_94
timestamp 1667941163
transform -1 0 160496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_95
timestamp 1667941163
transform -1 0 162848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_96
timestamp 1667941163
transform -1 0 163856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_97
timestamp 1667941163
transform -1 0 165536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_98
timestamp 1667941163
transform -1 0 167216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_99
timestamp 1667941163
transform -1 0 168896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_100
timestamp 1667941163
transform -1 0 170688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_101
timestamp 1667941163
transform -1 0 172256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_102
timestamp 1667941163
transform -1 0 173376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_103
timestamp 1667941163
transform -1 0 174608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_104
timestamp 1667941163
transform -1 0 175280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_105
timestamp 1667941163
transform -1 0 5040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_106
timestamp 1667941163
transform -1 0 9968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_107
timestamp 1667941163
transform -1 0 14448 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_108
timestamp 1667941163
transform -1 0 19152 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_109
timestamp 1667941163
transform -1 0 23856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_110
timestamp 1667941163
transform -1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_111
timestamp 1667941163
transform -1 0 33488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_112
timestamp 1667941163
transform -1 0 37968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_113
timestamp 1667941163
transform -1 0 42672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_114
timestamp 1667941163
transform -1 0 47376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_115
timestamp 1667941163
transform -1 0 52080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_116
timestamp 1667941163
transform -1 0 57008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_117
timestamp 1667941163
transform -1 0 61488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_118
timestamp 1667941163
transform -1 0 66192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_119
timestamp 1667941163
transform -1 0 70896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_120
timestamp 1667941163
transform -1 0 75600 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_121
timestamp 1667941163
transform -1 0 80528 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_122
timestamp 1667941163
transform -1 0 85008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_123
timestamp 1667941163
transform -1 0 89712 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_124
timestamp 1667941163
transform -1 0 94416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_125
timestamp 1667941163
transform -1 0 99120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_126
timestamp 1667941163
transform -1 0 104048 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_127
timestamp 1667941163
transform -1 0 108528 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_128
timestamp 1667941163
transform -1 0 113232 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_129
timestamp 1667941163
transform -1 0 117936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_130
timestamp 1667941163
transform -1 0 122640 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_131
timestamp 1667941163
transform -1 0 127568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_132
timestamp 1667941163
transform -1 0 132048 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_133
timestamp 1667941163
transform -1 0 136752 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_134
timestamp 1667941163
transform -1 0 141456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_135
timestamp 1667941163
transform -1 0 146160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_136
timestamp 1667941163
transform -1 0 151088 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_137
timestamp 1667941163
transform -1 0 155568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_138
timestamp 1667941163
transform -1 0 160272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_139
timestamp 1667941163
transform -1 0 164976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_140
timestamp 1667941163
transform -1 0 169680 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_141
timestamp 1667941163
transform -1 0 174608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_142
timestamp 1667941163
transform 1 0 177856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_143
timestamp 1667941163
transform -1 0 3472 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_144
timestamp 1667941163
transform -1 0 8176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_145
timestamp 1667941163
transform -1 0 12880 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_146
timestamp 1667941163
transform -1 0 17808 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_147
timestamp 1667941163
transform -1 0 22288 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_148
timestamp 1667941163
transform -1 0 26992 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_149
timestamp 1667941163
transform -1 0 31696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_150
timestamp 1667941163
transform -1 0 36400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_151
timestamp 1667941163
transform -1 0 41328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_152
timestamp 1667941163
transform -1 0 45808 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_153
timestamp 1667941163
transform -1 0 50512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_154
timestamp 1667941163
transform -1 0 55216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_155
timestamp 1667941163
transform -1 0 59920 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_156
timestamp 1667941163
transform -1 0 64848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_157
timestamp 1667941163
transform -1 0 69328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_158
timestamp 1667941163
transform -1 0 74032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_159
timestamp 1667941163
transform -1 0 78736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_160
timestamp 1667941163
transform -1 0 83440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_161
timestamp 1667941163
transform -1 0 88368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_162
timestamp 1667941163
transform -1 0 92848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_163
timestamp 1667941163
transform -1 0 97552 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_164
timestamp 1667941163
transform -1 0 102256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_165
timestamp 1667941163
transform -1 0 106960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_166
timestamp 1667941163
transform -1 0 111888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_167
timestamp 1667941163
transform -1 0 116368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_168
timestamp 1667941163
transform -1 0 121072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_169
timestamp 1667941163
transform -1 0 125776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_170
timestamp 1667941163
transform -1 0 130480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_171
timestamp 1667941163
transform -1 0 135408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_172
timestamp 1667941163
transform -1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_173
timestamp 1667941163
transform -1 0 144592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_174
timestamp 1667941163
transform -1 0 149296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_175
timestamp 1667941163
transform -1 0 154000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_176
timestamp 1667941163
transform -1 0 158928 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_177
timestamp 1667941163
transform -1 0 163408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_178
timestamp 1667941163
transform -1 0 168112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_179
timestamp 1667941163
transform -1 0 172816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_180
timestamp 1667941163
transform -1 0 177520 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_181
timestamp 1667941163
transform -1 0 7616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_182
timestamp 1667941163
transform -1 0 10976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_183
timestamp 1667941163
transform -1 0 13888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_184
timestamp 1667941163
transform -1 0 15456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_185
timestamp 1667941163
transform -1 0 17808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_186
timestamp 1667941163
transform -1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_187
timestamp 1667941163
transform -1 0 21728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_188
timestamp 1667941163
transform -1 0 23296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_189
timestamp 1667941163
transform -1 0 24752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_190
timestamp 1667941163
transform -1 0 26656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_191
timestamp 1667941163
transform -1 0 28336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_192
timestamp 1667941163
transform -1 0 30016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_193
timestamp 1667941163
transform -1 0 31696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_194
timestamp 1667941163
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_195
timestamp 1667941163
transform -1 0 36512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_196
timestamp 1667941163
transform -1 0 37408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_197
timestamp 1667941163
transform -1 0 38416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_198
timestamp 1667941163
transform -1 0 40096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_199
timestamp 1667941163
transform -1 0 41776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_200
timestamp 1667941163
transform -1 0 43456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_201
timestamp 1667941163
transform -1 0 45248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_202
timestamp 1667941163
transform -1 0 46816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_203
timestamp 1667941163
transform -1 0 49168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_204
timestamp 1667941163
transform -1 0 50176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_205
timestamp 1667941163
transform -1 0 51856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_206
timestamp 1667941163
transform -1 0 53536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_207
timestamp 1667941163
transform -1 0 55216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_208
timestamp 1667941163
transform -1 0 57008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_209
timestamp 1667941163
transform 1 0 57456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_210
timestamp 1667941163
transform -1 0 60928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_211
timestamp 1667941163
transform -1 0 61712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_212
timestamp 1667941163
transform 1 0 62608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_213
timestamp 1667941163
transform 1 0 62608 0 1 3136
box -86 -86 534 870
<< labels >>
flabel metal2 s 1344 19200 1456 20000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 48384 19200 48496 20000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 53088 19200 53200 20000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 57792 19200 57904 20000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 62496 19200 62608 20000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 67200 19200 67312 20000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 71904 19200 72016 20000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 76608 19200 76720 20000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 81312 19200 81424 20000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 86016 19200 86128 20000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 90720 19200 90832 20000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 6048 19200 6160 20000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 95424 19200 95536 20000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 100128 19200 100240 20000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 104832 19200 104944 20000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 109536 19200 109648 20000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 114240 19200 114352 20000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 118944 19200 119056 20000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 123648 19200 123760 20000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 128352 19200 128464 20000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 133056 19200 133168 20000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 137760 19200 137872 20000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 10752 19200 10864 20000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 142464 19200 142576 20000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 147168 19200 147280 20000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 151872 19200 151984 20000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 156576 19200 156688 20000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 161280 19200 161392 20000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 165984 19200 166096 20000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 170688 19200 170800 20000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 175392 19200 175504 20000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 15456 19200 15568 20000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 20160 19200 20272 20000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 24864 19200 24976 20000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 29568 19200 29680 20000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 34272 19200 34384 20000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 38976 19200 39088 20000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 43680 19200 43792 20000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 2912 19200 3024 20000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 49952 19200 50064 20000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 54656 19200 54768 20000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 59360 19200 59472 20000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 64064 19200 64176 20000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 68768 19200 68880 20000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 73472 19200 73584 20000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 78176 19200 78288 20000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 82880 19200 82992 20000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 87584 19200 87696 20000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 92288 19200 92400 20000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 7616 19200 7728 20000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 96992 19200 97104 20000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 101696 19200 101808 20000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 106400 19200 106512 20000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 111104 19200 111216 20000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 115808 19200 115920 20000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 120512 19200 120624 20000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 125216 19200 125328 20000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 129920 19200 130032 20000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 134624 19200 134736 20000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 139328 19200 139440 20000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 12320 19200 12432 20000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 144032 19200 144144 20000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 148736 19200 148848 20000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 153440 19200 153552 20000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 158144 19200 158256 20000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 162848 19200 162960 20000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 167552 19200 167664 20000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 172256 19200 172368 20000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 176960 19200 177072 20000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 17024 19200 17136 20000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 21728 19200 21840 20000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 26432 19200 26544 20000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 31136 19200 31248 20000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 35840 19200 35952 20000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 40544 19200 40656 20000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 45248 19200 45360 20000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4480 19200 4592 20000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 51520 19200 51632 20000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 56224 19200 56336 20000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 60928 19200 61040 20000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 65632 19200 65744 20000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 70336 19200 70448 20000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 75040 19200 75152 20000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 79744 19200 79856 20000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 84448 19200 84560 20000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 89152 19200 89264 20000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 93856 19200 93968 20000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 9184 19200 9296 20000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 98560 19200 98672 20000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 103264 19200 103376 20000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 107968 19200 108080 20000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 112672 19200 112784 20000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 117376 19200 117488 20000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 122080 19200 122192 20000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 126784 19200 126896 20000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 131488 19200 131600 20000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 136192 19200 136304 20000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 140896 19200 141008 20000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 13888 19200 14000 20000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 145600 19200 145712 20000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 150304 19200 150416 20000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 155008 19200 155120 20000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 159712 19200 159824 20000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 164416 19200 164528 20000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 169120 19200 169232 20000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 173824 19200 173936 20000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 178528 19200 178640 20000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 18592 19200 18704 20000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 23296 19200 23408 20000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 28000 19200 28112 20000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 32704 19200 32816 20000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 37408 19200 37520 20000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 42112 19200 42224 20000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 46816 19200 46928 20000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 172816 0 172928 800 0 FreeSans 448 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 173376 0 173488 800 0 FreeSans 448 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 173936 0 174048 800 0 FreeSans 448 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 65296 0 65408 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 82096 0 82208 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 118 nsew signal input
flabel metal2 s 83776 0 83888 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 119 nsew signal input
flabel metal2 s 85456 0 85568 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 120 nsew signal input
flabel metal2 s 87136 0 87248 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 121 nsew signal input
flabel metal2 s 88816 0 88928 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 122 nsew signal input
flabel metal2 s 90496 0 90608 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 123 nsew signal input
flabel metal2 s 92176 0 92288 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 124 nsew signal input
flabel metal2 s 93856 0 93968 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 125 nsew signal input
flabel metal2 s 95536 0 95648 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 126 nsew signal input
flabel metal2 s 97216 0 97328 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 127 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 128 nsew signal input
flabel metal2 s 98896 0 99008 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 129 nsew signal input
flabel metal2 s 100576 0 100688 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 130 nsew signal input
flabel metal2 s 102256 0 102368 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 131 nsew signal input
flabel metal2 s 103936 0 104048 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 132 nsew signal input
flabel metal2 s 105616 0 105728 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 133 nsew signal input
flabel metal2 s 107296 0 107408 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 134 nsew signal input
flabel metal2 s 108976 0 109088 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 135 nsew signal input
flabel metal2 s 110656 0 110768 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 136 nsew signal input
flabel metal2 s 112336 0 112448 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 137 nsew signal input
flabel metal2 s 114016 0 114128 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 138 nsew signal input
flabel metal2 s 68656 0 68768 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 139 nsew signal input
flabel metal2 s 115696 0 115808 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 140 nsew signal input
flabel metal2 s 117376 0 117488 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 141 nsew signal input
flabel metal2 s 119056 0 119168 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 142 nsew signal input
flabel metal2 s 120736 0 120848 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 143 nsew signal input
flabel metal2 s 122416 0 122528 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 144 nsew signal input
flabel metal2 s 124096 0 124208 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 145 nsew signal input
flabel metal2 s 125776 0 125888 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 146 nsew signal input
flabel metal2 s 127456 0 127568 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 147 nsew signal input
flabel metal2 s 129136 0 129248 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 148 nsew signal input
flabel metal2 s 130816 0 130928 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 149 nsew signal input
flabel metal2 s 70336 0 70448 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 150 nsew signal input
flabel metal2 s 132496 0 132608 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 151 nsew signal input
flabel metal2 s 134176 0 134288 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 152 nsew signal input
flabel metal2 s 135856 0 135968 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 153 nsew signal input
flabel metal2 s 137536 0 137648 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 154 nsew signal input
flabel metal2 s 139216 0 139328 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 155 nsew signal input
flabel metal2 s 140896 0 141008 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 156 nsew signal input
flabel metal2 s 142576 0 142688 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 157 nsew signal input
flabel metal2 s 144256 0 144368 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 158 nsew signal input
flabel metal2 s 145936 0 146048 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 159 nsew signal input
flabel metal2 s 147616 0 147728 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 160 nsew signal input
flabel metal2 s 72016 0 72128 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 161 nsew signal input
flabel metal2 s 149296 0 149408 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 162 nsew signal input
flabel metal2 s 150976 0 151088 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 163 nsew signal input
flabel metal2 s 152656 0 152768 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 164 nsew signal input
flabel metal2 s 154336 0 154448 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 165 nsew signal input
flabel metal2 s 156016 0 156128 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 166 nsew signal input
flabel metal2 s 157696 0 157808 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 167 nsew signal input
flabel metal2 s 159376 0 159488 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 168 nsew signal input
flabel metal2 s 161056 0 161168 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 169 nsew signal input
flabel metal2 s 162736 0 162848 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 170 nsew signal input
flabel metal2 s 164416 0 164528 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 171 nsew signal input
flabel metal2 s 73696 0 73808 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 172 nsew signal input
flabel metal2 s 166096 0 166208 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 173 nsew signal input
flabel metal2 s 167776 0 167888 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 174 nsew signal input
flabel metal2 s 169456 0 169568 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 175 nsew signal input
flabel metal2 s 171136 0 171248 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 176 nsew signal input
flabel metal2 s 75376 0 75488 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 177 nsew signal input
flabel metal2 s 77056 0 77168 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 178 nsew signal input
flabel metal2 s 78736 0 78848 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 179 nsew signal input
flabel metal2 s 80416 0 80528 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 180 nsew signal input
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_out[0]
port 181 nsew signal tristate
flabel metal2 s 82656 0 82768 800 0 FreeSans 448 90 0 0 la_data_out[10]
port 182 nsew signal tristate
flabel metal2 s 84336 0 84448 800 0 FreeSans 448 90 0 0 la_data_out[11]
port 183 nsew signal tristate
flabel metal2 s 86016 0 86128 800 0 FreeSans 448 90 0 0 la_data_out[12]
port 184 nsew signal tristate
flabel metal2 s 87696 0 87808 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 185 nsew signal tristate
flabel metal2 s 89376 0 89488 800 0 FreeSans 448 90 0 0 la_data_out[14]
port 186 nsew signal tristate
flabel metal2 s 91056 0 91168 800 0 FreeSans 448 90 0 0 la_data_out[15]
port 187 nsew signal tristate
flabel metal2 s 92736 0 92848 800 0 FreeSans 448 90 0 0 la_data_out[16]
port 188 nsew signal tristate
flabel metal2 s 94416 0 94528 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 189 nsew signal tristate
flabel metal2 s 96096 0 96208 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 190 nsew signal tristate
flabel metal2 s 97776 0 97888 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 191 nsew signal tristate
flabel metal2 s 67536 0 67648 800 0 FreeSans 448 90 0 0 la_data_out[1]
port 192 nsew signal tristate
flabel metal2 s 99456 0 99568 800 0 FreeSans 448 90 0 0 la_data_out[20]
port 193 nsew signal tristate
flabel metal2 s 101136 0 101248 800 0 FreeSans 448 90 0 0 la_data_out[21]
port 194 nsew signal tristate
flabel metal2 s 102816 0 102928 800 0 FreeSans 448 90 0 0 la_data_out[22]
port 195 nsew signal tristate
flabel metal2 s 104496 0 104608 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 196 nsew signal tristate
flabel metal2 s 106176 0 106288 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 197 nsew signal tristate
flabel metal2 s 107856 0 107968 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 198 nsew signal tristate
flabel metal2 s 109536 0 109648 800 0 FreeSans 448 90 0 0 la_data_out[26]
port 199 nsew signal tristate
flabel metal2 s 111216 0 111328 800 0 FreeSans 448 90 0 0 la_data_out[27]
port 200 nsew signal tristate
flabel metal2 s 112896 0 113008 800 0 FreeSans 448 90 0 0 la_data_out[28]
port 201 nsew signal tristate
flabel metal2 s 114576 0 114688 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 202 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_out[2]
port 203 nsew signal tristate
flabel metal2 s 116256 0 116368 800 0 FreeSans 448 90 0 0 la_data_out[30]
port 204 nsew signal tristate
flabel metal2 s 117936 0 118048 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 205 nsew signal tristate
flabel metal2 s 119616 0 119728 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 206 nsew signal tristate
flabel metal2 s 121296 0 121408 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 207 nsew signal tristate
flabel metal2 s 122976 0 123088 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 208 nsew signal tristate
flabel metal2 s 124656 0 124768 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 209 nsew signal tristate
flabel metal2 s 126336 0 126448 800 0 FreeSans 448 90 0 0 la_data_out[36]
port 210 nsew signal tristate
flabel metal2 s 128016 0 128128 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 211 nsew signal tristate
flabel metal2 s 129696 0 129808 800 0 FreeSans 448 90 0 0 la_data_out[38]
port 212 nsew signal tristate
flabel metal2 s 131376 0 131488 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 213 nsew signal tristate
flabel metal2 s 70896 0 71008 800 0 FreeSans 448 90 0 0 la_data_out[3]
port 214 nsew signal tristate
flabel metal2 s 133056 0 133168 800 0 FreeSans 448 90 0 0 la_data_out[40]
port 215 nsew signal tristate
flabel metal2 s 134736 0 134848 800 0 FreeSans 448 90 0 0 la_data_out[41]
port 216 nsew signal tristate
flabel metal2 s 136416 0 136528 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 217 nsew signal tristate
flabel metal2 s 138096 0 138208 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 218 nsew signal tristate
flabel metal2 s 139776 0 139888 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 219 nsew signal tristate
flabel metal2 s 141456 0 141568 800 0 FreeSans 448 90 0 0 la_data_out[45]
port 220 nsew signal tristate
flabel metal2 s 143136 0 143248 800 0 FreeSans 448 90 0 0 la_data_out[46]
port 221 nsew signal tristate
flabel metal2 s 144816 0 144928 800 0 FreeSans 448 90 0 0 la_data_out[47]
port 222 nsew signal tristate
flabel metal2 s 146496 0 146608 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 223 nsew signal tristate
flabel metal2 s 148176 0 148288 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 224 nsew signal tristate
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_out[4]
port 225 nsew signal tristate
flabel metal2 s 149856 0 149968 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 226 nsew signal tristate
flabel metal2 s 151536 0 151648 800 0 FreeSans 448 90 0 0 la_data_out[51]
port 227 nsew signal tristate
flabel metal2 s 153216 0 153328 800 0 FreeSans 448 90 0 0 la_data_out[52]
port 228 nsew signal tristate
flabel metal2 s 154896 0 155008 800 0 FreeSans 448 90 0 0 la_data_out[53]
port 229 nsew signal tristate
flabel metal2 s 156576 0 156688 800 0 FreeSans 448 90 0 0 la_data_out[54]
port 230 nsew signal tristate
flabel metal2 s 158256 0 158368 800 0 FreeSans 448 90 0 0 la_data_out[55]
port 231 nsew signal tristate
flabel metal2 s 159936 0 160048 800 0 FreeSans 448 90 0 0 la_data_out[56]
port 232 nsew signal tristate
flabel metal2 s 161616 0 161728 800 0 FreeSans 448 90 0 0 la_data_out[57]
port 233 nsew signal tristate
flabel metal2 s 163296 0 163408 800 0 FreeSans 448 90 0 0 la_data_out[58]
port 234 nsew signal tristate
flabel metal2 s 164976 0 165088 800 0 FreeSans 448 90 0 0 la_data_out[59]
port 235 nsew signal tristate
flabel metal2 s 74256 0 74368 800 0 FreeSans 448 90 0 0 la_data_out[5]
port 236 nsew signal tristate
flabel metal2 s 166656 0 166768 800 0 FreeSans 448 90 0 0 la_data_out[60]
port 237 nsew signal tristate
flabel metal2 s 168336 0 168448 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 238 nsew signal tristate
flabel metal2 s 170016 0 170128 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 239 nsew signal tristate
flabel metal2 s 171696 0 171808 800 0 FreeSans 448 90 0 0 la_data_out[63]
port 240 nsew signal tristate
flabel metal2 s 75936 0 76048 800 0 FreeSans 448 90 0 0 la_data_out[6]
port 241 nsew signal tristate
flabel metal2 s 77616 0 77728 800 0 FreeSans 448 90 0 0 la_data_out[7]
port 242 nsew signal tristate
flabel metal2 s 79296 0 79408 800 0 FreeSans 448 90 0 0 la_data_out[8]
port 243 nsew signal tristate
flabel metal2 s 80976 0 81088 800 0 FreeSans 448 90 0 0 la_data_out[9]
port 244 nsew signal tristate
flabel metal2 s 66416 0 66528 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 245 nsew signal input
flabel metal2 s 83216 0 83328 800 0 FreeSans 448 90 0 0 la_oenb[10]
port 246 nsew signal input
flabel metal2 s 84896 0 85008 800 0 FreeSans 448 90 0 0 la_oenb[11]
port 247 nsew signal input
flabel metal2 s 86576 0 86688 800 0 FreeSans 448 90 0 0 la_oenb[12]
port 248 nsew signal input
flabel metal2 s 88256 0 88368 800 0 FreeSans 448 90 0 0 la_oenb[13]
port 249 nsew signal input
flabel metal2 s 89936 0 90048 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 250 nsew signal input
flabel metal2 s 91616 0 91728 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 251 nsew signal input
flabel metal2 s 93296 0 93408 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 252 nsew signal input
flabel metal2 s 94976 0 95088 800 0 FreeSans 448 90 0 0 la_oenb[17]
port 253 nsew signal input
flabel metal2 s 96656 0 96768 800 0 FreeSans 448 90 0 0 la_oenb[18]
port 254 nsew signal input
flabel metal2 s 98336 0 98448 800 0 FreeSans 448 90 0 0 la_oenb[19]
port 255 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 256 nsew signal input
flabel metal2 s 100016 0 100128 800 0 FreeSans 448 90 0 0 la_oenb[20]
port 257 nsew signal input
flabel metal2 s 101696 0 101808 800 0 FreeSans 448 90 0 0 la_oenb[21]
port 258 nsew signal input
flabel metal2 s 103376 0 103488 800 0 FreeSans 448 90 0 0 la_oenb[22]
port 259 nsew signal input
flabel metal2 s 105056 0 105168 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 260 nsew signal input
flabel metal2 s 106736 0 106848 800 0 FreeSans 448 90 0 0 la_oenb[24]
port 261 nsew signal input
flabel metal2 s 108416 0 108528 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 262 nsew signal input
flabel metal2 s 110096 0 110208 800 0 FreeSans 448 90 0 0 la_oenb[26]
port 263 nsew signal input
flabel metal2 s 111776 0 111888 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 264 nsew signal input
flabel metal2 s 113456 0 113568 800 0 FreeSans 448 90 0 0 la_oenb[28]
port 265 nsew signal input
flabel metal2 s 115136 0 115248 800 0 FreeSans 448 90 0 0 la_oenb[29]
port 266 nsew signal input
flabel metal2 s 69776 0 69888 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 267 nsew signal input
flabel metal2 s 116816 0 116928 800 0 FreeSans 448 90 0 0 la_oenb[30]
port 268 nsew signal input
flabel metal2 s 118496 0 118608 800 0 FreeSans 448 90 0 0 la_oenb[31]
port 269 nsew signal input
flabel metal2 s 120176 0 120288 800 0 FreeSans 448 90 0 0 la_oenb[32]
port 270 nsew signal input
flabel metal2 s 121856 0 121968 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 271 nsew signal input
flabel metal2 s 123536 0 123648 800 0 FreeSans 448 90 0 0 la_oenb[34]
port 272 nsew signal input
flabel metal2 s 125216 0 125328 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 273 nsew signal input
flabel metal2 s 126896 0 127008 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 274 nsew signal input
flabel metal2 s 128576 0 128688 800 0 FreeSans 448 90 0 0 la_oenb[37]
port 275 nsew signal input
flabel metal2 s 130256 0 130368 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 276 nsew signal input
flabel metal2 s 131936 0 132048 800 0 FreeSans 448 90 0 0 la_oenb[39]
port 277 nsew signal input
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 278 nsew signal input
flabel metal2 s 133616 0 133728 800 0 FreeSans 448 90 0 0 la_oenb[40]
port 279 nsew signal input
flabel metal2 s 135296 0 135408 800 0 FreeSans 448 90 0 0 la_oenb[41]
port 280 nsew signal input
flabel metal2 s 136976 0 137088 800 0 FreeSans 448 90 0 0 la_oenb[42]
port 281 nsew signal input
flabel metal2 s 138656 0 138768 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 282 nsew signal input
flabel metal2 s 140336 0 140448 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 283 nsew signal input
flabel metal2 s 142016 0 142128 800 0 FreeSans 448 90 0 0 la_oenb[45]
port 284 nsew signal input
flabel metal2 s 143696 0 143808 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 285 nsew signal input
flabel metal2 s 145376 0 145488 800 0 FreeSans 448 90 0 0 la_oenb[47]
port 286 nsew signal input
flabel metal2 s 147056 0 147168 800 0 FreeSans 448 90 0 0 la_oenb[48]
port 287 nsew signal input
flabel metal2 s 148736 0 148848 800 0 FreeSans 448 90 0 0 la_oenb[49]
port 288 nsew signal input
flabel metal2 s 73136 0 73248 800 0 FreeSans 448 90 0 0 la_oenb[4]
port 289 nsew signal input
flabel metal2 s 150416 0 150528 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 290 nsew signal input
flabel metal2 s 152096 0 152208 800 0 FreeSans 448 90 0 0 la_oenb[51]
port 291 nsew signal input
flabel metal2 s 153776 0 153888 800 0 FreeSans 448 90 0 0 la_oenb[52]
port 292 nsew signal input
flabel metal2 s 155456 0 155568 800 0 FreeSans 448 90 0 0 la_oenb[53]
port 293 nsew signal input
flabel metal2 s 157136 0 157248 800 0 FreeSans 448 90 0 0 la_oenb[54]
port 294 nsew signal input
flabel metal2 s 158816 0 158928 800 0 FreeSans 448 90 0 0 la_oenb[55]
port 295 nsew signal input
flabel metal2 s 160496 0 160608 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 296 nsew signal input
flabel metal2 s 162176 0 162288 800 0 FreeSans 448 90 0 0 la_oenb[57]
port 297 nsew signal input
flabel metal2 s 163856 0 163968 800 0 FreeSans 448 90 0 0 la_oenb[58]
port 298 nsew signal input
flabel metal2 s 165536 0 165648 800 0 FreeSans 448 90 0 0 la_oenb[59]
port 299 nsew signal input
flabel metal2 s 74816 0 74928 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 300 nsew signal input
flabel metal2 s 167216 0 167328 800 0 FreeSans 448 90 0 0 la_oenb[60]
port 301 nsew signal input
flabel metal2 s 168896 0 169008 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 302 nsew signal input
flabel metal2 s 170576 0 170688 800 0 FreeSans 448 90 0 0 la_oenb[62]
port 303 nsew signal input
flabel metal2 s 172256 0 172368 800 0 FreeSans 448 90 0 0 la_oenb[63]
port 304 nsew signal input
flabel metal2 s 76496 0 76608 800 0 FreeSans 448 90 0 0 la_oenb[6]
port 305 nsew signal input
flabel metal2 s 78176 0 78288 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 306 nsew signal input
flabel metal2 s 79856 0 79968 800 0 FreeSans 448 90 0 0 la_oenb[8]
port 307 nsew signal input
flabel metal2 s 81536 0 81648 800 0 FreeSans 448 90 0 0 la_oenb[9]
port 308 nsew signal input
flabel metal4 s 23346 3076 23666 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 67670 3076 67990 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 111994 3076 112314 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 156318 3076 156638 16524 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 45508 3076 45828 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 89832 3076 90152 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 134156 3076 134476 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 178480 3076 178800 16524 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 wb_clk_i
port 311 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 wb_rst_i
port 312 nsew signal input
flabel metal2 s 7056 0 7168 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 313 nsew signal tristate
flabel metal2 s 9296 0 9408 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 314 nsew signal input
flabel metal2 s 28336 0 28448 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 315 nsew signal input
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 316 nsew signal input
flabel metal2 s 31696 0 31808 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 317 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 318 nsew signal input
flabel metal2 s 35056 0 35168 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 319 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 320 nsew signal input
flabel metal2 s 38416 0 38528 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 321 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 322 nsew signal input
flabel metal2 s 41776 0 41888 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 323 nsew signal input
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 324 nsew signal input
flabel metal2 s 11536 0 11648 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 325 nsew signal input
flabel metal2 s 45136 0 45248 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 326 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 327 nsew signal input
flabel metal2 s 48496 0 48608 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 328 nsew signal input
flabel metal2 s 50176 0 50288 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 329 nsew signal input
flabel metal2 s 51856 0 51968 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 330 nsew signal input
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 331 nsew signal input
flabel metal2 s 55216 0 55328 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 332 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 333 nsew signal input
flabel metal2 s 58576 0 58688 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 334 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 335 nsew signal input
flabel metal2 s 13776 0 13888 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 336 nsew signal input
flabel metal2 s 61936 0 62048 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 337 nsew signal input
flabel metal2 s 63616 0 63728 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 338 nsew signal input
flabel metal2 s 16016 0 16128 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 339 nsew signal input
flabel metal2 s 18256 0 18368 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 340 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 341 nsew signal input
flabel metal2 s 21616 0 21728 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 342 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 343 nsew signal input
flabel metal2 s 24976 0 25088 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 344 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 345 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 346 nsew signal input
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 347 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 348 nsew signal input
flabel metal2 s 30576 0 30688 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 349 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 350 nsew signal input
flabel metal2 s 33936 0 34048 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 351 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 352 nsew signal input
flabel metal2 s 37296 0 37408 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 353 nsew signal input
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 354 nsew signal input
flabel metal2 s 40656 0 40768 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 355 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 356 nsew signal input
flabel metal2 s 44016 0 44128 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 357 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 358 nsew signal input
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 359 nsew signal input
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 360 nsew signal input
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 361 nsew signal input
flabel metal2 s 50736 0 50848 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 362 nsew signal input
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 363 nsew signal input
flabel metal2 s 54096 0 54208 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 364 nsew signal input
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 365 nsew signal input
flabel metal2 s 57456 0 57568 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 366 nsew signal input
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 367 nsew signal input
flabel metal2 s 60816 0 60928 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 368 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 369 nsew signal input
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 370 nsew signal input
flabel metal2 s 64176 0 64288 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 371 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 372 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 373 nsew signal input
flabel metal2 s 20496 0 20608 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 374 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 375 nsew signal input
flabel metal2 s 23856 0 23968 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 376 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 377 nsew signal input
flabel metal2 s 27216 0 27328 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 378 nsew signal input
flabel metal2 s 10416 0 10528 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 379 nsew signal tristate
flabel metal2 s 29456 0 29568 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 380 nsew signal tristate
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 381 nsew signal tristate
flabel metal2 s 32816 0 32928 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 382 nsew signal tristate
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 383 nsew signal tristate
flabel metal2 s 36176 0 36288 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 384 nsew signal tristate
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 385 nsew signal tristate
flabel metal2 s 39536 0 39648 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 386 nsew signal tristate
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 387 nsew signal tristate
flabel metal2 s 42896 0 43008 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 388 nsew signal tristate
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 389 nsew signal tristate
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 390 nsew signal tristate
flabel metal2 s 46256 0 46368 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 391 nsew signal tristate
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 392 nsew signal tristate
flabel metal2 s 49616 0 49728 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 393 nsew signal tristate
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 394 nsew signal tristate
flabel metal2 s 52976 0 53088 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 395 nsew signal tristate
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 396 nsew signal tristate
flabel metal2 s 56336 0 56448 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 397 nsew signal tristate
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 398 nsew signal tristate
flabel metal2 s 59696 0 59808 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 399 nsew signal tristate
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 400 nsew signal tristate
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 401 nsew signal tristate
flabel metal2 s 63056 0 63168 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 402 nsew signal tristate
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 403 nsew signal tristate
flabel metal2 s 17136 0 17248 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 404 nsew signal tristate
flabel metal2 s 19376 0 19488 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 405 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 406 nsew signal tristate
flabel metal2 s 22736 0 22848 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 407 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 408 nsew signal tristate
flabel metal2 s 26096 0 26208 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 409 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 410 nsew signal tristate
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 411 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 412 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 413 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 414 nsew signal input
flabel metal2 s 8176 0 8288 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 415 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_we_i
port 416 nsew signal input
rlabel metal1 89992 16464 89992 16464 0 vdd
rlabel via1 90072 15680 90072 15680 0 vss
rlabel metal2 66472 3416 66472 3416 0 _000_
rlabel metal2 85960 5040 85960 5040 0 _001_
rlabel metal3 81648 4872 81648 4872 0 _002_
rlabel metal2 63784 3584 63784 3584 0 la_data_in[0]
rlabel metal2 67592 6160 67592 6160 0 la_data_in[1]
rlabel metal2 68936 3528 68936 3528 0 la_data_in[2]
rlabel metal2 70616 3528 70616 3528 0 la_data_in[3]
rlabel metal2 71960 4200 71960 4200 0 la_data_in[4]
rlabel metal2 73640 4200 73640 4200 0 la_data_in[5]
rlabel metal3 75880 3416 75880 3416 0 la_data_in[6]
rlabel metal2 77280 3416 77280 3416 0 la_data_in[7]
rlabel metal2 78792 2086 78792 2086 0 la_data_in[8]
rlabel metal2 80360 3416 80360 3416 0 la_data_in[9]
rlabel metal2 119672 1246 119672 1246 0 la_data_out[32]
rlabel metal2 121352 2086 121352 2086 0 la_data_out[33]
rlabel metal3 62776 3304 62776 3304 0 net1
rlabel metal3 27328 3528 27328 3528 0 net10
rlabel metal2 170072 2030 170072 2030 0 net100
rlabel metal2 171752 2030 171752 2030 0 net101
rlabel metal2 172872 2030 172872 2030 0 net102
rlabel metal2 173432 1246 173432 1246 0 net103
rlabel metal2 173992 2030 173992 2030 0 net104
rlabel metal2 4648 15960 4648 15960 0 net105
rlabel metal2 9688 16800 9688 16800 0 net106
rlabel metal2 14056 15960 14056 15960 0 net107
rlabel metal2 18760 15960 18760 15960 0 net108
rlabel metal2 23408 15960 23408 15960 0 net109
rlabel metal2 59864 4592 59864 4592 0 net11
rlabel metal2 28168 15960 28168 15960 0 net110
rlabel metal2 33208 16800 33208 16800 0 net111
rlabel metal2 37576 15960 37576 15960 0 net112
rlabel metal2 42280 15960 42280 15960 0 net113
rlabel metal2 46984 15960 46984 15960 0 net114
rlabel metal2 51688 15960 51688 15960 0 net115
rlabel metal2 56728 16800 56728 16800 0 net116
rlabel metal2 61096 15960 61096 15960 0 net117
rlabel metal2 65800 15960 65800 15960 0 net118
rlabel metal2 70504 15960 70504 15960 0 net119
rlabel metal2 51576 5488 51576 5488 0 net12
rlabel metal2 75208 15960 75208 15960 0 net120
rlabel metal2 80248 16800 80248 16800 0 net121
rlabel metal2 84616 15960 84616 15960 0 net122
rlabel metal2 89320 15960 89320 15960 0 net123
rlabel metal2 94024 15960 94024 15960 0 net124
rlabel metal2 98728 15960 98728 15960 0 net125
rlabel metal2 103768 16800 103768 16800 0 net126
rlabel metal2 108136 15960 108136 15960 0 net127
rlabel metal2 112840 15960 112840 15960 0 net128
rlabel metal2 117544 15960 117544 15960 0 net129
rlabel metal3 69776 4312 69776 4312 0 net13
rlabel metal2 122248 15960 122248 15960 0 net130
rlabel metal2 127288 16800 127288 16800 0 net131
rlabel metal2 131656 15960 131656 15960 0 net132
rlabel metal2 136360 15960 136360 15960 0 net133
rlabel metal2 141064 15960 141064 15960 0 net134
rlabel metal2 145768 15960 145768 15960 0 net135
rlabel metal2 150808 16800 150808 16800 0 net136
rlabel metal2 155176 15960 155176 15960 0 net137
rlabel metal2 159880 15960 159880 15960 0 net138
rlabel metal2 164584 15960 164584 15960 0 net139
rlabel metal2 60536 5880 60536 5880 0 net14
rlabel metal2 169288 15960 169288 15960 0 net140
rlabel metal2 174328 16800 174328 16800 0 net141
rlabel metal2 178136 16464 178136 16464 0 net142
rlabel metal2 3080 15960 3080 15960 0 net143
rlabel metal2 7784 15960 7784 15960 0 net144
rlabel metal2 12488 15960 12488 15960 0 net145
rlabel metal2 17528 16800 17528 16800 0 net146
rlabel metal2 22008 16296 22008 16296 0 net147
rlabel metal2 26600 15960 26600 15960 0 net148
rlabel metal2 31304 15960 31304 15960 0 net149
rlabel metal3 113288 5096 113288 5096 0 net15
rlabel metal2 36008 15960 36008 15960 0 net150
rlabel metal2 41048 16800 41048 16800 0 net151
rlabel metal2 45528 16296 45528 16296 0 net152
rlabel metal2 50120 15960 50120 15960 0 net153
rlabel metal2 54824 15960 54824 15960 0 net154
rlabel metal2 59528 15960 59528 15960 0 net155
rlabel metal2 64568 16800 64568 16800 0 net156
rlabel metal2 69048 16296 69048 16296 0 net157
rlabel metal2 73640 15960 73640 15960 0 net158
rlabel metal2 78344 15960 78344 15960 0 net159
rlabel metal2 96824 5040 96824 5040 0 net16
rlabel metal2 83048 15960 83048 15960 0 net160
rlabel metal2 88088 16800 88088 16800 0 net161
rlabel metal2 92568 16296 92568 16296 0 net162
rlabel metal2 97160 15960 97160 15960 0 net163
rlabel metal2 101864 15960 101864 15960 0 net164
rlabel metal2 106568 15960 106568 15960 0 net165
rlabel metal2 111608 16800 111608 16800 0 net166
rlabel metal2 116088 16296 116088 16296 0 net167
rlabel metal2 120680 15960 120680 15960 0 net168
rlabel metal2 125384 15960 125384 15960 0 net169
rlabel metal2 114632 4648 114632 4648 0 net17
rlabel metal2 130088 15960 130088 15960 0 net170
rlabel metal2 135128 16800 135128 16800 0 net171
rlabel metal2 139608 16296 139608 16296 0 net172
rlabel metal2 144200 15960 144200 15960 0 net173
rlabel metal2 148904 15960 148904 15960 0 net174
rlabel metal2 153608 15960 153608 15960 0 net175
rlabel metal2 158648 16800 158648 16800 0 net176
rlabel metal2 163128 16296 163128 16296 0 net177
rlabel metal2 167720 15960 167720 15960 0 net178
rlabel metal2 172424 15960 172424 15960 0 net179
rlabel metal2 97440 4984 97440 4984 0 net18
rlabel metal2 177128 15960 177128 15960 0 net180
rlabel metal2 7112 2030 7112 2030 0 net181
rlabel metal2 10472 2590 10472 2590 0 net182
rlabel metal2 12712 2030 12712 2030 0 net183
rlabel metal2 14952 2030 14952 2030 0 net184
rlabel metal2 17192 2030 17192 2030 0 net185
rlabel metal2 19432 2030 19432 2030 0 net186
rlabel metal2 21112 2030 21112 2030 0 net187
rlabel metal2 22792 2030 22792 2030 0 net188
rlabel metal2 24472 2030 24472 2030 0 net189
rlabel metal2 115640 5600 115640 5600 0 net19
rlabel metal2 26152 854 26152 854 0 net190
rlabel metal2 27832 2590 27832 2590 0 net191
rlabel metal2 29512 2030 29512 2030 0 net192
rlabel metal2 31192 2030 31192 2030 0 net193
rlabel metal2 32872 2030 32872 2030 0 net194
rlabel metal2 34552 2030 34552 2030 0 net195
rlabel metal2 36232 1246 36232 1246 0 net196
rlabel metal2 37912 2030 37912 2030 0 net197
rlabel metal2 39592 2030 39592 2030 0 net198
rlabel metal2 41272 2030 41272 2030 0 net199
rlabel metal3 54656 3640 54656 3640 0 net2
rlabel metal3 96880 4984 96880 4984 0 net20
rlabel metal2 42952 2030 42952 2030 0 net200
rlabel metal2 44632 2030 44632 2030 0 net201
rlabel metal2 46312 2030 46312 2030 0 net202
rlabel metal2 47992 2030 47992 2030 0 net203
rlabel metal2 49672 2030 49672 2030 0 net204
rlabel metal2 51352 2030 51352 2030 0 net205
rlabel metal2 53032 2590 53032 2590 0 net206
rlabel metal2 54712 2590 54712 2590 0 net207
rlabel metal2 56392 2030 56392 2030 0 net208
rlabel metal2 58072 2590 58072 2590 0 net209
rlabel metal2 115864 5544 115864 5544 0 net21
rlabel metal2 59752 2030 59752 2030 0 net210
rlabel metal2 61432 2030 61432 2030 0 net211
rlabel metal2 63112 2590 63112 2590 0 net212
rlabel metal2 64792 1190 64792 1190 0 net213
rlabel metal2 92456 5152 92456 5152 0 net214
rlabel metal2 92456 4256 92456 4256 0 net215
rlabel metal2 98056 5208 98056 5208 0 net22
rlabel metal3 112784 4536 112784 4536 0 net23
rlabel metal2 96544 3304 96544 3304 0 net24
rlabel metal2 113960 5208 113960 5208 0 net25
rlabel metal2 96096 4424 96096 4424 0 net26
rlabel metal2 113344 4984 113344 4984 0 net27
rlabel metal3 98000 4872 98000 4872 0 net28
rlabel metal2 115304 5208 115304 5208 0 net29
rlabel metal2 28728 3528 28728 3528 0 net3
rlabel metal3 96096 4536 96096 4536 0 net30
rlabel metal2 107688 5544 107688 5544 0 net31
rlabel metal2 107464 4592 107464 4592 0 net32
rlabel metal3 120792 4984 120792 4984 0 net33
rlabel metal2 120456 4368 120456 4368 0 net34
rlabel metal2 132888 3976 132888 3976 0 net35
rlabel metal2 132552 4312 132552 4312 0 net36
rlabel metal2 141064 4312 141064 4312 0 net37
rlabel metal2 141344 3528 141344 3528 0 net38
rlabel metal2 79072 4536 79072 4536 0 net39
rlabel metal2 70616 3136 70616 3136 0 net4
rlabel metal2 65912 2590 65912 2590 0 net40
rlabel metal2 67592 2030 67592 2030 0 net41
rlabel metal2 69272 1246 69272 1246 0 net42
rlabel metal2 70952 2590 70952 2590 0 net43
rlabel metal2 72632 1190 72632 1190 0 net44
rlabel metal2 74312 2086 74312 2086 0 net45
rlabel metal2 75992 2590 75992 2590 0 net46
rlabel metal2 77672 1246 77672 1246 0 net47
rlabel metal2 79352 1470 79352 1470 0 net48
rlabel metal2 81032 1246 81032 1246 0 net49
rlabel metal2 73416 4032 73416 4032 0 net5
rlabel metal2 82712 2030 82712 2030 0 net50
rlabel metal2 84392 2030 84392 2030 0 net51
rlabel metal2 86072 1246 86072 1246 0 net52
rlabel metal2 87752 2030 87752 2030 0 net53
rlabel metal2 89432 2030 89432 2030 0 net54
rlabel metal2 91112 2030 91112 2030 0 net55
rlabel metal2 92792 2086 92792 2086 0 net56
rlabel metal2 94472 2590 94472 2590 0 net57
rlabel metal2 96152 1246 96152 1246 0 net58
rlabel metal2 97832 2030 97832 2030 0 net59
rlabel metal2 89096 4032 89096 4032 0 net6
rlabel metal2 99512 2030 99512 2030 0 net60
rlabel metal2 101192 2030 101192 2030 0 net61
rlabel metal2 102872 1246 102872 1246 0 net62
rlabel metal2 104552 2030 104552 2030 0 net63
rlabel metal2 106232 2030 106232 2030 0 net64
rlabel metal2 107912 2590 107912 2590 0 net65
rlabel metal2 109592 2590 109592 2590 0 net66
rlabel metal2 111272 2030 111272 2030 0 net67
rlabel metal2 112952 2030 112952 2030 0 net68
rlabel metal2 114632 1246 114632 1246 0 net69
rlabel metal2 105560 3360 105560 3360 0 net7
rlabel metal2 116312 2030 116312 2030 0 net70
rlabel metal2 117992 2030 117992 2030 0 net71
rlabel metal2 123032 2030 123032 2030 0 net72
rlabel metal2 124712 2030 124712 2030 0 net73
rlabel metal2 126392 2030 126392 2030 0 net74
rlabel metal2 128072 2590 128072 2590 0 net75
rlabel metal2 129752 2590 129752 2590 0 net76
rlabel metal2 131432 2030 131432 2030 0 net77
rlabel metal2 133112 1246 133112 1246 0 net78
rlabel metal2 134792 2030 134792 2030 0 net79
rlabel metal2 77672 3080 77672 3080 0 net8
rlabel metal2 136472 2030 136472 2030 0 net80
rlabel metal2 138152 2030 138152 2030 0 net81
rlabel metal2 139832 2030 139832 2030 0 net82
rlabel metal2 141512 854 141512 854 0 net83
rlabel metal2 143192 2030 143192 2030 0 net84
rlabel metal2 144872 2030 144872 2030 0 net85
rlabel metal2 146552 2030 146552 2030 0 net86
rlabel metal2 148232 2030 148232 2030 0 net87
rlabel metal2 149912 2030 149912 2030 0 net88
rlabel metal2 151592 2590 151592 2590 0 net89
rlabel metal2 79352 3136 79352 3136 0 net9
rlabel metal2 153272 2590 153272 2590 0 net90
rlabel metal2 154952 2030 154952 2030 0 net91
rlabel metal2 156632 2030 156632 2030 0 net92
rlabel metal2 158312 2030 158312 2030 0 net93
rlabel metal2 159992 2030 159992 2030 0 net94
rlabel metal2 161672 1246 161672 1246 0 net95
rlabel metal2 163352 2030 163352 2030 0 net96
rlabel metal2 165032 2030 165032 2030 0 net97
rlabel metal2 166712 2030 166712 2030 0 net98
rlabel metal2 168392 2030 168392 2030 0 net99
rlabel metal2 70504 4144 70504 4144 0 u_inj.outn
rlabel metal2 49224 4760 49224 4760 0 u_inj.outp
rlabel metal3 79464 5208 79464 5208 0 u_inj.signal_n
rlabel metal2 105224 3920 105224 3920 0 u_inj.trim_n_r\[0\]
rlabel metal2 118216 3920 118216 3920 0 u_inj.trim_n_r\[1\]
rlabel metal3 130816 3640 130816 3640 0 u_inj.trim_n_r\[2\]
rlabel metal2 142632 3808 142632 3808 0 u_inj.trim_n_r\[3\]
rlabel metal2 49784 3976 49784 3976 0 u_inj.trim_p_r\[0\]
rlabel metal2 33656 4536 33656 4536 0 u_inj.trim_p_r\[1\]
rlabel metal2 30856 3976 30856 3976 0 u_inj.trim_p_r\[2\]
rlabel metal2 83720 3920 83720 3920 0 u_inj.trim_p_r\[3\]
<< properties >>
string FIXED_BBOX 0 0 180000 20000
<< end >>
